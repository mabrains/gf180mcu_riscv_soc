magic
tech gf180mcuD
magscale 1 5
timestamp 1700152632
<< metal1 >>
rect 672 8245 9296 8262
rect 672 8219 1685 8245
rect 1711 8219 1737 8245
rect 1763 8219 1789 8245
rect 1815 8219 3841 8245
rect 3867 8219 3893 8245
rect 3919 8219 3945 8245
rect 3971 8219 5997 8245
rect 6023 8219 6049 8245
rect 6075 8219 6101 8245
rect 6127 8219 8153 8245
rect 8179 8219 8205 8245
rect 8231 8219 8257 8245
rect 8283 8219 9296 8245
rect 672 8202 9296 8219
rect 4663 8161 4689 8167
rect 4663 8129 4689 8135
rect 1079 7993 1105 7999
rect 1079 7961 1105 7967
rect 1303 7993 1329 7999
rect 1303 7961 1329 7967
rect 3151 7993 3177 7999
rect 3151 7961 3177 7967
rect 3487 7993 3513 7999
rect 3487 7961 3513 7967
rect 3823 7993 3849 7999
rect 3823 7961 3849 7967
rect 4383 7993 4409 7999
rect 4383 7961 4409 7967
rect 5503 7993 5529 7999
rect 5503 7961 5529 7967
rect 5839 7993 5865 7999
rect 5839 7961 5865 7967
rect 6847 7993 6873 7999
rect 6847 7961 6873 7967
rect 7183 7993 7209 7999
rect 7183 7961 7209 7967
rect 7519 7993 7545 7999
rect 7519 7961 7545 7967
rect 855 7937 881 7943
rect 855 7905 881 7911
rect 5055 7937 5081 7943
rect 5055 7905 5081 7911
rect 9087 7937 9113 7943
rect 9087 7905 9113 7911
rect 672 7853 9376 7870
rect 672 7827 2763 7853
rect 2789 7827 2815 7853
rect 2841 7827 2867 7853
rect 2893 7827 4919 7853
rect 4945 7827 4971 7853
rect 4997 7827 5023 7853
rect 5049 7827 7075 7853
rect 7101 7827 7127 7853
rect 7153 7827 7179 7853
rect 7205 7827 9231 7853
rect 9257 7827 9283 7853
rect 9309 7827 9335 7853
rect 9361 7827 9376 7853
rect 672 7810 9376 7827
rect 4831 7769 4857 7775
rect 4831 7737 4857 7743
rect 855 7713 881 7719
rect 855 7681 881 7687
rect 9087 7713 9113 7719
rect 9087 7681 9113 7687
rect 672 7461 9296 7478
rect 672 7435 1685 7461
rect 1711 7435 1737 7461
rect 1763 7435 1789 7461
rect 1815 7435 3841 7461
rect 3867 7435 3893 7461
rect 3919 7435 3945 7461
rect 3971 7435 5997 7461
rect 6023 7435 6049 7461
rect 6075 7435 6101 7461
rect 6127 7435 8153 7461
rect 8179 7435 8205 7461
rect 8231 7435 8257 7461
rect 8283 7435 9296 7461
rect 672 7418 9296 7435
rect 855 7153 881 7159
rect 855 7121 881 7127
rect 9087 7153 9113 7159
rect 9087 7121 9113 7127
rect 672 7069 9376 7086
rect 672 7043 2763 7069
rect 2789 7043 2815 7069
rect 2841 7043 2867 7069
rect 2893 7043 4919 7069
rect 4945 7043 4971 7069
rect 4997 7043 5023 7069
rect 5049 7043 7075 7069
rect 7101 7043 7127 7069
rect 7153 7043 7179 7069
rect 7205 7043 9231 7069
rect 9257 7043 9283 7069
rect 9309 7043 9335 7069
rect 9361 7043 9376 7069
rect 672 7026 9376 7043
rect 5553 6847 5559 6873
rect 5585 6847 5591 6873
rect 911 6817 937 6823
rect 911 6785 937 6791
rect 3487 6817 3513 6823
rect 5889 6791 5895 6817
rect 5921 6791 5927 6817
rect 6953 6791 6959 6817
rect 6985 6791 6991 6817
rect 3487 6785 3513 6791
rect 3543 6761 3569 6767
rect 3543 6729 3569 6735
rect 672 6677 9296 6694
rect 672 6651 1685 6677
rect 1711 6651 1737 6677
rect 1763 6651 1789 6677
rect 1815 6651 3841 6677
rect 3867 6651 3893 6677
rect 3919 6651 3945 6677
rect 3971 6651 5997 6677
rect 6023 6651 6049 6677
rect 6075 6651 6101 6677
rect 6127 6651 8153 6677
rect 8179 6651 8205 6677
rect 8231 6651 8257 6677
rect 8283 6651 9296 6677
rect 672 6634 9296 6651
rect 4377 6511 4383 6537
rect 4409 6511 4415 6537
rect 6449 6511 6455 6537
rect 6481 6511 6487 6537
rect 8185 6511 8191 6537
rect 8217 6511 8223 6537
rect 2977 6455 2983 6481
rect 3009 6455 3015 6481
rect 5049 6455 5055 6481
rect 5081 6455 5087 6481
rect 7681 6455 7687 6481
rect 7713 6455 7719 6481
rect 8465 6455 8471 6481
rect 8497 6455 8503 6481
rect 855 6425 881 6431
rect 855 6393 881 6399
rect 1023 6425 1049 6431
rect 3313 6399 3319 6425
rect 3345 6399 3351 6425
rect 5385 6399 5391 6425
rect 5417 6399 5423 6425
rect 9025 6399 9031 6425
rect 9057 6399 9063 6425
rect 1023 6393 1049 6399
rect 1191 6369 1217 6375
rect 1191 6337 1217 6343
rect 672 6285 9376 6302
rect 672 6259 2763 6285
rect 2789 6259 2815 6285
rect 2841 6259 2867 6285
rect 2893 6259 4919 6285
rect 4945 6259 4971 6285
rect 4997 6259 5023 6285
rect 5049 6259 7075 6285
rect 7101 6259 7127 6285
rect 7153 6259 7179 6285
rect 7205 6259 9231 6285
rect 9257 6259 9283 6285
rect 9309 6259 9335 6285
rect 9361 6259 9376 6285
rect 672 6242 9376 6259
rect 3487 6201 3513 6207
rect 3487 6169 3513 6175
rect 3935 6201 3961 6207
rect 3935 6169 3961 6175
rect 3991 6201 4017 6207
rect 3991 6169 4017 6175
rect 4831 6201 4857 6207
rect 4831 6169 4857 6175
rect 5391 6201 5417 6207
rect 5391 6169 5417 6175
rect 855 6145 881 6151
rect 855 6113 881 6119
rect 3711 6145 3737 6151
rect 3711 6113 3737 6119
rect 4103 6145 4129 6151
rect 4103 6113 4129 6119
rect 8919 6145 8945 6151
rect 8919 6113 8945 6119
rect 3431 6089 3457 6095
rect 3431 6057 3457 6063
rect 3543 6089 3569 6095
rect 3543 6057 3569 6063
rect 3879 6089 3905 6095
rect 3879 6057 3905 6063
rect 4775 6089 4801 6095
rect 4775 6057 4801 6063
rect 4943 6089 4969 6095
rect 4943 6057 4969 6063
rect 5279 6089 5305 6095
rect 5279 6057 5305 6063
rect 5503 6089 5529 6095
rect 5503 6057 5529 6063
rect 5615 6089 5641 6095
rect 9087 6089 9113 6095
rect 5889 6063 5895 6089
rect 5921 6063 5927 6089
rect 5615 6057 5641 6063
rect 9087 6057 9113 6063
rect 5111 6033 5137 6039
rect 8807 6033 8833 6039
rect 7009 6007 7015 6033
rect 7041 6007 7047 6033
rect 5111 6001 5137 6007
rect 8807 6001 8833 6007
rect 672 5893 9296 5910
rect 672 5867 1685 5893
rect 1711 5867 1737 5893
rect 1763 5867 1789 5893
rect 1815 5867 3841 5893
rect 3867 5867 3893 5893
rect 3919 5867 3945 5893
rect 3971 5867 5997 5893
rect 6023 5867 6049 5893
rect 6075 5867 6101 5893
rect 6127 5867 8153 5893
rect 8179 5867 8205 5893
rect 8231 5867 8257 5893
rect 8283 5867 9296 5893
rect 672 5850 9296 5867
rect 6225 5783 6231 5809
rect 6257 5783 6263 5809
rect 6791 5753 6817 5759
rect 3537 5727 3543 5753
rect 3569 5727 3575 5753
rect 6791 5721 6817 5727
rect 7239 5753 7265 5759
rect 7239 5721 7265 5727
rect 6119 5697 6145 5703
rect 6735 5697 6761 5703
rect 1465 5671 1471 5697
rect 1497 5671 1503 5697
rect 5777 5671 5783 5697
rect 5809 5671 5815 5697
rect 6337 5671 6343 5697
rect 6369 5671 6375 5697
rect 6119 5665 6145 5671
rect 6735 5665 6761 5671
rect 6847 5697 6873 5703
rect 6847 5665 6873 5671
rect 7295 5697 7321 5703
rect 7295 5665 7321 5671
rect 7463 5697 7489 5703
rect 7463 5665 7489 5671
rect 7687 5697 7713 5703
rect 7687 5665 7713 5671
rect 7743 5697 7769 5703
rect 8465 5671 8471 5697
rect 8497 5671 8503 5697
rect 7743 5665 7769 5671
rect 5951 5641 5977 5647
rect 1017 5615 1023 5641
rect 1049 5615 1055 5641
rect 5951 5609 5977 5615
rect 7183 5641 7209 5647
rect 9025 5615 9031 5641
rect 9057 5615 9063 5641
rect 7183 5609 7209 5615
rect 6343 5585 6369 5591
rect 6343 5553 6369 5559
rect 6959 5585 6985 5591
rect 6959 5553 6985 5559
rect 7631 5585 7657 5591
rect 7631 5553 7657 5559
rect 7855 5585 7881 5591
rect 7855 5553 7881 5559
rect 672 5501 9376 5518
rect 672 5475 2763 5501
rect 2789 5475 2815 5501
rect 2841 5475 2867 5501
rect 2893 5475 4919 5501
rect 4945 5475 4971 5501
rect 4997 5475 5023 5501
rect 5049 5475 7075 5501
rect 7101 5475 7127 5501
rect 7153 5475 7179 5501
rect 7205 5475 9231 5501
rect 9257 5475 9283 5501
rect 9309 5475 9335 5501
rect 9361 5475 9376 5501
rect 672 5458 9376 5475
rect 1023 5361 1049 5367
rect 1023 5329 1049 5335
rect 4439 5361 4465 5367
rect 4439 5329 4465 5335
rect 4551 5361 4577 5367
rect 7911 5361 7937 5367
rect 5945 5335 5951 5361
rect 5977 5335 5983 5361
rect 4551 5329 4577 5335
rect 7911 5329 7937 5335
rect 8919 5361 8945 5367
rect 8919 5329 8945 5335
rect 855 5305 881 5311
rect 4383 5305 4409 5311
rect 9087 5305 9113 5311
rect 4041 5279 4047 5305
rect 4073 5279 4079 5305
rect 5105 5279 5111 5305
rect 5137 5279 5143 5305
rect 855 5273 881 5279
rect 4383 5273 4409 5279
rect 9087 5273 9113 5279
rect 1247 5249 1273 5255
rect 8807 5249 8833 5255
rect 2641 5223 2647 5249
rect 2673 5223 2679 5249
rect 3705 5223 3711 5249
rect 3737 5223 3743 5249
rect 7737 5223 7743 5249
rect 7769 5223 7775 5249
rect 1247 5217 1273 5223
rect 8807 5217 8833 5223
rect 672 5109 9296 5126
rect 672 5083 1685 5109
rect 1711 5083 1737 5109
rect 1763 5083 1789 5109
rect 1815 5083 3841 5109
rect 3867 5083 3893 5109
rect 3919 5083 3945 5109
rect 3971 5083 5997 5109
rect 6023 5083 6049 5109
rect 6075 5083 6101 5109
rect 6127 5083 8153 5109
rect 8179 5083 8205 5109
rect 8231 5083 8257 5109
rect 8283 5083 9296 5109
rect 672 5066 9296 5083
rect 6287 5025 6313 5031
rect 6287 4993 6313 4999
rect 6455 5025 6481 5031
rect 6455 4993 6481 4999
rect 3039 4969 3065 4975
rect 3039 4937 3065 4943
rect 3319 4969 3345 4975
rect 8465 4943 8471 4969
rect 8497 4943 8503 4969
rect 3319 4937 3345 4943
rect 3095 4913 3121 4919
rect 3095 4881 3121 4887
rect 3375 4913 3401 4919
rect 3375 4881 3401 4887
rect 3543 4913 3569 4919
rect 3543 4881 3569 4887
rect 3823 4913 3849 4919
rect 3823 4881 3849 4887
rect 3879 4913 3905 4919
rect 3879 4881 3905 4887
rect 4103 4913 4129 4919
rect 5279 4913 5305 4919
rect 6847 4913 6873 4919
rect 4209 4887 4215 4913
rect 4241 4887 4247 4913
rect 6449 4887 6455 4913
rect 6481 4887 6487 4913
rect 7009 4887 7015 4913
rect 7041 4887 7047 4913
rect 4103 4881 4129 4887
rect 5279 4881 5305 4887
rect 6847 4881 6873 4887
rect 855 4857 881 4863
rect 855 4825 881 4831
rect 3263 4857 3289 4863
rect 5503 4857 5529 4863
rect 8919 4857 8945 4863
rect 4265 4831 4271 4857
rect 4297 4831 4303 4857
rect 7401 4831 7407 4857
rect 7433 4831 7439 4857
rect 3263 4825 3289 4831
rect 5503 4825 5529 4831
rect 8919 4825 8945 4831
rect 9087 4857 9113 4863
rect 9087 4825 9113 4831
rect 1023 4801 1049 4807
rect 1023 4769 1049 4775
rect 1247 4801 1273 4807
rect 1247 4769 1273 4775
rect 3767 4801 3793 4807
rect 6679 4801 6705 4807
rect 4321 4775 4327 4801
rect 4353 4775 4359 4801
rect 3767 4769 3793 4775
rect 6679 4769 6705 4775
rect 6791 4801 6817 4807
rect 6791 4769 6817 4775
rect 8807 4801 8833 4807
rect 8807 4769 8833 4775
rect 672 4717 9376 4734
rect 672 4691 2763 4717
rect 2789 4691 2815 4717
rect 2841 4691 2867 4717
rect 2893 4691 4919 4717
rect 4945 4691 4971 4717
rect 4997 4691 5023 4717
rect 5049 4691 7075 4717
rect 7101 4691 7127 4717
rect 7153 4691 7179 4717
rect 7205 4691 9231 4717
rect 9257 4691 9283 4717
rect 9309 4691 9335 4717
rect 9361 4691 9376 4717
rect 672 4674 9376 4691
rect 7015 4633 7041 4639
rect 7015 4601 7041 4607
rect 1023 4577 1049 4583
rect 3991 4577 4017 4583
rect 2473 4551 2479 4577
rect 2505 4551 2511 4577
rect 2921 4551 2927 4577
rect 2953 4551 2959 4577
rect 5665 4551 5671 4577
rect 5697 4551 5703 4577
rect 6505 4551 6511 4577
rect 6537 4551 6543 4577
rect 6673 4551 6679 4577
rect 6705 4551 6711 4577
rect 8913 4551 8919 4577
rect 8945 4551 8951 4577
rect 1023 4545 1049 4551
rect 3991 4545 4017 4551
rect 855 4521 881 4527
rect 3935 4521 3961 4527
rect 6231 4521 6257 4527
rect 2249 4495 2255 4521
rect 2281 4495 2287 4521
rect 2977 4495 2983 4521
rect 3009 4495 3015 4521
rect 4321 4495 4327 4521
rect 4353 4495 4359 4521
rect 5217 4495 5223 4521
rect 5249 4495 5255 4521
rect 5441 4495 5447 4521
rect 5473 4495 5479 4521
rect 855 4489 881 4495
rect 3935 4489 3961 4495
rect 6231 4489 6257 4495
rect 6959 4521 6985 4527
rect 6959 4489 6985 4495
rect 7127 4521 7153 4527
rect 7127 4489 7153 4495
rect 7183 4521 7209 4527
rect 9087 4521 9113 4527
rect 7345 4495 7351 4521
rect 7377 4495 7383 4521
rect 7183 4489 7209 4495
rect 9087 4489 9113 4495
rect 1247 4465 1273 4471
rect 4439 4465 4465 4471
rect 6175 4465 6201 4471
rect 3817 4439 3823 4465
rect 3849 4439 3855 4465
rect 5497 4439 5503 4465
rect 5529 4439 5535 4465
rect 1247 4433 1273 4439
rect 4439 4433 4465 4439
rect 6175 4433 6201 4439
rect 8807 4465 8833 4471
rect 8807 4433 8833 4439
rect 3991 4409 4017 4415
rect 3991 4377 4017 4383
rect 4495 4409 4521 4415
rect 4495 4377 4521 4383
rect 672 4325 9296 4342
rect 672 4299 1685 4325
rect 1711 4299 1737 4325
rect 1763 4299 1789 4325
rect 1815 4299 3841 4325
rect 3867 4299 3893 4325
rect 3919 4299 3945 4325
rect 3971 4299 5997 4325
rect 6023 4299 6049 4325
rect 6075 4299 6101 4325
rect 6127 4299 8153 4325
rect 8179 4299 8205 4325
rect 8231 4299 8257 4325
rect 8283 4299 9296 4325
rect 672 4282 9296 4299
rect 2255 4241 2281 4247
rect 2255 4209 2281 4215
rect 6735 4241 6761 4247
rect 6735 4209 6761 4215
rect 5833 4159 5839 4185
rect 5865 4159 5871 4185
rect 6897 4159 6903 4185
rect 6929 4159 6935 4185
rect 7015 4129 7041 4135
rect 4321 4103 4327 4129
rect 4353 4103 4359 4129
rect 5329 4103 5335 4129
rect 5361 4103 5367 4129
rect 7015 4097 7041 4103
rect 855 4073 881 4079
rect 855 4041 881 4047
rect 1191 4073 1217 4079
rect 1191 4041 1217 4047
rect 1359 4073 1385 4079
rect 1359 4041 1385 4047
rect 2087 4073 2113 4079
rect 2087 4041 2113 4047
rect 4607 4073 4633 4079
rect 4607 4041 4633 4047
rect 5615 4073 5641 4079
rect 5615 4041 5641 4047
rect 6847 4073 6873 4079
rect 6847 4041 6873 4047
rect 7127 4073 7153 4079
rect 7127 4041 7153 4047
rect 7183 4073 7209 4079
rect 7183 4041 7209 4047
rect 8583 4073 8609 4079
rect 8583 4041 8609 4047
rect 8751 4073 8777 4079
rect 8751 4041 8777 4047
rect 9087 4073 9113 4079
rect 9087 4041 9113 4047
rect 1023 4017 1049 4023
rect 1023 3985 1049 3991
rect 1583 4017 1609 4023
rect 1583 3985 1609 3991
rect 2199 4017 2225 4023
rect 8913 3991 8919 4017
rect 8945 3991 8951 4017
rect 2199 3985 2225 3991
rect 672 3933 9376 3950
rect 672 3907 2763 3933
rect 2789 3907 2815 3933
rect 2841 3907 2867 3933
rect 2893 3907 4919 3933
rect 4945 3907 4971 3933
rect 4997 3907 5023 3933
rect 5049 3907 7075 3933
rect 7101 3907 7127 3933
rect 7153 3907 7179 3933
rect 7205 3907 9231 3933
rect 9257 3907 9283 3933
rect 9309 3907 9335 3933
rect 9361 3907 9376 3933
rect 672 3890 9376 3907
rect 1023 3849 1049 3855
rect 1023 3817 1049 3823
rect 1247 3849 1273 3855
rect 4103 3849 4129 3855
rect 2529 3823 2535 3849
rect 2561 3823 2567 3849
rect 1247 3817 1273 3823
rect 4103 3817 4129 3823
rect 4495 3849 4521 3855
rect 4495 3817 4521 3823
rect 4775 3849 4801 3855
rect 9143 3849 9169 3855
rect 5273 3823 5279 3849
rect 5305 3823 5311 3849
rect 5945 3823 5951 3849
rect 5977 3823 5983 3849
rect 4775 3817 4801 3823
rect 9143 3817 9169 3823
rect 3095 3793 3121 3799
rect 1857 3767 1863 3793
rect 1889 3767 1895 3793
rect 3095 3761 3121 3767
rect 4327 3793 4353 3799
rect 4327 3761 4353 3767
rect 4383 3793 4409 3799
rect 6455 3793 6481 3799
rect 5609 3767 5615 3793
rect 5641 3767 5647 3793
rect 4383 3761 4409 3767
rect 6455 3761 6481 3767
rect 7463 3793 7489 3799
rect 7463 3761 7489 3767
rect 855 3737 881 3743
rect 8863 3737 8889 3743
rect 1801 3711 1807 3737
rect 1833 3711 1839 3737
rect 2809 3711 2815 3737
rect 2841 3711 2847 3737
rect 5553 3711 5559 3737
rect 5585 3711 5591 3737
rect 6673 3711 6679 3737
rect 6705 3711 6711 3737
rect 7793 3711 7799 3737
rect 7825 3711 7831 3737
rect 855 3705 881 3711
rect 8863 3705 8889 3711
rect 1471 3681 1497 3687
rect 1471 3649 1497 3655
rect 4831 3681 4857 3687
rect 4831 3649 4857 3655
rect 3935 3625 3961 3631
rect 3935 3593 3961 3599
rect 4047 3625 4073 3631
rect 4047 3593 4073 3599
rect 4103 3625 4129 3631
rect 4103 3593 4129 3599
rect 672 3541 9296 3558
rect 672 3515 1685 3541
rect 1711 3515 1737 3541
rect 1763 3515 1789 3541
rect 1815 3515 3841 3541
rect 3867 3515 3893 3541
rect 3919 3515 3945 3541
rect 3971 3515 5997 3541
rect 6023 3515 6049 3541
rect 6075 3515 6101 3541
rect 6127 3515 8153 3541
rect 8179 3515 8205 3541
rect 8231 3515 8257 3541
rect 8283 3515 9296 3541
rect 672 3498 9296 3515
rect 4383 3345 4409 3351
rect 3313 3319 3319 3345
rect 3345 3319 3351 3345
rect 4383 3313 4409 3319
rect 855 3289 881 3295
rect 855 3257 881 3263
rect 1023 3289 1049 3295
rect 4663 3289 4689 3295
rect 3369 3263 3375 3289
rect 3401 3263 3407 3289
rect 1023 3257 1049 3263
rect 4663 3257 4689 3263
rect 1247 3233 1273 3239
rect 1247 3201 1273 3207
rect 1471 3233 1497 3239
rect 1471 3201 1497 3207
rect 1695 3233 1721 3239
rect 9087 3233 9113 3239
rect 4209 3207 4215 3233
rect 4241 3207 4247 3233
rect 1695 3201 1721 3207
rect 9087 3201 9113 3207
rect 672 3149 9376 3166
rect 672 3123 2763 3149
rect 2789 3123 2815 3149
rect 2841 3123 2867 3149
rect 2893 3123 4919 3149
rect 4945 3123 4971 3149
rect 4997 3123 5023 3149
rect 5049 3123 7075 3149
rect 7101 3123 7127 3149
rect 7153 3123 7179 3149
rect 7205 3123 9231 3149
rect 9257 3123 9283 3149
rect 9309 3123 9335 3149
rect 9361 3123 9376 3149
rect 672 3106 9376 3123
rect 4377 3039 4383 3065
rect 4409 3039 4415 3065
rect 5889 3039 5895 3065
rect 5921 3039 5927 3065
rect 1023 3009 1049 3015
rect 4159 3009 4185 3015
rect 2585 2983 2591 3009
rect 2617 2983 2623 3009
rect 1023 2977 1049 2983
rect 4159 2977 4185 2983
rect 6399 3009 6425 3015
rect 6399 2977 6425 2983
rect 7407 3009 7433 3015
rect 7407 2977 7433 2983
rect 855 2953 881 2959
rect 855 2921 881 2927
rect 3431 2953 3457 2959
rect 6679 2953 6705 2959
rect 3593 2927 3599 2953
rect 3625 2927 3631 2953
rect 7737 2927 7743 2953
rect 7769 2927 7775 2953
rect 3431 2921 3457 2927
rect 6679 2921 6705 2927
rect 1247 2897 1273 2903
rect 1247 2865 1273 2871
rect 1471 2897 1497 2903
rect 1471 2865 1497 2871
rect 1695 2897 1721 2903
rect 1695 2865 1721 2871
rect 1919 2897 1945 2903
rect 1919 2865 1945 2871
rect 2479 2897 2505 2903
rect 2479 2865 2505 2871
rect 5055 2897 5081 2903
rect 5055 2865 5081 2871
rect 5391 2897 5417 2903
rect 5391 2865 5417 2871
rect 5727 2897 5753 2903
rect 5727 2865 5753 2871
rect 8807 2897 8833 2903
rect 8807 2865 8833 2871
rect 9143 2897 9169 2903
rect 9143 2865 9169 2871
rect 672 2757 9296 2774
rect 672 2731 1685 2757
rect 1711 2731 1737 2757
rect 1763 2731 1789 2757
rect 1815 2731 3841 2757
rect 3867 2731 3893 2757
rect 3919 2731 3945 2757
rect 3971 2731 5997 2757
rect 6023 2731 6049 2757
rect 6075 2731 6101 2757
rect 6127 2731 8153 2757
rect 8179 2731 8205 2757
rect 8231 2731 8257 2757
rect 8283 2731 9296 2757
rect 672 2714 9296 2731
rect 2591 2617 2617 2623
rect 2591 2585 2617 2591
rect 1695 2561 1721 2567
rect 905 2535 911 2561
rect 937 2535 943 2561
rect 1695 2529 1721 2535
rect 3319 2561 3345 2567
rect 3319 2529 3345 2535
rect 3599 2561 3625 2567
rect 3599 2529 3625 2535
rect 3767 2561 3793 2567
rect 3767 2529 3793 2535
rect 4159 2561 4185 2567
rect 4159 2529 4185 2535
rect 5167 2561 5193 2567
rect 5167 2529 5193 2535
rect 6231 2561 6257 2567
rect 6231 2529 6257 2535
rect 7463 2561 7489 2567
rect 7463 2529 7489 2535
rect 8135 2561 8161 2567
rect 8135 2529 8161 2535
rect 8359 2561 8385 2567
rect 8359 2529 8385 2535
rect 8583 2561 8609 2567
rect 8583 2529 8609 2535
rect 9087 2561 9113 2567
rect 9087 2529 9113 2535
rect 1023 2505 1049 2511
rect 1023 2473 1049 2479
rect 3431 2505 3457 2511
rect 3431 2473 3457 2479
rect 3935 2505 3961 2511
rect 3935 2473 3961 2479
rect 4719 2505 4745 2511
rect 6001 2479 6007 2505
rect 6033 2479 6039 2505
rect 4719 2473 4745 2479
rect 1191 2449 1217 2455
rect 1191 2417 1217 2423
rect 1415 2449 1441 2455
rect 1415 2417 1441 2423
rect 1919 2449 1945 2455
rect 1919 2417 1945 2423
rect 2143 2449 2169 2455
rect 2143 2417 2169 2423
rect 3039 2449 3065 2455
rect 7799 2449 7825 2455
rect 5497 2423 5503 2449
rect 5529 2423 5535 2449
rect 3039 2417 3065 2423
rect 7799 2417 7825 2423
rect 8751 2449 8777 2455
rect 8751 2417 8777 2423
rect 8919 2449 8945 2455
rect 8919 2417 8945 2423
rect 672 2365 9376 2382
rect 672 2339 2763 2365
rect 2789 2339 2815 2365
rect 2841 2339 2867 2365
rect 2893 2339 4919 2365
rect 4945 2339 4971 2365
rect 4997 2339 5023 2365
rect 5049 2339 7075 2365
rect 7101 2339 7127 2365
rect 7153 2339 7179 2365
rect 7205 2339 9231 2365
rect 9257 2339 9283 2365
rect 9309 2339 9335 2365
rect 9361 2339 9376 2365
rect 672 2322 9376 2339
rect 1023 2281 1049 2287
rect 1023 2249 1049 2255
rect 1695 2281 1721 2287
rect 1695 2249 1721 2255
rect 7855 2281 7881 2287
rect 7855 2249 7881 2255
rect 8863 2281 8889 2287
rect 8863 2249 8889 2255
rect 1863 2225 1889 2231
rect 1353 2199 1359 2225
rect 1385 2199 1391 2225
rect 1863 2193 1889 2199
rect 2199 2225 2225 2231
rect 2199 2193 2225 2199
rect 2423 2225 2449 2231
rect 2423 2193 2449 2199
rect 3207 2225 3233 2231
rect 5111 2225 5137 2231
rect 4433 2199 4439 2225
rect 4465 2199 4471 2225
rect 3207 2193 3233 2199
rect 5111 2193 5137 2199
rect 6119 2225 6145 2231
rect 6119 2193 6145 2199
rect 8247 2225 8273 2231
rect 8247 2193 8273 2199
rect 855 2169 881 2175
rect 855 2137 881 2143
rect 1191 2169 1217 2175
rect 1191 2137 1217 2143
rect 1527 2169 1553 2175
rect 4831 2169 4857 2175
rect 8415 2169 8441 2175
rect 3481 2143 3487 2169
rect 3513 2143 3519 2169
rect 4489 2143 4495 2169
rect 4521 2143 4527 2169
rect 6673 2143 6679 2169
rect 6705 2143 6711 2169
rect 7961 2143 7967 2169
rect 7993 2143 7999 2169
rect 8969 2143 8975 2169
rect 9001 2143 9007 2169
rect 1527 2137 1553 2143
rect 4831 2137 4857 2143
rect 8415 2137 8441 2143
rect 6903 2113 6929 2119
rect 3537 2087 3543 2113
rect 3569 2087 3575 2113
rect 5049 2087 5055 2113
rect 5081 2087 5087 2113
rect 6903 2081 6929 2087
rect 7127 2113 7153 2119
rect 7127 2081 7153 2087
rect 7351 2113 7377 2119
rect 7351 2081 7377 2087
rect 7743 2113 7769 2119
rect 7743 2081 7769 2087
rect 672 1973 9296 1990
rect 672 1947 1685 1973
rect 1711 1947 1737 1973
rect 1763 1947 1789 1973
rect 1815 1947 3841 1973
rect 3867 1947 3893 1973
rect 3919 1947 3945 1973
rect 3971 1947 5997 1973
rect 6023 1947 6049 1973
rect 6075 1947 6101 1973
rect 6127 1947 8153 1973
rect 8179 1947 8205 1973
rect 8231 1947 8257 1973
rect 8283 1947 9296 1973
rect 672 1930 9296 1947
rect 4041 1807 4047 1833
rect 4073 1807 4079 1833
rect 1471 1777 1497 1783
rect 4831 1777 4857 1783
rect 2361 1751 2367 1777
rect 2393 1751 2399 1777
rect 3593 1751 3599 1777
rect 3625 1751 3631 1777
rect 4153 1751 4159 1777
rect 4185 1751 4191 1777
rect 5273 1751 5279 1777
rect 5305 1751 5311 1777
rect 5609 1751 5615 1777
rect 5641 1751 5647 1777
rect 5945 1751 5951 1777
rect 5977 1751 5983 1777
rect 6673 1751 6679 1777
rect 6705 1751 6711 1777
rect 7009 1751 7015 1777
rect 7041 1751 7047 1777
rect 7345 1751 7351 1777
rect 7377 1751 7383 1777
rect 7681 1751 7687 1777
rect 7713 1751 7719 1777
rect 8017 1751 8023 1777
rect 8049 1751 8055 1777
rect 8577 1751 8583 1777
rect 8609 1751 8615 1777
rect 8913 1751 8919 1777
rect 8945 1751 8951 1777
rect 1471 1745 1497 1751
rect 4831 1745 4857 1751
rect 1135 1721 1161 1727
rect 1135 1689 1161 1695
rect 1303 1721 1329 1727
rect 4999 1721 5025 1727
rect 1633 1695 1639 1721
rect 1665 1695 1671 1721
rect 1969 1695 1975 1721
rect 2001 1695 2007 1721
rect 2473 1695 2479 1721
rect 2505 1695 2511 1721
rect 3537 1695 3543 1721
rect 3569 1695 3575 1721
rect 4097 1695 4103 1721
rect 4129 1695 4135 1721
rect 1303 1689 1329 1695
rect 4999 1689 5025 1695
rect 5167 1721 5193 1727
rect 5167 1689 5193 1695
rect 5503 1721 5529 1727
rect 5503 1689 5529 1695
rect 5839 1721 5865 1727
rect 5839 1689 5865 1695
rect 6567 1721 6593 1727
rect 6567 1689 6593 1695
rect 7239 1721 7265 1727
rect 7239 1689 7265 1695
rect 7575 1721 7601 1727
rect 7575 1689 7601 1695
rect 7911 1721 7937 1727
rect 7911 1689 7937 1695
rect 8471 1721 8497 1727
rect 8471 1689 8497 1695
rect 855 1665 881 1671
rect 855 1633 881 1639
rect 1807 1665 1833 1671
rect 1807 1633 1833 1639
rect 6175 1665 6201 1671
rect 6175 1633 6201 1639
rect 6903 1665 6929 1671
rect 6903 1633 6929 1639
rect 8807 1665 8833 1671
rect 8807 1633 8833 1639
rect 672 1581 9376 1598
rect 672 1555 2763 1581
rect 2789 1555 2815 1581
rect 2841 1555 2867 1581
rect 2893 1555 4919 1581
rect 4945 1555 4971 1581
rect 4997 1555 5023 1581
rect 5049 1555 7075 1581
rect 7101 1555 7127 1581
rect 7153 1555 7179 1581
rect 7205 1555 9231 1581
rect 9257 1555 9283 1581
rect 9309 1555 9335 1581
rect 9361 1555 9376 1581
rect 672 1538 9376 1555
<< via1 >>
rect 1685 8219 1711 8245
rect 1737 8219 1763 8245
rect 1789 8219 1815 8245
rect 3841 8219 3867 8245
rect 3893 8219 3919 8245
rect 3945 8219 3971 8245
rect 5997 8219 6023 8245
rect 6049 8219 6075 8245
rect 6101 8219 6127 8245
rect 8153 8219 8179 8245
rect 8205 8219 8231 8245
rect 8257 8219 8283 8245
rect 4663 8135 4689 8161
rect 1079 7967 1105 7993
rect 1303 7967 1329 7993
rect 3151 7967 3177 7993
rect 3487 7967 3513 7993
rect 3823 7967 3849 7993
rect 4383 7967 4409 7993
rect 5503 7967 5529 7993
rect 5839 7967 5865 7993
rect 6847 7967 6873 7993
rect 7183 7967 7209 7993
rect 7519 7967 7545 7993
rect 855 7911 881 7937
rect 5055 7911 5081 7937
rect 9087 7911 9113 7937
rect 2763 7827 2789 7853
rect 2815 7827 2841 7853
rect 2867 7827 2893 7853
rect 4919 7827 4945 7853
rect 4971 7827 4997 7853
rect 5023 7827 5049 7853
rect 7075 7827 7101 7853
rect 7127 7827 7153 7853
rect 7179 7827 7205 7853
rect 9231 7827 9257 7853
rect 9283 7827 9309 7853
rect 9335 7827 9361 7853
rect 4831 7743 4857 7769
rect 855 7687 881 7713
rect 9087 7687 9113 7713
rect 1685 7435 1711 7461
rect 1737 7435 1763 7461
rect 1789 7435 1815 7461
rect 3841 7435 3867 7461
rect 3893 7435 3919 7461
rect 3945 7435 3971 7461
rect 5997 7435 6023 7461
rect 6049 7435 6075 7461
rect 6101 7435 6127 7461
rect 8153 7435 8179 7461
rect 8205 7435 8231 7461
rect 8257 7435 8283 7461
rect 855 7127 881 7153
rect 9087 7127 9113 7153
rect 2763 7043 2789 7069
rect 2815 7043 2841 7069
rect 2867 7043 2893 7069
rect 4919 7043 4945 7069
rect 4971 7043 4997 7069
rect 5023 7043 5049 7069
rect 7075 7043 7101 7069
rect 7127 7043 7153 7069
rect 7179 7043 7205 7069
rect 9231 7043 9257 7069
rect 9283 7043 9309 7069
rect 9335 7043 9361 7069
rect 5559 6847 5585 6873
rect 911 6791 937 6817
rect 3487 6791 3513 6817
rect 5895 6791 5921 6817
rect 6959 6791 6985 6817
rect 3543 6735 3569 6761
rect 1685 6651 1711 6677
rect 1737 6651 1763 6677
rect 1789 6651 1815 6677
rect 3841 6651 3867 6677
rect 3893 6651 3919 6677
rect 3945 6651 3971 6677
rect 5997 6651 6023 6677
rect 6049 6651 6075 6677
rect 6101 6651 6127 6677
rect 8153 6651 8179 6677
rect 8205 6651 8231 6677
rect 8257 6651 8283 6677
rect 4383 6511 4409 6537
rect 6455 6511 6481 6537
rect 8191 6511 8217 6537
rect 2983 6455 3009 6481
rect 5055 6455 5081 6481
rect 7687 6455 7713 6481
rect 8471 6455 8497 6481
rect 855 6399 881 6425
rect 1023 6399 1049 6425
rect 3319 6399 3345 6425
rect 5391 6399 5417 6425
rect 9031 6399 9057 6425
rect 1191 6343 1217 6369
rect 2763 6259 2789 6285
rect 2815 6259 2841 6285
rect 2867 6259 2893 6285
rect 4919 6259 4945 6285
rect 4971 6259 4997 6285
rect 5023 6259 5049 6285
rect 7075 6259 7101 6285
rect 7127 6259 7153 6285
rect 7179 6259 7205 6285
rect 9231 6259 9257 6285
rect 9283 6259 9309 6285
rect 9335 6259 9361 6285
rect 3487 6175 3513 6201
rect 3935 6175 3961 6201
rect 3991 6175 4017 6201
rect 4831 6175 4857 6201
rect 5391 6175 5417 6201
rect 855 6119 881 6145
rect 3711 6119 3737 6145
rect 4103 6119 4129 6145
rect 8919 6119 8945 6145
rect 3431 6063 3457 6089
rect 3543 6063 3569 6089
rect 3879 6063 3905 6089
rect 4775 6063 4801 6089
rect 4943 6063 4969 6089
rect 5279 6063 5305 6089
rect 5503 6063 5529 6089
rect 5615 6063 5641 6089
rect 5895 6063 5921 6089
rect 9087 6063 9113 6089
rect 5111 6007 5137 6033
rect 7015 6007 7041 6033
rect 8807 6007 8833 6033
rect 1685 5867 1711 5893
rect 1737 5867 1763 5893
rect 1789 5867 1815 5893
rect 3841 5867 3867 5893
rect 3893 5867 3919 5893
rect 3945 5867 3971 5893
rect 5997 5867 6023 5893
rect 6049 5867 6075 5893
rect 6101 5867 6127 5893
rect 8153 5867 8179 5893
rect 8205 5867 8231 5893
rect 8257 5867 8283 5893
rect 6231 5783 6257 5809
rect 3543 5727 3569 5753
rect 6791 5727 6817 5753
rect 7239 5727 7265 5753
rect 1471 5671 1497 5697
rect 5783 5671 5809 5697
rect 6119 5671 6145 5697
rect 6343 5671 6369 5697
rect 6735 5671 6761 5697
rect 6847 5671 6873 5697
rect 7295 5671 7321 5697
rect 7463 5671 7489 5697
rect 7687 5671 7713 5697
rect 7743 5671 7769 5697
rect 8471 5671 8497 5697
rect 1023 5615 1049 5641
rect 5951 5615 5977 5641
rect 7183 5615 7209 5641
rect 9031 5615 9057 5641
rect 6343 5559 6369 5585
rect 6959 5559 6985 5585
rect 7631 5559 7657 5585
rect 7855 5559 7881 5585
rect 2763 5475 2789 5501
rect 2815 5475 2841 5501
rect 2867 5475 2893 5501
rect 4919 5475 4945 5501
rect 4971 5475 4997 5501
rect 5023 5475 5049 5501
rect 7075 5475 7101 5501
rect 7127 5475 7153 5501
rect 7179 5475 7205 5501
rect 9231 5475 9257 5501
rect 9283 5475 9309 5501
rect 9335 5475 9361 5501
rect 1023 5335 1049 5361
rect 4439 5335 4465 5361
rect 4551 5335 4577 5361
rect 5951 5335 5977 5361
rect 7911 5335 7937 5361
rect 8919 5335 8945 5361
rect 855 5279 881 5305
rect 4047 5279 4073 5305
rect 4383 5279 4409 5305
rect 5111 5279 5137 5305
rect 9087 5279 9113 5305
rect 1247 5223 1273 5249
rect 2647 5223 2673 5249
rect 3711 5223 3737 5249
rect 7743 5223 7769 5249
rect 8807 5223 8833 5249
rect 1685 5083 1711 5109
rect 1737 5083 1763 5109
rect 1789 5083 1815 5109
rect 3841 5083 3867 5109
rect 3893 5083 3919 5109
rect 3945 5083 3971 5109
rect 5997 5083 6023 5109
rect 6049 5083 6075 5109
rect 6101 5083 6127 5109
rect 8153 5083 8179 5109
rect 8205 5083 8231 5109
rect 8257 5083 8283 5109
rect 6287 4999 6313 5025
rect 6455 4999 6481 5025
rect 3039 4943 3065 4969
rect 3319 4943 3345 4969
rect 8471 4943 8497 4969
rect 3095 4887 3121 4913
rect 3375 4887 3401 4913
rect 3543 4887 3569 4913
rect 3823 4887 3849 4913
rect 3879 4887 3905 4913
rect 4103 4887 4129 4913
rect 4215 4887 4241 4913
rect 5279 4887 5305 4913
rect 6455 4887 6481 4913
rect 6847 4887 6873 4913
rect 7015 4887 7041 4913
rect 855 4831 881 4857
rect 3263 4831 3289 4857
rect 4271 4831 4297 4857
rect 5503 4831 5529 4857
rect 7407 4831 7433 4857
rect 8919 4831 8945 4857
rect 9087 4831 9113 4857
rect 1023 4775 1049 4801
rect 1247 4775 1273 4801
rect 3767 4775 3793 4801
rect 4327 4775 4353 4801
rect 6679 4775 6705 4801
rect 6791 4775 6817 4801
rect 8807 4775 8833 4801
rect 2763 4691 2789 4717
rect 2815 4691 2841 4717
rect 2867 4691 2893 4717
rect 4919 4691 4945 4717
rect 4971 4691 4997 4717
rect 5023 4691 5049 4717
rect 7075 4691 7101 4717
rect 7127 4691 7153 4717
rect 7179 4691 7205 4717
rect 9231 4691 9257 4717
rect 9283 4691 9309 4717
rect 9335 4691 9361 4717
rect 7015 4607 7041 4633
rect 1023 4551 1049 4577
rect 2479 4551 2505 4577
rect 2927 4551 2953 4577
rect 3991 4551 4017 4577
rect 5671 4551 5697 4577
rect 6511 4551 6537 4577
rect 6679 4551 6705 4577
rect 8919 4551 8945 4577
rect 855 4495 881 4521
rect 2255 4495 2281 4521
rect 2983 4495 3009 4521
rect 3935 4495 3961 4521
rect 4327 4495 4353 4521
rect 5223 4495 5249 4521
rect 5447 4495 5473 4521
rect 6231 4495 6257 4521
rect 6959 4495 6985 4521
rect 7127 4495 7153 4521
rect 7183 4495 7209 4521
rect 7351 4495 7377 4521
rect 9087 4495 9113 4521
rect 1247 4439 1273 4465
rect 3823 4439 3849 4465
rect 4439 4439 4465 4465
rect 5503 4439 5529 4465
rect 6175 4439 6201 4465
rect 8807 4439 8833 4465
rect 3991 4383 4017 4409
rect 4495 4383 4521 4409
rect 1685 4299 1711 4325
rect 1737 4299 1763 4325
rect 1789 4299 1815 4325
rect 3841 4299 3867 4325
rect 3893 4299 3919 4325
rect 3945 4299 3971 4325
rect 5997 4299 6023 4325
rect 6049 4299 6075 4325
rect 6101 4299 6127 4325
rect 8153 4299 8179 4325
rect 8205 4299 8231 4325
rect 8257 4299 8283 4325
rect 2255 4215 2281 4241
rect 6735 4215 6761 4241
rect 5839 4159 5865 4185
rect 6903 4159 6929 4185
rect 4327 4103 4353 4129
rect 5335 4103 5361 4129
rect 7015 4103 7041 4129
rect 855 4047 881 4073
rect 1191 4047 1217 4073
rect 1359 4047 1385 4073
rect 2087 4047 2113 4073
rect 4607 4047 4633 4073
rect 5615 4047 5641 4073
rect 6847 4047 6873 4073
rect 7127 4047 7153 4073
rect 7183 4047 7209 4073
rect 8583 4047 8609 4073
rect 8751 4047 8777 4073
rect 9087 4047 9113 4073
rect 1023 3991 1049 4017
rect 1583 3991 1609 4017
rect 2199 3991 2225 4017
rect 8919 3991 8945 4017
rect 2763 3907 2789 3933
rect 2815 3907 2841 3933
rect 2867 3907 2893 3933
rect 4919 3907 4945 3933
rect 4971 3907 4997 3933
rect 5023 3907 5049 3933
rect 7075 3907 7101 3933
rect 7127 3907 7153 3933
rect 7179 3907 7205 3933
rect 9231 3907 9257 3933
rect 9283 3907 9309 3933
rect 9335 3907 9361 3933
rect 1023 3823 1049 3849
rect 1247 3823 1273 3849
rect 2535 3823 2561 3849
rect 4103 3823 4129 3849
rect 4495 3823 4521 3849
rect 4775 3823 4801 3849
rect 5279 3823 5305 3849
rect 5951 3823 5977 3849
rect 9143 3823 9169 3849
rect 1863 3767 1889 3793
rect 3095 3767 3121 3793
rect 4327 3767 4353 3793
rect 4383 3767 4409 3793
rect 5615 3767 5641 3793
rect 6455 3767 6481 3793
rect 7463 3767 7489 3793
rect 855 3711 881 3737
rect 1807 3711 1833 3737
rect 2815 3711 2841 3737
rect 5559 3711 5585 3737
rect 6679 3711 6705 3737
rect 7799 3711 7825 3737
rect 8863 3711 8889 3737
rect 1471 3655 1497 3681
rect 4831 3655 4857 3681
rect 3935 3599 3961 3625
rect 4047 3599 4073 3625
rect 4103 3599 4129 3625
rect 1685 3515 1711 3541
rect 1737 3515 1763 3541
rect 1789 3515 1815 3541
rect 3841 3515 3867 3541
rect 3893 3515 3919 3541
rect 3945 3515 3971 3541
rect 5997 3515 6023 3541
rect 6049 3515 6075 3541
rect 6101 3515 6127 3541
rect 8153 3515 8179 3541
rect 8205 3515 8231 3541
rect 8257 3515 8283 3541
rect 3319 3319 3345 3345
rect 4383 3319 4409 3345
rect 855 3263 881 3289
rect 1023 3263 1049 3289
rect 3375 3263 3401 3289
rect 4663 3263 4689 3289
rect 1247 3207 1273 3233
rect 1471 3207 1497 3233
rect 1695 3207 1721 3233
rect 4215 3207 4241 3233
rect 9087 3207 9113 3233
rect 2763 3123 2789 3149
rect 2815 3123 2841 3149
rect 2867 3123 2893 3149
rect 4919 3123 4945 3149
rect 4971 3123 4997 3149
rect 5023 3123 5049 3149
rect 7075 3123 7101 3149
rect 7127 3123 7153 3149
rect 7179 3123 7205 3149
rect 9231 3123 9257 3149
rect 9283 3123 9309 3149
rect 9335 3123 9361 3149
rect 4383 3039 4409 3065
rect 5895 3039 5921 3065
rect 1023 2983 1049 3009
rect 2591 2983 2617 3009
rect 4159 2983 4185 3009
rect 6399 2983 6425 3009
rect 7407 2983 7433 3009
rect 855 2927 881 2953
rect 3431 2927 3457 2953
rect 3599 2927 3625 2953
rect 6679 2927 6705 2953
rect 7743 2927 7769 2953
rect 1247 2871 1273 2897
rect 1471 2871 1497 2897
rect 1695 2871 1721 2897
rect 1919 2871 1945 2897
rect 2479 2871 2505 2897
rect 5055 2871 5081 2897
rect 5391 2871 5417 2897
rect 5727 2871 5753 2897
rect 8807 2871 8833 2897
rect 9143 2871 9169 2897
rect 1685 2731 1711 2757
rect 1737 2731 1763 2757
rect 1789 2731 1815 2757
rect 3841 2731 3867 2757
rect 3893 2731 3919 2757
rect 3945 2731 3971 2757
rect 5997 2731 6023 2757
rect 6049 2731 6075 2757
rect 6101 2731 6127 2757
rect 8153 2731 8179 2757
rect 8205 2731 8231 2757
rect 8257 2731 8283 2757
rect 2591 2591 2617 2617
rect 911 2535 937 2561
rect 1695 2535 1721 2561
rect 3319 2535 3345 2561
rect 3599 2535 3625 2561
rect 3767 2535 3793 2561
rect 4159 2535 4185 2561
rect 5167 2535 5193 2561
rect 6231 2535 6257 2561
rect 7463 2535 7489 2561
rect 8135 2535 8161 2561
rect 8359 2535 8385 2561
rect 8583 2535 8609 2561
rect 9087 2535 9113 2561
rect 1023 2479 1049 2505
rect 3431 2479 3457 2505
rect 3935 2479 3961 2505
rect 4719 2479 4745 2505
rect 6007 2479 6033 2505
rect 1191 2423 1217 2449
rect 1415 2423 1441 2449
rect 1919 2423 1945 2449
rect 2143 2423 2169 2449
rect 3039 2423 3065 2449
rect 5503 2423 5529 2449
rect 7799 2423 7825 2449
rect 8751 2423 8777 2449
rect 8919 2423 8945 2449
rect 2763 2339 2789 2365
rect 2815 2339 2841 2365
rect 2867 2339 2893 2365
rect 4919 2339 4945 2365
rect 4971 2339 4997 2365
rect 5023 2339 5049 2365
rect 7075 2339 7101 2365
rect 7127 2339 7153 2365
rect 7179 2339 7205 2365
rect 9231 2339 9257 2365
rect 9283 2339 9309 2365
rect 9335 2339 9361 2365
rect 1023 2255 1049 2281
rect 1695 2255 1721 2281
rect 7855 2255 7881 2281
rect 8863 2255 8889 2281
rect 1359 2199 1385 2225
rect 1863 2199 1889 2225
rect 2199 2199 2225 2225
rect 2423 2199 2449 2225
rect 3207 2199 3233 2225
rect 4439 2199 4465 2225
rect 5111 2199 5137 2225
rect 6119 2199 6145 2225
rect 8247 2199 8273 2225
rect 855 2143 881 2169
rect 1191 2143 1217 2169
rect 1527 2143 1553 2169
rect 3487 2143 3513 2169
rect 4495 2143 4521 2169
rect 4831 2143 4857 2169
rect 6679 2143 6705 2169
rect 7967 2143 7993 2169
rect 8415 2143 8441 2169
rect 8975 2143 9001 2169
rect 3543 2087 3569 2113
rect 5055 2087 5081 2113
rect 6903 2087 6929 2113
rect 7127 2087 7153 2113
rect 7351 2087 7377 2113
rect 7743 2087 7769 2113
rect 1685 1947 1711 1973
rect 1737 1947 1763 1973
rect 1789 1947 1815 1973
rect 3841 1947 3867 1973
rect 3893 1947 3919 1973
rect 3945 1947 3971 1973
rect 5997 1947 6023 1973
rect 6049 1947 6075 1973
rect 6101 1947 6127 1973
rect 8153 1947 8179 1973
rect 8205 1947 8231 1973
rect 8257 1947 8283 1973
rect 4047 1807 4073 1833
rect 1471 1751 1497 1777
rect 2367 1751 2393 1777
rect 3599 1751 3625 1777
rect 4159 1751 4185 1777
rect 4831 1751 4857 1777
rect 5279 1751 5305 1777
rect 5615 1751 5641 1777
rect 5951 1751 5977 1777
rect 6679 1751 6705 1777
rect 7015 1751 7041 1777
rect 7351 1751 7377 1777
rect 7687 1751 7713 1777
rect 8023 1751 8049 1777
rect 8583 1751 8609 1777
rect 8919 1751 8945 1777
rect 1135 1695 1161 1721
rect 1303 1695 1329 1721
rect 1639 1695 1665 1721
rect 1975 1695 2001 1721
rect 2479 1695 2505 1721
rect 3543 1695 3569 1721
rect 4103 1695 4129 1721
rect 4999 1695 5025 1721
rect 5167 1695 5193 1721
rect 5503 1695 5529 1721
rect 5839 1695 5865 1721
rect 6567 1695 6593 1721
rect 7239 1695 7265 1721
rect 7575 1695 7601 1721
rect 7911 1695 7937 1721
rect 8471 1695 8497 1721
rect 855 1639 881 1665
rect 1807 1639 1833 1665
rect 6175 1639 6201 1665
rect 6903 1639 6929 1665
rect 8807 1639 8833 1665
rect 2763 1555 2789 1581
rect 2815 1555 2841 1581
rect 2867 1555 2893 1581
rect 4919 1555 4945 1581
rect 4971 1555 4997 1581
rect 5023 1555 5049 1581
rect 7075 1555 7101 1581
rect 7127 1555 7153 1581
rect 7179 1555 7205 1581
rect 9231 1555 9257 1581
rect 9283 1555 9309 1581
rect 9335 1555 9361 1581
<< metal2 >>
rect 3024 9600 3080 10000
rect 3360 9600 3416 10000
rect 3696 9600 3752 10000
rect 4032 9600 4088 10000
rect 4368 9600 4424 10000
rect 4704 9600 4760 10000
rect 5376 9600 5432 10000
rect 5712 9600 5768 10000
rect 6720 9600 6776 10000
rect 7056 9600 7112 10000
rect 7392 9600 7448 10000
rect 1302 8386 1330 8391
rect 1078 8106 1106 8111
rect 1078 7993 1106 8078
rect 1078 7967 1079 7993
rect 1105 7967 1106 7993
rect 1078 7961 1106 7967
rect 1302 7993 1330 8358
rect 1684 8246 1816 8251
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1684 8213 1816 8218
rect 1302 7967 1303 7993
rect 1329 7967 1330 7993
rect 1302 7961 1330 7967
rect 3038 7994 3066 9600
rect 3150 7994 3178 7999
rect 3038 7993 3178 7994
rect 3038 7967 3151 7993
rect 3177 7967 3178 7993
rect 3038 7966 3178 7967
rect 3374 7994 3402 9600
rect 3486 7994 3514 7999
rect 3374 7993 3514 7994
rect 3374 7967 3487 7993
rect 3513 7967 3514 7993
rect 3374 7966 3514 7967
rect 3710 7994 3738 9600
rect 3840 8246 3972 8251
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3840 8213 3972 8218
rect 4046 8162 4074 9600
rect 4046 8129 4074 8134
rect 3822 7994 3850 7999
rect 3710 7993 3850 7994
rect 3710 7967 3823 7993
rect 3849 7967 3850 7993
rect 3710 7966 3850 7967
rect 3150 7961 3178 7966
rect 3486 7961 3514 7966
rect 3822 7961 3850 7966
rect 4382 7993 4410 9600
rect 4662 8162 4690 8167
rect 4662 8115 4690 8134
rect 4382 7967 4383 7993
rect 4409 7967 4410 7993
rect 4382 7961 4410 7967
rect 854 7938 882 7943
rect 854 7891 882 7910
rect 2762 7854 2894 7859
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2762 7821 2894 7826
rect 4718 7770 4746 9600
rect 5390 7994 5418 9600
rect 5502 7994 5530 7999
rect 5390 7993 5530 7994
rect 5390 7967 5503 7993
rect 5529 7967 5530 7993
rect 5390 7966 5530 7967
rect 5726 7994 5754 9600
rect 5996 8246 6128 8251
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 5996 8213 6128 8218
rect 5838 7994 5866 7999
rect 5726 7993 5866 7994
rect 5726 7967 5839 7993
rect 5865 7967 5866 7993
rect 5726 7966 5866 7967
rect 6734 7994 6762 9600
rect 6846 7994 6874 7999
rect 6734 7993 6874 7994
rect 6734 7967 6847 7993
rect 6873 7967 6874 7993
rect 6734 7966 6874 7967
rect 7070 7994 7098 9600
rect 7182 7994 7210 7999
rect 7070 7993 7210 7994
rect 7070 7967 7183 7993
rect 7209 7967 7210 7993
rect 7070 7966 7210 7967
rect 7406 7994 7434 9600
rect 8152 8246 8284 8251
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8152 8213 8284 8218
rect 7518 7994 7546 7999
rect 7406 7993 7546 7994
rect 7406 7967 7519 7993
rect 7545 7967 7546 7993
rect 7406 7966 7546 7967
rect 5502 7961 5530 7966
rect 5838 7961 5866 7966
rect 6846 7961 6874 7966
rect 7182 7961 7210 7966
rect 7518 7961 7546 7966
rect 5054 7938 5082 7943
rect 9086 7938 9114 7943
rect 5054 7937 5138 7938
rect 5054 7911 5055 7937
rect 5081 7911 5138 7937
rect 5054 7910 5138 7911
rect 5054 7905 5082 7910
rect 4918 7854 5050 7859
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 4918 7821 5050 7826
rect 4830 7770 4858 7775
rect 5110 7770 5138 7910
rect 9086 7937 9170 7938
rect 9086 7911 9087 7937
rect 9113 7911 9170 7937
rect 9086 7910 9170 7911
rect 9086 7905 9114 7910
rect 7074 7854 7206 7859
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7074 7821 7206 7826
rect 4718 7769 4858 7770
rect 4718 7743 4831 7769
rect 4857 7743 4858 7769
rect 4718 7742 4858 7743
rect 4830 7737 4858 7742
rect 4886 7742 5138 7770
rect 9142 7770 9170 7910
rect 9230 7854 9362 7859
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9230 7821 9362 7826
rect 854 7713 882 7719
rect 854 7687 855 7713
rect 881 7687 882 7713
rect 854 7602 882 7687
rect 854 7569 882 7574
rect 1684 7462 1816 7467
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1684 7429 1816 7434
rect 3840 7462 3972 7467
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3840 7429 3972 7434
rect 854 7154 882 7159
rect 4886 7154 4914 7742
rect 9142 7737 9170 7742
rect 9086 7713 9114 7719
rect 9086 7687 9087 7713
rect 9113 7687 9114 7713
rect 5996 7462 6128 7467
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 5996 7429 6128 7434
rect 8152 7462 8284 7467
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8152 7429 8284 7434
rect 9086 7434 9114 7687
rect 9086 7401 9114 7406
rect 854 7107 882 7126
rect 4830 7126 4914 7154
rect 9086 7154 9114 7159
rect 2762 7070 2894 7075
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2762 7037 2894 7042
rect 910 6817 938 6823
rect 910 6791 911 6817
rect 937 6791 938 6817
rect 854 6426 882 6431
rect 910 6426 938 6791
rect 3486 6817 3514 6823
rect 3486 6791 3487 6817
rect 3513 6791 3514 6817
rect 1684 6678 1816 6683
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1684 6645 1816 6650
rect 882 6398 938 6426
rect 1022 6594 1050 6599
rect 1022 6425 1050 6566
rect 3486 6594 3514 6791
rect 3486 6561 3514 6566
rect 3542 6761 3570 6767
rect 3542 6735 3543 6761
rect 3569 6735 3570 6761
rect 1022 6399 1023 6425
rect 1049 6399 1050 6425
rect 854 6379 882 6398
rect 1022 6393 1050 6399
rect 2982 6481 3010 6487
rect 2982 6455 2983 6481
rect 3009 6455 3010 6481
rect 1190 6369 1218 6375
rect 1190 6343 1191 6369
rect 1217 6343 1218 6369
rect 854 6145 882 6151
rect 854 6119 855 6145
rect 881 6119 882 6145
rect 854 5754 882 6119
rect 1190 6090 1218 6343
rect 2762 6286 2894 6291
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2762 6253 2894 6258
rect 1190 6057 1218 6062
rect 1684 5894 1816 5899
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1684 5861 1816 5866
rect 854 5721 882 5726
rect 2982 5754 3010 6455
rect 3318 6426 3346 6431
rect 3318 6425 3514 6426
rect 3318 6399 3319 6425
rect 3345 6399 3514 6425
rect 3318 6398 3514 6399
rect 3318 6393 3346 6398
rect 3486 6201 3514 6398
rect 3486 6175 3487 6201
rect 3513 6175 3514 6201
rect 3486 6169 3514 6175
rect 2982 5721 3010 5726
rect 3430 6089 3458 6095
rect 3430 6063 3431 6089
rect 3457 6063 3458 6089
rect 3430 5978 3458 6063
rect 3542 6089 3570 6735
rect 3840 6678 3972 6683
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3840 6645 3972 6650
rect 3990 6538 4018 6543
rect 3934 6202 3962 6207
rect 3710 6201 3962 6202
rect 3710 6175 3935 6201
rect 3961 6175 3962 6201
rect 3710 6174 3962 6175
rect 3710 6145 3738 6174
rect 3934 6169 3962 6174
rect 3990 6201 4018 6510
rect 4382 6538 4410 6543
rect 4382 6491 4410 6510
rect 4830 6538 4858 7126
rect 9086 7107 9114 7126
rect 4918 7070 5050 7075
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 4918 7037 5050 7042
rect 7074 7070 7206 7075
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7074 7037 7206 7042
rect 9230 7070 9362 7075
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9230 7037 9362 7042
rect 5558 6873 5586 6879
rect 5558 6847 5559 6873
rect 5585 6847 5586 6873
rect 3990 6175 3991 6201
rect 4017 6175 4018 6201
rect 3990 6169 4018 6175
rect 4830 6201 4858 6510
rect 5110 6762 5138 6767
rect 5054 6482 5082 6487
rect 5054 6435 5082 6454
rect 4918 6286 5050 6291
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 4918 6253 5050 6258
rect 4830 6175 4831 6201
rect 4857 6175 4858 6201
rect 4830 6169 4858 6175
rect 3710 6119 3711 6145
rect 3737 6119 3738 6145
rect 3710 6113 3738 6119
rect 4102 6145 4130 6151
rect 4102 6119 4103 6145
rect 4129 6119 4130 6145
rect 3542 6063 3543 6089
rect 3569 6063 3570 6089
rect 3542 6057 3570 6063
rect 3878 6089 3906 6095
rect 3878 6063 3879 6089
rect 3905 6063 3906 6089
rect 3878 5978 3906 6063
rect 3430 5950 3906 5978
rect 1470 5698 1498 5703
rect 1470 5651 1498 5670
rect 2646 5698 2674 5703
rect 1022 5641 1050 5647
rect 1022 5615 1023 5641
rect 1049 5615 1050 5641
rect 1022 5474 1050 5615
rect 1022 5441 1050 5446
rect 1022 5361 1050 5367
rect 1022 5335 1023 5361
rect 1049 5335 1050 5361
rect 854 5305 882 5311
rect 854 5279 855 5305
rect 881 5279 882 5305
rect 854 5082 882 5279
rect 854 5049 882 5054
rect 1022 4970 1050 5335
rect 1246 5249 1274 5255
rect 1246 5223 1247 5249
rect 1273 5223 1274 5249
rect 1246 5082 1274 5223
rect 2646 5250 2674 5670
rect 2762 5502 2894 5507
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2762 5469 2894 5474
rect 2646 5203 2674 5222
rect 1684 5110 1816 5115
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 3374 5082 3402 5087
rect 1684 5077 1816 5082
rect 1246 5049 1274 5054
rect 3318 5054 3374 5082
rect 1022 4937 1050 4942
rect 3038 4970 3066 4975
rect 3038 4923 3066 4942
rect 3318 4969 3346 5054
rect 3374 5049 3402 5054
rect 3318 4943 3319 4969
rect 3345 4943 3346 4969
rect 3318 4937 3346 4943
rect 3094 4914 3122 4919
rect 3094 4867 3122 4886
rect 3374 4914 3402 4919
rect 3374 4867 3402 4886
rect 854 4857 882 4863
rect 854 4831 855 4857
rect 881 4831 882 4857
rect 854 4746 882 4831
rect 3262 4857 3290 4863
rect 3262 4831 3263 4857
rect 3289 4831 3290 4857
rect 1022 4802 1050 4807
rect 1022 4801 1106 4802
rect 1022 4775 1023 4801
rect 1049 4775 1106 4801
rect 1022 4774 1106 4775
rect 1022 4769 1050 4774
rect 854 4713 882 4718
rect 1022 4577 1050 4583
rect 1022 4551 1023 4577
rect 1049 4551 1050 4577
rect 854 4521 882 4527
rect 854 4495 855 4521
rect 881 4495 882 4521
rect 854 4410 882 4495
rect 854 4377 882 4382
rect 1022 4214 1050 4551
rect 966 4186 1050 4214
rect 854 4074 882 4079
rect 854 4027 882 4046
rect 966 3850 994 4186
rect 1022 4018 1050 4037
rect 1022 3985 1050 3990
rect 966 3817 994 3822
rect 1022 3906 1050 3911
rect 1022 3849 1050 3878
rect 1022 3823 1023 3849
rect 1049 3823 1050 3849
rect 1022 3817 1050 3823
rect 854 3737 882 3743
rect 854 3711 855 3737
rect 881 3711 882 3737
rect 854 3682 882 3711
rect 1078 3738 1106 4774
rect 1246 4801 1274 4807
rect 1246 4775 1247 4801
rect 1273 4775 1274 4801
rect 1246 4746 1274 4775
rect 3262 4802 3290 4831
rect 3262 4769 3290 4774
rect 3430 4802 3458 5950
rect 3840 5894 3972 5899
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3840 5861 3972 5866
rect 3542 5754 3570 5759
rect 3542 5707 3570 5726
rect 4046 5754 4074 5759
rect 4046 5305 4074 5726
rect 4046 5279 4047 5305
rect 4073 5279 4074 5305
rect 4046 5273 4074 5279
rect 3710 5249 3738 5255
rect 3710 5223 3711 5249
rect 3737 5223 3738 5249
rect 3710 5082 3738 5223
rect 3710 5049 3738 5054
rect 3766 5250 3794 5255
rect 3766 5026 3794 5222
rect 3840 5110 3972 5115
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3840 5077 3972 5082
rect 3766 4998 3906 5026
rect 3542 4914 3570 4919
rect 3822 4914 3850 4919
rect 3542 4913 3850 4914
rect 3542 4887 3543 4913
rect 3569 4887 3823 4913
rect 3849 4887 3850 4913
rect 3542 4886 3850 4887
rect 3542 4881 3570 4886
rect 3822 4881 3850 4886
rect 3878 4913 3906 4998
rect 3878 4887 3879 4913
rect 3905 4887 3906 4913
rect 3878 4881 3906 4887
rect 4102 4914 4130 6119
rect 4774 6089 4802 6095
rect 4774 6063 4775 6089
rect 4801 6063 4802 6089
rect 4774 5754 4802 6063
rect 4942 6090 4970 6095
rect 4942 6043 4970 6062
rect 4382 5726 4802 5754
rect 5110 6033 5138 6734
rect 5558 6482 5586 6847
rect 5390 6425 5418 6431
rect 5390 6399 5391 6425
rect 5417 6399 5418 6425
rect 5390 6201 5418 6399
rect 5390 6175 5391 6201
rect 5417 6175 5418 6201
rect 5390 6169 5418 6175
rect 5278 6090 5306 6095
rect 5278 6043 5306 6062
rect 5502 6090 5530 6095
rect 5502 6043 5530 6062
rect 5110 6007 5111 6033
rect 5137 6007 5138 6033
rect 4382 5305 4410 5726
rect 4550 5642 4578 5647
rect 4438 5362 4466 5367
rect 4438 5315 4466 5334
rect 4550 5361 4578 5614
rect 4918 5502 5050 5507
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 4918 5469 5050 5474
rect 4550 5335 4551 5361
rect 4577 5335 4578 5361
rect 4550 5329 4578 5335
rect 4382 5279 4383 5305
rect 4409 5279 4410 5305
rect 4102 4867 4130 4886
rect 4214 4913 4242 4919
rect 4214 4887 4215 4913
rect 4241 4887 4242 4913
rect 3430 4769 3458 4774
rect 3766 4802 3794 4807
rect 1246 4713 1274 4718
rect 2762 4718 2894 4723
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2762 4685 2894 4690
rect 1358 4578 1386 4583
rect 1246 4465 1274 4471
rect 1246 4439 1247 4465
rect 1273 4439 1274 4465
rect 1246 4410 1274 4439
rect 1246 4377 1274 4382
rect 1190 4073 1218 4079
rect 1190 4047 1191 4073
rect 1217 4047 1218 4073
rect 1190 3794 1218 4047
rect 1246 4074 1274 4079
rect 1246 3849 1274 4046
rect 1358 4073 1386 4550
rect 2478 4577 2506 4583
rect 2478 4551 2479 4577
rect 2505 4551 2506 4577
rect 2254 4521 2282 4527
rect 2254 4495 2255 4521
rect 2281 4495 2282 4521
rect 1684 4326 1816 4331
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1684 4293 1816 4298
rect 2254 4241 2282 4495
rect 2254 4215 2255 4241
rect 2281 4215 2282 4241
rect 2254 4209 2282 4215
rect 2478 4214 2506 4551
rect 2926 4578 2954 4583
rect 2926 4531 2954 4550
rect 2982 4521 3010 4527
rect 2982 4495 2983 4521
rect 3009 4495 3010 4521
rect 2478 4186 2562 4214
rect 1358 4047 1359 4073
rect 1385 4047 1386 4073
rect 1358 4041 1386 4047
rect 2086 4073 2114 4079
rect 2086 4047 2087 4073
rect 2113 4047 2114 4073
rect 1246 3823 1247 3849
rect 1273 3823 1274 3849
rect 1246 3817 1274 3823
rect 1582 4017 1610 4023
rect 1582 3991 1583 4017
rect 1609 3991 1610 4017
rect 1190 3761 1218 3766
rect 1582 3794 1610 3991
rect 2086 3906 2114 4047
rect 2086 3873 2114 3878
rect 2198 4017 2226 4023
rect 2198 3991 2199 4017
rect 2225 3991 2226 4017
rect 1582 3761 1610 3766
rect 1862 3793 1890 3799
rect 1862 3767 1863 3793
rect 1889 3767 1890 3793
rect 1078 3705 1106 3710
rect 1806 3738 1834 3743
rect 1806 3691 1834 3710
rect 854 3402 882 3654
rect 1470 3682 1498 3687
rect 1470 3635 1498 3654
rect 854 3369 882 3374
rect 1022 3626 1050 3631
rect 854 3289 882 3295
rect 854 3263 855 3289
rect 881 3263 882 3289
rect 854 3066 882 3263
rect 1022 3289 1050 3598
rect 1684 3542 1816 3547
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1684 3509 1816 3514
rect 1134 3402 1162 3407
rect 1022 3263 1023 3289
rect 1049 3263 1050 3289
rect 1022 3257 1050 3263
rect 1078 3374 1134 3402
rect 854 3033 882 3038
rect 1022 3010 1050 3015
rect 1022 2963 1050 2982
rect 854 2953 882 2959
rect 854 2927 855 2953
rect 881 2927 882 2953
rect 854 2730 882 2927
rect 854 2697 882 2702
rect 966 2954 994 2959
rect 910 2561 938 2567
rect 910 2535 911 2561
rect 937 2535 938 2561
rect 910 2506 938 2535
rect 910 2473 938 2478
rect 966 2282 994 2926
rect 1078 2898 1106 3374
rect 1134 3369 1162 3374
rect 1862 3402 1890 3767
rect 2198 3626 2226 3991
rect 2534 3849 2562 4186
rect 2762 3934 2894 3939
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2762 3901 2894 3906
rect 2534 3823 2535 3849
rect 2561 3823 2562 3849
rect 2534 3817 2562 3823
rect 2814 3850 2842 3855
rect 2814 3737 2842 3822
rect 2814 3711 2815 3737
rect 2841 3711 2842 3737
rect 2814 3705 2842 3711
rect 2198 3593 2226 3598
rect 1862 3369 1890 3374
rect 2310 3346 2338 3351
rect 1190 3234 1218 3239
rect 1022 2870 1106 2898
rect 1134 3206 1190 3234
rect 1022 2505 1050 2870
rect 1134 2506 1162 3206
rect 1190 3201 1218 3206
rect 1246 3233 1274 3239
rect 1246 3207 1247 3233
rect 1273 3207 1274 3233
rect 1246 3066 1274 3207
rect 1470 3234 1498 3239
rect 1694 3234 1722 3239
rect 1470 3233 1554 3234
rect 1470 3207 1471 3233
rect 1497 3207 1554 3233
rect 1470 3206 1554 3207
rect 1470 3201 1498 3206
rect 1246 3033 1274 3038
rect 1246 2897 1274 2903
rect 1246 2871 1247 2897
rect 1273 2871 1274 2897
rect 1246 2730 1274 2871
rect 1470 2897 1498 2903
rect 1470 2871 1471 2897
rect 1497 2871 1498 2897
rect 1246 2697 1274 2702
rect 1302 2842 1330 2847
rect 1022 2479 1023 2505
rect 1049 2479 1050 2505
rect 1022 2473 1050 2479
rect 1078 2478 1162 2506
rect 1022 2282 1050 2287
rect 966 2281 1050 2282
rect 966 2255 1023 2281
rect 1049 2255 1050 2281
rect 966 2254 1050 2255
rect 1022 2249 1050 2254
rect 854 2170 882 2175
rect 798 2142 854 2170
rect 798 2114 826 2142
rect 854 2123 882 2142
rect 686 2086 826 2114
rect 14 1946 42 1951
rect 14 400 42 1918
rect 406 1890 434 1895
rect 350 1862 406 1890
rect 350 400 378 1862
rect 406 1857 434 1862
rect 686 400 714 2086
rect 854 2058 882 2063
rect 854 1665 882 2030
rect 1078 1722 1106 2478
rect 1190 2450 1218 2455
rect 1134 2449 1218 2450
rect 1134 2423 1191 2449
rect 1217 2423 1218 2449
rect 1134 2422 1218 2423
rect 1134 1834 1162 2422
rect 1190 2417 1218 2422
rect 1190 2282 1218 2287
rect 1190 2169 1218 2254
rect 1190 2143 1191 2169
rect 1217 2143 1218 2169
rect 1190 1946 1218 2143
rect 1190 1913 1218 1918
rect 1134 1801 1162 1806
rect 1134 1722 1162 1727
rect 854 1639 855 1665
rect 881 1639 882 1665
rect 854 1633 882 1639
rect 1022 1721 1162 1722
rect 1022 1695 1135 1721
rect 1161 1695 1162 1721
rect 1022 1694 1162 1695
rect 1022 400 1050 1694
rect 1134 1689 1162 1694
rect 1302 1721 1330 2814
rect 1470 2506 1498 2871
rect 1470 2473 1498 2478
rect 1414 2449 1442 2455
rect 1414 2423 1415 2449
rect 1441 2423 1442 2449
rect 1358 2226 1386 2231
rect 1358 2179 1386 2198
rect 1302 1695 1303 1721
rect 1329 1695 1330 1721
rect 1302 1689 1330 1695
rect 1414 1050 1442 2423
rect 1526 2282 1554 3206
rect 1694 3187 1722 3206
rect 1694 2897 1722 2903
rect 1694 2871 1695 2897
rect 1721 2871 1722 2897
rect 1694 2842 1722 2871
rect 1414 1017 1442 1022
rect 1470 2254 1554 2282
rect 1582 2814 1722 2842
rect 1918 2897 1946 2903
rect 1918 2871 1919 2897
rect 1945 2871 1946 2897
rect 1582 2282 1610 2814
rect 1684 2758 1816 2763
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1684 2725 1816 2730
rect 1694 2561 1722 2567
rect 1918 2562 1946 2871
rect 1694 2535 1695 2561
rect 1721 2535 1722 2561
rect 1694 2450 1722 2535
rect 1470 1777 1498 2254
rect 1582 2249 1610 2254
rect 1638 2422 1722 2450
rect 1806 2534 1946 2562
rect 1526 2170 1554 2175
rect 1638 2170 1666 2422
rect 1694 2282 1722 2287
rect 1694 2235 1722 2254
rect 1526 2169 1666 2170
rect 1526 2143 1527 2169
rect 1553 2143 1666 2169
rect 1526 2142 1666 2143
rect 1806 2170 1834 2534
rect 1918 2449 1946 2455
rect 1918 2423 1919 2449
rect 1945 2423 1946 2449
rect 1526 1890 1554 2142
rect 1806 2137 1834 2142
rect 1862 2225 1890 2231
rect 1862 2199 1863 2225
rect 1889 2199 1890 2225
rect 1684 1974 1816 1979
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1684 1941 1816 1946
rect 1526 1857 1554 1862
rect 1638 1890 1666 1895
rect 1862 1890 1890 2199
rect 1470 1751 1471 1777
rect 1497 1751 1498 1777
rect 1470 938 1498 1751
rect 1638 1721 1666 1862
rect 1638 1695 1639 1721
rect 1665 1695 1666 1721
rect 1638 1689 1666 1695
rect 1750 1862 1890 1890
rect 1750 1386 1778 1862
rect 1750 1353 1778 1358
rect 1806 1666 1834 1671
rect 1918 1666 1946 2423
rect 1974 2450 2002 2455
rect 2142 2450 2170 2455
rect 1974 1721 2002 2422
rect 1974 1695 1975 1721
rect 2001 1695 2002 1721
rect 1974 1689 2002 1695
rect 2030 2449 2170 2450
rect 2030 2423 2143 2449
rect 2169 2423 2170 2449
rect 2030 2422 2170 2423
rect 1806 1665 1946 1666
rect 1806 1639 1807 1665
rect 1833 1639 1946 1665
rect 1806 1638 1946 1639
rect 1806 1274 1834 1638
rect 1358 910 1498 938
rect 1694 1246 1834 1274
rect 1358 400 1386 910
rect 1694 400 1722 1246
rect 2030 400 2058 2422
rect 2142 2417 2170 2422
rect 2198 2226 2226 2231
rect 2198 2225 2282 2226
rect 2198 2199 2199 2225
rect 2225 2199 2282 2225
rect 2198 2198 2282 2199
rect 2198 2193 2226 2198
rect 2254 490 2282 2198
rect 2310 1666 2338 3318
rect 2762 3150 2894 3155
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2762 3117 2894 3122
rect 2590 3009 2618 3015
rect 2590 2983 2591 3009
rect 2617 2983 2618 3009
rect 2478 2898 2506 2903
rect 2366 2897 2506 2898
rect 2366 2871 2479 2897
rect 2505 2871 2506 2897
rect 2366 2870 2506 2871
rect 2366 1778 2394 2870
rect 2478 2865 2506 2870
rect 2590 2842 2618 2983
rect 2982 3010 3010 4495
rect 3766 4242 3794 4774
rect 3934 4662 4130 4690
rect 3934 4521 3962 4662
rect 3934 4495 3935 4521
rect 3961 4495 3962 4521
rect 3934 4489 3962 4495
rect 3990 4577 4018 4583
rect 3990 4551 3991 4577
rect 4017 4551 4018 4577
rect 3990 4522 4018 4551
rect 3990 4489 4018 4494
rect 4046 4578 4074 4583
rect 3822 4466 3850 4471
rect 3822 4419 3850 4438
rect 3990 4410 4018 4415
rect 4046 4410 4074 4550
rect 3990 4409 4074 4410
rect 3990 4383 3991 4409
rect 4017 4383 4074 4409
rect 3990 4382 4074 4383
rect 3990 4377 4018 4382
rect 3840 4326 3972 4331
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3840 4293 3972 4298
rect 3766 4209 3794 4214
rect 3094 4018 3122 4023
rect 3094 3793 3122 3990
rect 4102 3850 4130 4662
rect 4158 4522 4186 4527
rect 4158 4074 4186 4494
rect 4214 4466 4242 4887
rect 4270 4857 4298 4863
rect 4270 4831 4271 4857
rect 4297 4831 4298 4857
rect 4270 4578 4298 4831
rect 4270 4545 4298 4550
rect 4326 4802 4354 4807
rect 4382 4802 4410 5279
rect 5110 5305 5138 6007
rect 5558 6034 5586 6454
rect 5894 6817 5922 6823
rect 5894 6791 5895 6817
rect 5921 6791 5922 6817
rect 5894 6202 5922 6791
rect 6958 6817 6986 6823
rect 6958 6791 6959 6817
rect 6985 6791 6986 6817
rect 5996 6678 6128 6683
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 5996 6645 6128 6650
rect 6454 6538 6482 6543
rect 6454 6491 6482 6510
rect 6846 6538 6874 6543
rect 5894 6169 5922 6174
rect 5558 6001 5586 6006
rect 5614 6089 5642 6095
rect 5614 6063 5615 6089
rect 5641 6063 5642 6089
rect 5614 5754 5642 6063
rect 5614 5721 5642 5726
rect 5894 6089 5922 6095
rect 5894 6063 5895 6089
rect 5921 6063 5922 6089
rect 5782 5697 5810 5703
rect 5782 5671 5783 5697
rect 5809 5671 5810 5697
rect 5782 5362 5810 5671
rect 5894 5362 5922 6063
rect 5996 5894 6128 5899
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 5996 5861 6128 5866
rect 6230 5810 6258 5815
rect 6230 5809 6314 5810
rect 6230 5783 6231 5809
rect 6257 5783 6314 5809
rect 6230 5782 6314 5783
rect 6230 5777 6258 5782
rect 6118 5697 6146 5703
rect 6118 5671 6119 5697
rect 6145 5671 6146 5697
rect 5950 5642 5978 5647
rect 5950 5641 6034 5642
rect 5950 5615 5951 5641
rect 5977 5615 6034 5641
rect 5950 5614 6034 5615
rect 5950 5609 5978 5614
rect 5950 5362 5978 5367
rect 5782 5361 5978 5362
rect 5782 5335 5951 5361
rect 5977 5335 5978 5361
rect 5782 5334 5978 5335
rect 5950 5329 5978 5334
rect 5110 5279 5111 5305
rect 5137 5279 5138 5305
rect 5110 5273 5138 5279
rect 6006 5194 6034 5614
rect 5894 5166 6034 5194
rect 6118 5194 6146 5671
rect 4326 4801 4410 4802
rect 4326 4775 4327 4801
rect 4353 4775 4410 4801
rect 4326 4774 4410 4775
rect 5278 4913 5306 4919
rect 5278 4887 5279 4913
rect 5305 4887 5306 4913
rect 4326 4521 4354 4774
rect 4918 4718 5050 4723
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 4918 4685 5050 4690
rect 4326 4495 4327 4521
rect 4353 4495 4354 4521
rect 4326 4489 4354 4495
rect 5222 4521 5250 4527
rect 5222 4495 5223 4521
rect 5249 4495 5250 4521
rect 4214 4214 4242 4438
rect 4438 4466 4466 4471
rect 4438 4419 4466 4438
rect 4494 4410 4522 4415
rect 4494 4363 4522 4382
rect 4214 4186 4354 4214
rect 4158 4041 4186 4046
rect 4102 3803 4130 3822
rect 3094 3767 3095 3793
rect 3121 3767 3122 3793
rect 3094 3761 3122 3767
rect 3934 3626 3962 3631
rect 3766 3625 3962 3626
rect 3766 3599 3935 3625
rect 3961 3599 3962 3625
rect 3766 3598 3962 3599
rect 3318 3345 3346 3351
rect 3318 3319 3319 3345
rect 3345 3319 3346 3345
rect 3318 3290 3346 3319
rect 3318 3122 3346 3262
rect 3374 3290 3402 3295
rect 3766 3290 3794 3598
rect 3934 3593 3962 3598
rect 4046 3625 4074 3631
rect 4046 3599 4047 3625
rect 4073 3599 4074 3625
rect 3840 3542 3972 3547
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3840 3509 3972 3514
rect 3374 3289 3794 3290
rect 3374 3263 3375 3289
rect 3401 3263 3794 3289
rect 3374 3262 3794 3263
rect 4046 3290 4074 3599
rect 4102 3625 4130 3631
rect 4102 3599 4103 3625
rect 4129 3599 4130 3625
rect 4102 3346 4130 3599
rect 4102 3313 4130 3318
rect 3374 3257 3402 3262
rect 3430 3122 3458 3262
rect 4046 3257 4074 3262
rect 4214 3233 4242 3239
rect 4214 3207 4215 3233
rect 4241 3207 4242 3233
rect 3318 3094 3402 3122
rect 3430 3094 3514 3122
rect 2982 2977 3010 2982
rect 2590 2809 2618 2814
rect 2590 2618 2618 2623
rect 2590 2571 2618 2590
rect 3318 2562 3346 2567
rect 3318 2515 3346 2534
rect 3038 2449 3066 2455
rect 3038 2423 3039 2449
rect 3065 2423 3066 2449
rect 2762 2366 2894 2371
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2762 2333 2894 2338
rect 2422 2226 2450 2231
rect 2422 2225 2674 2226
rect 2422 2199 2423 2225
rect 2449 2199 2674 2225
rect 2422 2198 2674 2199
rect 2422 2193 2450 2198
rect 2366 1731 2394 1750
rect 2478 1722 2506 1727
rect 2422 1721 2506 1722
rect 2422 1695 2479 1721
rect 2505 1695 2506 1721
rect 2422 1694 2506 1695
rect 2422 1666 2450 1694
rect 2478 1689 2506 1694
rect 2310 1638 2450 1666
rect 2646 490 2674 2198
rect 2762 1582 2894 1587
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2762 1549 2894 1554
rect 2254 462 2394 490
rect 2646 462 2730 490
rect 2366 400 2394 462
rect 2702 400 2730 462
rect 3038 400 3066 2423
rect 3206 2225 3234 2231
rect 3206 2199 3207 2225
rect 3233 2199 3234 2225
rect 3206 1722 3234 2199
rect 3374 2226 3402 3094
rect 3430 2953 3458 2959
rect 3430 2927 3431 2953
rect 3457 2927 3458 2953
rect 3430 2505 3458 2927
rect 3430 2479 3431 2505
rect 3457 2479 3458 2505
rect 3430 2473 3458 2479
rect 3486 2394 3514 3094
rect 4158 3010 4186 3015
rect 4046 3009 4186 3010
rect 4046 2983 4159 3009
rect 4185 2983 4186 3009
rect 4046 2982 4186 2983
rect 3598 2954 3626 2959
rect 3598 2907 3626 2926
rect 3840 2758 3972 2763
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3840 2725 3972 2730
rect 4046 2674 4074 2982
rect 4158 2977 4186 2982
rect 4214 2674 4242 3207
rect 4270 3010 4298 4186
rect 4326 4129 4354 4186
rect 4326 4103 4327 4129
rect 4353 4103 4354 4129
rect 4326 4097 4354 4103
rect 4606 4074 4634 4079
rect 4494 4073 4634 4074
rect 4494 4047 4607 4073
rect 4633 4047 4634 4073
rect 4494 4046 4634 4047
rect 4326 3850 4354 3855
rect 4326 3793 4354 3822
rect 4494 3849 4522 4046
rect 4606 4041 4634 4046
rect 4774 4074 4802 4079
rect 4494 3823 4495 3849
rect 4521 3823 4522 3849
rect 4494 3817 4522 3823
rect 4774 3849 4802 4046
rect 4918 3934 5050 3939
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 4918 3901 5050 3906
rect 4774 3823 4775 3849
rect 4801 3823 4802 3849
rect 4774 3817 4802 3823
rect 4326 3767 4327 3793
rect 4353 3767 4354 3793
rect 4326 3761 4354 3767
rect 4382 3794 4410 3799
rect 4382 3793 4466 3794
rect 4382 3767 4383 3793
rect 4409 3767 4466 3793
rect 4382 3766 4466 3767
rect 4382 3761 4410 3766
rect 4326 3402 4354 3407
rect 4326 3066 4354 3374
rect 4382 3346 4410 3351
rect 4382 3299 4410 3318
rect 4438 3290 4466 3766
rect 4830 3681 4858 3687
rect 4830 3655 4831 3681
rect 4857 3655 4858 3681
rect 4830 3514 4858 3655
rect 4662 3486 4858 3514
rect 4662 3290 4690 3486
rect 4438 3289 4690 3290
rect 4438 3263 4663 3289
rect 4689 3263 4690 3289
rect 4438 3262 4690 3263
rect 4382 3066 4410 3071
rect 4326 3065 4410 3066
rect 4326 3039 4383 3065
rect 4409 3039 4410 3065
rect 4326 3038 4410 3039
rect 4270 2982 4354 3010
rect 3934 2646 4074 2674
rect 4102 2646 4242 2674
rect 3598 2618 3626 2623
rect 3598 2562 3626 2590
rect 3766 2562 3794 2567
rect 3598 2561 3738 2562
rect 3598 2535 3599 2561
rect 3625 2535 3738 2561
rect 3598 2534 3738 2535
rect 3598 2529 3626 2534
rect 3374 2193 3402 2198
rect 3430 2366 3514 2394
rect 3542 2506 3570 2511
rect 3374 1890 3402 1895
rect 3430 1890 3458 2366
rect 3486 2170 3514 2175
rect 3486 2123 3514 2142
rect 3402 1862 3458 1890
rect 3542 2113 3570 2478
rect 3542 2087 3543 2113
rect 3569 2087 3570 2113
rect 3374 1857 3402 1862
rect 3206 1689 3234 1694
rect 3374 1778 3402 1783
rect 3374 400 3402 1750
rect 3542 1721 3570 2087
rect 3598 2114 3626 2119
rect 3598 1777 3626 2086
rect 3598 1751 3599 1777
rect 3625 1751 3626 1777
rect 3598 1745 3626 1751
rect 3542 1695 3543 1721
rect 3569 1695 3570 1721
rect 3542 1689 3570 1695
rect 3710 400 3738 2534
rect 3766 1666 3794 2534
rect 3934 2505 3962 2646
rect 3934 2479 3935 2505
rect 3961 2479 3962 2505
rect 3934 2473 3962 2479
rect 4046 2562 4074 2567
rect 3840 1974 3972 1979
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3840 1941 3972 1946
rect 4046 1833 4074 2534
rect 4046 1807 4047 1833
rect 4073 1807 4074 1833
rect 4046 1801 4074 1807
rect 4102 1721 4130 2646
rect 4158 2562 4186 2567
rect 4326 2562 4354 2982
rect 4158 2561 4354 2562
rect 4158 2535 4159 2561
rect 4185 2535 4354 2561
rect 4158 2534 4354 2535
rect 4158 2529 4186 2534
rect 4382 2506 4410 3038
rect 4214 2478 4410 2506
rect 4214 2338 4242 2478
rect 4662 2450 4690 3262
rect 4718 3346 4746 3351
rect 4718 2505 4746 3318
rect 4918 3150 5050 3155
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 4918 3117 5050 3122
rect 5054 2897 5082 2903
rect 5054 2871 5055 2897
rect 5081 2871 5082 2897
rect 4718 2479 4719 2505
rect 4745 2479 4746 2505
rect 4718 2473 4746 2479
rect 4774 2618 4802 2623
rect 4662 2417 4690 2422
rect 4158 2310 4242 2338
rect 4158 1777 4186 2310
rect 4438 2225 4466 2231
rect 4438 2199 4439 2225
rect 4465 2199 4466 2225
rect 4438 2002 4466 2199
rect 4438 1969 4466 1974
rect 4494 2169 4522 2175
rect 4494 2143 4495 2169
rect 4521 2143 4522 2169
rect 4494 1890 4522 2143
rect 4494 1857 4522 1862
rect 4158 1751 4159 1777
rect 4185 1751 4186 1777
rect 4158 1745 4186 1751
rect 4382 1778 4410 1783
rect 4774 1778 4802 2590
rect 5054 2450 5082 2871
rect 5166 2562 5194 2567
rect 5222 2562 5250 4495
rect 5278 4130 5306 4887
rect 5502 4857 5530 4863
rect 5502 4831 5503 4857
rect 5529 4831 5530 4857
rect 5446 4521 5474 4527
rect 5446 4495 5447 4521
rect 5473 4495 5474 4521
rect 5334 4130 5362 4135
rect 5278 4129 5362 4130
rect 5278 4103 5335 4129
rect 5361 4103 5362 4129
rect 5278 4102 5362 4103
rect 5278 3849 5306 4102
rect 5334 4097 5362 4102
rect 5278 3823 5279 3849
rect 5305 3823 5306 3849
rect 5278 3346 5306 3823
rect 5278 3313 5306 3318
rect 5390 2897 5418 2903
rect 5390 2871 5391 2897
rect 5417 2871 5418 2897
rect 5222 2534 5306 2562
rect 5166 2515 5194 2534
rect 5278 2506 5306 2534
rect 5278 2473 5306 2478
rect 5054 2422 5250 2450
rect 4918 2366 5050 2371
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 4918 2333 5050 2338
rect 5110 2226 5138 2231
rect 5110 2225 5194 2226
rect 5110 2199 5111 2225
rect 5137 2199 5194 2225
rect 5110 2198 5194 2199
rect 5110 2193 5138 2198
rect 4830 2170 4858 2175
rect 4830 2169 5026 2170
rect 4830 2143 4831 2169
rect 4857 2143 5026 2169
rect 4830 2142 5026 2143
rect 4830 2137 4858 2142
rect 4830 1778 4858 1783
rect 4102 1695 4103 1721
rect 4129 1695 4130 1721
rect 4102 1689 4130 1695
rect 3766 1638 4074 1666
rect 4046 400 4074 1638
rect 4382 400 4410 1750
rect 4718 1777 4858 1778
rect 4718 1751 4831 1777
rect 4857 1751 4858 1777
rect 4718 1750 4858 1751
rect 4718 400 4746 1750
rect 4830 1745 4858 1750
rect 4998 1721 5026 2142
rect 5054 2114 5082 2119
rect 5054 2067 5082 2086
rect 4998 1695 4999 1721
rect 5025 1695 5026 1721
rect 4998 1689 5026 1695
rect 5166 1721 5194 2198
rect 5222 1778 5250 2422
rect 5278 1778 5306 1783
rect 5222 1777 5306 1778
rect 5222 1751 5279 1777
rect 5305 1751 5306 1777
rect 5222 1750 5306 1751
rect 5166 1695 5167 1721
rect 5193 1695 5194 1721
rect 5166 1689 5194 1695
rect 4918 1582 5050 1587
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 4918 1549 5050 1554
rect 5278 1498 5306 1750
rect 5054 1470 5306 1498
rect 5390 1554 5418 2871
rect 5446 2114 5474 4495
rect 5502 4466 5530 4831
rect 5670 4577 5698 4583
rect 5670 4551 5671 4577
rect 5697 4551 5698 4577
rect 5502 4465 5642 4466
rect 5502 4439 5503 4465
rect 5529 4439 5642 4465
rect 5502 4438 5642 4439
rect 5502 4433 5530 4438
rect 5502 4242 5530 4247
rect 5502 2449 5530 4214
rect 5614 4073 5642 4438
rect 5614 4047 5615 4073
rect 5641 4047 5642 4073
rect 5614 4041 5642 4047
rect 5558 3850 5586 3855
rect 5558 3737 5586 3822
rect 5558 3711 5559 3737
rect 5585 3711 5586 3737
rect 5558 3705 5586 3711
rect 5614 3793 5642 3799
rect 5614 3767 5615 3793
rect 5641 3767 5642 3793
rect 5614 3066 5642 3767
rect 5670 3402 5698 4551
rect 5838 4410 5866 4415
rect 5894 4410 5922 5166
rect 6118 5161 6146 5166
rect 5996 5110 6128 5115
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 5996 5077 6128 5082
rect 6286 5025 6314 5782
rect 6790 5754 6818 5759
rect 6790 5707 6818 5726
rect 6342 5698 6370 5703
rect 6454 5698 6482 5703
rect 6342 5697 6426 5698
rect 6342 5671 6343 5697
rect 6369 5671 6426 5697
rect 6342 5670 6426 5671
rect 6342 5665 6370 5670
rect 6342 5586 6370 5591
rect 6342 5539 6370 5558
rect 6286 4999 6287 5025
rect 6313 4999 6314 5025
rect 6286 4634 6314 4999
rect 6398 4914 6426 5670
rect 6454 5025 6482 5670
rect 6734 5698 6762 5703
rect 6734 5651 6762 5670
rect 6846 5697 6874 6510
rect 6958 6482 6986 6791
rect 8152 6678 8284 6683
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8152 6645 8284 6650
rect 8190 6537 8218 6543
rect 8190 6511 8191 6537
rect 8217 6511 8218 6537
rect 6958 6449 6986 6454
rect 7686 6482 7714 6487
rect 7714 6454 7770 6482
rect 7686 6435 7714 6454
rect 7074 6286 7206 6291
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7074 6253 7206 6258
rect 7238 6202 7266 6207
rect 6846 5671 6847 5697
rect 6873 5671 6874 5697
rect 6846 5665 6874 5671
rect 6902 6090 6930 6095
rect 6454 4999 6455 5025
rect 6481 4999 6482 5025
rect 6454 4993 6482 4999
rect 6454 4914 6482 4919
rect 6398 4913 6482 4914
rect 6398 4887 6455 4913
rect 6481 4887 6482 4913
rect 6398 4886 6482 4887
rect 6286 4601 6314 4606
rect 6230 4522 6258 4527
rect 6230 4475 6258 4494
rect 6454 4522 6482 4886
rect 6846 4914 6874 4919
rect 6846 4867 6874 4886
rect 6678 4802 6706 4807
rect 6678 4801 6762 4802
rect 6678 4775 6679 4801
rect 6705 4775 6762 4801
rect 6678 4774 6762 4775
rect 6678 4769 6706 4774
rect 6454 4489 6482 4494
rect 6510 4577 6538 4583
rect 6510 4551 6511 4577
rect 6537 4551 6538 4577
rect 5866 4382 5922 4410
rect 6174 4465 6202 4471
rect 6174 4439 6175 4465
rect 6201 4439 6202 4465
rect 5838 4185 5866 4382
rect 5996 4326 6128 4331
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 5996 4293 6128 4298
rect 6174 4214 6202 4439
rect 6174 4186 6258 4214
rect 5838 4159 5839 4185
rect 5865 4159 5866 4185
rect 5838 4153 5866 4159
rect 5950 3850 5978 3855
rect 5950 3803 5978 3822
rect 5996 3542 6128 3547
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 5996 3509 6128 3514
rect 5670 3369 5698 3374
rect 5894 3066 5922 3071
rect 5614 3065 5922 3066
rect 5614 3039 5895 3065
rect 5921 3039 5922 3065
rect 5614 3038 5922 3039
rect 5894 3033 5922 3038
rect 5502 2423 5503 2449
rect 5529 2423 5530 2449
rect 5502 2417 5530 2423
rect 5726 2897 5754 2903
rect 5726 2871 5727 2897
rect 5753 2871 5754 2897
rect 5446 2081 5474 2086
rect 5614 1777 5642 1783
rect 5614 1751 5615 1777
rect 5641 1751 5642 1777
rect 5502 1722 5530 1727
rect 5502 1675 5530 1694
rect 5614 1554 5642 1751
rect 5726 1778 5754 2871
rect 5996 2758 6128 2763
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 5996 2725 6128 2730
rect 6230 2674 6258 4186
rect 6510 4074 6538 4551
rect 6678 4577 6706 4583
rect 6678 4551 6679 4577
rect 6705 4551 6706 4577
rect 6678 4130 6706 4551
rect 6734 4241 6762 4774
rect 6734 4215 6735 4241
rect 6761 4215 6762 4241
rect 6734 4209 6762 4215
rect 6790 4801 6818 4807
rect 6790 4775 6791 4801
rect 6817 4775 6818 4801
rect 6790 4130 6818 4775
rect 6902 4634 6930 6062
rect 7014 6034 7042 6039
rect 6958 5585 6986 5591
rect 6958 5559 6959 5585
rect 6985 5559 6986 5585
rect 6958 5250 6986 5559
rect 6958 4914 6986 5222
rect 6958 4881 6986 4886
rect 7014 4913 7042 6006
rect 7238 5753 7266 6174
rect 7238 5727 7239 5753
rect 7265 5727 7266 5753
rect 7238 5721 7266 5727
rect 7294 5697 7322 5703
rect 7294 5671 7295 5697
rect 7321 5671 7322 5697
rect 7182 5642 7210 5647
rect 7182 5595 7210 5614
rect 7294 5586 7322 5671
rect 7462 5698 7490 5703
rect 7686 5698 7714 5703
rect 7462 5697 7714 5698
rect 7462 5671 7463 5697
rect 7489 5671 7687 5697
rect 7713 5671 7714 5697
rect 7462 5670 7714 5671
rect 7462 5665 7490 5670
rect 7686 5665 7714 5670
rect 7742 5697 7770 6454
rect 8190 6090 8218 6511
rect 8470 6538 8498 6543
rect 8470 6481 8498 6510
rect 8470 6455 8471 6481
rect 8497 6455 8498 6481
rect 8470 6449 8498 6455
rect 9030 6426 9058 6431
rect 9030 6379 9058 6398
rect 9230 6286 9362 6291
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9230 6253 9362 6258
rect 8918 6146 8946 6151
rect 8190 6057 8218 6062
rect 8750 6145 8946 6146
rect 8750 6119 8919 6145
rect 8945 6119 8946 6145
rect 8750 6118 8946 6119
rect 8152 5894 8284 5899
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8152 5861 8284 5866
rect 7742 5671 7743 5697
rect 7769 5671 7770 5697
rect 7742 5665 7770 5671
rect 8470 5697 8498 5703
rect 8470 5671 8471 5697
rect 8497 5671 8498 5697
rect 7294 5553 7322 5558
rect 7630 5586 7658 5591
rect 7630 5539 7658 5558
rect 7854 5585 7882 5591
rect 7854 5559 7855 5585
rect 7881 5559 7882 5585
rect 7074 5502 7206 5507
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7074 5469 7206 5474
rect 7742 5250 7770 5255
rect 7854 5250 7882 5559
rect 7910 5362 7938 5367
rect 7910 5315 7938 5334
rect 7770 5222 7882 5250
rect 7742 5203 7770 5222
rect 8152 5110 8284 5115
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8152 5077 8284 5082
rect 8470 4969 8498 5671
rect 8470 4943 8471 4969
rect 8497 4943 8498 4969
rect 8470 4937 8498 4943
rect 7014 4887 7015 4913
rect 7041 4887 7042 4913
rect 7014 4881 7042 4887
rect 7406 4857 7434 4863
rect 7406 4831 7407 4857
rect 7433 4831 7434 4857
rect 7074 4718 7206 4723
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7074 4685 7206 4690
rect 7014 4634 7042 4639
rect 6902 4633 7042 4634
rect 6902 4607 7015 4633
rect 7041 4607 7042 4633
rect 6902 4606 7042 4607
rect 7014 4601 7042 4606
rect 7182 4634 7210 4639
rect 7126 4578 7154 4583
rect 6958 4521 6986 4527
rect 6958 4495 6959 4521
rect 6985 4495 6986 4521
rect 6678 4102 6818 4130
rect 6510 4041 6538 4046
rect 6790 4018 6818 4102
rect 6846 4466 6874 4471
rect 6846 4073 6874 4438
rect 6958 4410 6986 4495
rect 7126 4521 7154 4550
rect 7126 4495 7127 4521
rect 7153 4495 7154 4521
rect 7126 4489 7154 4495
rect 7182 4521 7210 4606
rect 7182 4495 7183 4521
rect 7209 4495 7210 4521
rect 6958 4377 6986 4382
rect 6958 4298 6986 4303
rect 6958 4214 6986 4270
rect 7182 4214 7210 4495
rect 7350 4522 7378 4527
rect 7350 4475 7378 4494
rect 7406 4298 7434 4831
rect 8750 4578 8778 6118
rect 8918 6113 8946 6118
rect 9086 6089 9114 6095
rect 9086 6063 9087 6089
rect 9113 6063 9114 6089
rect 8806 6034 8834 6039
rect 9086 6034 9114 6063
rect 8806 6033 9114 6034
rect 8806 6007 8807 6033
rect 8833 6007 9114 6033
rect 8806 6006 9114 6007
rect 8806 6001 8834 6006
rect 9086 5754 9114 6006
rect 9086 5721 9114 5726
rect 9030 5641 9058 5647
rect 9030 5615 9031 5641
rect 9057 5615 9058 5641
rect 9030 5418 9058 5615
rect 9230 5502 9362 5507
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9230 5469 9362 5474
rect 9030 5385 9058 5390
rect 8918 5362 8946 5367
rect 8918 5315 8946 5334
rect 9086 5305 9114 5311
rect 9086 5279 9087 5305
rect 9113 5279 9114 5305
rect 8806 5250 8834 5255
rect 9086 5250 9114 5279
rect 8806 5249 9114 5250
rect 8806 5223 8807 5249
rect 8833 5223 9114 5249
rect 8806 5222 9114 5223
rect 8806 5217 8834 5222
rect 8918 5138 8946 5143
rect 8918 4857 8946 5110
rect 9086 5082 9114 5222
rect 9086 5049 9114 5054
rect 8918 4831 8919 4857
rect 8945 4831 8946 4857
rect 8918 4825 8946 4831
rect 9086 4857 9114 4863
rect 9086 4831 9087 4857
rect 9113 4831 9114 4857
rect 8806 4802 8834 4807
rect 8806 4755 8834 4774
rect 9086 4802 9114 4831
rect 9086 4769 9114 4774
rect 9230 4718 9362 4723
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9230 4685 9362 4690
rect 8750 4545 8778 4550
rect 8918 4577 8946 4583
rect 8918 4551 8919 4577
rect 8945 4551 8946 4577
rect 8918 4522 8946 4551
rect 8918 4489 8946 4494
rect 9086 4521 9114 4527
rect 9086 4495 9087 4521
rect 9113 4495 9114 4521
rect 8806 4465 8834 4471
rect 8806 4439 8807 4465
rect 8833 4439 8834 4465
rect 8806 4410 8834 4439
rect 8806 4377 8834 4382
rect 9086 4410 9114 4495
rect 9086 4377 9114 4382
rect 8152 4326 8284 4331
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8152 4293 8284 4298
rect 7406 4265 7434 4270
rect 6902 4186 6986 4214
rect 7014 4186 7210 4214
rect 6902 4185 6930 4186
rect 6902 4159 6903 4185
rect 6929 4159 6930 4185
rect 6902 4153 6930 4159
rect 7014 4129 7042 4186
rect 7014 4103 7015 4129
rect 7041 4103 7042 4129
rect 7014 4097 7042 4103
rect 6846 4047 6847 4073
rect 6873 4047 6874 4073
rect 6846 4041 6874 4047
rect 7126 4074 7154 4079
rect 7126 4027 7154 4046
rect 7182 4073 7210 4079
rect 7182 4047 7183 4073
rect 7209 4047 7210 4073
rect 6790 3985 6818 3990
rect 7182 4018 7210 4047
rect 8582 4074 8610 4079
rect 8582 4027 8610 4046
rect 8750 4073 8778 4079
rect 8750 4047 8751 4073
rect 8777 4047 8778 4073
rect 7182 3985 7210 3990
rect 7074 3934 7206 3939
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7074 3901 7206 3906
rect 6454 3794 6482 3799
rect 6454 3747 6482 3766
rect 7462 3794 7490 3799
rect 8470 3794 8498 3799
rect 7462 3793 7546 3794
rect 7462 3767 7463 3793
rect 7489 3767 7546 3793
rect 7462 3766 7546 3767
rect 7462 3761 7490 3766
rect 6678 3738 6706 3743
rect 6566 3737 6706 3738
rect 6566 3711 6679 3737
rect 6705 3711 6706 3737
rect 6566 3710 6706 3711
rect 6006 2646 6258 2674
rect 6398 3009 6426 3015
rect 6398 2983 6399 3009
rect 6425 2983 6426 3009
rect 6006 2505 6034 2646
rect 6230 2562 6258 2567
rect 6230 2515 6258 2534
rect 6006 2479 6007 2505
rect 6033 2479 6034 2505
rect 6006 2473 6034 2479
rect 6398 2282 6426 2983
rect 6398 2249 6426 2254
rect 6118 2226 6146 2231
rect 6118 2179 6146 2198
rect 5726 1745 5754 1750
rect 5838 2002 5866 2007
rect 5838 1721 5866 1974
rect 5996 1974 6128 1979
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 5996 1941 6128 1946
rect 5950 1778 5978 1783
rect 5950 1731 5978 1750
rect 6398 1778 6426 1783
rect 5838 1695 5839 1721
rect 5865 1695 5866 1721
rect 5838 1689 5866 1695
rect 6062 1722 6090 1727
rect 5390 1526 5642 1554
rect 5726 1666 5754 1671
rect 5054 400 5082 1470
rect 5390 400 5418 1526
rect 5726 400 5754 1638
rect 6062 400 6090 1694
rect 6174 1666 6202 1671
rect 6174 1619 6202 1638
rect 6398 400 6426 1750
rect 6566 1721 6594 3710
rect 6678 3705 6706 3710
rect 7074 3150 7206 3155
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7074 3117 7206 3122
rect 7406 3009 7434 3015
rect 7406 2983 7407 3009
rect 7433 2983 7434 3009
rect 6678 2953 6706 2959
rect 6678 2927 6679 2953
rect 6705 2927 6706 2953
rect 6678 2338 6706 2927
rect 7074 2366 7206 2371
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 6678 2310 6986 2338
rect 7074 2333 7206 2338
rect 6678 2169 6706 2175
rect 6678 2143 6679 2169
rect 6705 2143 6706 2169
rect 6678 2114 6706 2143
rect 6678 2081 6706 2086
rect 6902 2113 6930 2119
rect 6902 2087 6903 2113
rect 6929 2087 6930 2113
rect 6566 1695 6567 1721
rect 6593 1695 6594 1721
rect 6566 1689 6594 1695
rect 6678 1778 6706 1783
rect 6902 1778 6930 2087
rect 6678 1777 6930 1778
rect 6678 1751 6679 1777
rect 6705 1751 6930 1777
rect 6678 1750 6930 1751
rect 6678 1722 6706 1750
rect 6958 1722 6986 2310
rect 7238 2282 7266 2287
rect 7406 2282 7434 2983
rect 7518 2730 7546 3766
rect 7798 3737 7826 3743
rect 7798 3711 7799 3737
rect 7825 3711 7826 3737
rect 7742 2953 7770 2959
rect 7742 2927 7743 2953
rect 7769 2927 7770 2953
rect 7518 2702 7602 2730
rect 7462 2562 7490 2567
rect 7462 2561 7546 2562
rect 7462 2535 7463 2561
rect 7489 2535 7546 2561
rect 7462 2534 7546 2535
rect 7462 2529 7490 2534
rect 7462 2282 7490 2287
rect 7406 2254 7462 2282
rect 7126 2113 7154 2119
rect 7126 2087 7127 2113
rect 7153 2087 7154 2113
rect 7014 1778 7042 1783
rect 7126 1778 7154 2087
rect 7042 1750 7154 1778
rect 7014 1731 7042 1750
rect 6678 1689 6706 1694
rect 6902 1694 6986 1722
rect 7238 1721 7266 2254
rect 7462 2249 7490 2254
rect 7238 1695 7239 1721
rect 7265 1695 7266 1721
rect 6902 1665 6930 1694
rect 7238 1689 7266 1695
rect 7350 2113 7378 2119
rect 7350 2087 7351 2113
rect 7377 2087 7378 2113
rect 7350 1777 7378 2087
rect 7350 1751 7351 1777
rect 7377 1751 7378 1777
rect 6902 1639 6903 1665
rect 6929 1639 6930 1665
rect 6902 1633 6930 1639
rect 7074 1582 7206 1587
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7074 1549 7206 1554
rect 7350 1274 7378 1751
rect 6734 1246 7378 1274
rect 7406 1722 7434 1727
rect 7518 1722 7546 2534
rect 7434 1694 7546 1722
rect 7574 1721 7602 2702
rect 7742 2506 7770 2927
rect 7798 2674 7826 3711
rect 8152 3542 8284 3547
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8152 3509 8284 3514
rect 8152 2758 8284 2763
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8152 2725 8284 2730
rect 7798 2646 8050 2674
rect 7742 2473 7770 2478
rect 7798 2449 7826 2455
rect 7798 2423 7799 2449
rect 7825 2423 7826 2449
rect 7798 2226 7826 2423
rect 7854 2282 7882 2287
rect 7854 2235 7882 2254
rect 7574 1695 7575 1721
rect 7601 1695 7602 1721
rect 6734 400 6762 1246
rect 7406 1162 7434 1694
rect 7574 1689 7602 1695
rect 7630 2198 7826 2226
rect 7630 1778 7658 2198
rect 7966 2169 7994 2175
rect 7966 2143 7967 2169
rect 7993 2143 7994 2169
rect 7742 2114 7770 2119
rect 7966 2114 7994 2143
rect 7742 2113 7994 2114
rect 7742 2087 7743 2113
rect 7769 2087 7994 2113
rect 7742 2086 7994 2087
rect 7630 1610 7658 1750
rect 7686 1777 7714 1783
rect 7686 1751 7687 1777
rect 7713 1751 7714 1777
rect 7686 1722 7714 1751
rect 7686 1689 7714 1694
rect 7070 1134 7434 1162
rect 7518 1582 7658 1610
rect 7070 400 7098 1134
rect 7518 1106 7546 1582
rect 7406 1078 7546 1106
rect 7406 400 7434 1078
rect 7742 400 7770 2086
rect 8022 2058 8050 2646
rect 8134 2562 8162 2567
rect 7910 2030 8050 2058
rect 8078 2561 8162 2562
rect 8078 2535 8135 2561
rect 8161 2535 8162 2561
rect 8078 2534 8162 2535
rect 7910 1721 7938 2030
rect 8078 1890 8106 2534
rect 8134 2529 8162 2534
rect 8358 2561 8386 2567
rect 8358 2535 8359 2561
rect 8385 2535 8386 2561
rect 8358 2450 8386 2535
rect 8358 2417 8386 2422
rect 8246 2226 8274 2231
rect 8246 2179 8274 2198
rect 8414 2170 8442 2175
rect 8414 2123 8442 2142
rect 8152 1974 8284 1979
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8152 1941 8284 1946
rect 8078 1862 8162 1890
rect 8022 1778 8050 1783
rect 8022 1731 8050 1750
rect 7910 1695 7911 1721
rect 7937 1695 7938 1721
rect 7910 1689 7938 1695
rect 8134 1722 8162 1862
rect 8134 1610 8162 1694
rect 8470 1721 8498 3766
rect 8750 3738 8778 4047
rect 9086 4074 9114 4079
rect 9114 4046 9170 4074
rect 9086 4027 9114 4046
rect 8918 4018 8946 4023
rect 8918 3971 8946 3990
rect 9142 3849 9170 4046
rect 9230 3934 9362 3939
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9230 3901 9362 3906
rect 9142 3823 9143 3849
rect 9169 3823 9170 3849
rect 9142 3817 9170 3823
rect 8862 3738 8890 3743
rect 8750 3710 8862 3738
rect 8862 3691 8890 3710
rect 9086 3233 9114 3239
rect 9086 3207 9087 3233
rect 9113 3207 9114 3233
rect 9086 3066 9114 3207
rect 9230 3150 9362 3155
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9230 3117 9362 3122
rect 9086 3033 9114 3038
rect 8806 2897 8834 2903
rect 8806 2871 8807 2897
rect 8833 2871 8834 2897
rect 8582 2561 8610 2567
rect 8582 2535 8583 2561
rect 8609 2535 8610 2561
rect 8582 2170 8610 2535
rect 8582 2137 8610 2142
rect 8750 2449 8778 2455
rect 8750 2423 8751 2449
rect 8777 2423 8778 2449
rect 8750 2058 8778 2423
rect 8750 2025 8778 2030
rect 8750 1890 8778 1895
rect 8470 1695 8471 1721
rect 8497 1695 8498 1721
rect 8470 1689 8498 1695
rect 8582 1777 8610 1783
rect 8582 1751 8583 1777
rect 8609 1751 8610 1777
rect 8582 1722 8610 1751
rect 8750 1722 8778 1862
rect 8806 1778 8834 2871
rect 9142 2897 9170 2903
rect 9142 2871 9143 2897
rect 9169 2871 9170 2897
rect 9086 2562 9114 2567
rect 9142 2562 9170 2871
rect 9086 2561 9170 2562
rect 9086 2535 9087 2561
rect 9113 2535 9170 2561
rect 9086 2534 9170 2535
rect 8862 2506 8890 2511
rect 8862 2281 8890 2478
rect 8862 2255 8863 2281
rect 8889 2255 8890 2281
rect 8862 2249 8890 2255
rect 8918 2449 8946 2455
rect 8918 2423 8919 2449
rect 8945 2423 8946 2449
rect 8918 2114 8946 2423
rect 8918 2081 8946 2086
rect 8974 2450 9002 2455
rect 8974 2169 9002 2422
rect 8974 2143 8975 2169
rect 9001 2143 9002 2169
rect 8918 1778 8946 1783
rect 8806 1777 8946 1778
rect 8806 1751 8919 1777
rect 8945 1751 8946 1777
rect 8806 1750 8946 1751
rect 8750 1694 8834 1722
rect 8582 1689 8610 1694
rect 8806 1665 8834 1694
rect 8806 1639 8807 1665
rect 8833 1639 8834 1665
rect 8806 1633 8834 1639
rect 8078 1582 8162 1610
rect 8078 400 8106 1582
rect 8918 1554 8946 1750
rect 8414 1526 8946 1554
rect 8414 400 8442 1526
rect 8974 1442 9002 2143
rect 8750 1414 9002 1442
rect 9030 2170 9058 2175
rect 9030 1442 9058 2142
rect 9086 1834 9114 2534
rect 9230 2366 9362 2371
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9230 2333 9362 2338
rect 9086 1806 9450 1834
rect 9230 1582 9362 1587
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9230 1549 9362 1554
rect 9030 1414 9114 1442
rect 8750 400 8778 1414
rect 9086 400 9114 1414
rect 9422 400 9450 1806
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 5376 0 5432 400
rect 5712 0 5768 400
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
<< via2 >>
rect 1302 8358 1330 8386
rect 1078 8078 1106 8106
rect 1684 8245 1712 8246
rect 1684 8219 1685 8245
rect 1685 8219 1711 8245
rect 1711 8219 1712 8245
rect 1684 8218 1712 8219
rect 1736 8245 1764 8246
rect 1736 8219 1737 8245
rect 1737 8219 1763 8245
rect 1763 8219 1764 8245
rect 1736 8218 1764 8219
rect 1788 8245 1816 8246
rect 1788 8219 1789 8245
rect 1789 8219 1815 8245
rect 1815 8219 1816 8245
rect 1788 8218 1816 8219
rect 3840 8245 3868 8246
rect 3840 8219 3841 8245
rect 3841 8219 3867 8245
rect 3867 8219 3868 8245
rect 3840 8218 3868 8219
rect 3892 8245 3920 8246
rect 3892 8219 3893 8245
rect 3893 8219 3919 8245
rect 3919 8219 3920 8245
rect 3892 8218 3920 8219
rect 3944 8245 3972 8246
rect 3944 8219 3945 8245
rect 3945 8219 3971 8245
rect 3971 8219 3972 8245
rect 3944 8218 3972 8219
rect 4046 8134 4074 8162
rect 4662 8161 4690 8162
rect 4662 8135 4663 8161
rect 4663 8135 4689 8161
rect 4689 8135 4690 8161
rect 4662 8134 4690 8135
rect 854 7937 882 7938
rect 854 7911 855 7937
rect 855 7911 881 7937
rect 881 7911 882 7937
rect 854 7910 882 7911
rect 2762 7853 2790 7854
rect 2762 7827 2763 7853
rect 2763 7827 2789 7853
rect 2789 7827 2790 7853
rect 2762 7826 2790 7827
rect 2814 7853 2842 7854
rect 2814 7827 2815 7853
rect 2815 7827 2841 7853
rect 2841 7827 2842 7853
rect 2814 7826 2842 7827
rect 2866 7853 2894 7854
rect 2866 7827 2867 7853
rect 2867 7827 2893 7853
rect 2893 7827 2894 7853
rect 2866 7826 2894 7827
rect 5996 8245 6024 8246
rect 5996 8219 5997 8245
rect 5997 8219 6023 8245
rect 6023 8219 6024 8245
rect 5996 8218 6024 8219
rect 6048 8245 6076 8246
rect 6048 8219 6049 8245
rect 6049 8219 6075 8245
rect 6075 8219 6076 8245
rect 6048 8218 6076 8219
rect 6100 8245 6128 8246
rect 6100 8219 6101 8245
rect 6101 8219 6127 8245
rect 6127 8219 6128 8245
rect 6100 8218 6128 8219
rect 8152 8245 8180 8246
rect 8152 8219 8153 8245
rect 8153 8219 8179 8245
rect 8179 8219 8180 8245
rect 8152 8218 8180 8219
rect 8204 8245 8232 8246
rect 8204 8219 8205 8245
rect 8205 8219 8231 8245
rect 8231 8219 8232 8245
rect 8204 8218 8232 8219
rect 8256 8245 8284 8246
rect 8256 8219 8257 8245
rect 8257 8219 8283 8245
rect 8283 8219 8284 8245
rect 8256 8218 8284 8219
rect 4918 7853 4946 7854
rect 4918 7827 4919 7853
rect 4919 7827 4945 7853
rect 4945 7827 4946 7853
rect 4918 7826 4946 7827
rect 4970 7853 4998 7854
rect 4970 7827 4971 7853
rect 4971 7827 4997 7853
rect 4997 7827 4998 7853
rect 4970 7826 4998 7827
rect 5022 7853 5050 7854
rect 5022 7827 5023 7853
rect 5023 7827 5049 7853
rect 5049 7827 5050 7853
rect 5022 7826 5050 7827
rect 7074 7853 7102 7854
rect 7074 7827 7075 7853
rect 7075 7827 7101 7853
rect 7101 7827 7102 7853
rect 7074 7826 7102 7827
rect 7126 7853 7154 7854
rect 7126 7827 7127 7853
rect 7127 7827 7153 7853
rect 7153 7827 7154 7853
rect 7126 7826 7154 7827
rect 7178 7853 7206 7854
rect 7178 7827 7179 7853
rect 7179 7827 7205 7853
rect 7205 7827 7206 7853
rect 7178 7826 7206 7827
rect 9230 7853 9258 7854
rect 9230 7827 9231 7853
rect 9231 7827 9257 7853
rect 9257 7827 9258 7853
rect 9230 7826 9258 7827
rect 9282 7853 9310 7854
rect 9282 7827 9283 7853
rect 9283 7827 9309 7853
rect 9309 7827 9310 7853
rect 9282 7826 9310 7827
rect 9334 7853 9362 7854
rect 9334 7827 9335 7853
rect 9335 7827 9361 7853
rect 9361 7827 9362 7853
rect 9334 7826 9362 7827
rect 9142 7742 9170 7770
rect 854 7574 882 7602
rect 1684 7461 1712 7462
rect 1684 7435 1685 7461
rect 1685 7435 1711 7461
rect 1711 7435 1712 7461
rect 1684 7434 1712 7435
rect 1736 7461 1764 7462
rect 1736 7435 1737 7461
rect 1737 7435 1763 7461
rect 1763 7435 1764 7461
rect 1736 7434 1764 7435
rect 1788 7461 1816 7462
rect 1788 7435 1789 7461
rect 1789 7435 1815 7461
rect 1815 7435 1816 7461
rect 1788 7434 1816 7435
rect 3840 7461 3868 7462
rect 3840 7435 3841 7461
rect 3841 7435 3867 7461
rect 3867 7435 3868 7461
rect 3840 7434 3868 7435
rect 3892 7461 3920 7462
rect 3892 7435 3893 7461
rect 3893 7435 3919 7461
rect 3919 7435 3920 7461
rect 3892 7434 3920 7435
rect 3944 7461 3972 7462
rect 3944 7435 3945 7461
rect 3945 7435 3971 7461
rect 3971 7435 3972 7461
rect 3944 7434 3972 7435
rect 5996 7461 6024 7462
rect 5996 7435 5997 7461
rect 5997 7435 6023 7461
rect 6023 7435 6024 7461
rect 5996 7434 6024 7435
rect 6048 7461 6076 7462
rect 6048 7435 6049 7461
rect 6049 7435 6075 7461
rect 6075 7435 6076 7461
rect 6048 7434 6076 7435
rect 6100 7461 6128 7462
rect 6100 7435 6101 7461
rect 6101 7435 6127 7461
rect 6127 7435 6128 7461
rect 6100 7434 6128 7435
rect 8152 7461 8180 7462
rect 8152 7435 8153 7461
rect 8153 7435 8179 7461
rect 8179 7435 8180 7461
rect 8152 7434 8180 7435
rect 8204 7461 8232 7462
rect 8204 7435 8205 7461
rect 8205 7435 8231 7461
rect 8231 7435 8232 7461
rect 8204 7434 8232 7435
rect 8256 7461 8284 7462
rect 8256 7435 8257 7461
rect 8257 7435 8283 7461
rect 8283 7435 8284 7461
rect 8256 7434 8284 7435
rect 9086 7406 9114 7434
rect 854 7153 882 7154
rect 854 7127 855 7153
rect 855 7127 881 7153
rect 881 7127 882 7153
rect 854 7126 882 7127
rect 9086 7153 9114 7154
rect 9086 7127 9087 7153
rect 9087 7127 9113 7153
rect 9113 7127 9114 7153
rect 9086 7126 9114 7127
rect 2762 7069 2790 7070
rect 2762 7043 2763 7069
rect 2763 7043 2789 7069
rect 2789 7043 2790 7069
rect 2762 7042 2790 7043
rect 2814 7069 2842 7070
rect 2814 7043 2815 7069
rect 2815 7043 2841 7069
rect 2841 7043 2842 7069
rect 2814 7042 2842 7043
rect 2866 7069 2894 7070
rect 2866 7043 2867 7069
rect 2867 7043 2893 7069
rect 2893 7043 2894 7069
rect 2866 7042 2894 7043
rect 1684 6677 1712 6678
rect 1684 6651 1685 6677
rect 1685 6651 1711 6677
rect 1711 6651 1712 6677
rect 1684 6650 1712 6651
rect 1736 6677 1764 6678
rect 1736 6651 1737 6677
rect 1737 6651 1763 6677
rect 1763 6651 1764 6677
rect 1736 6650 1764 6651
rect 1788 6677 1816 6678
rect 1788 6651 1789 6677
rect 1789 6651 1815 6677
rect 1815 6651 1816 6677
rect 1788 6650 1816 6651
rect 854 6425 882 6426
rect 854 6399 855 6425
rect 855 6399 881 6425
rect 881 6399 882 6425
rect 854 6398 882 6399
rect 1022 6566 1050 6594
rect 3486 6566 3514 6594
rect 2762 6285 2790 6286
rect 2762 6259 2763 6285
rect 2763 6259 2789 6285
rect 2789 6259 2790 6285
rect 2762 6258 2790 6259
rect 2814 6285 2842 6286
rect 2814 6259 2815 6285
rect 2815 6259 2841 6285
rect 2841 6259 2842 6285
rect 2814 6258 2842 6259
rect 2866 6285 2894 6286
rect 2866 6259 2867 6285
rect 2867 6259 2893 6285
rect 2893 6259 2894 6285
rect 2866 6258 2894 6259
rect 1190 6062 1218 6090
rect 1684 5893 1712 5894
rect 1684 5867 1685 5893
rect 1685 5867 1711 5893
rect 1711 5867 1712 5893
rect 1684 5866 1712 5867
rect 1736 5893 1764 5894
rect 1736 5867 1737 5893
rect 1737 5867 1763 5893
rect 1763 5867 1764 5893
rect 1736 5866 1764 5867
rect 1788 5893 1816 5894
rect 1788 5867 1789 5893
rect 1789 5867 1815 5893
rect 1815 5867 1816 5893
rect 1788 5866 1816 5867
rect 854 5726 882 5754
rect 2982 5726 3010 5754
rect 3840 6677 3868 6678
rect 3840 6651 3841 6677
rect 3841 6651 3867 6677
rect 3867 6651 3868 6677
rect 3840 6650 3868 6651
rect 3892 6677 3920 6678
rect 3892 6651 3893 6677
rect 3893 6651 3919 6677
rect 3919 6651 3920 6677
rect 3892 6650 3920 6651
rect 3944 6677 3972 6678
rect 3944 6651 3945 6677
rect 3945 6651 3971 6677
rect 3971 6651 3972 6677
rect 3944 6650 3972 6651
rect 3990 6510 4018 6538
rect 4382 6537 4410 6538
rect 4382 6511 4383 6537
rect 4383 6511 4409 6537
rect 4409 6511 4410 6537
rect 4382 6510 4410 6511
rect 4918 7069 4946 7070
rect 4918 7043 4919 7069
rect 4919 7043 4945 7069
rect 4945 7043 4946 7069
rect 4918 7042 4946 7043
rect 4970 7069 4998 7070
rect 4970 7043 4971 7069
rect 4971 7043 4997 7069
rect 4997 7043 4998 7069
rect 4970 7042 4998 7043
rect 5022 7069 5050 7070
rect 5022 7043 5023 7069
rect 5023 7043 5049 7069
rect 5049 7043 5050 7069
rect 5022 7042 5050 7043
rect 7074 7069 7102 7070
rect 7074 7043 7075 7069
rect 7075 7043 7101 7069
rect 7101 7043 7102 7069
rect 7074 7042 7102 7043
rect 7126 7069 7154 7070
rect 7126 7043 7127 7069
rect 7127 7043 7153 7069
rect 7153 7043 7154 7069
rect 7126 7042 7154 7043
rect 7178 7069 7206 7070
rect 7178 7043 7179 7069
rect 7179 7043 7205 7069
rect 7205 7043 7206 7069
rect 7178 7042 7206 7043
rect 9230 7069 9258 7070
rect 9230 7043 9231 7069
rect 9231 7043 9257 7069
rect 9257 7043 9258 7069
rect 9230 7042 9258 7043
rect 9282 7069 9310 7070
rect 9282 7043 9283 7069
rect 9283 7043 9309 7069
rect 9309 7043 9310 7069
rect 9282 7042 9310 7043
rect 9334 7069 9362 7070
rect 9334 7043 9335 7069
rect 9335 7043 9361 7069
rect 9361 7043 9362 7069
rect 9334 7042 9362 7043
rect 4830 6510 4858 6538
rect 5110 6734 5138 6762
rect 5054 6481 5082 6482
rect 5054 6455 5055 6481
rect 5055 6455 5081 6481
rect 5081 6455 5082 6481
rect 5054 6454 5082 6455
rect 4918 6285 4946 6286
rect 4918 6259 4919 6285
rect 4919 6259 4945 6285
rect 4945 6259 4946 6285
rect 4918 6258 4946 6259
rect 4970 6285 4998 6286
rect 4970 6259 4971 6285
rect 4971 6259 4997 6285
rect 4997 6259 4998 6285
rect 4970 6258 4998 6259
rect 5022 6285 5050 6286
rect 5022 6259 5023 6285
rect 5023 6259 5049 6285
rect 5049 6259 5050 6285
rect 5022 6258 5050 6259
rect 1470 5697 1498 5698
rect 1470 5671 1471 5697
rect 1471 5671 1497 5697
rect 1497 5671 1498 5697
rect 1470 5670 1498 5671
rect 2646 5670 2674 5698
rect 1022 5446 1050 5474
rect 854 5054 882 5082
rect 2762 5501 2790 5502
rect 2762 5475 2763 5501
rect 2763 5475 2789 5501
rect 2789 5475 2790 5501
rect 2762 5474 2790 5475
rect 2814 5501 2842 5502
rect 2814 5475 2815 5501
rect 2815 5475 2841 5501
rect 2841 5475 2842 5501
rect 2814 5474 2842 5475
rect 2866 5501 2894 5502
rect 2866 5475 2867 5501
rect 2867 5475 2893 5501
rect 2893 5475 2894 5501
rect 2866 5474 2894 5475
rect 2646 5249 2674 5250
rect 2646 5223 2647 5249
rect 2647 5223 2673 5249
rect 2673 5223 2674 5249
rect 2646 5222 2674 5223
rect 1246 5054 1274 5082
rect 1684 5109 1712 5110
rect 1684 5083 1685 5109
rect 1685 5083 1711 5109
rect 1711 5083 1712 5109
rect 1684 5082 1712 5083
rect 1736 5109 1764 5110
rect 1736 5083 1737 5109
rect 1737 5083 1763 5109
rect 1763 5083 1764 5109
rect 1736 5082 1764 5083
rect 1788 5109 1816 5110
rect 1788 5083 1789 5109
rect 1789 5083 1815 5109
rect 1815 5083 1816 5109
rect 1788 5082 1816 5083
rect 3374 5054 3402 5082
rect 1022 4942 1050 4970
rect 3038 4969 3066 4970
rect 3038 4943 3039 4969
rect 3039 4943 3065 4969
rect 3065 4943 3066 4969
rect 3038 4942 3066 4943
rect 3094 4913 3122 4914
rect 3094 4887 3095 4913
rect 3095 4887 3121 4913
rect 3121 4887 3122 4913
rect 3094 4886 3122 4887
rect 3374 4913 3402 4914
rect 3374 4887 3375 4913
rect 3375 4887 3401 4913
rect 3401 4887 3402 4913
rect 3374 4886 3402 4887
rect 854 4718 882 4746
rect 854 4382 882 4410
rect 854 4073 882 4074
rect 854 4047 855 4073
rect 855 4047 881 4073
rect 881 4047 882 4073
rect 854 4046 882 4047
rect 1022 4017 1050 4018
rect 1022 3991 1023 4017
rect 1023 3991 1049 4017
rect 1049 3991 1050 4017
rect 1022 3990 1050 3991
rect 966 3822 994 3850
rect 1022 3878 1050 3906
rect 3262 4774 3290 4802
rect 3840 5893 3868 5894
rect 3840 5867 3841 5893
rect 3841 5867 3867 5893
rect 3867 5867 3868 5893
rect 3840 5866 3868 5867
rect 3892 5893 3920 5894
rect 3892 5867 3893 5893
rect 3893 5867 3919 5893
rect 3919 5867 3920 5893
rect 3892 5866 3920 5867
rect 3944 5893 3972 5894
rect 3944 5867 3945 5893
rect 3945 5867 3971 5893
rect 3971 5867 3972 5893
rect 3944 5866 3972 5867
rect 3542 5753 3570 5754
rect 3542 5727 3543 5753
rect 3543 5727 3569 5753
rect 3569 5727 3570 5753
rect 3542 5726 3570 5727
rect 4046 5726 4074 5754
rect 3710 5054 3738 5082
rect 3766 5222 3794 5250
rect 3840 5109 3868 5110
rect 3840 5083 3841 5109
rect 3841 5083 3867 5109
rect 3867 5083 3868 5109
rect 3840 5082 3868 5083
rect 3892 5109 3920 5110
rect 3892 5083 3893 5109
rect 3893 5083 3919 5109
rect 3919 5083 3920 5109
rect 3892 5082 3920 5083
rect 3944 5109 3972 5110
rect 3944 5083 3945 5109
rect 3945 5083 3971 5109
rect 3971 5083 3972 5109
rect 3944 5082 3972 5083
rect 4942 6089 4970 6090
rect 4942 6063 4943 6089
rect 4943 6063 4969 6089
rect 4969 6063 4970 6089
rect 4942 6062 4970 6063
rect 5558 6454 5586 6482
rect 5278 6089 5306 6090
rect 5278 6063 5279 6089
rect 5279 6063 5305 6089
rect 5305 6063 5306 6089
rect 5278 6062 5306 6063
rect 5502 6089 5530 6090
rect 5502 6063 5503 6089
rect 5503 6063 5529 6089
rect 5529 6063 5530 6089
rect 5502 6062 5530 6063
rect 4550 5614 4578 5642
rect 4438 5361 4466 5362
rect 4438 5335 4439 5361
rect 4439 5335 4465 5361
rect 4465 5335 4466 5361
rect 4438 5334 4466 5335
rect 4918 5501 4946 5502
rect 4918 5475 4919 5501
rect 4919 5475 4945 5501
rect 4945 5475 4946 5501
rect 4918 5474 4946 5475
rect 4970 5501 4998 5502
rect 4970 5475 4971 5501
rect 4971 5475 4997 5501
rect 4997 5475 4998 5501
rect 4970 5474 4998 5475
rect 5022 5501 5050 5502
rect 5022 5475 5023 5501
rect 5023 5475 5049 5501
rect 5049 5475 5050 5501
rect 5022 5474 5050 5475
rect 4102 4913 4130 4914
rect 4102 4887 4103 4913
rect 4103 4887 4129 4913
rect 4129 4887 4130 4913
rect 4102 4886 4130 4887
rect 3430 4774 3458 4802
rect 3766 4801 3794 4802
rect 3766 4775 3767 4801
rect 3767 4775 3793 4801
rect 3793 4775 3794 4801
rect 3766 4774 3794 4775
rect 1246 4718 1274 4746
rect 2762 4717 2790 4718
rect 2762 4691 2763 4717
rect 2763 4691 2789 4717
rect 2789 4691 2790 4717
rect 2762 4690 2790 4691
rect 2814 4717 2842 4718
rect 2814 4691 2815 4717
rect 2815 4691 2841 4717
rect 2841 4691 2842 4717
rect 2814 4690 2842 4691
rect 2866 4717 2894 4718
rect 2866 4691 2867 4717
rect 2867 4691 2893 4717
rect 2893 4691 2894 4717
rect 2866 4690 2894 4691
rect 1358 4550 1386 4578
rect 1246 4382 1274 4410
rect 1246 4046 1274 4074
rect 1684 4325 1712 4326
rect 1684 4299 1685 4325
rect 1685 4299 1711 4325
rect 1711 4299 1712 4325
rect 1684 4298 1712 4299
rect 1736 4325 1764 4326
rect 1736 4299 1737 4325
rect 1737 4299 1763 4325
rect 1763 4299 1764 4325
rect 1736 4298 1764 4299
rect 1788 4325 1816 4326
rect 1788 4299 1789 4325
rect 1789 4299 1815 4325
rect 1815 4299 1816 4325
rect 1788 4298 1816 4299
rect 2926 4577 2954 4578
rect 2926 4551 2927 4577
rect 2927 4551 2953 4577
rect 2953 4551 2954 4577
rect 2926 4550 2954 4551
rect 1190 3766 1218 3794
rect 2086 3878 2114 3906
rect 1582 3766 1610 3794
rect 1078 3710 1106 3738
rect 1806 3737 1834 3738
rect 1806 3711 1807 3737
rect 1807 3711 1833 3737
rect 1833 3711 1834 3737
rect 1806 3710 1834 3711
rect 854 3654 882 3682
rect 1470 3681 1498 3682
rect 1470 3655 1471 3681
rect 1471 3655 1497 3681
rect 1497 3655 1498 3681
rect 1470 3654 1498 3655
rect 854 3374 882 3402
rect 1022 3598 1050 3626
rect 1684 3541 1712 3542
rect 1684 3515 1685 3541
rect 1685 3515 1711 3541
rect 1711 3515 1712 3541
rect 1684 3514 1712 3515
rect 1736 3541 1764 3542
rect 1736 3515 1737 3541
rect 1737 3515 1763 3541
rect 1763 3515 1764 3541
rect 1736 3514 1764 3515
rect 1788 3541 1816 3542
rect 1788 3515 1789 3541
rect 1789 3515 1815 3541
rect 1815 3515 1816 3541
rect 1788 3514 1816 3515
rect 1134 3374 1162 3402
rect 854 3038 882 3066
rect 1022 3009 1050 3010
rect 1022 2983 1023 3009
rect 1023 2983 1049 3009
rect 1049 2983 1050 3009
rect 1022 2982 1050 2983
rect 854 2702 882 2730
rect 966 2926 994 2954
rect 910 2478 938 2506
rect 2762 3933 2790 3934
rect 2762 3907 2763 3933
rect 2763 3907 2789 3933
rect 2789 3907 2790 3933
rect 2762 3906 2790 3907
rect 2814 3933 2842 3934
rect 2814 3907 2815 3933
rect 2815 3907 2841 3933
rect 2841 3907 2842 3933
rect 2814 3906 2842 3907
rect 2866 3933 2894 3934
rect 2866 3907 2867 3933
rect 2867 3907 2893 3933
rect 2893 3907 2894 3933
rect 2866 3906 2894 3907
rect 2814 3822 2842 3850
rect 2198 3598 2226 3626
rect 1862 3374 1890 3402
rect 2310 3318 2338 3346
rect 1190 3206 1218 3234
rect 1246 3038 1274 3066
rect 1246 2702 1274 2730
rect 1302 2814 1330 2842
rect 854 2169 882 2170
rect 854 2143 855 2169
rect 855 2143 881 2169
rect 881 2143 882 2169
rect 854 2142 882 2143
rect 14 1918 42 1946
rect 406 1862 434 1890
rect 854 2030 882 2058
rect 1190 2254 1218 2282
rect 1190 1918 1218 1946
rect 1134 1806 1162 1834
rect 1470 2478 1498 2506
rect 1358 2225 1386 2226
rect 1358 2199 1359 2225
rect 1359 2199 1385 2225
rect 1385 2199 1386 2225
rect 1358 2198 1386 2199
rect 1694 3233 1722 3234
rect 1694 3207 1695 3233
rect 1695 3207 1721 3233
rect 1721 3207 1722 3233
rect 1694 3206 1722 3207
rect 1414 1022 1442 1050
rect 1684 2757 1712 2758
rect 1684 2731 1685 2757
rect 1685 2731 1711 2757
rect 1711 2731 1712 2757
rect 1684 2730 1712 2731
rect 1736 2757 1764 2758
rect 1736 2731 1737 2757
rect 1737 2731 1763 2757
rect 1763 2731 1764 2757
rect 1736 2730 1764 2731
rect 1788 2757 1816 2758
rect 1788 2731 1789 2757
rect 1789 2731 1815 2757
rect 1815 2731 1816 2757
rect 1788 2730 1816 2731
rect 1582 2254 1610 2282
rect 1694 2281 1722 2282
rect 1694 2255 1695 2281
rect 1695 2255 1721 2281
rect 1721 2255 1722 2281
rect 1694 2254 1722 2255
rect 1806 2142 1834 2170
rect 1684 1973 1712 1974
rect 1684 1947 1685 1973
rect 1685 1947 1711 1973
rect 1711 1947 1712 1973
rect 1684 1946 1712 1947
rect 1736 1973 1764 1974
rect 1736 1947 1737 1973
rect 1737 1947 1763 1973
rect 1763 1947 1764 1973
rect 1736 1946 1764 1947
rect 1788 1973 1816 1974
rect 1788 1947 1789 1973
rect 1789 1947 1815 1973
rect 1815 1947 1816 1973
rect 1788 1946 1816 1947
rect 1526 1862 1554 1890
rect 1638 1862 1666 1890
rect 1750 1358 1778 1386
rect 1974 2422 2002 2450
rect 2762 3149 2790 3150
rect 2762 3123 2763 3149
rect 2763 3123 2789 3149
rect 2789 3123 2790 3149
rect 2762 3122 2790 3123
rect 2814 3149 2842 3150
rect 2814 3123 2815 3149
rect 2815 3123 2841 3149
rect 2841 3123 2842 3149
rect 2814 3122 2842 3123
rect 2866 3149 2894 3150
rect 2866 3123 2867 3149
rect 2867 3123 2893 3149
rect 2893 3123 2894 3149
rect 2866 3122 2894 3123
rect 3990 4494 4018 4522
rect 4046 4550 4074 4578
rect 3822 4465 3850 4466
rect 3822 4439 3823 4465
rect 3823 4439 3849 4465
rect 3849 4439 3850 4465
rect 3822 4438 3850 4439
rect 3840 4325 3868 4326
rect 3840 4299 3841 4325
rect 3841 4299 3867 4325
rect 3867 4299 3868 4325
rect 3840 4298 3868 4299
rect 3892 4325 3920 4326
rect 3892 4299 3893 4325
rect 3893 4299 3919 4325
rect 3919 4299 3920 4325
rect 3892 4298 3920 4299
rect 3944 4325 3972 4326
rect 3944 4299 3945 4325
rect 3945 4299 3971 4325
rect 3971 4299 3972 4325
rect 3944 4298 3972 4299
rect 3766 4214 3794 4242
rect 3094 3990 3122 4018
rect 4158 4494 4186 4522
rect 4270 4550 4298 4578
rect 5996 6677 6024 6678
rect 5996 6651 5997 6677
rect 5997 6651 6023 6677
rect 6023 6651 6024 6677
rect 5996 6650 6024 6651
rect 6048 6677 6076 6678
rect 6048 6651 6049 6677
rect 6049 6651 6075 6677
rect 6075 6651 6076 6677
rect 6048 6650 6076 6651
rect 6100 6677 6128 6678
rect 6100 6651 6101 6677
rect 6101 6651 6127 6677
rect 6127 6651 6128 6677
rect 6100 6650 6128 6651
rect 6454 6537 6482 6538
rect 6454 6511 6455 6537
rect 6455 6511 6481 6537
rect 6481 6511 6482 6537
rect 6454 6510 6482 6511
rect 6846 6510 6874 6538
rect 5894 6174 5922 6202
rect 5558 6006 5586 6034
rect 5614 5726 5642 5754
rect 5996 5893 6024 5894
rect 5996 5867 5997 5893
rect 5997 5867 6023 5893
rect 6023 5867 6024 5893
rect 5996 5866 6024 5867
rect 6048 5893 6076 5894
rect 6048 5867 6049 5893
rect 6049 5867 6075 5893
rect 6075 5867 6076 5893
rect 6048 5866 6076 5867
rect 6100 5893 6128 5894
rect 6100 5867 6101 5893
rect 6101 5867 6127 5893
rect 6127 5867 6128 5893
rect 6100 5866 6128 5867
rect 6118 5166 6146 5194
rect 4918 4717 4946 4718
rect 4918 4691 4919 4717
rect 4919 4691 4945 4717
rect 4945 4691 4946 4717
rect 4918 4690 4946 4691
rect 4970 4717 4998 4718
rect 4970 4691 4971 4717
rect 4971 4691 4997 4717
rect 4997 4691 4998 4717
rect 4970 4690 4998 4691
rect 5022 4717 5050 4718
rect 5022 4691 5023 4717
rect 5023 4691 5049 4717
rect 5049 4691 5050 4717
rect 5022 4690 5050 4691
rect 4214 4438 4242 4466
rect 4438 4465 4466 4466
rect 4438 4439 4439 4465
rect 4439 4439 4465 4465
rect 4465 4439 4466 4465
rect 4438 4438 4466 4439
rect 4494 4409 4522 4410
rect 4494 4383 4495 4409
rect 4495 4383 4521 4409
rect 4521 4383 4522 4409
rect 4494 4382 4522 4383
rect 4158 4046 4186 4074
rect 4102 3849 4130 3850
rect 4102 3823 4103 3849
rect 4103 3823 4129 3849
rect 4129 3823 4130 3849
rect 4102 3822 4130 3823
rect 3318 3262 3346 3290
rect 3840 3541 3868 3542
rect 3840 3515 3841 3541
rect 3841 3515 3867 3541
rect 3867 3515 3868 3541
rect 3840 3514 3868 3515
rect 3892 3541 3920 3542
rect 3892 3515 3893 3541
rect 3893 3515 3919 3541
rect 3919 3515 3920 3541
rect 3892 3514 3920 3515
rect 3944 3541 3972 3542
rect 3944 3515 3945 3541
rect 3945 3515 3971 3541
rect 3971 3515 3972 3541
rect 3944 3514 3972 3515
rect 4102 3318 4130 3346
rect 4046 3262 4074 3290
rect 2982 2982 3010 3010
rect 2590 2814 2618 2842
rect 2590 2617 2618 2618
rect 2590 2591 2591 2617
rect 2591 2591 2617 2617
rect 2617 2591 2618 2617
rect 2590 2590 2618 2591
rect 3318 2561 3346 2562
rect 3318 2535 3319 2561
rect 3319 2535 3345 2561
rect 3345 2535 3346 2561
rect 3318 2534 3346 2535
rect 2762 2365 2790 2366
rect 2762 2339 2763 2365
rect 2763 2339 2789 2365
rect 2789 2339 2790 2365
rect 2762 2338 2790 2339
rect 2814 2365 2842 2366
rect 2814 2339 2815 2365
rect 2815 2339 2841 2365
rect 2841 2339 2842 2365
rect 2814 2338 2842 2339
rect 2866 2365 2894 2366
rect 2866 2339 2867 2365
rect 2867 2339 2893 2365
rect 2893 2339 2894 2365
rect 2866 2338 2894 2339
rect 2366 1777 2394 1778
rect 2366 1751 2367 1777
rect 2367 1751 2393 1777
rect 2393 1751 2394 1777
rect 2366 1750 2394 1751
rect 2762 1581 2790 1582
rect 2762 1555 2763 1581
rect 2763 1555 2789 1581
rect 2789 1555 2790 1581
rect 2762 1554 2790 1555
rect 2814 1581 2842 1582
rect 2814 1555 2815 1581
rect 2815 1555 2841 1581
rect 2841 1555 2842 1581
rect 2814 1554 2842 1555
rect 2866 1581 2894 1582
rect 2866 1555 2867 1581
rect 2867 1555 2893 1581
rect 2893 1555 2894 1581
rect 2866 1554 2894 1555
rect 3598 2953 3626 2954
rect 3598 2927 3599 2953
rect 3599 2927 3625 2953
rect 3625 2927 3626 2953
rect 3598 2926 3626 2927
rect 3840 2757 3868 2758
rect 3840 2731 3841 2757
rect 3841 2731 3867 2757
rect 3867 2731 3868 2757
rect 3840 2730 3868 2731
rect 3892 2757 3920 2758
rect 3892 2731 3893 2757
rect 3893 2731 3919 2757
rect 3919 2731 3920 2757
rect 3892 2730 3920 2731
rect 3944 2757 3972 2758
rect 3944 2731 3945 2757
rect 3945 2731 3971 2757
rect 3971 2731 3972 2757
rect 3944 2730 3972 2731
rect 4326 3822 4354 3850
rect 4774 4046 4802 4074
rect 4918 3933 4946 3934
rect 4918 3907 4919 3933
rect 4919 3907 4945 3933
rect 4945 3907 4946 3933
rect 4918 3906 4946 3907
rect 4970 3933 4998 3934
rect 4970 3907 4971 3933
rect 4971 3907 4997 3933
rect 4997 3907 4998 3933
rect 4970 3906 4998 3907
rect 5022 3933 5050 3934
rect 5022 3907 5023 3933
rect 5023 3907 5049 3933
rect 5049 3907 5050 3933
rect 5022 3906 5050 3907
rect 4326 3374 4354 3402
rect 4382 3345 4410 3346
rect 4382 3319 4383 3345
rect 4383 3319 4409 3345
rect 4409 3319 4410 3345
rect 4382 3318 4410 3319
rect 3598 2590 3626 2618
rect 3374 2198 3402 2226
rect 3542 2478 3570 2506
rect 3486 2169 3514 2170
rect 3486 2143 3487 2169
rect 3487 2143 3513 2169
rect 3513 2143 3514 2169
rect 3486 2142 3514 2143
rect 3374 1862 3402 1890
rect 3206 1694 3234 1722
rect 3374 1750 3402 1778
rect 3598 2086 3626 2114
rect 3766 2561 3794 2562
rect 3766 2535 3767 2561
rect 3767 2535 3793 2561
rect 3793 2535 3794 2561
rect 3766 2534 3794 2535
rect 4046 2534 4074 2562
rect 3840 1973 3868 1974
rect 3840 1947 3841 1973
rect 3841 1947 3867 1973
rect 3867 1947 3868 1973
rect 3840 1946 3868 1947
rect 3892 1973 3920 1974
rect 3892 1947 3893 1973
rect 3893 1947 3919 1973
rect 3919 1947 3920 1973
rect 3892 1946 3920 1947
rect 3944 1973 3972 1974
rect 3944 1947 3945 1973
rect 3945 1947 3971 1973
rect 3971 1947 3972 1973
rect 3944 1946 3972 1947
rect 4718 3318 4746 3346
rect 4918 3149 4946 3150
rect 4918 3123 4919 3149
rect 4919 3123 4945 3149
rect 4945 3123 4946 3149
rect 4918 3122 4946 3123
rect 4970 3149 4998 3150
rect 4970 3123 4971 3149
rect 4971 3123 4997 3149
rect 4997 3123 4998 3149
rect 4970 3122 4998 3123
rect 5022 3149 5050 3150
rect 5022 3123 5023 3149
rect 5023 3123 5049 3149
rect 5049 3123 5050 3149
rect 5022 3122 5050 3123
rect 4774 2590 4802 2618
rect 4662 2422 4690 2450
rect 4438 1974 4466 2002
rect 4494 1862 4522 1890
rect 5166 2561 5194 2562
rect 5166 2535 5167 2561
rect 5167 2535 5193 2561
rect 5193 2535 5194 2561
rect 5166 2534 5194 2535
rect 5278 3318 5306 3346
rect 5278 2478 5306 2506
rect 4918 2365 4946 2366
rect 4918 2339 4919 2365
rect 4919 2339 4945 2365
rect 4945 2339 4946 2365
rect 4918 2338 4946 2339
rect 4970 2365 4998 2366
rect 4970 2339 4971 2365
rect 4971 2339 4997 2365
rect 4997 2339 4998 2365
rect 4970 2338 4998 2339
rect 5022 2365 5050 2366
rect 5022 2339 5023 2365
rect 5023 2339 5049 2365
rect 5049 2339 5050 2365
rect 5022 2338 5050 2339
rect 4382 1750 4410 1778
rect 5054 2113 5082 2114
rect 5054 2087 5055 2113
rect 5055 2087 5081 2113
rect 5081 2087 5082 2113
rect 5054 2086 5082 2087
rect 4918 1581 4946 1582
rect 4918 1555 4919 1581
rect 4919 1555 4945 1581
rect 4945 1555 4946 1581
rect 4918 1554 4946 1555
rect 4970 1581 4998 1582
rect 4970 1555 4971 1581
rect 4971 1555 4997 1581
rect 4997 1555 4998 1581
rect 4970 1554 4998 1555
rect 5022 1581 5050 1582
rect 5022 1555 5023 1581
rect 5023 1555 5049 1581
rect 5049 1555 5050 1581
rect 5022 1554 5050 1555
rect 5502 4214 5530 4242
rect 5558 3822 5586 3850
rect 5996 5109 6024 5110
rect 5996 5083 5997 5109
rect 5997 5083 6023 5109
rect 6023 5083 6024 5109
rect 5996 5082 6024 5083
rect 6048 5109 6076 5110
rect 6048 5083 6049 5109
rect 6049 5083 6075 5109
rect 6075 5083 6076 5109
rect 6048 5082 6076 5083
rect 6100 5109 6128 5110
rect 6100 5083 6101 5109
rect 6101 5083 6127 5109
rect 6127 5083 6128 5109
rect 6100 5082 6128 5083
rect 6790 5753 6818 5754
rect 6790 5727 6791 5753
rect 6791 5727 6817 5753
rect 6817 5727 6818 5753
rect 6790 5726 6818 5727
rect 6342 5585 6370 5586
rect 6342 5559 6343 5585
rect 6343 5559 6369 5585
rect 6369 5559 6370 5585
rect 6342 5558 6370 5559
rect 6454 5670 6482 5698
rect 6734 5697 6762 5698
rect 6734 5671 6735 5697
rect 6735 5671 6761 5697
rect 6761 5671 6762 5697
rect 6734 5670 6762 5671
rect 8152 6677 8180 6678
rect 8152 6651 8153 6677
rect 8153 6651 8179 6677
rect 8179 6651 8180 6677
rect 8152 6650 8180 6651
rect 8204 6677 8232 6678
rect 8204 6651 8205 6677
rect 8205 6651 8231 6677
rect 8231 6651 8232 6677
rect 8204 6650 8232 6651
rect 8256 6677 8284 6678
rect 8256 6651 8257 6677
rect 8257 6651 8283 6677
rect 8283 6651 8284 6677
rect 8256 6650 8284 6651
rect 6958 6454 6986 6482
rect 7686 6481 7714 6482
rect 7686 6455 7687 6481
rect 7687 6455 7713 6481
rect 7713 6455 7714 6481
rect 7686 6454 7714 6455
rect 7074 6285 7102 6286
rect 7074 6259 7075 6285
rect 7075 6259 7101 6285
rect 7101 6259 7102 6285
rect 7074 6258 7102 6259
rect 7126 6285 7154 6286
rect 7126 6259 7127 6285
rect 7127 6259 7153 6285
rect 7153 6259 7154 6285
rect 7126 6258 7154 6259
rect 7178 6285 7206 6286
rect 7178 6259 7179 6285
rect 7179 6259 7205 6285
rect 7205 6259 7206 6285
rect 7178 6258 7206 6259
rect 7238 6174 7266 6202
rect 6902 6062 6930 6090
rect 6286 4606 6314 4634
rect 6230 4521 6258 4522
rect 6230 4495 6231 4521
rect 6231 4495 6257 4521
rect 6257 4495 6258 4521
rect 6230 4494 6258 4495
rect 6846 4913 6874 4914
rect 6846 4887 6847 4913
rect 6847 4887 6873 4913
rect 6873 4887 6874 4913
rect 6846 4886 6874 4887
rect 6454 4494 6482 4522
rect 5838 4382 5866 4410
rect 5996 4325 6024 4326
rect 5996 4299 5997 4325
rect 5997 4299 6023 4325
rect 6023 4299 6024 4325
rect 5996 4298 6024 4299
rect 6048 4325 6076 4326
rect 6048 4299 6049 4325
rect 6049 4299 6075 4325
rect 6075 4299 6076 4325
rect 6048 4298 6076 4299
rect 6100 4325 6128 4326
rect 6100 4299 6101 4325
rect 6101 4299 6127 4325
rect 6127 4299 6128 4325
rect 6100 4298 6128 4299
rect 5950 3849 5978 3850
rect 5950 3823 5951 3849
rect 5951 3823 5977 3849
rect 5977 3823 5978 3849
rect 5950 3822 5978 3823
rect 5996 3541 6024 3542
rect 5996 3515 5997 3541
rect 5997 3515 6023 3541
rect 6023 3515 6024 3541
rect 5996 3514 6024 3515
rect 6048 3541 6076 3542
rect 6048 3515 6049 3541
rect 6049 3515 6075 3541
rect 6075 3515 6076 3541
rect 6048 3514 6076 3515
rect 6100 3541 6128 3542
rect 6100 3515 6101 3541
rect 6101 3515 6127 3541
rect 6127 3515 6128 3541
rect 6100 3514 6128 3515
rect 5670 3374 5698 3402
rect 5446 2086 5474 2114
rect 5502 1721 5530 1722
rect 5502 1695 5503 1721
rect 5503 1695 5529 1721
rect 5529 1695 5530 1721
rect 5502 1694 5530 1695
rect 5996 2757 6024 2758
rect 5996 2731 5997 2757
rect 5997 2731 6023 2757
rect 6023 2731 6024 2757
rect 5996 2730 6024 2731
rect 6048 2757 6076 2758
rect 6048 2731 6049 2757
rect 6049 2731 6075 2757
rect 6075 2731 6076 2757
rect 6048 2730 6076 2731
rect 6100 2757 6128 2758
rect 6100 2731 6101 2757
rect 6101 2731 6127 2757
rect 6127 2731 6128 2757
rect 6100 2730 6128 2731
rect 7014 6033 7042 6034
rect 7014 6007 7015 6033
rect 7015 6007 7041 6033
rect 7041 6007 7042 6033
rect 7014 6006 7042 6007
rect 6958 5222 6986 5250
rect 6958 4886 6986 4914
rect 7182 5641 7210 5642
rect 7182 5615 7183 5641
rect 7183 5615 7209 5641
rect 7209 5615 7210 5641
rect 7182 5614 7210 5615
rect 8470 6510 8498 6538
rect 9030 6425 9058 6426
rect 9030 6399 9031 6425
rect 9031 6399 9057 6425
rect 9057 6399 9058 6425
rect 9030 6398 9058 6399
rect 9230 6285 9258 6286
rect 9230 6259 9231 6285
rect 9231 6259 9257 6285
rect 9257 6259 9258 6285
rect 9230 6258 9258 6259
rect 9282 6285 9310 6286
rect 9282 6259 9283 6285
rect 9283 6259 9309 6285
rect 9309 6259 9310 6285
rect 9282 6258 9310 6259
rect 9334 6285 9362 6286
rect 9334 6259 9335 6285
rect 9335 6259 9361 6285
rect 9361 6259 9362 6285
rect 9334 6258 9362 6259
rect 8190 6062 8218 6090
rect 8152 5893 8180 5894
rect 8152 5867 8153 5893
rect 8153 5867 8179 5893
rect 8179 5867 8180 5893
rect 8152 5866 8180 5867
rect 8204 5893 8232 5894
rect 8204 5867 8205 5893
rect 8205 5867 8231 5893
rect 8231 5867 8232 5893
rect 8204 5866 8232 5867
rect 8256 5893 8284 5894
rect 8256 5867 8257 5893
rect 8257 5867 8283 5893
rect 8283 5867 8284 5893
rect 8256 5866 8284 5867
rect 7294 5558 7322 5586
rect 7630 5585 7658 5586
rect 7630 5559 7631 5585
rect 7631 5559 7657 5585
rect 7657 5559 7658 5585
rect 7630 5558 7658 5559
rect 7074 5501 7102 5502
rect 7074 5475 7075 5501
rect 7075 5475 7101 5501
rect 7101 5475 7102 5501
rect 7074 5474 7102 5475
rect 7126 5501 7154 5502
rect 7126 5475 7127 5501
rect 7127 5475 7153 5501
rect 7153 5475 7154 5501
rect 7126 5474 7154 5475
rect 7178 5501 7206 5502
rect 7178 5475 7179 5501
rect 7179 5475 7205 5501
rect 7205 5475 7206 5501
rect 7178 5474 7206 5475
rect 7910 5361 7938 5362
rect 7910 5335 7911 5361
rect 7911 5335 7937 5361
rect 7937 5335 7938 5361
rect 7910 5334 7938 5335
rect 7742 5249 7770 5250
rect 7742 5223 7743 5249
rect 7743 5223 7769 5249
rect 7769 5223 7770 5249
rect 7742 5222 7770 5223
rect 8152 5109 8180 5110
rect 8152 5083 8153 5109
rect 8153 5083 8179 5109
rect 8179 5083 8180 5109
rect 8152 5082 8180 5083
rect 8204 5109 8232 5110
rect 8204 5083 8205 5109
rect 8205 5083 8231 5109
rect 8231 5083 8232 5109
rect 8204 5082 8232 5083
rect 8256 5109 8284 5110
rect 8256 5083 8257 5109
rect 8257 5083 8283 5109
rect 8283 5083 8284 5109
rect 8256 5082 8284 5083
rect 7074 4717 7102 4718
rect 7074 4691 7075 4717
rect 7075 4691 7101 4717
rect 7101 4691 7102 4717
rect 7074 4690 7102 4691
rect 7126 4717 7154 4718
rect 7126 4691 7127 4717
rect 7127 4691 7153 4717
rect 7153 4691 7154 4717
rect 7126 4690 7154 4691
rect 7178 4717 7206 4718
rect 7178 4691 7179 4717
rect 7179 4691 7205 4717
rect 7205 4691 7206 4717
rect 7178 4690 7206 4691
rect 7182 4606 7210 4634
rect 7126 4550 7154 4578
rect 6510 4046 6538 4074
rect 6846 4438 6874 4466
rect 6958 4382 6986 4410
rect 6958 4270 6986 4298
rect 7350 4521 7378 4522
rect 7350 4495 7351 4521
rect 7351 4495 7377 4521
rect 7377 4495 7378 4521
rect 7350 4494 7378 4495
rect 9086 5726 9114 5754
rect 9230 5501 9258 5502
rect 9230 5475 9231 5501
rect 9231 5475 9257 5501
rect 9257 5475 9258 5501
rect 9230 5474 9258 5475
rect 9282 5501 9310 5502
rect 9282 5475 9283 5501
rect 9283 5475 9309 5501
rect 9309 5475 9310 5501
rect 9282 5474 9310 5475
rect 9334 5501 9362 5502
rect 9334 5475 9335 5501
rect 9335 5475 9361 5501
rect 9361 5475 9362 5501
rect 9334 5474 9362 5475
rect 9030 5390 9058 5418
rect 8918 5361 8946 5362
rect 8918 5335 8919 5361
rect 8919 5335 8945 5361
rect 8945 5335 8946 5361
rect 8918 5334 8946 5335
rect 8918 5110 8946 5138
rect 9086 5054 9114 5082
rect 8806 4801 8834 4802
rect 8806 4775 8807 4801
rect 8807 4775 8833 4801
rect 8833 4775 8834 4801
rect 8806 4774 8834 4775
rect 9086 4774 9114 4802
rect 9230 4717 9258 4718
rect 9230 4691 9231 4717
rect 9231 4691 9257 4717
rect 9257 4691 9258 4717
rect 9230 4690 9258 4691
rect 9282 4717 9310 4718
rect 9282 4691 9283 4717
rect 9283 4691 9309 4717
rect 9309 4691 9310 4717
rect 9282 4690 9310 4691
rect 9334 4717 9362 4718
rect 9334 4691 9335 4717
rect 9335 4691 9361 4717
rect 9361 4691 9362 4717
rect 9334 4690 9362 4691
rect 8750 4550 8778 4578
rect 8918 4494 8946 4522
rect 8806 4382 8834 4410
rect 9086 4382 9114 4410
rect 7406 4270 7434 4298
rect 8152 4325 8180 4326
rect 8152 4299 8153 4325
rect 8153 4299 8179 4325
rect 8179 4299 8180 4325
rect 8152 4298 8180 4299
rect 8204 4325 8232 4326
rect 8204 4299 8205 4325
rect 8205 4299 8231 4325
rect 8231 4299 8232 4325
rect 8204 4298 8232 4299
rect 8256 4325 8284 4326
rect 8256 4299 8257 4325
rect 8257 4299 8283 4325
rect 8283 4299 8284 4325
rect 8256 4298 8284 4299
rect 7126 4073 7154 4074
rect 7126 4047 7127 4073
rect 7127 4047 7153 4073
rect 7153 4047 7154 4073
rect 7126 4046 7154 4047
rect 6790 3990 6818 4018
rect 8582 4073 8610 4074
rect 8582 4047 8583 4073
rect 8583 4047 8609 4073
rect 8609 4047 8610 4073
rect 8582 4046 8610 4047
rect 7182 3990 7210 4018
rect 7074 3933 7102 3934
rect 7074 3907 7075 3933
rect 7075 3907 7101 3933
rect 7101 3907 7102 3933
rect 7074 3906 7102 3907
rect 7126 3933 7154 3934
rect 7126 3907 7127 3933
rect 7127 3907 7153 3933
rect 7153 3907 7154 3933
rect 7126 3906 7154 3907
rect 7178 3933 7206 3934
rect 7178 3907 7179 3933
rect 7179 3907 7205 3933
rect 7205 3907 7206 3933
rect 7178 3906 7206 3907
rect 6454 3793 6482 3794
rect 6454 3767 6455 3793
rect 6455 3767 6481 3793
rect 6481 3767 6482 3793
rect 6454 3766 6482 3767
rect 6230 2561 6258 2562
rect 6230 2535 6231 2561
rect 6231 2535 6257 2561
rect 6257 2535 6258 2561
rect 6230 2534 6258 2535
rect 6398 2254 6426 2282
rect 6118 2225 6146 2226
rect 6118 2199 6119 2225
rect 6119 2199 6145 2225
rect 6145 2199 6146 2225
rect 6118 2198 6146 2199
rect 5726 1750 5754 1778
rect 5838 1974 5866 2002
rect 5996 1973 6024 1974
rect 5996 1947 5997 1973
rect 5997 1947 6023 1973
rect 6023 1947 6024 1973
rect 5996 1946 6024 1947
rect 6048 1973 6076 1974
rect 6048 1947 6049 1973
rect 6049 1947 6075 1973
rect 6075 1947 6076 1973
rect 6048 1946 6076 1947
rect 6100 1973 6128 1974
rect 6100 1947 6101 1973
rect 6101 1947 6127 1973
rect 6127 1947 6128 1973
rect 6100 1946 6128 1947
rect 5950 1777 5978 1778
rect 5950 1751 5951 1777
rect 5951 1751 5977 1777
rect 5977 1751 5978 1777
rect 5950 1750 5978 1751
rect 6398 1750 6426 1778
rect 6062 1694 6090 1722
rect 5726 1638 5754 1666
rect 6174 1665 6202 1666
rect 6174 1639 6175 1665
rect 6175 1639 6201 1665
rect 6201 1639 6202 1665
rect 6174 1638 6202 1639
rect 7074 3149 7102 3150
rect 7074 3123 7075 3149
rect 7075 3123 7101 3149
rect 7101 3123 7102 3149
rect 7074 3122 7102 3123
rect 7126 3149 7154 3150
rect 7126 3123 7127 3149
rect 7127 3123 7153 3149
rect 7153 3123 7154 3149
rect 7126 3122 7154 3123
rect 7178 3149 7206 3150
rect 7178 3123 7179 3149
rect 7179 3123 7205 3149
rect 7205 3123 7206 3149
rect 7178 3122 7206 3123
rect 7074 2365 7102 2366
rect 7074 2339 7075 2365
rect 7075 2339 7101 2365
rect 7101 2339 7102 2365
rect 7074 2338 7102 2339
rect 7126 2365 7154 2366
rect 7126 2339 7127 2365
rect 7127 2339 7153 2365
rect 7153 2339 7154 2365
rect 7126 2338 7154 2339
rect 7178 2365 7206 2366
rect 7178 2339 7179 2365
rect 7179 2339 7205 2365
rect 7205 2339 7206 2365
rect 7178 2338 7206 2339
rect 6678 2086 6706 2114
rect 7238 2254 7266 2282
rect 8470 3766 8498 3794
rect 7462 2254 7490 2282
rect 7014 1777 7042 1778
rect 7014 1751 7015 1777
rect 7015 1751 7041 1777
rect 7041 1751 7042 1777
rect 7014 1750 7042 1751
rect 6678 1694 6706 1722
rect 7074 1581 7102 1582
rect 7074 1555 7075 1581
rect 7075 1555 7101 1581
rect 7101 1555 7102 1581
rect 7074 1554 7102 1555
rect 7126 1581 7154 1582
rect 7126 1555 7127 1581
rect 7127 1555 7153 1581
rect 7153 1555 7154 1581
rect 7126 1554 7154 1555
rect 7178 1581 7206 1582
rect 7178 1555 7179 1581
rect 7179 1555 7205 1581
rect 7205 1555 7206 1581
rect 7178 1554 7206 1555
rect 7406 1694 7434 1722
rect 8152 3541 8180 3542
rect 8152 3515 8153 3541
rect 8153 3515 8179 3541
rect 8179 3515 8180 3541
rect 8152 3514 8180 3515
rect 8204 3541 8232 3542
rect 8204 3515 8205 3541
rect 8205 3515 8231 3541
rect 8231 3515 8232 3541
rect 8204 3514 8232 3515
rect 8256 3541 8284 3542
rect 8256 3515 8257 3541
rect 8257 3515 8283 3541
rect 8283 3515 8284 3541
rect 8256 3514 8284 3515
rect 8152 2757 8180 2758
rect 8152 2731 8153 2757
rect 8153 2731 8179 2757
rect 8179 2731 8180 2757
rect 8152 2730 8180 2731
rect 8204 2757 8232 2758
rect 8204 2731 8205 2757
rect 8205 2731 8231 2757
rect 8231 2731 8232 2757
rect 8204 2730 8232 2731
rect 8256 2757 8284 2758
rect 8256 2731 8257 2757
rect 8257 2731 8283 2757
rect 8283 2731 8284 2757
rect 8256 2730 8284 2731
rect 7742 2478 7770 2506
rect 7854 2281 7882 2282
rect 7854 2255 7855 2281
rect 7855 2255 7881 2281
rect 7881 2255 7882 2281
rect 7854 2254 7882 2255
rect 7630 1750 7658 1778
rect 7686 1694 7714 1722
rect 8358 2422 8386 2450
rect 8246 2225 8274 2226
rect 8246 2199 8247 2225
rect 8247 2199 8273 2225
rect 8273 2199 8274 2225
rect 8246 2198 8274 2199
rect 8414 2169 8442 2170
rect 8414 2143 8415 2169
rect 8415 2143 8441 2169
rect 8441 2143 8442 2169
rect 8414 2142 8442 2143
rect 8152 1973 8180 1974
rect 8152 1947 8153 1973
rect 8153 1947 8179 1973
rect 8179 1947 8180 1973
rect 8152 1946 8180 1947
rect 8204 1973 8232 1974
rect 8204 1947 8205 1973
rect 8205 1947 8231 1973
rect 8231 1947 8232 1973
rect 8204 1946 8232 1947
rect 8256 1973 8284 1974
rect 8256 1947 8257 1973
rect 8257 1947 8283 1973
rect 8283 1947 8284 1973
rect 8256 1946 8284 1947
rect 8022 1777 8050 1778
rect 8022 1751 8023 1777
rect 8023 1751 8049 1777
rect 8049 1751 8050 1777
rect 8022 1750 8050 1751
rect 8134 1694 8162 1722
rect 9086 4073 9114 4074
rect 9086 4047 9087 4073
rect 9087 4047 9113 4073
rect 9113 4047 9114 4073
rect 9086 4046 9114 4047
rect 8918 4017 8946 4018
rect 8918 3991 8919 4017
rect 8919 3991 8945 4017
rect 8945 3991 8946 4017
rect 8918 3990 8946 3991
rect 9230 3933 9258 3934
rect 9230 3907 9231 3933
rect 9231 3907 9257 3933
rect 9257 3907 9258 3933
rect 9230 3906 9258 3907
rect 9282 3933 9310 3934
rect 9282 3907 9283 3933
rect 9283 3907 9309 3933
rect 9309 3907 9310 3933
rect 9282 3906 9310 3907
rect 9334 3933 9362 3934
rect 9334 3907 9335 3933
rect 9335 3907 9361 3933
rect 9361 3907 9362 3933
rect 9334 3906 9362 3907
rect 8862 3737 8890 3738
rect 8862 3711 8863 3737
rect 8863 3711 8889 3737
rect 8889 3711 8890 3737
rect 8862 3710 8890 3711
rect 9230 3149 9258 3150
rect 9230 3123 9231 3149
rect 9231 3123 9257 3149
rect 9257 3123 9258 3149
rect 9230 3122 9258 3123
rect 9282 3149 9310 3150
rect 9282 3123 9283 3149
rect 9283 3123 9309 3149
rect 9309 3123 9310 3149
rect 9282 3122 9310 3123
rect 9334 3149 9362 3150
rect 9334 3123 9335 3149
rect 9335 3123 9361 3149
rect 9361 3123 9362 3149
rect 9334 3122 9362 3123
rect 9086 3038 9114 3066
rect 8582 2142 8610 2170
rect 8750 2030 8778 2058
rect 8750 1862 8778 1890
rect 8582 1694 8610 1722
rect 8862 2478 8890 2506
rect 8918 2086 8946 2114
rect 8974 2422 9002 2450
rect 9030 2142 9058 2170
rect 9230 2365 9258 2366
rect 9230 2339 9231 2365
rect 9231 2339 9257 2365
rect 9257 2339 9258 2365
rect 9230 2338 9258 2339
rect 9282 2365 9310 2366
rect 9282 2339 9283 2365
rect 9283 2339 9309 2365
rect 9309 2339 9310 2365
rect 9282 2338 9310 2339
rect 9334 2365 9362 2366
rect 9334 2339 9335 2365
rect 9335 2339 9361 2365
rect 9361 2339 9362 2365
rect 9334 2338 9362 2339
rect 9230 1581 9258 1582
rect 9230 1555 9231 1581
rect 9231 1555 9257 1581
rect 9257 1555 9258 1581
rect 9230 1554 9258 1555
rect 9282 1581 9310 1582
rect 9282 1555 9283 1581
rect 9283 1555 9309 1581
rect 9309 1555 9310 1581
rect 9282 1554 9310 1555
rect 9334 1581 9362 1582
rect 9334 1555 9335 1581
rect 9335 1555 9361 1581
rect 9361 1555 9362 1581
rect 9334 1554 9362 1555
<< metal3 >>
rect 0 8442 400 8456
rect 0 8414 1330 8442
rect 0 8400 400 8414
rect 1302 8386 1330 8414
rect 1297 8358 1302 8386
rect 1330 8358 1335 8386
rect 1679 8218 1684 8246
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1816 8218 1821 8246
rect 3835 8218 3840 8246
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3972 8218 3977 8246
rect 5991 8218 5996 8246
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 6128 8218 6133 8246
rect 8147 8218 8152 8246
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8284 8218 8289 8246
rect 4041 8134 4046 8162
rect 4074 8134 4662 8162
rect 4690 8134 4695 8162
rect 0 8106 400 8120
rect 0 8078 1078 8106
rect 1106 8078 1111 8106
rect 0 8064 400 8078
rect 849 7910 854 7938
rect 882 7910 887 7938
rect 854 7826 882 7910
rect 2757 7826 2762 7854
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2894 7826 2899 7854
rect 4913 7826 4918 7854
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 5050 7826 5055 7854
rect 7069 7826 7074 7854
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7206 7826 7211 7854
rect 9225 7826 9230 7854
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9362 7826 9367 7854
rect 462 7798 882 7826
rect 0 7770 400 7784
rect 462 7770 490 7798
rect 9600 7770 10000 7784
rect 0 7742 490 7770
rect 9137 7742 9142 7770
rect 9170 7742 10000 7770
rect 0 7728 400 7742
rect 9600 7728 10000 7742
rect 849 7574 854 7602
rect 882 7574 887 7602
rect 0 7434 400 7448
rect 854 7434 882 7574
rect 1679 7434 1684 7462
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1816 7434 1821 7462
rect 3835 7434 3840 7462
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3972 7434 3977 7462
rect 5991 7434 5996 7462
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 6128 7434 6133 7462
rect 8147 7434 8152 7462
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8284 7434 8289 7462
rect 9600 7434 10000 7448
rect 0 7406 882 7434
rect 9081 7406 9086 7434
rect 9114 7406 10000 7434
rect 0 7392 400 7406
rect 9600 7392 10000 7406
rect 849 7126 854 7154
rect 882 7126 887 7154
rect 9081 7126 9086 7154
rect 9114 7126 9450 7154
rect 0 7098 400 7112
rect 854 7098 882 7126
rect 0 7070 882 7098
rect 9422 7098 9450 7126
rect 9600 7098 10000 7112
rect 9422 7070 10000 7098
rect 0 7056 400 7070
rect 2757 7042 2762 7070
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2894 7042 2899 7070
rect 4913 7042 4918 7070
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 5050 7042 5055 7070
rect 7069 7042 7074 7070
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7206 7042 7211 7070
rect 9225 7042 9230 7070
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9362 7042 9367 7070
rect 9600 7056 10000 7070
rect 0 6762 400 6776
rect 0 6734 5110 6762
rect 5138 6734 5143 6762
rect 0 6720 400 6734
rect 1679 6650 1684 6678
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1816 6650 1821 6678
rect 3835 6650 3840 6678
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3972 6650 3977 6678
rect 5991 6650 5996 6678
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 6128 6650 6133 6678
rect 8147 6650 8152 6678
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8284 6650 8289 6678
rect 1017 6566 1022 6594
rect 1050 6566 3486 6594
rect 3514 6566 3519 6594
rect 3985 6510 3990 6538
rect 4018 6510 4382 6538
rect 4410 6510 4830 6538
rect 4858 6510 4863 6538
rect 6449 6510 6454 6538
rect 6482 6510 6846 6538
rect 6874 6510 8470 6538
rect 8498 6510 8503 6538
rect 5049 6454 5054 6482
rect 5082 6454 5558 6482
rect 5586 6454 5591 6482
rect 6953 6454 6958 6482
rect 6986 6454 7686 6482
rect 7714 6454 7719 6482
rect 0 6426 400 6440
rect 9600 6426 10000 6440
rect 0 6398 854 6426
rect 882 6398 887 6426
rect 9025 6398 9030 6426
rect 9058 6398 10000 6426
rect 0 6384 400 6398
rect 9600 6384 10000 6398
rect 2757 6258 2762 6286
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2894 6258 2899 6286
rect 4913 6258 4918 6286
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 5050 6258 5055 6286
rect 7069 6258 7074 6286
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7206 6258 7211 6286
rect 9225 6258 9230 6286
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9362 6258 9367 6286
rect 5889 6174 5894 6202
rect 5922 6174 7238 6202
rect 7266 6174 7271 6202
rect 0 6090 400 6104
rect 9600 6090 10000 6104
rect 0 6062 1190 6090
rect 1218 6062 1223 6090
rect 4937 6062 4942 6090
rect 4970 6062 5278 6090
rect 5306 6062 5311 6090
rect 5497 6062 5502 6090
rect 5530 6062 6902 6090
rect 6930 6062 6935 6090
rect 8185 6062 8190 6090
rect 8218 6062 10000 6090
rect 0 6048 400 6062
rect 9600 6048 10000 6062
rect 5553 6006 5558 6034
rect 5586 6006 7014 6034
rect 7042 6006 7047 6034
rect 1679 5866 1684 5894
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1816 5866 1821 5894
rect 3835 5866 3840 5894
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3972 5866 3977 5894
rect 5991 5866 5996 5894
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 6128 5866 6133 5894
rect 8147 5866 8152 5894
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8284 5866 8289 5894
rect 0 5754 400 5768
rect 9600 5754 10000 5768
rect 0 5726 854 5754
rect 882 5726 887 5754
rect 2977 5726 2982 5754
rect 3010 5726 3542 5754
rect 3570 5726 4046 5754
rect 4074 5726 4079 5754
rect 5609 5726 5614 5754
rect 5642 5726 6790 5754
rect 6818 5726 6823 5754
rect 9081 5726 9086 5754
rect 9114 5726 10000 5754
rect 0 5712 400 5726
rect 9600 5712 10000 5726
rect 1465 5670 1470 5698
rect 1498 5670 2646 5698
rect 2674 5670 2679 5698
rect 6449 5670 6454 5698
rect 6482 5670 6734 5698
rect 6762 5670 7658 5698
rect 4545 5614 4550 5642
rect 4578 5614 7182 5642
rect 7210 5614 7215 5642
rect 7630 5586 7658 5670
rect 6337 5558 6342 5586
rect 6370 5558 7294 5586
rect 7322 5558 7327 5586
rect 7625 5558 7630 5586
rect 7658 5558 7663 5586
rect 2757 5474 2762 5502
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2894 5474 2899 5502
rect 4913 5474 4918 5502
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 5050 5474 5055 5502
rect 7069 5474 7074 5502
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7206 5474 7211 5502
rect 9225 5474 9230 5502
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9362 5474 9367 5502
rect 1017 5446 1022 5474
rect 1050 5446 1055 5474
rect 0 5418 400 5432
rect 1022 5418 1050 5446
rect 9600 5418 10000 5432
rect 0 5390 1050 5418
rect 9025 5390 9030 5418
rect 9058 5390 10000 5418
rect 0 5376 400 5390
rect 9600 5376 10000 5390
rect 4186 5334 4438 5362
rect 4466 5334 4471 5362
rect 7905 5334 7910 5362
rect 7938 5334 8918 5362
rect 8946 5334 8951 5362
rect 4186 5250 4214 5334
rect 2641 5222 2646 5250
rect 2674 5222 3766 5250
rect 3794 5222 4214 5250
rect 6953 5222 6958 5250
rect 6986 5222 7742 5250
rect 7770 5222 7775 5250
rect 6113 5166 6118 5194
rect 6146 5166 8946 5194
rect 8918 5138 8946 5166
rect 8913 5110 8918 5138
rect 8946 5110 8951 5138
rect 0 5082 400 5096
rect 1679 5082 1684 5110
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1816 5082 1821 5110
rect 3835 5082 3840 5110
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3972 5082 3977 5110
rect 5991 5082 5996 5110
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 6128 5082 6133 5110
rect 8147 5082 8152 5110
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8284 5082 8289 5110
rect 9600 5082 10000 5096
rect 0 5054 854 5082
rect 882 5054 1246 5082
rect 1274 5054 1279 5082
rect 3369 5054 3374 5082
rect 3402 5054 3710 5082
rect 3738 5054 3743 5082
rect 9081 5054 9086 5082
rect 9114 5054 10000 5082
rect 0 5040 400 5054
rect 9600 5040 10000 5054
rect 1017 4942 1022 4970
rect 1050 4942 3038 4970
rect 3066 4942 3071 4970
rect 3089 4886 3094 4914
rect 3122 4886 3374 4914
rect 3402 4886 3407 4914
rect 4097 4886 4102 4914
rect 4130 4886 6846 4914
rect 6874 4886 6958 4914
rect 6986 4886 6991 4914
rect 3257 4774 3262 4802
rect 3290 4774 3430 4802
rect 3458 4774 3766 4802
rect 3794 4774 3799 4802
rect 8801 4774 8806 4802
rect 8834 4774 9086 4802
rect 9114 4774 9450 4802
rect 0 4746 400 4760
rect 9422 4746 9450 4774
rect 9600 4746 10000 4760
rect 0 4718 854 4746
rect 882 4718 1246 4746
rect 1274 4718 1279 4746
rect 9422 4718 10000 4746
rect 0 4704 400 4718
rect 2757 4690 2762 4718
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2894 4690 2899 4718
rect 4913 4690 4918 4718
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 5050 4690 5055 4718
rect 7069 4690 7074 4718
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7206 4690 7211 4718
rect 9225 4690 9230 4718
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9362 4690 9367 4718
rect 9600 4704 10000 4718
rect 6281 4606 6286 4634
rect 6314 4606 7182 4634
rect 7210 4606 7215 4634
rect 1353 4550 1358 4578
rect 1386 4550 2926 4578
rect 2954 4550 2959 4578
rect 4041 4550 4046 4578
rect 4074 4550 4270 4578
rect 4298 4550 4303 4578
rect 7121 4550 7126 4578
rect 7154 4550 8750 4578
rect 8778 4550 8783 4578
rect 3985 4494 3990 4522
rect 4018 4494 4158 4522
rect 4186 4494 4191 4522
rect 6225 4494 6230 4522
rect 6258 4494 6454 4522
rect 6482 4494 7350 4522
rect 7378 4494 8918 4522
rect 8946 4494 8951 4522
rect 3817 4438 3822 4466
rect 3850 4438 4214 4466
rect 4242 4438 4247 4466
rect 4433 4438 4438 4466
rect 4466 4438 6846 4466
rect 6874 4438 6879 4466
rect 0 4410 400 4424
rect 9600 4410 10000 4424
rect 0 4382 854 4410
rect 882 4382 1246 4410
rect 1274 4382 1279 4410
rect 4489 4382 4494 4410
rect 4522 4382 5838 4410
rect 5866 4382 6958 4410
rect 6986 4382 6991 4410
rect 8801 4382 8806 4410
rect 8834 4382 9086 4410
rect 9114 4382 10000 4410
rect 0 4368 400 4382
rect 9600 4368 10000 4382
rect 1679 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1821 4326
rect 3835 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3977 4326
rect 5991 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6133 4326
rect 8147 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8289 4326
rect 6953 4270 6958 4298
rect 6986 4270 7406 4298
rect 7434 4270 7439 4298
rect 3761 4214 3766 4242
rect 3794 4214 5502 4242
rect 5530 4214 5535 4242
rect 0 4074 400 4088
rect 9600 4074 10000 4088
rect 0 4046 854 4074
rect 882 4046 1246 4074
rect 1274 4046 1279 4074
rect 4153 4046 4158 4074
rect 4186 4046 4774 4074
rect 4802 4046 4807 4074
rect 6505 4046 6510 4074
rect 6538 4046 7126 4074
rect 7154 4046 8582 4074
rect 8610 4046 8615 4074
rect 9081 4046 9086 4074
rect 9114 4046 10000 4074
rect 0 4032 400 4046
rect 9600 4032 10000 4046
rect 1017 3990 1022 4018
rect 1050 3990 3094 4018
rect 3122 3990 3127 4018
rect 6785 3990 6790 4018
rect 6818 3990 7182 4018
rect 7210 3990 8918 4018
rect 8946 3990 8951 4018
rect 2757 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2899 3934
rect 4913 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5055 3934
rect 7069 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7211 3934
rect 9225 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9367 3934
rect 1017 3878 1022 3906
rect 1050 3878 2086 3906
rect 2114 3878 2119 3906
rect 961 3822 966 3850
rect 994 3822 2814 3850
rect 2842 3822 2847 3850
rect 4097 3822 4102 3850
rect 4130 3822 4326 3850
rect 4354 3822 4359 3850
rect 5553 3822 5558 3850
rect 5586 3822 5950 3850
rect 5978 3822 5983 3850
rect 910 3766 1190 3794
rect 1218 3766 1582 3794
rect 1610 3766 1615 3794
rect 6449 3766 6454 3794
rect 6482 3766 8470 3794
rect 8498 3766 8503 3794
rect 0 3738 400 3752
rect 910 3738 938 3766
rect 9600 3738 10000 3752
rect 0 3710 938 3738
rect 1073 3710 1078 3738
rect 1106 3710 1806 3738
rect 1834 3710 1839 3738
rect 8857 3710 8862 3738
rect 8890 3710 10000 3738
rect 0 3696 400 3710
rect 9600 3696 10000 3710
rect 849 3654 854 3682
rect 882 3654 1470 3682
rect 1498 3654 1503 3682
rect 1017 3598 1022 3626
rect 1050 3598 2198 3626
rect 2226 3598 2231 3626
rect 1679 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1821 3542
rect 3835 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3977 3542
rect 5991 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6133 3542
rect 8147 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8289 3542
rect 0 3402 400 3416
rect 0 3374 854 3402
rect 882 3374 887 3402
rect 1129 3374 1134 3402
rect 1162 3374 1862 3402
rect 1890 3374 1895 3402
rect 4321 3374 4326 3402
rect 4354 3374 5670 3402
rect 5698 3374 5703 3402
rect 0 3360 400 3374
rect 2305 3318 2310 3346
rect 2338 3318 4102 3346
rect 4130 3318 4382 3346
rect 4410 3318 4415 3346
rect 4713 3318 4718 3346
rect 4746 3318 5278 3346
rect 5306 3318 5311 3346
rect 3313 3262 3318 3290
rect 3346 3262 4046 3290
rect 4074 3262 4079 3290
rect 1185 3206 1190 3234
rect 1218 3206 1694 3234
rect 1722 3206 1727 3234
rect 2757 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2899 3150
rect 4913 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5055 3150
rect 7069 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7211 3150
rect 9225 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9367 3150
rect 0 3066 400 3080
rect 9600 3066 10000 3080
rect 0 3038 854 3066
rect 882 3038 1246 3066
rect 1274 3038 1279 3066
rect 9081 3038 9086 3066
rect 9114 3038 10000 3066
rect 0 3024 400 3038
rect 9600 3024 10000 3038
rect 1017 2982 1022 3010
rect 1050 2982 2982 3010
rect 3010 2982 3015 3010
rect 961 2926 966 2954
rect 994 2926 3598 2954
rect 3626 2926 3631 2954
rect 1297 2814 1302 2842
rect 1330 2814 2590 2842
rect 2618 2814 2623 2842
rect 0 2730 400 2744
rect 1679 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1821 2758
rect 3835 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3977 2758
rect 5991 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6133 2758
rect 8147 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8289 2758
rect 0 2702 854 2730
rect 882 2702 1246 2730
rect 1274 2702 1279 2730
rect 0 2688 400 2702
rect 2585 2590 2590 2618
rect 2618 2590 3598 2618
rect 3626 2590 3631 2618
rect 4769 2590 4774 2618
rect 4802 2590 6258 2618
rect 6230 2562 6258 2590
rect 3313 2534 3318 2562
rect 3346 2534 3766 2562
rect 3794 2534 3799 2562
rect 4041 2534 4046 2562
rect 4074 2534 5166 2562
rect 5194 2534 5199 2562
rect 6225 2534 6230 2562
rect 6258 2534 6263 2562
rect 905 2478 910 2506
rect 938 2478 1470 2506
rect 1498 2478 1503 2506
rect 3537 2478 3542 2506
rect 3570 2478 5278 2506
rect 5306 2478 5311 2506
rect 7737 2478 7742 2506
rect 7770 2478 8862 2506
rect 8890 2478 8895 2506
rect 0 2394 400 2408
rect 910 2394 938 2478
rect 1969 2422 1974 2450
rect 2002 2422 4662 2450
rect 4690 2422 4695 2450
rect 8353 2422 8358 2450
rect 8386 2422 8974 2450
rect 9002 2422 9007 2450
rect 0 2366 938 2394
rect 0 2352 400 2366
rect 2757 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2899 2366
rect 4913 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5055 2366
rect 7069 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7211 2366
rect 9225 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9367 2366
rect 1185 2254 1190 2282
rect 1218 2254 1582 2282
rect 1610 2254 1615 2282
rect 1689 2254 1694 2282
rect 1722 2254 4214 2282
rect 6393 2254 6398 2282
rect 6426 2254 7238 2282
rect 7266 2254 7271 2282
rect 7457 2254 7462 2282
rect 7490 2254 7854 2282
rect 7882 2254 7887 2282
rect 4186 2226 4214 2254
rect 1353 2198 1358 2226
rect 1386 2198 3374 2226
rect 3402 2198 3407 2226
rect 4186 2198 6118 2226
rect 6146 2198 6151 2226
rect 8241 2198 8246 2226
rect 8274 2198 8279 2226
rect 8246 2170 8274 2198
rect 849 2142 854 2170
rect 882 2142 1806 2170
rect 1834 2142 1839 2170
rect 3481 2142 3486 2170
rect 3514 2142 8274 2170
rect 8409 2142 8414 2170
rect 8442 2142 8582 2170
rect 8610 2142 9030 2170
rect 9058 2142 9063 2170
rect 3593 2086 3598 2114
rect 3626 2086 5054 2114
rect 5082 2086 5446 2114
rect 5474 2086 5479 2114
rect 6673 2086 6678 2114
rect 6706 2086 8918 2114
rect 8946 2086 8951 2114
rect 0 2058 400 2072
rect 9600 2058 10000 2072
rect 0 2030 854 2058
rect 882 2030 887 2058
rect 8745 2030 8750 2058
rect 8778 2030 10000 2058
rect 0 2016 400 2030
rect 9600 2016 10000 2030
rect 4433 1974 4438 2002
rect 4466 1974 5838 2002
rect 5866 1974 5871 2002
rect 1679 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1821 1974
rect 3835 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3977 1974
rect 5991 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6133 1974
rect 8147 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8289 1974
rect 9 1918 14 1946
rect 42 1918 1190 1946
rect 1218 1918 1223 1946
rect 401 1862 406 1890
rect 434 1862 1526 1890
rect 1554 1862 1559 1890
rect 1633 1862 1638 1890
rect 1666 1862 3374 1890
rect 3402 1862 3407 1890
rect 4489 1862 4494 1890
rect 4522 1862 8750 1890
rect 8778 1862 8783 1890
rect 1129 1806 1134 1834
rect 1162 1806 1167 1834
rect 0 1722 400 1736
rect 1134 1722 1162 1806
rect 2361 1750 2366 1778
rect 2394 1750 3374 1778
rect 3402 1750 3407 1778
rect 4377 1750 4382 1778
rect 4410 1750 5726 1778
rect 5754 1750 5950 1778
rect 5978 1750 5983 1778
rect 6393 1750 6398 1778
rect 6426 1750 7014 1778
rect 7042 1750 7047 1778
rect 7625 1750 7630 1778
rect 7658 1750 8022 1778
rect 8050 1750 8055 1778
rect 0 1694 1162 1722
rect 3201 1694 3206 1722
rect 3234 1694 5502 1722
rect 5530 1694 5535 1722
rect 6057 1694 6062 1722
rect 6090 1694 6678 1722
rect 6706 1694 6711 1722
rect 7401 1694 7406 1722
rect 7434 1694 7686 1722
rect 7714 1694 7719 1722
rect 8129 1694 8134 1722
rect 8162 1694 8582 1722
rect 8610 1694 8615 1722
rect 0 1680 400 1694
rect 5721 1638 5726 1666
rect 5754 1638 6174 1666
rect 6202 1638 6207 1666
rect 2757 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2899 1582
rect 4913 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5055 1582
rect 7069 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7211 1582
rect 9225 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9367 1582
rect 0 1386 400 1400
rect 0 1358 1750 1386
rect 1778 1358 1783 1386
rect 0 1344 400 1358
rect 0 1050 400 1064
rect 0 1022 1414 1050
rect 1442 1022 1447 1050
rect 0 1008 400 1022
<< via3 >>
rect 1684 8218 1712 8246
rect 1736 8218 1764 8246
rect 1788 8218 1816 8246
rect 3840 8218 3868 8246
rect 3892 8218 3920 8246
rect 3944 8218 3972 8246
rect 5996 8218 6024 8246
rect 6048 8218 6076 8246
rect 6100 8218 6128 8246
rect 8152 8218 8180 8246
rect 8204 8218 8232 8246
rect 8256 8218 8284 8246
rect 2762 7826 2790 7854
rect 2814 7826 2842 7854
rect 2866 7826 2894 7854
rect 4918 7826 4946 7854
rect 4970 7826 4998 7854
rect 5022 7826 5050 7854
rect 7074 7826 7102 7854
rect 7126 7826 7154 7854
rect 7178 7826 7206 7854
rect 9230 7826 9258 7854
rect 9282 7826 9310 7854
rect 9334 7826 9362 7854
rect 1684 7434 1712 7462
rect 1736 7434 1764 7462
rect 1788 7434 1816 7462
rect 3840 7434 3868 7462
rect 3892 7434 3920 7462
rect 3944 7434 3972 7462
rect 5996 7434 6024 7462
rect 6048 7434 6076 7462
rect 6100 7434 6128 7462
rect 8152 7434 8180 7462
rect 8204 7434 8232 7462
rect 8256 7434 8284 7462
rect 2762 7042 2790 7070
rect 2814 7042 2842 7070
rect 2866 7042 2894 7070
rect 4918 7042 4946 7070
rect 4970 7042 4998 7070
rect 5022 7042 5050 7070
rect 7074 7042 7102 7070
rect 7126 7042 7154 7070
rect 7178 7042 7206 7070
rect 9230 7042 9258 7070
rect 9282 7042 9310 7070
rect 9334 7042 9362 7070
rect 1684 6650 1712 6678
rect 1736 6650 1764 6678
rect 1788 6650 1816 6678
rect 3840 6650 3868 6678
rect 3892 6650 3920 6678
rect 3944 6650 3972 6678
rect 5996 6650 6024 6678
rect 6048 6650 6076 6678
rect 6100 6650 6128 6678
rect 8152 6650 8180 6678
rect 8204 6650 8232 6678
rect 8256 6650 8284 6678
rect 2762 6258 2790 6286
rect 2814 6258 2842 6286
rect 2866 6258 2894 6286
rect 4918 6258 4946 6286
rect 4970 6258 4998 6286
rect 5022 6258 5050 6286
rect 7074 6258 7102 6286
rect 7126 6258 7154 6286
rect 7178 6258 7206 6286
rect 9230 6258 9258 6286
rect 9282 6258 9310 6286
rect 9334 6258 9362 6286
rect 1684 5866 1712 5894
rect 1736 5866 1764 5894
rect 1788 5866 1816 5894
rect 3840 5866 3868 5894
rect 3892 5866 3920 5894
rect 3944 5866 3972 5894
rect 5996 5866 6024 5894
rect 6048 5866 6076 5894
rect 6100 5866 6128 5894
rect 8152 5866 8180 5894
rect 8204 5866 8232 5894
rect 8256 5866 8284 5894
rect 2762 5474 2790 5502
rect 2814 5474 2842 5502
rect 2866 5474 2894 5502
rect 4918 5474 4946 5502
rect 4970 5474 4998 5502
rect 5022 5474 5050 5502
rect 7074 5474 7102 5502
rect 7126 5474 7154 5502
rect 7178 5474 7206 5502
rect 9230 5474 9258 5502
rect 9282 5474 9310 5502
rect 9334 5474 9362 5502
rect 1684 5082 1712 5110
rect 1736 5082 1764 5110
rect 1788 5082 1816 5110
rect 3840 5082 3868 5110
rect 3892 5082 3920 5110
rect 3944 5082 3972 5110
rect 5996 5082 6024 5110
rect 6048 5082 6076 5110
rect 6100 5082 6128 5110
rect 8152 5082 8180 5110
rect 8204 5082 8232 5110
rect 8256 5082 8284 5110
rect 2762 4690 2790 4718
rect 2814 4690 2842 4718
rect 2866 4690 2894 4718
rect 4918 4690 4946 4718
rect 4970 4690 4998 4718
rect 5022 4690 5050 4718
rect 7074 4690 7102 4718
rect 7126 4690 7154 4718
rect 7178 4690 7206 4718
rect 9230 4690 9258 4718
rect 9282 4690 9310 4718
rect 9334 4690 9362 4718
rect 1684 4298 1712 4326
rect 1736 4298 1764 4326
rect 1788 4298 1816 4326
rect 3840 4298 3868 4326
rect 3892 4298 3920 4326
rect 3944 4298 3972 4326
rect 5996 4298 6024 4326
rect 6048 4298 6076 4326
rect 6100 4298 6128 4326
rect 8152 4298 8180 4326
rect 8204 4298 8232 4326
rect 8256 4298 8284 4326
rect 2762 3906 2790 3934
rect 2814 3906 2842 3934
rect 2866 3906 2894 3934
rect 4918 3906 4946 3934
rect 4970 3906 4998 3934
rect 5022 3906 5050 3934
rect 7074 3906 7102 3934
rect 7126 3906 7154 3934
rect 7178 3906 7206 3934
rect 9230 3906 9258 3934
rect 9282 3906 9310 3934
rect 9334 3906 9362 3934
rect 1684 3514 1712 3542
rect 1736 3514 1764 3542
rect 1788 3514 1816 3542
rect 3840 3514 3868 3542
rect 3892 3514 3920 3542
rect 3944 3514 3972 3542
rect 5996 3514 6024 3542
rect 6048 3514 6076 3542
rect 6100 3514 6128 3542
rect 8152 3514 8180 3542
rect 8204 3514 8232 3542
rect 8256 3514 8284 3542
rect 2762 3122 2790 3150
rect 2814 3122 2842 3150
rect 2866 3122 2894 3150
rect 4918 3122 4946 3150
rect 4970 3122 4998 3150
rect 5022 3122 5050 3150
rect 7074 3122 7102 3150
rect 7126 3122 7154 3150
rect 7178 3122 7206 3150
rect 9230 3122 9258 3150
rect 9282 3122 9310 3150
rect 9334 3122 9362 3150
rect 1684 2730 1712 2758
rect 1736 2730 1764 2758
rect 1788 2730 1816 2758
rect 3840 2730 3868 2758
rect 3892 2730 3920 2758
rect 3944 2730 3972 2758
rect 5996 2730 6024 2758
rect 6048 2730 6076 2758
rect 6100 2730 6128 2758
rect 8152 2730 8180 2758
rect 8204 2730 8232 2758
rect 8256 2730 8284 2758
rect 2762 2338 2790 2366
rect 2814 2338 2842 2366
rect 2866 2338 2894 2366
rect 4918 2338 4946 2366
rect 4970 2338 4998 2366
rect 5022 2338 5050 2366
rect 7074 2338 7102 2366
rect 7126 2338 7154 2366
rect 7178 2338 7206 2366
rect 9230 2338 9258 2366
rect 9282 2338 9310 2366
rect 9334 2338 9362 2366
rect 1684 1946 1712 1974
rect 1736 1946 1764 1974
rect 1788 1946 1816 1974
rect 3840 1946 3868 1974
rect 3892 1946 3920 1974
rect 3944 1946 3972 1974
rect 5996 1946 6024 1974
rect 6048 1946 6076 1974
rect 6100 1946 6128 1974
rect 8152 1946 8180 1974
rect 8204 1946 8232 1974
rect 8256 1946 8284 1974
rect 2762 1554 2790 1582
rect 2814 1554 2842 1582
rect 2866 1554 2894 1582
rect 4918 1554 4946 1582
rect 4970 1554 4998 1582
rect 5022 1554 5050 1582
rect 7074 1554 7102 1582
rect 7126 1554 7154 1582
rect 7178 1554 7206 1582
rect 9230 1554 9258 1582
rect 9282 1554 9310 1582
rect 9334 1554 9362 1582
<< metal4 >>
rect 1670 8246 1830 8262
rect 1670 8218 1684 8246
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1816 8218 1830 8246
rect 1670 7462 1830 8218
rect 1670 7434 1684 7462
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1816 7434 1830 7462
rect 1670 6678 1830 7434
rect 1670 6650 1684 6678
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1816 6650 1830 6678
rect 1670 5894 1830 6650
rect 1670 5866 1684 5894
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1816 5866 1830 5894
rect 1670 5110 1830 5866
rect 1670 5082 1684 5110
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1816 5082 1830 5110
rect 1670 4326 1830 5082
rect 1670 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1830 4326
rect 1670 3542 1830 4298
rect 1670 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1830 3542
rect 1670 2758 1830 3514
rect 1670 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1830 2758
rect 1670 1974 1830 2730
rect 1670 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1830 1974
rect 1670 1538 1830 1946
rect 2748 7854 2908 8262
rect 2748 7826 2762 7854
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2894 7826 2908 7854
rect 2748 7070 2908 7826
rect 2748 7042 2762 7070
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2894 7042 2908 7070
rect 2748 6286 2908 7042
rect 2748 6258 2762 6286
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2894 6258 2908 6286
rect 2748 5502 2908 6258
rect 2748 5474 2762 5502
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2894 5474 2908 5502
rect 2748 4718 2908 5474
rect 2748 4690 2762 4718
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2894 4690 2908 4718
rect 2748 3934 2908 4690
rect 2748 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2908 3934
rect 2748 3150 2908 3906
rect 2748 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2908 3150
rect 2748 2366 2908 3122
rect 2748 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2908 2366
rect 2748 1582 2908 2338
rect 2748 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2908 1582
rect 2748 1538 2908 1554
rect 3826 8246 3986 8262
rect 3826 8218 3840 8246
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3972 8218 3986 8246
rect 3826 7462 3986 8218
rect 3826 7434 3840 7462
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3972 7434 3986 7462
rect 3826 6678 3986 7434
rect 3826 6650 3840 6678
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3972 6650 3986 6678
rect 3826 5894 3986 6650
rect 3826 5866 3840 5894
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3972 5866 3986 5894
rect 3826 5110 3986 5866
rect 3826 5082 3840 5110
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3972 5082 3986 5110
rect 3826 4326 3986 5082
rect 3826 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3986 4326
rect 3826 3542 3986 4298
rect 3826 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3986 3542
rect 3826 2758 3986 3514
rect 3826 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3986 2758
rect 3826 1974 3986 2730
rect 3826 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3986 1974
rect 3826 1538 3986 1946
rect 4904 7854 5064 8262
rect 4904 7826 4918 7854
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 5050 7826 5064 7854
rect 4904 7070 5064 7826
rect 4904 7042 4918 7070
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 5050 7042 5064 7070
rect 4904 6286 5064 7042
rect 4904 6258 4918 6286
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 5050 6258 5064 6286
rect 4904 5502 5064 6258
rect 4904 5474 4918 5502
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 5050 5474 5064 5502
rect 4904 4718 5064 5474
rect 4904 4690 4918 4718
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 5050 4690 5064 4718
rect 4904 3934 5064 4690
rect 4904 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5064 3934
rect 4904 3150 5064 3906
rect 4904 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5064 3150
rect 4904 2366 5064 3122
rect 4904 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5064 2366
rect 4904 1582 5064 2338
rect 4904 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5064 1582
rect 4904 1538 5064 1554
rect 5982 8246 6142 8262
rect 5982 8218 5996 8246
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 6128 8218 6142 8246
rect 5982 7462 6142 8218
rect 5982 7434 5996 7462
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 6128 7434 6142 7462
rect 5982 6678 6142 7434
rect 5982 6650 5996 6678
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 6128 6650 6142 6678
rect 5982 5894 6142 6650
rect 5982 5866 5996 5894
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 6128 5866 6142 5894
rect 5982 5110 6142 5866
rect 5982 5082 5996 5110
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 6128 5082 6142 5110
rect 5982 4326 6142 5082
rect 5982 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6142 4326
rect 5982 3542 6142 4298
rect 5982 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6142 3542
rect 5982 2758 6142 3514
rect 5982 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6142 2758
rect 5982 1974 6142 2730
rect 5982 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6142 1974
rect 5982 1538 6142 1946
rect 7060 7854 7220 8262
rect 7060 7826 7074 7854
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7206 7826 7220 7854
rect 7060 7070 7220 7826
rect 7060 7042 7074 7070
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7206 7042 7220 7070
rect 7060 6286 7220 7042
rect 7060 6258 7074 6286
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7206 6258 7220 6286
rect 7060 5502 7220 6258
rect 7060 5474 7074 5502
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7206 5474 7220 5502
rect 7060 4718 7220 5474
rect 7060 4690 7074 4718
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7206 4690 7220 4718
rect 7060 3934 7220 4690
rect 7060 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7220 3934
rect 7060 3150 7220 3906
rect 7060 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7220 3150
rect 7060 2366 7220 3122
rect 7060 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7220 2366
rect 7060 1582 7220 2338
rect 7060 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7220 1582
rect 7060 1538 7220 1554
rect 8138 8246 8298 8262
rect 8138 8218 8152 8246
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8284 8218 8298 8246
rect 8138 7462 8298 8218
rect 8138 7434 8152 7462
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8284 7434 8298 7462
rect 8138 6678 8298 7434
rect 8138 6650 8152 6678
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8284 6650 8298 6678
rect 8138 5894 8298 6650
rect 8138 5866 8152 5894
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8284 5866 8298 5894
rect 8138 5110 8298 5866
rect 8138 5082 8152 5110
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8284 5082 8298 5110
rect 8138 4326 8298 5082
rect 8138 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8298 4326
rect 8138 3542 8298 4298
rect 8138 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8298 3542
rect 8138 2758 8298 3514
rect 8138 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8298 2758
rect 8138 1974 8298 2730
rect 8138 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8298 1974
rect 8138 1538 8298 1946
rect 9216 7854 9376 8262
rect 9216 7826 9230 7854
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9362 7826 9376 7854
rect 9216 7070 9376 7826
rect 9216 7042 9230 7070
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9362 7042 9376 7070
rect 9216 6286 9376 7042
rect 9216 6258 9230 6286
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9362 6258 9376 6286
rect 9216 5502 9376 6258
rect 9216 5474 9230 5502
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9362 5474 9376 5502
rect 9216 4718 9376 5474
rect 9216 4690 9230 4718
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9362 4690 9376 4718
rect 9216 3934 9376 4690
rect 9216 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9376 3934
rect 9216 3150 9376 3906
rect 9216 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9376 3150
rect 9216 2366 9376 3122
rect 9216 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9376 2366
rect 9216 1582 9376 2338
rect 9216 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9376 1582
rect 9216 1538 9376 1554
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _040_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2968 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _041_
timestamp 1698431365
transform 1 0 3416 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _042_
timestamp 1698431365
transform -1 0 4928 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _043_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8008 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _044_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4592 0 -1 2352
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _045_
timestamp 1698431365
transform -1 0 6776 0 -1 2352
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _046_
timestamp 1698431365
transform 1 0 2520 0 -1 3136
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _047_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6160 0 -1 4704
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _048_
timestamp 1698431365
transform 1 0 5824 0 -1 3920
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _049_
timestamp 1698431365
transform 1 0 5768 0 -1 3136
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _050_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4928 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _051_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _052_
timestamp 1698431365
transform 1 0 1736 0 -1 3920
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _053_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2072 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _054_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4256 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _055_
timestamp 1698431365
transform -1 0 5320 0 1 3136
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _056_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3864 0 -1 4704
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _057_
timestamp 1698431365
transform 1 0 4144 0 1 4704
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _058_
timestamp 1698431365
transform 1 0 4256 0 -1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _059_
timestamp 1698431365
transform 1 0 4256 0 1 3920
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _060_
timestamp 1698431365
transform -1 0 4592 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _061_
timestamp 1698431365
transform -1 0 6944 0 1 4704
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _062_
timestamp 1698431365
transform 1 0 6664 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _063_
timestamp 1698431365
transform -1 0 7280 0 1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _064_
timestamp 1698431365
transform 1 0 6216 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _065_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6888 0 -1 4704
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _066_
timestamp 1698431365
transform 1 0 4704 0 -1 6272
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _067_
timestamp 1698431365
transform -1 0 4480 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _068_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6664 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _069_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5264 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _070_
timestamp 1698431365
transform 1 0 5880 0 1 5488
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _071_
timestamp 1698431365
transform 1 0 4312 0 -1 5488
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _072_
timestamp 1698431365
transform 1 0 7560 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _073_
timestamp 1698431365
transform 1 0 7112 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _074_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6160 0 -1 4704
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _075_
timestamp 1698431365
transform -1 0 6104 0 1 2352
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _076_
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _077_
timestamp 1698431365
transform 1 0 3360 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _078_
timestamp 1698431365
transform 1 0 3696 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _079_
timestamp 1698431365
transform 1 0 3192 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _080_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6944 0 1 4704
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _081_
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _082_
timestamp 1698431365
transform 1 0 5432 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _083_
timestamp 1698431365
transform 1 0 2856 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _084_
timestamp 1698431365
transform -1 0 4200 0 -1 5488
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5096 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 8848 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 8848 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 1680 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 1680 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 9184 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 8624 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 5432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 5768 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 8848 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 8400 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 7784 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 7336 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 7112 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 1456 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 7840 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 7504 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 8176 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 6888 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 1232 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 1232 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 1456 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 1232 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 1232 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 1568 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 1904 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 1456 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 1232 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 2520 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 1904 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 3360 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 1680 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 6216 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 5096 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 8848 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 896 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 1232 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 9184 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 8848 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 8848 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4872 0 -1 5488
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 5880 0 1 5488
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 5712 0 -1 6272
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_6 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1008 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_25 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2072 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_27
timestamp 1698431365
transform 1 0 2184 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_72
timestamp 1698431365
transform 1 0 4704 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 6328 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_134
timestamp 1698431365
transform 1 0 8176 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_150
timestamp 1698431365
transform 1 0 9072 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_24
timestamp 1698431365
transform 1 0 2016 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_109
timestamp 1698431365
transform 1 0 6776 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_113
timestamp 1698431365
transform 1 0 7000 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_117
timestamp 1698431365
transform 1 0 7224 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_121 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7448 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_133
timestamp 1698431365
transform 1 0 8120 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698431365
transform 1 0 8736 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_151
timestamp 1698431365
transform 1 0 9128 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_16
timestamp 1698431365
transform 1 0 1568 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_20
timestamp 1698431365
transform 1 0 1792 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_24
timestamp 1698431365
transform 1 0 2016 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_29
timestamp 1698431365
transform 1 0 2296 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 2744 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_39
timestamp 1698431365
transform 1 0 2856 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_44
timestamp 1698431365
transform 1 0 3136 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_97
timestamp 1698431365
transform 1 0 6104 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_107 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6664 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_115
timestamp 1698431365
transform 1 0 7112 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_119
timestamp 1698431365
transform 1 0 7336 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_122
timestamp 1698431365
transform 1 0 7504 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_128
timestamp 1698431365
transform 1 0 7840 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_134
timestamp 1698431365
transform 1 0 8176 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_138
timestamp 1698431365
transform 1 0 8400 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_8
timestamp 1698431365
transform 1 0 1120 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_12
timestamp 1698431365
transform 1 0 1344 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_16
timestamp 1698431365
transform 1 0 1568 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_20
timestamp 1698431365
transform 1 0 1792 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_24
timestamp 1698431365
transform 1 0 2016 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_28
timestamp 1698431365
transform 1 0 2240 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_30
timestamp 1698431365
transform 1 0 2352 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_72
timestamp 1698431365
transform 1 0 4704 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_76
timestamp 1698431365
transform 1 0 4928 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_79
timestamp 1698431365
transform 1 0 5096 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_85
timestamp 1698431365
transform 1 0 5432 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_128
timestamp 1698431365
transform 1 0 7840 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 8624 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_146
timestamp 1698431365
transform 1 0 8848 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_8
timestamp 1698431365
transform 1 0 1120 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_12
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_16
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_20
timestamp 1698431365
transform 1 0 1792 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_28
timestamp 1698431365
transform 1 0 2240 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_37
timestamp 1698431365
transform 1 0 2744 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_45
timestamp 1698431365
transform 1 0 3192 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_83 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5320 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_99
timestamp 1698431365
transform 1 0 6216 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 6440 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_107 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6664 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_139
timestamp 1698431365
transform 1 0 8456 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_147
timestamp 1698431365
transform 1 0 8904 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_8
timestamp 1698431365
transform 1 0 1120 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_12
timestamp 1698431365
transform 1 0 1344 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_16
timestamp 1698431365
transform 1 0 1568 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_18
timestamp 1698431365
transform 1 0 1680 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 4536 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_129
timestamp 1698431365
transform 1 0 7896 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_137
timestamp 1698431365
transform 1 0 8344 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 8456 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_142
timestamp 1698431365
transform 1 0 8624 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_148
timestamp 1698431365
transform 1 0 8960 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_14
timestamp 1698431365
transform 1 0 1456 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_18
timestamp 1698431365
transform 1 0 1680 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_22
timestamp 1698431365
transform 1 0 1904 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_30
timestamp 1698431365
transform 1 0 2352 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_37
timestamp 1698431365
transform 1 0 2744 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_53
timestamp 1698431365
transform 1 0 3640 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_61
timestamp 1698431365
transform 1 0 4088 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_63
timestamp 1698431365
transform 1 0 4200 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_118
timestamp 1698431365
transform 1 0 7280 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_134
timestamp 1698431365
transform 1 0 8176 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_138
timestamp 1698431365
transform 1 0 8400 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 1120 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_12
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_20
timestamp 1698431365
transform 1 0 1792 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_24
timestamp 1698431365
transform 1 0 2016 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_62
timestamp 1698431365
transform 1 0 4144 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_121
timestamp 1698431365
transform 1 0 7448 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 8344 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 8456 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698431365
transform 1 0 1120 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_37
timestamp 1698431365
transform 1 0 2744 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_53
timestamp 1698431365
transform 1 0 3640 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_141
timestamp 1698431365
transform 1 0 8568 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_143
timestamp 1698431365
transform 1 0 8680 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_8
timestamp 1698431365
transform 1 0 1120 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_12
timestamp 1698431365
transform 1 0 1344 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_28
timestamp 1698431365
transform 1 0 2240 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_32
timestamp 1698431365
transform 1 0 2464 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_63
timestamp 1698431365
transform 1 0 4200 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 4704 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_74
timestamp 1698431365
transform 1 0 4816 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_131
timestamp 1698431365
transform 1 0 8008 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 8456 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 8624 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_16
timestamp 1698431365
transform 1 0 1568 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 2464 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_37
timestamp 1698431365
transform 1 0 2744 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_41
timestamp 1698431365
transform 1 0 2968 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 6440 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_131
timestamp 1698431365
transform 1 0 8008 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_135
timestamp 1698431365
transform 1 0 8232 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_137
timestamp 1698431365
transform 1 0 8344 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_6
timestamp 1698431365
transform 1 0 1008 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_38
timestamp 1698431365
transform 1 0 2800 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_46
timestamp 1698431365
transform 1 0 3248 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_64
timestamp 1698431365
transform 1 0 4256 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_77
timestamp 1698431365
transform 1 0 4984 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_81
timestamp 1698431365
transform 1 0 5208 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698431365
transform 1 0 2240 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 2744 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_68
timestamp 1698431365
transform 1 0 4480 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698431365
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_123
timestamp 1698431365
transform 1 0 7560 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_2
timestamp 1698431365
transform 1 0 784 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_6
timestamp 1698431365
transform 1 0 1008 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_38
timestamp 1698431365
transform 1 0 2800 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_46
timestamp 1698431365
transform 1 0 3248 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_48
timestamp 1698431365
transform 1 0 3360 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_53
timestamp 1698431365
transform 1 0 3640 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 4536 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698431365
transform 1 0 4704 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_80
timestamp 1698431365
transform 1 0 5152 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_84
timestamp 1698431365
transform 1 0 5376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_114
timestamp 1698431365
transform 1 0 7056 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_130
timestamp 1698431365
transform 1 0 7952 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 8400 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 8624 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 9072 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_6
timestamp 1698431365
transform 1 0 1008 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_22
timestamp 1698431365
transform 1 0 1904 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_30
timestamp 1698431365
transform 1 0 2352 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698431365
transform 1 0 6664 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_139
timestamp 1698431365
transform 1 0 8456 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_147
timestamp 1698431365
transform 1 0 8904 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_6
timestamp 1698431365
transform 1 0 1008 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_72
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_77
timestamp 1698431365
transform 1 0 4984 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_109
timestamp 1698431365
transform 1 0 6776 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_125
timestamp 1698431365
transform 1 0 7672 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698431365
transform 1 0 8120 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 8344 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 8456 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698431365
transform 1 0 8848 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_14
timestamp 1698431365
transform 1 0 1456 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_30
timestamp 1698431365
transform 1 0 2352 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_36
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_40
timestamp 1698431365
transform 1 0 2912 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_42
timestamp 1698431365
transform 1 0 3024 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_47
timestamp 1698431365
transform 1 0 3304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_53
timestamp 1698431365
transform 1 0 3640 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_59
timestamp 1698431365
transform 1 0 3976 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_63
timestamp 1698431365
transform 1 0 4200 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_80
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_84
timestamp 1698431365
transform 1 0 5376 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_89
timestamp 1698431365
transform 1 0 5656 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_95
timestamp 1698431365
transform 1 0 5992 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_99
timestamp 1698431365
transform 1 0 6216 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_101
timestamp 1698431365
transform 1 0 6328 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_104
timestamp 1698431365
transform 1 0 6496 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_108
timestamp 1698431365
transform 1 0 6720 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_113
timestamp 1698431365
transform 1 0 7000 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698431365
transform 1 0 7336 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_125
timestamp 1698431365
transform 1 0 7672 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_133
timestamp 1698431365
transform 1 0 8120 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_135
timestamp 1698431365
transform 1 0 8232 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_138
timestamp 1698431365
transform 1 0 8400 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_146
timestamp 1698431365
transform 1 0 8848 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 9184 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1120 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 1456 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 9184 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 8512 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 5768 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 6104 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 9072 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 9128 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 8120 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 7504 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 7168 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1698431365
transform 1 0 1400 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 8176 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 7840 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 8736 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 6832 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 784 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 784 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 784 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 784 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 784 0 -1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 1120 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698431365
transform 1 0 1736 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 784 0 -1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 784 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input28
timestamp 1698431365
transform 1 0 2240 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 784 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 3696 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 1064 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 3696 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 4760 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 5432 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 8848 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 784 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 784 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input38
timestamp 1698431365
transform -1 0 9184 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input39
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform -1 0 9184 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output41 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5152 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output42 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 1568 0 1 5488
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output43 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8400 0 1 5488
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output44
timestamp 1698431365
transform 1 0 8400 0 1 6272
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output45
timestamp 1698431365
transform 1 0 7616 0 1 6272
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_17 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 9296 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_18
timestamp 1698431365
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_19
timestamp 1698431365
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 9296 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_20
timestamp 1698431365
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 9296 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_21
timestamp 1698431365
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 9296 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_22
timestamp 1698431365
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 9296 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_23
timestamp 1698431365
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 9296 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_24
timestamp 1698431365
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 9296 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_25
timestamp 1698431365
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 9296 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_26
timestamp 1698431365
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 9296 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_27
timestamp 1698431365
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 9296 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_28
timestamp 1698431365
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 9296 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_29
timestamp 1698431365
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 9296 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_30
timestamp 1698431365
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 9296 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_31
timestamp 1698431365
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 9296 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_32
timestamp 1698431365
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 9296 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_33
timestamp 1698431365
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 9296 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1698431365
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_38
timestamp 1698431365
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1698431365
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_40
timestamp 1698431365
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_41
timestamp 1698431365
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_42
timestamp 1698431365
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_43
timestamp 1698431365
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_44
timestamp 1698431365
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_45
timestamp 1698431365
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_46
timestamp 1698431365
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_47
timestamp 1698431365
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_48
timestamp 1698431365
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_49
timestamp 1698431365
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_50
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_51
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_52
timestamp 1698431365
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_53
timestamp 1698431365
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_54
timestamp 1698431365
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_55
timestamp 1698431365
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_56
timestamp 1698431365
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_57
timestamp 1698431365
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_58
timestamp 1698431365
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_59
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_60
timestamp 1698431365
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_61
timestamp 1698431365
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_62
timestamp 1698431365
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_63
timestamp 1698431365
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_64
timestamp 1698431365
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_65
timestamp 1698431365
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_66
timestamp 1698431365
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_67
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_68
timestamp 1698431365
transform 1 0 2576 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_69
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_70
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_71
timestamp 1698431365
transform 1 0 8288 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_46 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2296 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_47
timestamp 1698431365
transform -1 0 5656 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_48
timestamp 1698431365
transform -1 0 7000 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_49
timestamp 1698431365
transform -1 0 7336 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_50
timestamp 1698431365
transform -1 0 1008 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_51
timestamp 1698431365
transform -1 0 1232 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_52
timestamp 1698431365
transform -1 0 1008 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_53
timestamp 1698431365
transform -1 0 5992 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_54
timestamp 1698431365
transform -1 0 2296 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_55
timestamp 1698431365
transform -1 0 1344 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_56
timestamp 1698431365
transform -1 0 1568 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_57
timestamp 1698431365
transform 1 0 8624 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_58
timestamp 1698431365
transform -1 0 4984 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_59
timestamp 1698431365
transform -1 0 1456 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_60
timestamp 1698431365
transform -1 0 3304 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_61
timestamp 1698431365
transform -1 0 3976 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_62
timestamp 1698431365
transform -1 0 1008 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_63
timestamp 1698431365
transform 1 0 2912 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_64
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_65
timestamp 1698431365
transform 1 0 2072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_66
timestamp 1698431365
transform 1 0 8960 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_67
timestamp 1698431365
transform -1 0 7672 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_68
timestamp 1698431365
transform -1 0 1008 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_69
timestamp 1698431365
transform -1 0 3640 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_70
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_71
timestamp 1698431365
transform -1 0 2016 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_72
timestamp 1698431365
transform -1 0 6328 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_73
timestamp 1698431365
transform -1 0 1344 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_74
timestamp 1698431365
transform 1 0 8960 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_75
timestamp 1698431365
transform -1 0 1008 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_76
timestamp 1698431365
transform 1 0 4256 0 1 7840
box -43 -43 267 435
<< labels >>
flabel metal4 s 1670 1538 1830 8262 0 FreeSans 640 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 3826 1538 3986 8262 0 FreeSans 640 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 5982 1538 6142 8262 0 FreeSans 640 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 8138 1538 8298 8262 0 FreeSans 640 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 2748 1538 2908 8262 0 FreeSans 640 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 4904 1538 5064 8262 0 FreeSans 640 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 7060 1538 7220 8262 0 FreeSans 640 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 9216 1538 9376 8262 0 FreeSans 640 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 s 9600 5712 10000 5768 0 FreeSans 224 0 0 0 buttons[0]
port 2 nsew signal input
flabel metal3 s 9600 4704 10000 4760 0 FreeSans 224 0 0 0 buttons[1]
port 3 nsew signal input
flabel metal3 s 0 6720 400 6776 0 FreeSans 224 0 0 0 clk
port 4 nsew signal input
flabel metal2 s 0 0 56 400 0 FreeSans 224 90 0 0 i_wb_addr[0]
port 5 nsew signal input
flabel metal2 s 336 0 392 400 0 FreeSans 224 90 0 0 i_wb_addr[10]
port 6 nsew signal input
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 i_wb_addr[11]
port 7 nsew signal input
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 i_wb_addr[12]
port 8 nsew signal input
flabel metal2 s 5376 0 5432 400 0 FreeSans 224 90 0 0 i_wb_addr[13]
port 9 nsew signal input
flabel metal2 s 4368 0 4424 400 0 FreeSans 224 90 0 0 i_wb_addr[14]
port 10 nsew signal input
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 i_wb_addr[15]
port 11 nsew signal input
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 i_wb_addr[16]
port 12 nsew signal input
flabel metal2 s 7728 0 7784 400 0 FreeSans 224 90 0 0 i_wb_addr[17]
port 13 nsew signal input
flabel metal2 s 6720 0 6776 400 0 FreeSans 224 90 0 0 i_wb_addr[18]
port 14 nsew signal input
flabel metal2 s 6384 0 6440 400 0 FreeSans 224 90 0 0 i_wb_addr[19]
port 15 nsew signal input
flabel metal2 s 1344 0 1400 400 0 FreeSans 224 90 0 0 i_wb_addr[1]
port 16 nsew signal input
flabel metal2 s 7392 0 7448 400 0 FreeSans 224 90 0 0 i_wb_addr[20]
port 17 nsew signal input
flabel metal2 s 7056 0 7112 400 0 FreeSans 224 90 0 0 i_wb_addr[21]
port 18 nsew signal input
flabel metal2 s 8064 0 8120 400 0 FreeSans 224 90 0 0 i_wb_addr[22]
port 19 nsew signal input
flabel metal2 s 6048 0 6104 400 0 FreeSans 224 90 0 0 i_wb_addr[23]
port 20 nsew signal input
flabel metal3 s 0 4368 400 4424 0 FreeSans 224 0 0 0 i_wb_addr[24]
port 21 nsew signal input
flabel metal3 s 0 4032 400 4088 0 FreeSans 224 0 0 0 i_wb_addr[25]
port 22 nsew signal input
flabel metal3 s 0 2352 400 2408 0 FreeSans 224 0 0 0 i_wb_addr[26]
port 23 nsew signal input
flabel metal3 s 0 4704 400 4760 0 FreeSans 224 0 0 0 i_wb_addr[27]
port 24 nsew signal input
flabel metal3 s 0 2688 400 2744 0 FreeSans 224 0 0 0 i_wb_addr[28]
port 25 nsew signal input
flabel metal3 s 0 3696 400 3752 0 FreeSans 224 0 0 0 i_wb_addr[29]
port 26 nsew signal input
flabel metal2 s 1680 0 1736 400 0 FreeSans 224 90 0 0 i_wb_addr[2]
port 27 nsew signal input
flabel metal3 s 0 3360 400 3416 0 FreeSans 224 0 0 0 i_wb_addr[30]
port 28 nsew signal input
flabel metal3 s 0 3024 400 3080 0 FreeSans 224 0 0 0 i_wb_addr[31]
port 29 nsew signal input
flabel metal2 s 3360 0 3416 400 0 FreeSans 224 90 0 0 i_wb_addr[3]
port 30 nsew signal input
flabel metal2 s 672 0 728 400 0 FreeSans 224 90 0 0 i_wb_addr[4]
port 31 nsew signal input
flabel metal2 s 4032 0 4088 400 0 FreeSans 224 90 0 0 i_wb_addr[5]
port 32 nsew signal input
flabel metal2 s 1008 0 1064 400 0 FreeSans 224 90 0 0 i_wb_addr[6]
port 33 nsew signal input
flabel metal2 s 3696 0 3752 400 0 FreeSans 224 90 0 0 i_wb_addr[7]
port 34 nsew signal input
flabel metal2 s 4704 0 4760 400 0 FreeSans 224 90 0 0 i_wb_addr[8]
port 35 nsew signal input
flabel metal2 s 5040 0 5096 400 0 FreeSans 224 90 0 0 i_wb_addr[9]
port 36 nsew signal input
flabel metal3 s 9600 3696 10000 3752 0 FreeSans 224 0 0 0 i_wb_cyc
port 37 nsew signal input
flabel metal3 s 0 6384 400 6440 0 FreeSans 224 0 0 0 i_wb_data[0]
port 38 nsew signal input
flabel metal3 s 0 5040 400 5096 0 FreeSans 224 0 0 0 i_wb_data[1]
port 39 nsew signal input
flabel metal3 s 9600 4032 10000 4088 0 FreeSans 224 0 0 0 i_wb_stb
port 40 nsew signal input
flabel metal3 s 9600 4368 10000 4424 0 FreeSans 224 0 0 0 i_wb_we
port 41 nsew signal input
flabel metal2 s 4032 9600 4088 10000 0 FreeSans 224 90 0 0 leds[0]
port 42 nsew signal tristate
flabel metal3 s 0 5376 400 5432 0 FreeSans 224 0 0 0 leds[1]
port 43 nsew signal tristate
flabel metal3 s 9600 5376 10000 5432 0 FreeSans 224 0 0 0 o_wb_ack
port 44 nsew signal tristate
flabel metal3 s 9600 6384 10000 6440 0 FreeSans 224 0 0 0 o_wb_data[0]
port 45 nsew signal tristate
flabel metal2 s 2016 0 2072 400 0 FreeSans 224 90 0 0 o_wb_data[10]
port 46 nsew signal tristate
flabel metal3 s 0 6048 400 6104 0 FreeSans 224 0 0 0 o_wb_data[11]
port 47 nsew signal tristate
flabel metal3 s 0 1008 400 1064 0 FreeSans 224 0 0 0 o_wb_data[12]
port 48 nsew signal tristate
flabel metal3 s 9600 2016 10000 2072 0 FreeSans 224 0 0 0 o_wb_data[13]
port 49 nsew signal tristate
flabel metal2 s 4704 9600 4760 10000 0 FreeSans 224 90 0 0 o_wb_data[14]
port 50 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 o_wb_data[15]
port 51 nsew signal tristate
flabel metal2 s 3024 9600 3080 10000 0 FreeSans 224 90 0 0 o_wb_data[16]
port 52 nsew signal tristate
flabel metal2 s 3696 9600 3752 10000 0 FreeSans 224 90 0 0 o_wb_data[17]
port 53 nsew signal tristate
flabel metal3 s 0 7392 400 7448 0 FreeSans 224 0 0 0 o_wb_data[18]
port 54 nsew signal tristate
flabel metal2 s 3024 0 3080 400 0 FreeSans 224 90 0 0 o_wb_data[19]
port 55 nsew signal tristate
flabel metal3 s 9600 6048 10000 6104 0 FreeSans 224 0 0 0 o_wb_data[1]
port 56 nsew signal tristate
flabel metal3 s 9600 3024 10000 3080 0 FreeSans 224 0 0 0 o_wb_data[20]
port 57 nsew signal tristate
flabel metal2 s 2352 0 2408 400 0 FreeSans 224 90 0 0 o_wb_data[21]
port 58 nsew signal tristate
flabel metal3 s 9600 7728 10000 7784 0 FreeSans 224 0 0 0 o_wb_data[22]
port 59 nsew signal tristate
flabel metal2 s 7392 9600 7448 10000 0 FreeSans 224 90 0 0 o_wb_data[23]
port 60 nsew signal tristate
flabel metal3 s 0 7728 400 7784 0 FreeSans 224 0 0 0 o_wb_data[24]
port 61 nsew signal tristate
flabel metal2 s 3360 9600 3416 10000 0 FreeSans 224 90 0 0 o_wb_data[25]
port 62 nsew signal tristate
flabel metal3 s 9600 7392 10000 7448 0 FreeSans 224 0 0 0 o_wb_data[26]
port 63 nsew signal tristate
flabel metal3 s 0 1344 400 1400 0 FreeSans 224 0 0 0 o_wb_data[27]
port 64 nsew signal tristate
flabel metal2 s 5712 0 5768 400 0 FreeSans 224 90 0 0 o_wb_data[28]
port 65 nsew signal tristate
flabel metal3 s 0 1680 400 1736 0 FreeSans 224 0 0 0 o_wb_data[29]
port 66 nsew signal tristate
flabel metal2 s 2688 0 2744 400 0 FreeSans 224 90 0 0 o_wb_data[2]
port 67 nsew signal tristate
flabel metal3 s 9600 7056 10000 7112 0 FreeSans 224 0 0 0 o_wb_data[30]
port 68 nsew signal tristate
flabel metal3 s 0 2016 400 2072 0 FreeSans 224 0 0 0 o_wb_data[31]
port 69 nsew signal tristate
flabel metal2 s 5376 9600 5432 10000 0 FreeSans 224 90 0 0 o_wb_data[3]
port 70 nsew signal tristate
flabel metal2 s 6720 9600 6776 10000 0 FreeSans 224 90 0 0 o_wb_data[4]
port 71 nsew signal tristate
flabel metal2 s 7056 9600 7112 10000 0 FreeSans 224 90 0 0 o_wb_data[5]
port 72 nsew signal tristate
flabel metal3 s 0 5712 400 5768 0 FreeSans 224 0 0 0 o_wb_data[6]
port 73 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 o_wb_data[7]
port 74 nsew signal tristate
flabel metal3 s 0 7056 400 7112 0 FreeSans 224 0 0 0 o_wb_data[8]
port 75 nsew signal tristate
flabel metal2 s 5712 9600 5768 10000 0 FreeSans 224 90 0 0 o_wb_data[9]
port 76 nsew signal tristate
flabel metal2 s 4368 9600 4424 10000 0 FreeSans 224 90 0 0 o_wb_stall
port 77 nsew signal tristate
flabel metal3 s 9600 5040 10000 5096 0 FreeSans 224 0 0 0 reset
port 78 nsew signal input
rlabel metal1 4984 8232 4984 8232 0 VDD
rlabel via1 5024 7840 5024 7840 0 VSS
rlabel metal2 6916 4186 6916 4186 0 _000_
rlabel metal2 5404 6300 5404 6300 0 _001_
rlabel metal2 7252 5964 7252 5964 0 _002_
rlabel metal2 3500 6300 3500 6300 0 _003_
rlabel metal2 3332 5012 3332 5012 0 _004_
rlabel metal3 3248 4900 3248 4900 0 _005_
rlabel metal2 3556 6412 3556 6412 0 _006_
rlabel metal3 4088 4508 4088 4508 0 _007_
rlabel metal2 4116 5516 4116 5516 0 _008_
rlabel metal2 3556 1904 3556 1904 0 _009_
rlabel metal2 3612 1932 3612 1932 0 _010_
rlabel metal2 4172 2044 4172 2044 0 _011_
rlabel metal2 5516 4648 5516 4648 0 _012_
rlabel metal2 5572 3780 5572 3780 0 _013_
rlabel metal2 5628 3416 5628 3416 0 _014_
rlabel metal2 5320 4116 5320 4116 0 _015_
rlabel metal2 2268 4368 2268 4368 0 _016_
rlabel metal2 2548 4018 2548 4018 0 _017_
rlabel metal2 4340 2772 4340 2772 0 _018_
rlabel metal2 4032 4676 4032 4676 0 _019_
rlabel metal2 4116 2184 4116 2184 0 _020_
rlabel metal2 4032 4396 4032 4396 0 _021_
rlabel metal2 4340 4648 4340 4648 0 _022_
rlabel metal2 4508 3948 4508 3948 0 _023_
rlabel metal3 5180 4396 5180 4396 0 _024_
rlabel metal3 5656 4452 5656 4452 0 _025_
rlabel metal2 6748 4508 6748 4508 0 _026_
rlabel metal2 7028 4158 7028 4158 0 _027_
rlabel metal3 7196 5684 7196 5684 0 _028_
rlabel metal3 6216 6076 6216 6076 0 _029_
rlabel metal3 5124 6076 5124 6076 0 _030_
rlabel metal2 4060 2184 4060 2184 0 _031_
rlabel metal3 6216 5740 6216 5740 0 _032_
rlabel metal2 7308 5628 7308 5628 0 _033_
rlabel metal2 4564 5488 4564 5488 0 _034_
rlabel metal2 7588 5684 7588 5684 0 _035_
rlabel metal2 6020 2576 6020 2576 0 _036_
rlabel metal2 3780 4508 3780 4508 0 _037_
rlabel metal2 3724 6160 3724 6160 0 _038_
rlabel metal2 3696 4900 3696 4900 0 _039_
rlabel metal2 9100 5908 9100 5908 0 buttons[0]
rlabel metal2 9100 4816 9100 4816 0 buttons[1]
rlabel metal2 5124 5656 5124 5656 0 clk
rlabel metal2 5796 5516 5796 5516 0 clknet_0_clk
rlabel metal3 3276 5740 3276 5740 0 clknet_1_0__leaf_clk
rlabel metal2 7028 5460 7028 5460 0 clknet_1_1__leaf_clk
rlabel metal2 1204 2044 1204 2044 0 i_wb_addr[0]
rlabel metal2 1540 2016 1540 2016 0 i_wb_addr[10]
rlabel metal2 9100 2184 9100 2184 0 i_wb_addr[11]
rlabel metal3 8736 2156 8736 2156 0 i_wb_addr[12]
rlabel metal2 5628 1652 5628 1652 0 i_wb_addr[13]
rlabel metal3 5180 1764 5180 1764 0 i_wb_addr[14]
rlabel metal2 8932 1652 8932 1652 0 i_wb_addr[15]
rlabel metal2 8988 1792 8988 1792 0 i_wb_addr[16]
rlabel metal2 7756 1239 7756 1239 0 i_wb_addr[17]
rlabel metal2 7364 1512 7364 1512 0 i_wb_addr[18]
rlabel metal3 6720 1764 6720 1764 0 i_wb_addr[19]
rlabel metal2 1484 2016 1484 2016 0 i_wb_addr[1]
rlabel metal3 7840 1764 7840 1764 0 i_wb_addr[20]
rlabel metal2 7700 1736 7700 1736 0 i_wb_addr[21]
rlabel metal2 8596 1736 8596 1736 0 i_wb_addr[22]
rlabel metal2 6692 1736 6692 1736 0 i_wb_addr[23]
rlabel metal2 868 4452 868 4452 0 i_wb_addr[24]
rlabel metal3 623 4060 623 4060 0 i_wb_addr[25]
rlabel metal2 924 2520 924 2520 0 i_wb_addr[26]
rlabel metal2 868 4788 868 4788 0 i_wb_addr[27]
rlabel metal2 868 2828 868 2828 0 i_wb_addr[28]
rlabel metal2 1204 3920 1204 3920 0 i_wb_addr[29]
rlabel metal2 1820 1456 1820 1456 0 i_wb_addr[2]
rlabel metal2 868 3556 868 3556 0 i_wb_addr[30]
rlabel metal2 868 3164 868 3164 0 i_wb_addr[31]
rlabel metal3 2884 1764 2884 1764 0 i_wb_addr[3]
rlabel metal2 840 2156 840 2156 0 i_wb_addr[4]
rlabel metal2 3780 2100 3780 2100 0 i_wb_addr[5]
rlabel metal2 1120 1708 1120 1708 0 i_wb_addr[6]
rlabel metal2 3668 2548 3668 2548 0 i_wb_addr[7]
rlabel metal2 4816 1764 4816 1764 0 i_wb_addr[8]
rlabel metal2 5292 1624 5292 1624 0 i_wb_addr[9]
rlabel metal3 9261 3724 9261 3724 0 i_wb_cyc
rlabel metal3 623 6412 623 6412 0 i_wb_data[0]
rlabel metal2 868 5180 868 5180 0 i_wb_data[1]
rlabel metal3 9373 4060 9373 4060 0 i_wb_stb
rlabel metal2 9100 4452 9100 4452 0 i_wb_we
rlabel metal2 4060 8897 4060 8897 0 leds[0]
rlabel metal3 707 5404 707 5404 0 leds[1]
rlabel metal2 7140 4536 7140 4536 0 net1
rlabel metal2 7756 2716 7756 2716 0 net10
rlabel metal2 7420 2632 7420 2632 0 net11
rlabel metal2 7252 1988 7252 1988 0 net12
rlabel metal2 6692 2632 6692 2632 0 net13
rlabel metal2 3416 3276 3416 3276 0 net14
rlabel metal2 7812 3192 7812 3192 0 net15
rlabel metal2 7588 2212 7588 2212 0 net16
rlabel metal2 8484 2744 8484 2744 0 net17
rlabel metal2 6580 2716 6580 2716 0 net18
rlabel metal3 1904 3836 1904 3836 0 net19
rlabel metal2 8932 4984 8932 4984 0 net2
rlabel metal3 2072 4004 2072 4004 0 net20
rlabel metal2 1036 2688 1036 2688 0 net21
rlabel metal3 1456 3724 1456 3724 0 net22
rlabel metal3 2016 2996 2016 2996 0 net23
rlabel metal3 2156 4564 2156 4564 0 net24
rlabel metal2 1988 2072 1988 2072 0 net25
rlabel metal2 1036 3864 1036 3864 0 net26
rlabel metal2 1036 3444 1036 3444 0 net27
rlabel metal2 2324 2492 2324 2492 0 net28
rlabel metal2 1008 2268 1008 2268 0 net29
rlabel metal2 3332 3220 3332 3220 0 net3
rlabel metal2 3948 2576 3948 2576 0 net30
rlabel metal2 1316 2268 1316 2268 0 net31
rlabel metal2 3444 2716 3444 2716 0 net32
rlabel metal2 5012 1932 5012 1932 0 net33
rlabel metal2 5180 1960 5180 1960 0 net34
rlabel metal3 7868 4060 7868 4060 0 net35
rlabel metal2 1036 6496 1036 6496 0 net36
rlabel metal3 2044 4956 2044 4956 0 net37
rlabel metal2 7196 4032 7196 4032 0 net38
rlabel metal3 8148 4508 8148 4508 0 net39
rlabel metal3 2954 2268 2954 2268 0 net4
rlabel metal3 8428 5348 8428 5348 0 net40
rlabel metal2 4004 6356 4004 6356 0 net41
rlabel metal2 2660 5460 2660 5460 0 net42
rlabel metal2 8484 5320 8484 5320 0 net43
rlabel metal3 7476 6524 7476 6524 0 net44
rlabel metal3 7336 6468 7336 6468 0 net45
rlabel metal2 2716 427 2716 427 0 net46
rlabel metal2 5460 7980 5460 7980 0 net47
rlabel metal2 6804 7980 6804 7980 0 net48
rlabel metal2 7140 7980 7140 7980 0 net49
rlabel metal2 6692 2128 6692 2128 0 net5
rlabel metal3 623 5740 623 5740 0 net50
rlabel metal2 1092 8036 1092 8036 0 net51
rlabel metal3 623 7084 623 7084 0 net52
rlabel metal2 5796 7980 5796 7980 0 net53
rlabel metal2 2044 1407 2044 1407 0 net54
rlabel metal3 791 6076 791 6076 0 net55
rlabel metal3 903 1036 903 1036 0 net56
rlabel metal2 8764 2240 8764 2240 0 net57
rlabel metal2 4788 7756 4788 7756 0 net58
rlabel metal2 1316 8176 1316 8176 0 net59
rlabel metal3 8260 2184 8260 2184 0 net6
rlabel metal2 3108 7980 3108 7980 0 net60
rlabel metal2 3780 7980 3780 7980 0 net61
rlabel metal3 623 7420 623 7420 0 net62
rlabel metal2 3052 1407 3052 1407 0 net63
rlabel metal2 9100 3136 9100 3136 0 net64
rlabel metal2 2380 427 2380 427 0 net65
rlabel metal2 9128 7924 9128 7924 0 net66
rlabel metal2 7476 7980 7476 7980 0 net67
rlabel metal3 427 7756 427 7756 0 net68
rlabel metal2 3444 7980 3444 7980 0 net69
rlabel metal2 3220 1960 3220 1960 0 net7
rlabel metal2 9100 7560 9100 7560 0 net70
rlabel metal3 1071 1372 1071 1372 0 net71
rlabel metal2 5740 1015 5740 1015 0 net72
rlabel metal3 763 1708 763 1708 0 net73
rlabel metal3 9268 7140 9268 7140 0 net74
rlabel metal2 868 1848 868 1848 0 net75
rlabel metal2 4396 8813 4396 8813 0 net76
rlabel metal2 4452 2100 4452 2100 0 net8
rlabel metal2 4508 2016 4508 2016 0 net9
rlabel metal3 9345 5404 9345 5404 0 o_wb_ack
rlabel metal3 9345 6412 9345 6412 0 o_wb_data[0]
rlabel metal2 8204 6300 8204 6300 0 o_wb_data[1]
rlabel metal2 9100 5180 9100 5180 0 reset
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>
