magic
tech gf180mcuD
magscale 1 5
timestamp 1700745744
<< obsm1 >>
rect 672 1538 254296 173294
<< metal2 >>
rect 127344 174600 127400 175000
rect 127008 0 127064 400
rect 127344 0 127400 400
<< obsm2 >>
rect 2238 174570 127314 174600
rect 127430 174570 248130 174600
rect 2238 430 248130 174570
rect 2238 400 126978 430
rect 127094 400 127314 430
rect 127430 400 248130 430
<< obsm3 >>
rect 2233 1554 248135 173278
<< metal4 >>
rect 2224 1538 2384 173294
rect 9904 1538 10064 173294
rect 17584 1538 17744 173294
rect 25264 1538 25424 173294
rect 32944 1538 33104 173294
rect 40624 1538 40784 173294
rect 48304 1538 48464 173294
rect 55984 1538 56144 173294
rect 63664 1538 63824 173294
rect 71344 1538 71504 173294
rect 79024 1538 79184 173294
rect 86704 1538 86864 173294
rect 94384 1538 94544 173294
rect 102064 1538 102224 173294
rect 109744 1538 109904 173294
rect 117424 1538 117584 173294
rect 125104 1538 125264 173294
rect 132784 1538 132944 173294
rect 140464 1538 140624 173294
rect 148144 1538 148304 173294
rect 155824 1538 155984 173294
rect 163504 1538 163664 173294
rect 171184 1538 171344 173294
rect 178864 1538 179024 173294
rect 186544 1538 186704 173294
rect 194224 1538 194384 173294
rect 201904 1538 202064 173294
rect 209584 1538 209744 173294
rect 217264 1538 217424 173294
rect 224944 1538 225104 173294
rect 232624 1538 232784 173294
rect 240304 1538 240464 173294
rect 247984 1538 248144 173294
<< labels >>
rlabel metal2 s 127344 0 127400 400 6 in1
port 1 nsew signal input
rlabel metal2 s 127008 0 127064 400 6 in2
port 2 nsew signal input
rlabel metal2 s 127344 174600 127400 175000 6 out
port 3 nsew signal output
rlabel metal4 s 2224 1538 2384 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 173294 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 173294 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 173294 6 vss
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 255000 175000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5138800
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/analog_wrapper/runs/23_11_23_15_21/results/signoff/analog_wrapper.magic.gds
string GDS_START 3112
<< end >>

