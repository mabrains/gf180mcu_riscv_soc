magic
tech gf180mcuD
magscale 1 10
timestamp 1700703346
<< metal1 >>
rect 1344 96458 38640 96492
rect 1344 96406 4024 96458
rect 4076 96406 4148 96458
rect 4200 96406 4272 96458
rect 4324 96406 4396 96458
rect 4448 96406 4520 96458
rect 4572 96406 4644 96458
rect 4696 96406 4768 96458
rect 4820 96406 4892 96458
rect 4944 96406 5016 96458
rect 5068 96406 5140 96458
rect 5192 96406 24024 96458
rect 24076 96406 24148 96458
rect 24200 96406 24272 96458
rect 24324 96406 24396 96458
rect 24448 96406 24520 96458
rect 24572 96406 24644 96458
rect 24696 96406 24768 96458
rect 24820 96406 24892 96458
rect 24944 96406 25016 96458
rect 25068 96406 25140 96458
rect 25192 96406 38640 96458
rect 1344 96372 38640 96406
rect 30258 96014 30270 96066
rect 30322 96014 30334 96066
rect 30046 95954 30098 95966
rect 30046 95890 30098 95902
rect 1710 95842 1762 95854
rect 1710 95778 1762 95790
rect 29822 95842 29874 95854
rect 29822 95778 29874 95790
rect 1344 95674 38640 95708
rect 1344 95622 14024 95674
rect 14076 95622 14148 95674
rect 14200 95622 14272 95674
rect 14324 95622 14396 95674
rect 14448 95622 14520 95674
rect 14572 95622 14644 95674
rect 14696 95622 14768 95674
rect 14820 95622 14892 95674
rect 14944 95622 15016 95674
rect 15068 95622 15140 95674
rect 15192 95622 34024 95674
rect 34076 95622 34148 95674
rect 34200 95622 34272 95674
rect 34324 95622 34396 95674
rect 34448 95622 34520 95674
rect 34572 95622 34644 95674
rect 34696 95622 34768 95674
rect 34820 95622 34892 95674
rect 34944 95622 35016 95674
rect 35068 95622 35140 95674
rect 35192 95622 38640 95674
rect 1344 95588 38640 95622
rect 1344 94890 38640 94924
rect 1344 94838 4024 94890
rect 4076 94838 4148 94890
rect 4200 94838 4272 94890
rect 4324 94838 4396 94890
rect 4448 94838 4520 94890
rect 4572 94838 4644 94890
rect 4696 94838 4768 94890
rect 4820 94838 4892 94890
rect 4944 94838 5016 94890
rect 5068 94838 5140 94890
rect 5192 94838 24024 94890
rect 24076 94838 24148 94890
rect 24200 94838 24272 94890
rect 24324 94838 24396 94890
rect 24448 94838 24520 94890
rect 24572 94838 24644 94890
rect 24696 94838 24768 94890
rect 24820 94838 24892 94890
rect 24944 94838 25016 94890
rect 25068 94838 25140 94890
rect 25192 94838 38640 94890
rect 1344 94804 38640 94838
rect 1710 94274 1762 94286
rect 1710 94210 1762 94222
rect 1344 94106 38640 94140
rect 1344 94054 14024 94106
rect 14076 94054 14148 94106
rect 14200 94054 14272 94106
rect 14324 94054 14396 94106
rect 14448 94054 14520 94106
rect 14572 94054 14644 94106
rect 14696 94054 14768 94106
rect 14820 94054 14892 94106
rect 14944 94054 15016 94106
rect 15068 94054 15140 94106
rect 15192 94054 34024 94106
rect 34076 94054 34148 94106
rect 34200 94054 34272 94106
rect 34324 94054 34396 94106
rect 34448 94054 34520 94106
rect 34572 94054 34644 94106
rect 34696 94054 34768 94106
rect 34820 94054 34892 94106
rect 34944 94054 35016 94106
rect 35068 94054 35140 94106
rect 35192 94054 38640 94106
rect 1344 94020 38640 94054
rect 1710 93826 1762 93838
rect 1710 93762 1762 93774
rect 1344 93322 38640 93356
rect 1344 93270 4024 93322
rect 4076 93270 4148 93322
rect 4200 93270 4272 93322
rect 4324 93270 4396 93322
rect 4448 93270 4520 93322
rect 4572 93270 4644 93322
rect 4696 93270 4768 93322
rect 4820 93270 4892 93322
rect 4944 93270 5016 93322
rect 5068 93270 5140 93322
rect 5192 93270 24024 93322
rect 24076 93270 24148 93322
rect 24200 93270 24272 93322
rect 24324 93270 24396 93322
rect 24448 93270 24520 93322
rect 24572 93270 24644 93322
rect 24696 93270 24768 93322
rect 24820 93270 24892 93322
rect 24944 93270 25016 93322
rect 25068 93270 25140 93322
rect 25192 93270 38640 93322
rect 1344 93236 38640 93270
rect 1344 92538 38640 92572
rect 1344 92486 14024 92538
rect 14076 92486 14148 92538
rect 14200 92486 14272 92538
rect 14324 92486 14396 92538
rect 14448 92486 14520 92538
rect 14572 92486 14644 92538
rect 14696 92486 14768 92538
rect 14820 92486 14892 92538
rect 14944 92486 15016 92538
rect 15068 92486 15140 92538
rect 15192 92486 34024 92538
rect 34076 92486 34148 92538
rect 34200 92486 34272 92538
rect 34324 92486 34396 92538
rect 34448 92486 34520 92538
rect 34572 92486 34644 92538
rect 34696 92486 34768 92538
rect 34820 92486 34892 92538
rect 34944 92486 35016 92538
rect 35068 92486 35140 92538
rect 35192 92486 38640 92538
rect 1344 92452 38640 92486
rect 1710 92258 1762 92270
rect 1710 92194 1762 92206
rect 1344 91754 38640 91788
rect 1344 91702 4024 91754
rect 4076 91702 4148 91754
rect 4200 91702 4272 91754
rect 4324 91702 4396 91754
rect 4448 91702 4520 91754
rect 4572 91702 4644 91754
rect 4696 91702 4768 91754
rect 4820 91702 4892 91754
rect 4944 91702 5016 91754
rect 5068 91702 5140 91754
rect 5192 91702 24024 91754
rect 24076 91702 24148 91754
rect 24200 91702 24272 91754
rect 24324 91702 24396 91754
rect 24448 91702 24520 91754
rect 24572 91702 24644 91754
rect 24696 91702 24768 91754
rect 24820 91702 24892 91754
rect 24944 91702 25016 91754
rect 25068 91702 25140 91754
rect 25192 91702 38640 91754
rect 1344 91668 38640 91702
rect 1710 91138 1762 91150
rect 1710 91074 1762 91086
rect 1344 90970 38640 91004
rect 1344 90918 14024 90970
rect 14076 90918 14148 90970
rect 14200 90918 14272 90970
rect 14324 90918 14396 90970
rect 14448 90918 14520 90970
rect 14572 90918 14644 90970
rect 14696 90918 14768 90970
rect 14820 90918 14892 90970
rect 14944 90918 15016 90970
rect 15068 90918 15140 90970
rect 15192 90918 34024 90970
rect 34076 90918 34148 90970
rect 34200 90918 34272 90970
rect 34324 90918 34396 90970
rect 34448 90918 34520 90970
rect 34572 90918 34644 90970
rect 34696 90918 34768 90970
rect 34820 90918 34892 90970
rect 34944 90918 35016 90970
rect 35068 90918 35140 90970
rect 35192 90918 38640 90970
rect 1344 90884 38640 90918
rect 1344 90186 38640 90220
rect 1344 90134 4024 90186
rect 4076 90134 4148 90186
rect 4200 90134 4272 90186
rect 4324 90134 4396 90186
rect 4448 90134 4520 90186
rect 4572 90134 4644 90186
rect 4696 90134 4768 90186
rect 4820 90134 4892 90186
rect 4944 90134 5016 90186
rect 5068 90134 5140 90186
rect 5192 90134 24024 90186
rect 24076 90134 24148 90186
rect 24200 90134 24272 90186
rect 24324 90134 24396 90186
rect 24448 90134 24520 90186
rect 24572 90134 24644 90186
rect 24696 90134 24768 90186
rect 24820 90134 24892 90186
rect 24944 90134 25016 90186
rect 25068 90134 25140 90186
rect 25192 90134 38640 90186
rect 1344 90100 38640 90134
rect 1710 89682 1762 89694
rect 1710 89618 1762 89630
rect 13694 89570 13746 89582
rect 13694 89506 13746 89518
rect 1344 89402 38640 89436
rect 1344 89350 14024 89402
rect 14076 89350 14148 89402
rect 14200 89350 14272 89402
rect 14324 89350 14396 89402
rect 14448 89350 14520 89402
rect 14572 89350 14644 89402
rect 14696 89350 14768 89402
rect 14820 89350 14892 89402
rect 14944 89350 15016 89402
rect 15068 89350 15140 89402
rect 15192 89350 34024 89402
rect 34076 89350 34148 89402
rect 34200 89350 34272 89402
rect 34324 89350 34396 89402
rect 34448 89350 34520 89402
rect 34572 89350 34644 89402
rect 34696 89350 34768 89402
rect 34820 89350 34892 89402
rect 34944 89350 35016 89402
rect 35068 89350 35140 89402
rect 35192 89350 38640 89402
rect 1344 89316 38640 89350
rect 1710 89122 1762 89134
rect 1710 89058 1762 89070
rect 12350 89122 12402 89134
rect 12350 89058 12402 89070
rect 9438 89010 9490 89022
rect 9986 88958 9998 89010
rect 10050 88958 10062 89010
rect 9438 88946 9490 88958
rect 8542 88898 8594 88910
rect 8542 88834 8594 88846
rect 8990 88898 9042 88910
rect 8990 88834 9042 88846
rect 13582 88898 13634 88910
rect 13582 88834 13634 88846
rect 13918 88898 13970 88910
rect 13918 88834 13970 88846
rect 13134 88786 13186 88798
rect 13134 88722 13186 88734
rect 1344 88618 38640 88652
rect 1344 88566 4024 88618
rect 4076 88566 4148 88618
rect 4200 88566 4272 88618
rect 4324 88566 4396 88618
rect 4448 88566 4520 88618
rect 4572 88566 4644 88618
rect 4696 88566 4768 88618
rect 4820 88566 4892 88618
rect 4944 88566 5016 88618
rect 5068 88566 5140 88618
rect 5192 88566 24024 88618
rect 24076 88566 24148 88618
rect 24200 88566 24272 88618
rect 24324 88566 24396 88618
rect 24448 88566 24520 88618
rect 24572 88566 24644 88618
rect 24696 88566 24768 88618
rect 24820 88566 24892 88618
rect 24944 88566 25016 88618
rect 25068 88566 25140 88618
rect 25192 88566 38640 88618
rect 1344 88532 38640 88566
rect 9102 88226 9154 88238
rect 13918 88226 13970 88238
rect 9762 88174 9774 88226
rect 9826 88174 9838 88226
rect 9102 88162 9154 88174
rect 13918 88162 13970 88174
rect 14130 88062 14142 88114
rect 14194 88062 14206 88114
rect 14690 88062 14702 88114
rect 14754 88062 14766 88114
rect 1710 88002 1762 88014
rect 1710 87938 1762 87950
rect 8430 88002 8482 88014
rect 8430 87938 8482 87950
rect 8878 88002 8930 88014
rect 12798 88002 12850 88014
rect 12002 87950 12014 88002
rect 12066 87950 12078 88002
rect 8878 87938 8930 87950
rect 12798 87938 12850 87950
rect 13582 88002 13634 88014
rect 13582 87938 13634 87950
rect 1344 87834 38640 87868
rect 1344 87782 14024 87834
rect 14076 87782 14148 87834
rect 14200 87782 14272 87834
rect 14324 87782 14396 87834
rect 14448 87782 14520 87834
rect 14572 87782 14644 87834
rect 14696 87782 14768 87834
rect 14820 87782 14892 87834
rect 14944 87782 15016 87834
rect 15068 87782 15140 87834
rect 15192 87782 34024 87834
rect 34076 87782 34148 87834
rect 34200 87782 34272 87834
rect 34324 87782 34396 87834
rect 34448 87782 34520 87834
rect 34572 87782 34644 87834
rect 34696 87782 34768 87834
rect 34820 87782 34892 87834
rect 34944 87782 35016 87834
rect 35068 87782 35140 87834
rect 35192 87782 38640 87834
rect 1344 87748 38640 87782
rect 9886 87666 9938 87678
rect 8418 87614 8430 87666
rect 8482 87614 8494 87666
rect 9886 87602 9938 87614
rect 10334 87666 10386 87678
rect 16382 87666 16434 87678
rect 15026 87614 15038 87666
rect 15090 87614 15102 87666
rect 20402 87614 20414 87666
rect 20466 87614 20478 87666
rect 10334 87602 10386 87614
rect 16382 87602 16434 87614
rect 10882 87502 10894 87554
rect 10946 87502 10958 87554
rect 11442 87502 11454 87554
rect 11506 87502 11518 87554
rect 5630 87442 5682 87454
rect 9102 87442 9154 87454
rect 6066 87390 6078 87442
rect 6130 87390 6142 87442
rect 5630 87378 5682 87390
rect 9102 87378 9154 87390
rect 12126 87442 12178 87454
rect 20974 87442 21026 87454
rect 12562 87390 12574 87442
rect 12626 87390 12638 87442
rect 17378 87390 17390 87442
rect 17442 87390 17454 87442
rect 17938 87390 17950 87442
rect 18002 87390 18014 87442
rect 12126 87378 12178 87390
rect 20974 87378 21026 87390
rect 21310 87442 21362 87454
rect 21310 87378 21362 87390
rect 16046 87330 16098 87342
rect 16046 87266 16098 87278
rect 16942 87330 16994 87342
rect 16942 87266 16994 87278
rect 10670 87218 10722 87230
rect 10670 87154 10722 87166
rect 15598 87218 15650 87230
rect 16034 87166 16046 87218
rect 16098 87215 16110 87218
rect 16930 87215 16942 87218
rect 16098 87169 16942 87215
rect 16098 87166 16110 87169
rect 16930 87166 16942 87169
rect 16994 87166 17006 87218
rect 15598 87154 15650 87166
rect 1344 87050 38640 87084
rect 1344 86998 4024 87050
rect 4076 86998 4148 87050
rect 4200 86998 4272 87050
rect 4324 86998 4396 87050
rect 4448 86998 4520 87050
rect 4572 86998 4644 87050
rect 4696 86998 4768 87050
rect 4820 86998 4892 87050
rect 4944 86998 5016 87050
rect 5068 86998 5140 87050
rect 5192 86998 24024 87050
rect 24076 86998 24148 87050
rect 24200 86998 24272 87050
rect 24324 86998 24396 87050
rect 24448 86998 24520 87050
rect 24572 86998 24644 87050
rect 24696 86998 24768 87050
rect 24820 86998 24892 87050
rect 24944 86998 25016 87050
rect 25068 86998 25140 87050
rect 25192 86998 38640 87050
rect 1344 86964 38640 86998
rect 7646 86882 7698 86894
rect 18398 86882 18450 86894
rect 12226 86830 12238 86882
rect 12290 86879 12302 86882
rect 13010 86879 13022 86882
rect 12290 86833 13022 86879
rect 12290 86830 12302 86833
rect 13010 86830 13022 86833
rect 13074 86830 13086 86882
rect 7646 86818 7698 86830
rect 18398 86818 18450 86830
rect 9998 86770 10050 86782
rect 9998 86706 10050 86718
rect 12014 86770 12066 86782
rect 12014 86706 12066 86718
rect 12910 86770 12962 86782
rect 12910 86706 12962 86718
rect 7982 86658 8034 86670
rect 9326 86658 9378 86670
rect 8754 86606 8766 86658
rect 8818 86606 8830 86658
rect 7982 86594 8034 86606
rect 9326 86594 9378 86606
rect 9886 86658 9938 86670
rect 9886 86594 9938 86606
rect 10334 86658 10386 86670
rect 10334 86594 10386 86606
rect 10894 86658 10946 86670
rect 10894 86594 10946 86606
rect 12462 86658 12514 86670
rect 14366 86658 14418 86670
rect 18734 86658 18786 86670
rect 13570 86606 13582 86658
rect 13634 86606 13646 86658
rect 15026 86606 15038 86658
rect 15090 86606 15102 86658
rect 12462 86594 12514 86606
rect 14366 86594 14418 86606
rect 18734 86594 18786 86606
rect 7310 86546 7362 86558
rect 10222 86546 10274 86558
rect 8530 86494 8542 86546
rect 8594 86494 8606 86546
rect 7310 86482 7362 86494
rect 10222 86482 10274 86494
rect 11902 86546 11954 86558
rect 11902 86482 11954 86494
rect 14030 86546 14082 86558
rect 18946 86494 18958 86546
rect 19010 86494 19022 86546
rect 19394 86494 19406 86546
rect 19458 86494 19470 86546
rect 14030 86482 14082 86494
rect 1710 86434 1762 86446
rect 18062 86434 18114 86446
rect 17266 86382 17278 86434
rect 17330 86382 17342 86434
rect 1710 86370 1762 86382
rect 18062 86370 18114 86382
rect 1344 86266 38640 86300
rect 1344 86214 14024 86266
rect 14076 86214 14148 86266
rect 14200 86214 14272 86266
rect 14324 86214 14396 86266
rect 14448 86214 14520 86266
rect 14572 86214 14644 86266
rect 14696 86214 14768 86266
rect 14820 86214 14892 86266
rect 14944 86214 15016 86266
rect 15068 86214 15140 86266
rect 15192 86214 34024 86266
rect 34076 86214 34148 86266
rect 34200 86214 34272 86266
rect 34324 86214 34396 86266
rect 34448 86214 34520 86266
rect 34572 86214 34644 86266
rect 34696 86214 34768 86266
rect 34820 86214 34892 86266
rect 34944 86214 35016 86266
rect 35068 86214 35140 86266
rect 35192 86214 38640 86266
rect 1344 86180 38640 86214
rect 9662 86098 9714 86110
rect 9662 86034 9714 86046
rect 10222 86098 10274 86110
rect 10222 86034 10274 86046
rect 10782 86098 10834 86110
rect 10782 86034 10834 86046
rect 13582 86098 13634 86110
rect 13582 86034 13634 86046
rect 15374 86098 15426 86110
rect 23090 86046 23102 86098
rect 23154 86046 23166 86098
rect 15374 86034 15426 86046
rect 1710 85986 1762 85998
rect 1710 85922 1762 85934
rect 9998 85986 10050 85998
rect 9998 85922 10050 85934
rect 15710 85986 15762 85998
rect 15710 85922 15762 85934
rect 16606 85986 16658 85998
rect 16606 85922 16658 85934
rect 14142 85874 14194 85886
rect 14142 85810 14194 85822
rect 15038 85874 15090 85886
rect 15038 85810 15090 85822
rect 15374 85874 15426 85886
rect 24558 85874 24610 85886
rect 20066 85822 20078 85874
rect 20130 85822 20142 85874
rect 20626 85822 20638 85874
rect 20690 85822 20702 85874
rect 15374 85810 15426 85822
rect 24558 85810 24610 85822
rect 7422 85762 7474 85774
rect 14814 85762 14866 85774
rect 10322 85710 10334 85762
rect 10386 85710 10398 85762
rect 7422 85698 7474 85710
rect 14814 85698 14866 85710
rect 16158 85762 16210 85774
rect 16830 85762 16882 85774
rect 16482 85710 16494 85762
rect 16546 85710 16558 85762
rect 16158 85698 16210 85710
rect 16830 85698 16882 85710
rect 18174 85762 18226 85774
rect 18174 85698 18226 85710
rect 18622 85762 18674 85774
rect 18622 85698 18674 85710
rect 23662 85762 23714 85774
rect 23662 85698 23714 85710
rect 23998 85762 24050 85774
rect 23998 85698 24050 85710
rect 1344 85482 38640 85516
rect 1344 85430 4024 85482
rect 4076 85430 4148 85482
rect 4200 85430 4272 85482
rect 4324 85430 4396 85482
rect 4448 85430 4520 85482
rect 4572 85430 4644 85482
rect 4696 85430 4768 85482
rect 4820 85430 4892 85482
rect 4944 85430 5016 85482
rect 5068 85430 5140 85482
rect 5192 85430 24024 85482
rect 24076 85430 24148 85482
rect 24200 85430 24272 85482
rect 24324 85430 24396 85482
rect 24448 85430 24520 85482
rect 24572 85430 24644 85482
rect 24696 85430 24768 85482
rect 24820 85430 24892 85482
rect 24944 85430 25016 85482
rect 25068 85430 25140 85482
rect 25192 85430 38640 85482
rect 1344 85396 38640 85430
rect 21422 85314 21474 85326
rect 21422 85250 21474 85262
rect 4846 85202 4898 85214
rect 4846 85138 4898 85150
rect 14366 85202 14418 85214
rect 14366 85138 14418 85150
rect 6526 85090 6578 85102
rect 10782 85090 10834 85102
rect 6962 85038 6974 85090
rect 7026 85038 7038 85090
rect 6526 85026 6578 85038
rect 10782 85026 10834 85038
rect 14254 85090 14306 85102
rect 14254 85026 14306 85038
rect 21758 85090 21810 85102
rect 21758 85026 21810 85038
rect 9214 84978 9266 84990
rect 9214 84914 9266 84926
rect 13918 84978 13970 84990
rect 13918 84914 13970 84926
rect 14478 84978 14530 84990
rect 14478 84914 14530 84926
rect 20750 84978 20802 84990
rect 21970 84926 21982 84978
rect 22034 84926 22046 84978
rect 22530 84926 22542 84978
rect 22594 84926 22606 84978
rect 20750 84914 20802 84926
rect 5854 84866 5906 84878
rect 5854 84802 5906 84814
rect 9998 84866 10050 84878
rect 9998 84802 10050 84814
rect 10334 84866 10386 84878
rect 10334 84802 10386 84814
rect 12574 84866 12626 84878
rect 12574 84802 12626 84814
rect 13022 84866 13074 84878
rect 13022 84802 13074 84814
rect 13694 84866 13746 84878
rect 13694 84802 13746 84814
rect 18174 84866 18226 84878
rect 18174 84802 18226 84814
rect 1344 84698 38640 84732
rect 1344 84646 14024 84698
rect 14076 84646 14148 84698
rect 14200 84646 14272 84698
rect 14324 84646 14396 84698
rect 14448 84646 14520 84698
rect 14572 84646 14644 84698
rect 14696 84646 14768 84698
rect 14820 84646 14892 84698
rect 14944 84646 15016 84698
rect 15068 84646 15140 84698
rect 15192 84646 34024 84698
rect 34076 84646 34148 84698
rect 34200 84646 34272 84698
rect 34324 84646 34396 84698
rect 34448 84646 34520 84698
rect 34572 84646 34644 84698
rect 34696 84646 34768 84698
rect 34820 84646 34892 84698
rect 34944 84646 35016 84698
rect 35068 84646 35140 84698
rect 35192 84646 38640 84698
rect 1344 84612 38640 84646
rect 8318 84530 8370 84542
rect 6738 84478 6750 84530
rect 6802 84478 6814 84530
rect 8318 84466 8370 84478
rect 9662 84530 9714 84542
rect 9662 84466 9714 84478
rect 12238 84530 12290 84542
rect 12238 84466 12290 84478
rect 12686 84530 12738 84542
rect 12686 84466 12738 84478
rect 18734 84530 18786 84542
rect 18734 84466 18786 84478
rect 22094 84530 22146 84542
rect 22094 84466 22146 84478
rect 1710 84418 1762 84430
rect 1710 84354 1762 84366
rect 8542 84418 8594 84430
rect 8542 84354 8594 84366
rect 9774 84418 9826 84430
rect 9774 84354 9826 84366
rect 13358 84418 13410 84430
rect 13358 84354 13410 84366
rect 13582 84418 13634 84430
rect 13582 84354 13634 84366
rect 14478 84418 14530 84430
rect 14478 84354 14530 84366
rect 14590 84418 14642 84430
rect 14590 84354 14642 84366
rect 15038 84418 15090 84430
rect 19282 84366 19294 84418
rect 19346 84366 19358 84418
rect 19618 84366 19630 84418
rect 19682 84366 19694 84418
rect 21074 84366 21086 84418
rect 21138 84366 21150 84418
rect 15038 84354 15090 84366
rect 3838 84306 3890 84318
rect 8094 84306 8146 84318
rect 4162 84254 4174 84306
rect 4226 84254 4238 84306
rect 3838 84242 3890 84254
rect 8094 84242 8146 84254
rect 8766 84306 8818 84318
rect 8766 84242 8818 84254
rect 12574 84306 12626 84318
rect 12574 84242 12626 84254
rect 12798 84306 12850 84318
rect 12798 84242 12850 84254
rect 13246 84306 13298 84318
rect 13246 84242 13298 84254
rect 13694 84306 13746 84318
rect 13694 84242 13746 84254
rect 20526 84306 20578 84318
rect 20962 84254 20974 84306
rect 21026 84254 21038 84306
rect 20526 84242 20578 84254
rect 7870 84194 7922 84206
rect 7870 84130 7922 84142
rect 11790 84194 11842 84206
rect 11790 84130 11842 84142
rect 17502 84194 17554 84206
rect 17502 84130 17554 84142
rect 18286 84194 18338 84206
rect 18286 84130 18338 84142
rect 7310 84082 7362 84094
rect 7310 84018 7362 84030
rect 14478 84082 14530 84094
rect 14478 84018 14530 84030
rect 19070 84082 19122 84094
rect 19070 84018 19122 84030
rect 21758 84082 21810 84094
rect 21758 84018 21810 84030
rect 1344 83914 38640 83948
rect 1344 83862 4024 83914
rect 4076 83862 4148 83914
rect 4200 83862 4272 83914
rect 4324 83862 4396 83914
rect 4448 83862 4520 83914
rect 4572 83862 4644 83914
rect 4696 83862 4768 83914
rect 4820 83862 4892 83914
rect 4944 83862 5016 83914
rect 5068 83862 5140 83914
rect 5192 83862 24024 83914
rect 24076 83862 24148 83914
rect 24200 83862 24272 83914
rect 24324 83862 24396 83914
rect 24448 83862 24520 83914
rect 24572 83862 24644 83914
rect 24696 83862 24768 83914
rect 24820 83862 24892 83914
rect 24944 83862 25016 83914
rect 25068 83862 25140 83914
rect 25192 83862 38640 83914
rect 1344 83828 38640 83862
rect 5966 83746 6018 83758
rect 5966 83682 6018 83694
rect 6302 83746 6354 83758
rect 6302 83682 6354 83694
rect 8766 83746 8818 83758
rect 12114 83694 12126 83746
rect 12178 83694 12190 83746
rect 8766 83682 8818 83694
rect 20302 83634 20354 83646
rect 12562 83582 12574 83634
rect 12626 83582 12638 83634
rect 20302 83570 20354 83582
rect 3726 83522 3778 83534
rect 17614 83522 17666 83534
rect 4274 83470 4286 83522
rect 4338 83470 4350 83522
rect 7074 83470 7086 83522
rect 7138 83470 7150 83522
rect 8754 83470 8766 83522
rect 8818 83470 8830 83522
rect 12450 83470 12462 83522
rect 12514 83470 12526 83522
rect 13458 83470 13470 83522
rect 13522 83470 13534 83522
rect 14018 83470 14030 83522
rect 14082 83470 14094 83522
rect 3726 83458 3778 83470
rect 17614 83458 17666 83470
rect 17838 83522 17890 83534
rect 17838 83458 17890 83470
rect 18286 83522 18338 83534
rect 18286 83458 18338 83470
rect 18958 83522 19010 83534
rect 18958 83458 19010 83470
rect 19182 83522 19234 83534
rect 22990 83522 23042 83534
rect 19394 83470 19406 83522
rect 19458 83470 19470 83522
rect 19182 83458 19234 83470
rect 22990 83458 23042 83470
rect 8206 83410 8258 83422
rect 4498 83358 4510 83410
rect 4562 83358 4574 83410
rect 6850 83358 6862 83410
rect 6914 83358 6926 83410
rect 8206 83346 8258 83358
rect 8430 83410 8482 83422
rect 8430 83346 8482 83358
rect 18398 83410 18450 83422
rect 18398 83346 18450 83358
rect 18734 83410 18786 83422
rect 18734 83346 18786 83358
rect 19070 83410 19122 83422
rect 19070 83346 19122 83358
rect 1710 83298 1762 83310
rect 1710 83234 1762 83246
rect 3390 83298 3442 83310
rect 3390 83234 3442 83246
rect 5070 83298 5122 83310
rect 5070 83234 5122 83246
rect 7646 83298 7698 83310
rect 7646 83234 7698 83246
rect 9214 83298 9266 83310
rect 17054 83298 17106 83310
rect 16482 83246 16494 83298
rect 16546 83246 16558 83298
rect 9214 83234 9266 83246
rect 17054 83234 17106 83246
rect 17502 83298 17554 83310
rect 17502 83234 17554 83246
rect 22542 83298 22594 83310
rect 22542 83234 22594 83246
rect 22654 83298 22706 83310
rect 22654 83234 22706 83246
rect 22878 83298 22930 83310
rect 22878 83234 22930 83246
rect 1344 83130 38640 83164
rect 1344 83078 14024 83130
rect 14076 83078 14148 83130
rect 14200 83078 14272 83130
rect 14324 83078 14396 83130
rect 14448 83078 14520 83130
rect 14572 83078 14644 83130
rect 14696 83078 14768 83130
rect 14820 83078 14892 83130
rect 14944 83078 15016 83130
rect 15068 83078 15140 83130
rect 15192 83078 34024 83130
rect 34076 83078 34148 83130
rect 34200 83078 34272 83130
rect 34324 83078 34396 83130
rect 34448 83078 34520 83130
rect 34572 83078 34644 83130
rect 34696 83078 34768 83130
rect 34820 83078 34892 83130
rect 34944 83078 35016 83130
rect 35068 83078 35140 83130
rect 35192 83078 38640 83130
rect 1344 83044 38640 83078
rect 5294 82962 5346 82974
rect 4722 82910 4734 82962
rect 4786 82910 4798 82962
rect 5294 82898 5346 82910
rect 5630 82962 5682 82974
rect 5630 82898 5682 82910
rect 6190 82962 6242 82974
rect 6190 82898 6242 82910
rect 11118 82962 11170 82974
rect 11118 82898 11170 82910
rect 12910 82962 12962 82974
rect 12910 82898 12962 82910
rect 15934 82962 15986 82974
rect 15934 82898 15986 82910
rect 16718 82962 16770 82974
rect 16718 82898 16770 82910
rect 25342 82962 25394 82974
rect 25342 82898 25394 82910
rect 5518 82850 5570 82862
rect 5518 82786 5570 82798
rect 13022 82850 13074 82862
rect 13022 82786 13074 82798
rect 13582 82850 13634 82862
rect 13582 82786 13634 82798
rect 14366 82850 14418 82862
rect 14366 82786 14418 82798
rect 16270 82850 16322 82862
rect 16270 82786 16322 82798
rect 17390 82850 17442 82862
rect 17390 82786 17442 82798
rect 21870 82850 21922 82862
rect 21870 82786 21922 82798
rect 1822 82738 1874 82750
rect 6302 82738 6354 82750
rect 2258 82686 2270 82738
rect 2322 82686 2334 82738
rect 1822 82674 1874 82686
rect 6302 82674 6354 82686
rect 10670 82738 10722 82750
rect 10670 82674 10722 82686
rect 10894 82738 10946 82750
rect 10894 82674 10946 82686
rect 11342 82738 11394 82750
rect 11342 82674 11394 82686
rect 14142 82738 14194 82750
rect 14142 82674 14194 82686
rect 14478 82738 14530 82750
rect 16830 82738 16882 82750
rect 24558 82738 24610 82750
rect 16482 82686 16494 82738
rect 16546 82686 16558 82738
rect 17602 82686 17614 82738
rect 17666 82686 17678 82738
rect 17826 82686 17838 82738
rect 17890 82686 17902 82738
rect 24098 82686 24110 82738
rect 24162 82686 24174 82738
rect 14478 82674 14530 82686
rect 16830 82674 16882 82686
rect 24558 82674 24610 82686
rect 25790 82738 25842 82750
rect 25790 82674 25842 82686
rect 6750 82626 6802 82638
rect 6750 82562 6802 82574
rect 7198 82626 7250 82638
rect 7198 82562 7250 82574
rect 7646 82626 7698 82638
rect 7646 82562 7698 82574
rect 11230 82626 11282 82638
rect 11230 82562 11282 82574
rect 12574 82626 12626 82638
rect 12574 82562 12626 82574
rect 13358 82626 13410 82638
rect 15486 82626 15538 82638
rect 13682 82574 13694 82626
rect 13746 82574 13758 82626
rect 13358 82562 13410 82574
rect 15486 82562 15538 82574
rect 18846 82626 18898 82638
rect 18846 82562 18898 82574
rect 5630 82514 5682 82526
rect 5630 82450 5682 82462
rect 6190 82514 6242 82526
rect 21086 82514 21138 82526
rect 15474 82462 15486 82514
rect 15538 82511 15550 82514
rect 16034 82511 16046 82514
rect 15538 82465 16046 82511
rect 15538 82462 15550 82465
rect 16034 82462 16046 82465
rect 16098 82462 16110 82514
rect 6190 82450 6242 82462
rect 21086 82450 21138 82462
rect 1344 82346 38640 82380
rect 1344 82294 4024 82346
rect 4076 82294 4148 82346
rect 4200 82294 4272 82346
rect 4324 82294 4396 82346
rect 4448 82294 4520 82346
rect 4572 82294 4644 82346
rect 4696 82294 4768 82346
rect 4820 82294 4892 82346
rect 4944 82294 5016 82346
rect 5068 82294 5140 82346
rect 5192 82294 24024 82346
rect 24076 82294 24148 82346
rect 24200 82294 24272 82346
rect 24324 82294 24396 82346
rect 24448 82294 24520 82346
rect 24572 82294 24644 82346
rect 24696 82294 24768 82346
rect 24820 82294 24892 82346
rect 24944 82294 25016 82346
rect 25068 82294 25140 82346
rect 25192 82294 38640 82346
rect 1344 82260 38640 82294
rect 20638 82178 20690 82190
rect 20638 82114 20690 82126
rect 4510 82066 4562 82078
rect 4510 82002 4562 82014
rect 5966 82066 6018 82078
rect 5966 82002 6018 82014
rect 6414 82066 6466 82078
rect 6414 82002 6466 82014
rect 9438 82066 9490 82078
rect 14478 82066 14530 82078
rect 10434 82014 10446 82066
rect 10498 82014 10510 82066
rect 9438 82002 9490 82014
rect 14478 82002 14530 82014
rect 21422 82066 21474 82078
rect 21422 82002 21474 82014
rect 22430 82066 22482 82078
rect 22430 82002 22482 82014
rect 10110 81954 10162 81966
rect 10110 81890 10162 81902
rect 10334 81954 10386 81966
rect 11118 81954 11170 81966
rect 10546 81902 10558 81954
rect 10610 81902 10622 81954
rect 10334 81890 10386 81902
rect 11118 81890 11170 81902
rect 11342 81954 11394 81966
rect 11342 81890 11394 81902
rect 11454 81954 11506 81966
rect 11454 81890 11506 81902
rect 11790 81954 11842 81966
rect 15038 81954 15090 81966
rect 12114 81902 12126 81954
rect 12178 81902 12190 81954
rect 11790 81890 11842 81902
rect 15038 81890 15090 81902
rect 15262 81954 15314 81966
rect 15262 81890 15314 81902
rect 16158 81954 16210 81966
rect 16158 81890 16210 81902
rect 16270 81954 16322 81966
rect 16270 81890 16322 81902
rect 16606 81954 16658 81966
rect 16606 81890 16658 81902
rect 16942 81954 16994 81966
rect 17490 81902 17502 81954
rect 17554 81902 17566 81954
rect 16942 81890 16994 81902
rect 1710 81842 1762 81854
rect 1710 81778 1762 81790
rect 4846 81842 4898 81854
rect 4846 81778 4898 81790
rect 9886 81842 9938 81854
rect 9886 81778 9938 81790
rect 10894 81842 10946 81854
rect 10894 81778 10946 81790
rect 12350 81842 12402 81854
rect 12350 81778 12402 81790
rect 13694 81842 13746 81854
rect 13694 81778 13746 81790
rect 13806 81842 13858 81854
rect 13806 81778 13858 81790
rect 14814 81842 14866 81854
rect 14814 81778 14866 81790
rect 15486 81842 15538 81854
rect 15486 81778 15538 81790
rect 22766 81842 22818 81854
rect 22766 81778 22818 81790
rect 4398 81730 4450 81742
rect 4398 81666 4450 81678
rect 4622 81730 4674 81742
rect 4622 81666 4674 81678
rect 11230 81730 11282 81742
rect 11230 81666 11282 81678
rect 12462 81730 12514 81742
rect 12462 81666 12514 81678
rect 14702 81730 14754 81742
rect 14702 81666 14754 81678
rect 16382 81730 16434 81742
rect 16382 81666 16434 81678
rect 16494 81730 16546 81742
rect 21982 81730 22034 81742
rect 20066 81678 20078 81730
rect 20130 81678 20142 81730
rect 16494 81666 16546 81678
rect 21982 81666 22034 81678
rect 22318 81730 22370 81742
rect 22318 81666 22370 81678
rect 22542 81730 22594 81742
rect 22542 81666 22594 81678
rect 1344 81562 38640 81596
rect 1344 81510 14024 81562
rect 14076 81510 14148 81562
rect 14200 81510 14272 81562
rect 14324 81510 14396 81562
rect 14448 81510 14520 81562
rect 14572 81510 14644 81562
rect 14696 81510 14768 81562
rect 14820 81510 14892 81562
rect 14944 81510 15016 81562
rect 15068 81510 15140 81562
rect 15192 81510 34024 81562
rect 34076 81510 34148 81562
rect 34200 81510 34272 81562
rect 34324 81510 34396 81562
rect 34448 81510 34520 81562
rect 34572 81510 34644 81562
rect 34696 81510 34768 81562
rect 34820 81510 34892 81562
rect 34944 81510 35016 81562
rect 35068 81510 35140 81562
rect 35192 81510 38640 81562
rect 1344 81476 38640 81510
rect 15374 81394 15426 81406
rect 15374 81330 15426 81342
rect 1710 81282 1762 81294
rect 1710 81218 1762 81230
rect 8318 81282 8370 81294
rect 8318 81218 8370 81230
rect 10894 81282 10946 81294
rect 10894 81218 10946 81230
rect 15262 81282 15314 81294
rect 15262 81218 15314 81230
rect 15934 81282 15986 81294
rect 15934 81218 15986 81230
rect 5630 81170 5682 81182
rect 10334 81170 10386 81182
rect 6066 81118 6078 81170
rect 6130 81118 6142 81170
rect 9650 81118 9662 81170
rect 9714 81118 9726 81170
rect 5630 81106 5682 81118
rect 10334 81106 10386 81118
rect 10446 81170 10498 81182
rect 11678 81170 11730 81182
rect 10546 81118 10558 81170
rect 10610 81118 10622 81170
rect 10446 81106 10498 81118
rect 11678 81106 11730 81118
rect 11902 81170 11954 81182
rect 11902 81106 11954 81118
rect 12350 81170 12402 81182
rect 15486 81170 15538 81182
rect 14802 81118 14814 81170
rect 14866 81118 14878 81170
rect 15026 81118 15038 81170
rect 15090 81118 15102 81170
rect 12350 81106 12402 81118
rect 15486 81106 15538 81118
rect 16046 81170 16098 81182
rect 16046 81106 16098 81118
rect 16494 81170 16546 81182
rect 16494 81106 16546 81118
rect 16718 81170 16770 81182
rect 16718 81106 16770 81118
rect 17390 81170 17442 81182
rect 18274 81118 18286 81170
rect 18338 81118 18350 81170
rect 19282 81118 19294 81170
rect 19346 81118 19358 81170
rect 22530 81118 22542 81170
rect 22594 81118 22606 81170
rect 17390 81106 17442 81118
rect 5182 81058 5234 81070
rect 12126 81058 12178 81070
rect 9874 81006 9886 81058
rect 9938 81006 9950 81058
rect 5182 80994 5234 81006
rect 12126 80994 12178 81006
rect 13470 81058 13522 81070
rect 13470 80994 13522 81006
rect 13918 81058 13970 81070
rect 13918 80994 13970 81006
rect 14366 81058 14418 81070
rect 20078 81058 20130 81070
rect 16258 81006 16270 81058
rect 16322 81006 16334 81058
rect 18050 81006 18062 81058
rect 18114 81006 18126 81058
rect 19170 81006 19182 81058
rect 19234 81006 19246 81058
rect 14366 80994 14418 81006
rect 20078 80994 20130 81006
rect 20526 81058 20578 81070
rect 20526 80994 20578 81006
rect 22206 81058 22258 81070
rect 23662 81058 23714 81070
rect 22306 81006 22318 81058
rect 22370 81006 22382 81058
rect 22206 80994 22258 81006
rect 23662 80994 23714 81006
rect 9102 80946 9154 80958
rect 9102 80882 9154 80894
rect 11118 80946 11170 80958
rect 11118 80882 11170 80894
rect 11230 80946 11282 80958
rect 11230 80882 11282 80894
rect 12798 80946 12850 80958
rect 18946 80894 18958 80946
rect 19010 80894 19022 80946
rect 12798 80882 12850 80894
rect 1344 80778 38640 80812
rect 1344 80726 4024 80778
rect 4076 80726 4148 80778
rect 4200 80726 4272 80778
rect 4324 80726 4396 80778
rect 4448 80726 4520 80778
rect 4572 80726 4644 80778
rect 4696 80726 4768 80778
rect 4820 80726 4892 80778
rect 4944 80726 5016 80778
rect 5068 80726 5140 80778
rect 5192 80726 24024 80778
rect 24076 80726 24148 80778
rect 24200 80726 24272 80778
rect 24324 80726 24396 80778
rect 24448 80726 24520 80778
rect 24572 80726 24644 80778
rect 24696 80726 24768 80778
rect 24820 80726 24892 80778
rect 24944 80726 25016 80778
rect 25068 80726 25140 80778
rect 25192 80726 38640 80778
rect 1344 80692 38640 80726
rect 5966 80610 6018 80622
rect 5966 80546 6018 80558
rect 6078 80610 6130 80622
rect 6078 80546 6130 80558
rect 6750 80610 6802 80622
rect 7982 80610 8034 80622
rect 6962 80558 6974 80610
rect 7026 80607 7038 80610
rect 7746 80607 7758 80610
rect 7026 80561 7758 80607
rect 7026 80558 7038 80561
rect 7746 80558 7758 80561
rect 7810 80558 7822 80610
rect 6750 80546 6802 80558
rect 7982 80546 8034 80558
rect 10334 80610 10386 80622
rect 19406 80610 19458 80622
rect 15138 80558 15150 80610
rect 15202 80558 15214 80610
rect 10334 80546 10386 80558
rect 19406 80546 19458 80558
rect 9774 80498 9826 80510
rect 9774 80434 9826 80446
rect 10110 80498 10162 80510
rect 19966 80498 20018 80510
rect 11666 80446 11678 80498
rect 11730 80446 11742 80498
rect 10110 80434 10162 80446
rect 19966 80434 20018 80446
rect 6078 80386 6130 80398
rect 6078 80322 6130 80334
rect 6526 80386 6578 80398
rect 6526 80322 6578 80334
rect 7310 80386 7362 80398
rect 7310 80322 7362 80334
rect 9886 80386 9938 80398
rect 14142 80386 14194 80398
rect 11890 80334 11902 80386
rect 11954 80334 11966 80386
rect 9886 80322 9938 80334
rect 14142 80322 14194 80334
rect 14478 80386 14530 80398
rect 14478 80322 14530 80334
rect 14590 80386 14642 80398
rect 14590 80322 14642 80334
rect 14702 80386 14754 80398
rect 15810 80334 15822 80386
rect 15874 80334 15886 80386
rect 16258 80334 16270 80386
rect 16322 80334 16334 80386
rect 14702 80322 14754 80334
rect 8318 80274 8370 80286
rect 8318 80210 8370 80222
rect 8654 80274 8706 80286
rect 8654 80210 8706 80222
rect 8766 80274 8818 80286
rect 8766 80210 8818 80222
rect 9214 80274 9266 80286
rect 9214 80210 9266 80222
rect 11230 80274 11282 80286
rect 11230 80210 11282 80222
rect 13806 80274 13858 80286
rect 13806 80210 13858 80222
rect 1710 80162 1762 80174
rect 1710 80098 1762 80110
rect 8094 80162 8146 80174
rect 8094 80098 8146 80110
rect 9662 80162 9714 80174
rect 9662 80098 9714 80110
rect 11454 80162 11506 80174
rect 11454 80098 11506 80110
rect 11678 80162 11730 80174
rect 11678 80098 11730 80110
rect 12910 80162 12962 80174
rect 12910 80098 12962 80110
rect 13918 80162 13970 80174
rect 18834 80110 18846 80162
rect 18898 80110 18910 80162
rect 13918 80098 13970 80110
rect 1344 79994 38640 80028
rect 1344 79942 14024 79994
rect 14076 79942 14148 79994
rect 14200 79942 14272 79994
rect 14324 79942 14396 79994
rect 14448 79942 14520 79994
rect 14572 79942 14644 79994
rect 14696 79942 14768 79994
rect 14820 79942 14892 79994
rect 14944 79942 15016 79994
rect 15068 79942 15140 79994
rect 15192 79942 34024 79994
rect 34076 79942 34148 79994
rect 34200 79942 34272 79994
rect 34324 79942 34396 79994
rect 34448 79942 34520 79994
rect 34572 79942 34644 79994
rect 34696 79942 34768 79994
rect 34820 79942 34892 79994
rect 34944 79942 35016 79994
rect 35068 79942 35140 79994
rect 35192 79942 38640 79994
rect 1344 79908 38640 79942
rect 5854 79826 5906 79838
rect 4722 79774 4734 79826
rect 4786 79774 4798 79826
rect 5854 79762 5906 79774
rect 6302 79826 6354 79838
rect 6302 79762 6354 79774
rect 6750 79826 6802 79838
rect 6750 79762 6802 79774
rect 17502 79826 17554 79838
rect 17502 79762 17554 79774
rect 7422 79714 7474 79726
rect 7422 79650 7474 79662
rect 7534 79714 7586 79726
rect 14130 79662 14142 79714
rect 14194 79662 14206 79714
rect 15138 79662 15150 79714
rect 15202 79662 15214 79714
rect 7534 79650 7586 79662
rect 1822 79602 1874 79614
rect 5406 79602 5458 79614
rect 8654 79602 8706 79614
rect 13246 79602 13298 79614
rect 2258 79550 2270 79602
rect 2322 79550 2334 79602
rect 8306 79550 8318 79602
rect 8370 79550 8382 79602
rect 10994 79550 11006 79602
rect 11058 79550 11070 79602
rect 11554 79550 11566 79602
rect 11618 79550 11630 79602
rect 12002 79550 12014 79602
rect 12066 79550 12078 79602
rect 13010 79550 13022 79602
rect 13074 79550 13086 79602
rect 13682 79550 13694 79602
rect 13746 79550 13758 79602
rect 15250 79550 15262 79602
rect 15314 79550 15326 79602
rect 22082 79550 22094 79602
rect 22146 79550 22158 79602
rect 1822 79538 1874 79550
rect 5406 79538 5458 79550
rect 8654 79538 8706 79550
rect 13246 79538 13298 79550
rect 20638 79490 20690 79502
rect 13794 79438 13806 79490
rect 13858 79438 13870 79490
rect 20638 79426 20690 79438
rect 20974 79490 21026 79502
rect 22654 79490 22706 79502
rect 22194 79438 22206 79490
rect 22258 79438 22270 79490
rect 20974 79426 21026 79438
rect 22654 79426 22706 79438
rect 12910 79378 12962 79390
rect 7970 79326 7982 79378
rect 8034 79326 8046 79378
rect 20626 79326 20638 79378
rect 20690 79375 20702 79378
rect 21410 79375 21422 79378
rect 20690 79329 21422 79375
rect 20690 79326 20702 79329
rect 21410 79326 21422 79329
rect 21474 79326 21486 79378
rect 12910 79314 12962 79326
rect 1344 79210 38640 79244
rect 1344 79158 4024 79210
rect 4076 79158 4148 79210
rect 4200 79158 4272 79210
rect 4324 79158 4396 79210
rect 4448 79158 4520 79210
rect 4572 79158 4644 79210
rect 4696 79158 4768 79210
rect 4820 79158 4892 79210
rect 4944 79158 5016 79210
rect 5068 79158 5140 79210
rect 5192 79158 24024 79210
rect 24076 79158 24148 79210
rect 24200 79158 24272 79210
rect 24324 79158 24396 79210
rect 24448 79158 24520 79210
rect 24572 79158 24644 79210
rect 24696 79158 24768 79210
rect 24820 79158 24892 79210
rect 24944 79158 25016 79210
rect 25068 79158 25140 79210
rect 25192 79158 38640 79210
rect 1344 79124 38640 79158
rect 3278 79042 3330 79054
rect 3278 78978 3330 78990
rect 13918 79042 13970 79054
rect 13918 78978 13970 78990
rect 3390 78930 3442 78942
rect 12014 78930 12066 78942
rect 4498 78878 4510 78930
rect 4562 78878 4574 78930
rect 6514 78878 6526 78930
rect 6578 78878 6590 78930
rect 15922 78878 15934 78930
rect 15986 78878 15998 78930
rect 19954 78878 19966 78930
rect 20018 78878 20030 78930
rect 23314 78878 23326 78930
rect 23378 78878 23390 78930
rect 3390 78866 3442 78878
rect 12014 78866 12066 78878
rect 4622 78818 4674 78830
rect 7534 78818 7586 78830
rect 11230 78818 11282 78830
rect 6066 78766 6078 78818
rect 6130 78766 6142 78818
rect 8194 78766 8206 78818
rect 8258 78766 8270 78818
rect 4622 78754 4674 78766
rect 7534 78754 7586 78766
rect 11230 78754 11282 78766
rect 11566 78818 11618 78830
rect 22206 78818 22258 78830
rect 13906 78766 13918 78818
rect 13970 78766 13982 78818
rect 14242 78766 14254 78818
rect 14306 78766 14318 78818
rect 15586 78766 15598 78818
rect 15650 78766 15662 78818
rect 16034 78766 16046 78818
rect 16098 78766 16110 78818
rect 20290 78766 20302 78818
rect 20354 78766 20366 78818
rect 11566 78754 11618 78766
rect 22206 78754 22258 78766
rect 5070 78706 5122 78718
rect 5070 78642 5122 78654
rect 5630 78706 5682 78718
rect 5630 78642 5682 78654
rect 13582 78706 13634 78718
rect 20750 78706 20802 78718
rect 22990 78706 23042 78718
rect 15474 78654 15486 78706
rect 15538 78654 15550 78706
rect 16258 78654 16270 78706
rect 16322 78654 16334 78706
rect 21410 78654 21422 78706
rect 21474 78654 21486 78706
rect 21858 78654 21870 78706
rect 21922 78654 21934 78706
rect 13582 78642 13634 78654
rect 20750 78642 20802 78654
rect 22990 78642 23042 78654
rect 23214 78706 23266 78718
rect 23214 78642 23266 78654
rect 1710 78594 1762 78606
rect 1710 78530 1762 78542
rect 4174 78594 4226 78606
rect 4174 78530 4226 78542
rect 4510 78594 4562 78606
rect 4510 78530 4562 78542
rect 4846 78594 4898 78606
rect 4846 78530 4898 78542
rect 7086 78594 7138 78606
rect 11454 78594 11506 78606
rect 10658 78542 10670 78594
rect 10722 78542 10734 78594
rect 7086 78530 7138 78542
rect 11454 78530 11506 78542
rect 22542 78594 22594 78606
rect 22542 78530 22594 78542
rect 1344 78426 38640 78460
rect 1344 78374 14024 78426
rect 14076 78374 14148 78426
rect 14200 78374 14272 78426
rect 14324 78374 14396 78426
rect 14448 78374 14520 78426
rect 14572 78374 14644 78426
rect 14696 78374 14768 78426
rect 14820 78374 14892 78426
rect 14944 78374 15016 78426
rect 15068 78374 15140 78426
rect 15192 78374 34024 78426
rect 34076 78374 34148 78426
rect 34200 78374 34272 78426
rect 34324 78374 34396 78426
rect 34448 78374 34520 78426
rect 34572 78374 34644 78426
rect 34696 78374 34768 78426
rect 34820 78374 34892 78426
rect 34944 78374 35016 78426
rect 35068 78374 35140 78426
rect 35192 78374 38640 78426
rect 1344 78340 38640 78374
rect 5294 78258 5346 78270
rect 4722 78206 4734 78258
rect 4786 78206 4798 78258
rect 5294 78194 5346 78206
rect 9886 78258 9938 78270
rect 9886 78194 9938 78206
rect 15262 78258 15314 78270
rect 15262 78194 15314 78206
rect 20302 78258 20354 78270
rect 24334 78258 24386 78270
rect 20962 78206 20974 78258
rect 21026 78206 21038 78258
rect 20302 78194 20354 78206
rect 24334 78194 24386 78206
rect 25342 78258 25394 78270
rect 25342 78194 25394 78206
rect 7310 78146 7362 78158
rect 6178 78094 6190 78146
rect 6242 78094 6254 78146
rect 6738 78094 6750 78146
rect 6802 78094 6814 78146
rect 7310 78082 7362 78094
rect 8878 78146 8930 78158
rect 8878 78082 8930 78094
rect 1822 78034 1874 78046
rect 5966 78034 6018 78046
rect 2258 77982 2270 78034
rect 2322 77982 2334 78034
rect 1822 77970 1874 77982
rect 5966 77970 6018 77982
rect 7198 78034 7250 78046
rect 7198 77970 7250 77982
rect 7758 78034 7810 78046
rect 7758 77970 7810 77982
rect 9550 78034 9602 78046
rect 9550 77970 9602 77982
rect 9886 78034 9938 78046
rect 9886 77970 9938 77982
rect 10110 78034 10162 78046
rect 10110 77970 10162 77982
rect 10558 78034 10610 78046
rect 15150 78034 15202 78046
rect 12450 77982 12462 78034
rect 12514 77982 12526 78034
rect 10558 77970 10610 77982
rect 15150 77970 15202 77982
rect 15374 78034 15426 78046
rect 15374 77970 15426 77982
rect 15822 78034 15874 78046
rect 23314 77982 23326 78034
rect 23378 77982 23390 78034
rect 23874 77982 23886 78034
rect 23938 77982 23950 78034
rect 15822 77970 15874 77982
rect 8318 77922 8370 77934
rect 11342 77922 11394 77934
rect 15598 77922 15650 77934
rect 8978 77870 8990 77922
rect 9042 77870 9054 77922
rect 13570 77870 13582 77922
rect 13634 77870 13646 77922
rect 8318 77858 8370 77870
rect 11342 77858 11394 77870
rect 15598 77858 15650 77870
rect 16382 77922 16434 77934
rect 16382 77858 16434 77870
rect 5630 77810 5682 77822
rect 5630 77746 5682 77758
rect 7310 77810 7362 77822
rect 7310 77746 7362 77758
rect 7870 77810 7922 77822
rect 7870 77746 7922 77758
rect 8654 77810 8706 77822
rect 8654 77746 8706 77758
rect 1344 77642 38640 77676
rect 1344 77590 4024 77642
rect 4076 77590 4148 77642
rect 4200 77590 4272 77642
rect 4324 77590 4396 77642
rect 4448 77590 4520 77642
rect 4572 77590 4644 77642
rect 4696 77590 4768 77642
rect 4820 77590 4892 77642
rect 4944 77590 5016 77642
rect 5068 77590 5140 77642
rect 5192 77590 24024 77642
rect 24076 77590 24148 77642
rect 24200 77590 24272 77642
rect 24324 77590 24396 77642
rect 24448 77590 24520 77642
rect 24572 77590 24644 77642
rect 24696 77590 24768 77642
rect 24820 77590 24892 77642
rect 24944 77590 25016 77642
rect 25068 77590 25140 77642
rect 25192 77590 38640 77642
rect 1344 77556 38640 77590
rect 3278 77474 3330 77486
rect 3278 77410 3330 77422
rect 3614 77474 3666 77486
rect 3614 77410 3666 77422
rect 25678 77362 25730 77374
rect 25678 77298 25730 77310
rect 5070 77250 5122 77262
rect 5070 77186 5122 77198
rect 5742 77250 5794 77262
rect 5742 77186 5794 77198
rect 6638 77250 6690 77262
rect 6638 77186 6690 77198
rect 6974 77250 7026 77262
rect 21198 77250 21250 77262
rect 25230 77250 25282 77262
rect 9650 77198 9662 77250
rect 9714 77198 9726 77250
rect 10098 77198 10110 77250
rect 10162 77198 10174 77250
rect 13794 77198 13806 77250
rect 13858 77198 13870 77250
rect 14578 77198 14590 77250
rect 14642 77198 14654 77250
rect 15474 77198 15486 77250
rect 15538 77198 15550 77250
rect 24210 77198 24222 77250
rect 24274 77198 24286 77250
rect 24770 77198 24782 77250
rect 24834 77198 24846 77250
rect 6974 77186 7026 77198
rect 21198 77186 21250 77198
rect 25230 77186 25282 77198
rect 1710 77138 1762 77150
rect 5966 77138 6018 77150
rect 3826 77086 3838 77138
rect 3890 77086 3902 77138
rect 4274 77086 4286 77138
rect 4338 77086 4350 77138
rect 1710 77074 1762 77086
rect 5966 77074 6018 77086
rect 6302 77138 6354 77150
rect 6302 77074 6354 77086
rect 6750 77138 6802 77150
rect 10558 77138 10610 77150
rect 21982 77138 22034 77150
rect 7970 77086 7982 77138
rect 8034 77086 8046 77138
rect 14690 77086 14702 77138
rect 14754 77086 14766 77138
rect 15362 77086 15374 77138
rect 15426 77086 15438 77138
rect 6750 77074 6802 77086
rect 10558 77074 10610 77086
rect 21982 77074 22034 77086
rect 6078 77026 6130 77038
rect 6078 76962 6130 76974
rect 7534 77026 7586 77038
rect 7534 76962 7586 76974
rect 8430 77026 8482 77038
rect 15138 76974 15150 77026
rect 15202 76974 15214 77026
rect 8430 76962 8482 76974
rect 1344 76858 38640 76892
rect 1344 76806 14024 76858
rect 14076 76806 14148 76858
rect 14200 76806 14272 76858
rect 14324 76806 14396 76858
rect 14448 76806 14520 76858
rect 14572 76806 14644 76858
rect 14696 76806 14768 76858
rect 14820 76806 14892 76858
rect 14944 76806 15016 76858
rect 15068 76806 15140 76858
rect 15192 76806 34024 76858
rect 34076 76806 34148 76858
rect 34200 76806 34272 76858
rect 34324 76806 34396 76858
rect 34448 76806 34520 76858
rect 34572 76806 34644 76858
rect 34696 76806 34768 76858
rect 34820 76806 34892 76858
rect 34944 76806 35016 76858
rect 35068 76806 35140 76858
rect 35192 76806 38640 76858
rect 1344 76772 38640 76806
rect 4734 76690 4786 76702
rect 4734 76626 4786 76638
rect 5406 76690 5458 76702
rect 5406 76626 5458 76638
rect 9774 76690 9826 76702
rect 16830 76690 16882 76702
rect 13794 76638 13806 76690
rect 13858 76638 13870 76690
rect 9774 76626 9826 76638
rect 16830 76626 16882 76638
rect 18734 76690 18786 76702
rect 18734 76626 18786 76638
rect 20302 76690 20354 76702
rect 20302 76626 20354 76638
rect 22318 76690 22370 76702
rect 22318 76626 22370 76638
rect 1710 76578 1762 76590
rect 1710 76514 1762 76526
rect 14590 76578 14642 76590
rect 17390 76578 17442 76590
rect 15250 76526 15262 76578
rect 15314 76526 15326 76578
rect 15810 76526 15822 76578
rect 15874 76526 15886 76578
rect 14590 76514 14642 76526
rect 17390 76514 17442 76526
rect 17726 76578 17778 76590
rect 21298 76526 21310 76578
rect 21362 76526 21374 76578
rect 21746 76526 21758 76578
rect 21810 76526 21822 76578
rect 17726 76514 17778 76526
rect 11118 76466 11170 76478
rect 16382 76466 16434 76478
rect 11554 76414 11566 76466
rect 11618 76414 11630 76466
rect 15922 76414 15934 76466
rect 15986 76414 15998 76466
rect 11118 76402 11170 76414
rect 16382 76402 16434 76414
rect 17838 76466 17890 76478
rect 17838 76402 17890 76414
rect 18398 76466 18450 76478
rect 18398 76402 18450 76414
rect 18846 76466 18898 76478
rect 18846 76402 18898 76414
rect 21982 76466 22034 76478
rect 21982 76402 22034 76414
rect 6526 76354 6578 76366
rect 6526 76290 6578 76302
rect 10222 76354 10274 76366
rect 10222 76290 10274 76302
rect 10670 76354 10722 76366
rect 10670 76290 10722 76302
rect 14702 76354 14754 76366
rect 14702 76290 14754 76302
rect 17502 76354 17554 76366
rect 17502 76290 17554 76302
rect 18286 76354 18338 76366
rect 18286 76290 18338 76302
rect 20750 76354 20802 76366
rect 20750 76290 20802 76302
rect 1344 76074 38640 76108
rect 1344 76022 4024 76074
rect 4076 76022 4148 76074
rect 4200 76022 4272 76074
rect 4324 76022 4396 76074
rect 4448 76022 4520 76074
rect 4572 76022 4644 76074
rect 4696 76022 4768 76074
rect 4820 76022 4892 76074
rect 4944 76022 5016 76074
rect 5068 76022 5140 76074
rect 5192 76022 24024 76074
rect 24076 76022 24148 76074
rect 24200 76022 24272 76074
rect 24324 76022 24396 76074
rect 24448 76022 24520 76074
rect 24572 76022 24644 76074
rect 24696 76022 24768 76074
rect 24820 76022 24892 76074
rect 24944 76022 25016 76074
rect 25068 76022 25140 76074
rect 25192 76022 38640 76074
rect 1344 75988 38640 76022
rect 11006 75906 11058 75918
rect 11006 75842 11058 75854
rect 11678 75906 11730 75918
rect 11678 75842 11730 75854
rect 12014 75906 12066 75918
rect 12014 75842 12066 75854
rect 20190 75906 20242 75918
rect 20190 75842 20242 75854
rect 4398 75794 4450 75806
rect 6750 75794 6802 75806
rect 14478 75794 14530 75806
rect 5842 75742 5854 75794
rect 5906 75742 5918 75794
rect 9650 75742 9662 75794
rect 9714 75742 9726 75794
rect 4398 75730 4450 75742
rect 6750 75730 6802 75742
rect 14478 75730 14530 75742
rect 14926 75794 14978 75806
rect 14926 75730 14978 75742
rect 15374 75794 15426 75806
rect 15374 75730 15426 75742
rect 6078 75682 6130 75694
rect 10894 75682 10946 75694
rect 15710 75682 15762 75694
rect 5618 75630 5630 75682
rect 5682 75630 5694 75682
rect 6290 75630 6302 75682
rect 6354 75630 6366 75682
rect 8530 75630 8542 75682
rect 8594 75630 8606 75682
rect 12786 75630 12798 75682
rect 12850 75630 12862 75682
rect 6078 75618 6130 75630
rect 10894 75618 10946 75630
rect 15710 75618 15762 75630
rect 16046 75682 16098 75694
rect 16046 75618 16098 75630
rect 16494 75682 16546 75694
rect 17154 75630 17166 75682
rect 17218 75630 17230 75682
rect 16494 75618 16546 75630
rect 5854 75570 5906 75582
rect 16270 75570 16322 75582
rect 12562 75518 12574 75570
rect 12626 75518 12638 75570
rect 5854 75506 5906 75518
rect 16270 75506 16322 75518
rect 1710 75458 1762 75470
rect 1710 75394 1762 75406
rect 4286 75458 4338 75470
rect 4286 75394 4338 75406
rect 15934 75458 15986 75470
rect 20526 75458 20578 75470
rect 19394 75406 19406 75458
rect 19458 75406 19470 75458
rect 15934 75394 15986 75406
rect 20526 75394 20578 75406
rect 1344 75290 38640 75324
rect 1344 75238 14024 75290
rect 14076 75238 14148 75290
rect 14200 75238 14272 75290
rect 14324 75238 14396 75290
rect 14448 75238 14520 75290
rect 14572 75238 14644 75290
rect 14696 75238 14768 75290
rect 14820 75238 14892 75290
rect 14944 75238 15016 75290
rect 15068 75238 15140 75290
rect 15192 75238 34024 75290
rect 34076 75238 34148 75290
rect 34200 75238 34272 75290
rect 34324 75238 34396 75290
rect 34448 75238 34520 75290
rect 34572 75238 34644 75290
rect 34696 75238 34768 75290
rect 34820 75238 34892 75290
rect 34944 75238 35016 75290
rect 35068 75238 35140 75290
rect 35192 75238 38640 75290
rect 1344 75204 38640 75238
rect 6974 75122 7026 75134
rect 6066 75070 6078 75122
rect 6130 75070 6142 75122
rect 6974 75058 7026 75070
rect 8878 75122 8930 75134
rect 8878 75058 8930 75070
rect 13358 75122 13410 75134
rect 13358 75058 13410 75070
rect 14254 75122 14306 75134
rect 14254 75058 14306 75070
rect 15710 75122 15762 75134
rect 15710 75058 15762 75070
rect 16158 75122 16210 75134
rect 16158 75058 16210 75070
rect 17838 75122 17890 75134
rect 17838 75058 17890 75070
rect 9886 75010 9938 75022
rect 9886 74946 9938 74958
rect 9998 75010 10050 75022
rect 9998 74946 10050 74958
rect 11678 75010 11730 75022
rect 11678 74946 11730 74958
rect 12686 75010 12738 75022
rect 12686 74946 12738 74958
rect 16606 75010 16658 75022
rect 16606 74946 16658 74958
rect 16830 75010 16882 75022
rect 16830 74946 16882 74958
rect 17726 75010 17778 75022
rect 17726 74946 17778 74958
rect 17950 75010 18002 75022
rect 17950 74946 18002 74958
rect 3166 74898 3218 74910
rect 7982 74898 8034 74910
rect 3602 74846 3614 74898
rect 3666 74846 3678 74898
rect 3166 74834 3218 74846
rect 7982 74834 8034 74846
rect 8990 74898 9042 74910
rect 8990 74834 9042 74846
rect 10222 74898 10274 74910
rect 12238 74898 12290 74910
rect 10770 74846 10782 74898
rect 10834 74846 10846 74898
rect 10222 74834 10274 74846
rect 12238 74834 12290 74846
rect 12910 74898 12962 74910
rect 12910 74834 12962 74846
rect 14366 74898 14418 74910
rect 14366 74834 14418 74846
rect 7422 74786 7474 74798
rect 7422 74722 7474 74734
rect 8542 74786 8594 74798
rect 12462 74786 12514 74798
rect 10882 74734 10894 74786
rect 10946 74734 10958 74786
rect 8542 74722 8594 74734
rect 12462 74722 12514 74734
rect 15262 74786 15314 74798
rect 18510 74786 18562 74798
rect 16482 74734 16494 74786
rect 16546 74734 16558 74786
rect 15262 74722 15314 74734
rect 18510 74722 18562 74734
rect 6638 74674 6690 74686
rect 8878 74674 8930 74686
rect 7410 74622 7422 74674
rect 7474 74671 7486 74674
rect 8306 74671 8318 74674
rect 7474 74625 8318 74671
rect 7474 74622 7486 74625
rect 8306 74622 8318 74625
rect 8370 74622 8382 74674
rect 15250 74622 15262 74674
rect 15314 74671 15326 74674
rect 16146 74671 16158 74674
rect 15314 74625 16158 74671
rect 15314 74622 15326 74625
rect 16146 74622 16158 74625
rect 16210 74622 16222 74674
rect 6638 74610 6690 74622
rect 8878 74610 8930 74622
rect 1344 74506 38640 74540
rect 1344 74454 4024 74506
rect 4076 74454 4148 74506
rect 4200 74454 4272 74506
rect 4324 74454 4396 74506
rect 4448 74454 4520 74506
rect 4572 74454 4644 74506
rect 4696 74454 4768 74506
rect 4820 74454 4892 74506
rect 4944 74454 5016 74506
rect 5068 74454 5140 74506
rect 5192 74454 24024 74506
rect 24076 74454 24148 74506
rect 24200 74454 24272 74506
rect 24324 74454 24396 74506
rect 24448 74454 24520 74506
rect 24572 74454 24644 74506
rect 24696 74454 24768 74506
rect 24820 74454 24892 74506
rect 24944 74454 25016 74506
rect 25068 74454 25140 74506
rect 25192 74454 38640 74506
rect 1344 74420 38640 74454
rect 10894 74338 10946 74350
rect 10894 74274 10946 74286
rect 12574 74338 12626 74350
rect 12574 74274 12626 74286
rect 12910 74338 12962 74350
rect 12910 74274 12962 74286
rect 19518 74338 19570 74350
rect 19518 74274 19570 74286
rect 5742 74226 5794 74238
rect 5742 74162 5794 74174
rect 6190 74226 6242 74238
rect 6190 74162 6242 74174
rect 6638 74226 6690 74238
rect 6638 74162 6690 74174
rect 11230 74226 11282 74238
rect 11230 74162 11282 74174
rect 11790 74226 11842 74238
rect 11790 74162 11842 74174
rect 3838 74114 3890 74126
rect 3838 74050 3890 74062
rect 7198 74114 7250 74126
rect 12238 74114 12290 74126
rect 7858 74062 7870 74114
rect 7922 74062 7934 74114
rect 7198 74050 7250 74062
rect 12238 74050 12290 74062
rect 15822 74114 15874 74126
rect 16370 74062 16382 74114
rect 16434 74062 16446 74114
rect 15822 74050 15874 74062
rect 3502 74002 3554 74014
rect 12798 74002 12850 74014
rect 4050 73950 4062 74002
rect 4114 73950 4126 74002
rect 4610 73950 4622 74002
rect 4674 73950 4686 74002
rect 3502 73938 3554 73950
rect 12798 73938 12850 73950
rect 1710 73890 1762 73902
rect 1710 73826 1762 73838
rect 2158 73890 2210 73902
rect 15598 73890 15650 73902
rect 19854 73890 19906 73902
rect 10098 73838 10110 73890
rect 10162 73838 10174 73890
rect 18722 73838 18734 73890
rect 18786 73838 18798 73890
rect 2158 73826 2210 73838
rect 15598 73826 15650 73838
rect 19854 73826 19906 73838
rect 1344 73722 38640 73756
rect 1344 73670 14024 73722
rect 14076 73670 14148 73722
rect 14200 73670 14272 73722
rect 14324 73670 14396 73722
rect 14448 73670 14520 73722
rect 14572 73670 14644 73722
rect 14696 73670 14768 73722
rect 14820 73670 14892 73722
rect 14944 73670 15016 73722
rect 15068 73670 15140 73722
rect 15192 73670 34024 73722
rect 34076 73670 34148 73722
rect 34200 73670 34272 73722
rect 34324 73670 34396 73722
rect 34448 73670 34520 73722
rect 34572 73670 34644 73722
rect 34696 73670 34768 73722
rect 34820 73670 34892 73722
rect 34944 73670 35016 73722
rect 35068 73670 35140 73722
rect 35192 73670 38640 73722
rect 1344 73636 38640 73670
rect 5294 73554 5346 73566
rect 4722 73502 4734 73554
rect 4786 73502 4798 73554
rect 5294 73490 5346 73502
rect 9102 73554 9154 73566
rect 9102 73490 9154 73502
rect 9662 73554 9714 73566
rect 15150 73554 15202 73566
rect 14354 73502 14366 73554
rect 14418 73502 14430 73554
rect 9662 73490 9714 73502
rect 15150 73490 15202 73502
rect 15934 73554 15986 73566
rect 15934 73490 15986 73502
rect 8318 73442 8370 73454
rect 8318 73378 8370 73390
rect 20638 73442 20690 73454
rect 20638 73378 20690 73390
rect 1822 73330 1874 73342
rect 5630 73330 5682 73342
rect 9550 73330 9602 73342
rect 2258 73278 2270 73330
rect 2322 73278 2334 73330
rect 6066 73278 6078 73330
rect 6130 73278 6142 73330
rect 1822 73266 1874 73278
rect 5630 73266 5682 73278
rect 9550 73266 9602 73278
rect 9774 73330 9826 73342
rect 9774 73266 9826 73278
rect 10222 73330 10274 73342
rect 10222 73266 10274 73278
rect 11006 73330 11058 73342
rect 11006 73266 11058 73278
rect 11454 73330 11506 73342
rect 12114 73278 12126 73330
rect 12178 73278 12190 73330
rect 22866 73278 22878 73330
rect 22930 73278 22942 73330
rect 23426 73278 23438 73330
rect 23490 73278 23502 73330
rect 11454 73266 11506 73278
rect 10558 73218 10610 73230
rect 10558 73154 10610 73166
rect 15486 73218 15538 73230
rect 15486 73154 15538 73166
rect 23886 73218 23938 73230
rect 23886 73154 23938 73166
rect 24334 73218 24386 73230
rect 24334 73154 24386 73166
rect 19854 73106 19906 73118
rect 10770 73054 10782 73106
rect 10834 73103 10846 73106
rect 11330 73103 11342 73106
rect 10834 73057 11342 73103
rect 10834 73054 10846 73057
rect 11330 73054 11342 73057
rect 11394 73054 11406 73106
rect 19854 73042 19906 73054
rect 1344 72938 38640 72972
rect 1344 72886 4024 72938
rect 4076 72886 4148 72938
rect 4200 72886 4272 72938
rect 4324 72886 4396 72938
rect 4448 72886 4520 72938
rect 4572 72886 4644 72938
rect 4696 72886 4768 72938
rect 4820 72886 4892 72938
rect 4944 72886 5016 72938
rect 5068 72886 5140 72938
rect 5192 72886 24024 72938
rect 24076 72886 24148 72938
rect 24200 72886 24272 72938
rect 24324 72886 24396 72938
rect 24448 72886 24520 72938
rect 24572 72886 24644 72938
rect 24696 72886 24768 72938
rect 24820 72886 24892 72938
rect 24944 72886 25016 72938
rect 25068 72886 25140 72938
rect 25192 72886 38640 72938
rect 1344 72852 38640 72886
rect 3838 72770 3890 72782
rect 3838 72706 3890 72718
rect 21534 72770 21586 72782
rect 21534 72706 21586 72718
rect 7758 72658 7810 72670
rect 7758 72594 7810 72606
rect 9550 72658 9602 72670
rect 9550 72594 9602 72606
rect 4174 72546 4226 72558
rect 5966 72546 6018 72558
rect 4722 72494 4734 72546
rect 4786 72494 4798 72546
rect 4174 72482 4226 72494
rect 5966 72482 6018 72494
rect 6078 72546 6130 72558
rect 6078 72482 6130 72494
rect 7870 72546 7922 72558
rect 23538 72494 23550 72546
rect 23602 72494 23614 72546
rect 7870 72482 7922 72494
rect 8094 72434 8146 72446
rect 4946 72382 4958 72434
rect 5010 72382 5022 72434
rect 8094 72370 8146 72382
rect 1710 72322 1762 72334
rect 1710 72258 1762 72270
rect 7646 72322 7698 72334
rect 7646 72258 7698 72270
rect 8654 72322 8706 72334
rect 8654 72258 8706 72270
rect 9886 72322 9938 72334
rect 9886 72258 9938 72270
rect 24334 72322 24386 72334
rect 24334 72258 24386 72270
rect 1344 72154 38640 72188
rect 1344 72102 14024 72154
rect 14076 72102 14148 72154
rect 14200 72102 14272 72154
rect 14324 72102 14396 72154
rect 14448 72102 14520 72154
rect 14572 72102 14644 72154
rect 14696 72102 14768 72154
rect 14820 72102 14892 72154
rect 14944 72102 15016 72154
rect 15068 72102 15140 72154
rect 15192 72102 34024 72154
rect 34076 72102 34148 72154
rect 34200 72102 34272 72154
rect 34324 72102 34396 72154
rect 34448 72102 34520 72154
rect 34572 72102 34644 72154
rect 34696 72102 34768 72154
rect 34820 72102 34892 72154
rect 34944 72102 35016 72154
rect 35068 72102 35140 72154
rect 35192 72102 38640 72154
rect 1344 72068 38640 72102
rect 21758 71986 21810 71998
rect 18274 71934 18286 71986
rect 18338 71934 18350 71986
rect 21758 71922 21810 71934
rect 35534 71986 35586 71998
rect 35534 71922 35586 71934
rect 22306 71822 22318 71874
rect 22370 71822 22382 71874
rect 22642 71822 22654 71874
rect 22706 71822 22718 71874
rect 21198 71762 21250 71774
rect 35870 71762 35922 71774
rect 20738 71710 20750 71762
rect 20802 71710 20814 71762
rect 27794 71710 27806 71762
rect 27858 71710 27870 71762
rect 21198 71698 21250 71710
rect 35870 71698 35922 71710
rect 36094 71762 36146 71774
rect 36094 71698 36146 71710
rect 36318 71762 36370 71774
rect 36318 71698 36370 71710
rect 5294 71650 5346 71662
rect 5294 71586 5346 71598
rect 23438 71650 23490 71662
rect 23438 71586 23490 71598
rect 27470 71650 27522 71662
rect 35086 71650 35138 71662
rect 30146 71598 30158 71650
rect 30210 71598 30222 71650
rect 27470 71586 27522 71598
rect 35086 71586 35138 71598
rect 35982 71650 36034 71662
rect 35982 71586 36034 71598
rect 17726 71538 17778 71550
rect 17726 71474 17778 71486
rect 22094 71538 22146 71550
rect 22094 71474 22146 71486
rect 34974 71538 35026 71550
rect 34974 71474 35026 71486
rect 1344 71370 38640 71404
rect 1344 71318 4024 71370
rect 4076 71318 4148 71370
rect 4200 71318 4272 71370
rect 4324 71318 4396 71370
rect 4448 71318 4520 71370
rect 4572 71318 4644 71370
rect 4696 71318 4768 71370
rect 4820 71318 4892 71370
rect 4944 71318 5016 71370
rect 5068 71318 5140 71370
rect 5192 71318 24024 71370
rect 24076 71318 24148 71370
rect 24200 71318 24272 71370
rect 24324 71318 24396 71370
rect 24448 71318 24520 71370
rect 24572 71318 24644 71370
rect 24696 71318 24768 71370
rect 24820 71318 24892 71370
rect 24944 71318 25016 71370
rect 25068 71318 25140 71370
rect 25192 71318 38640 71370
rect 1344 71284 38640 71318
rect 20302 71202 20354 71214
rect 21522 71150 21534 71202
rect 21586 71199 21598 71202
rect 22306 71199 22318 71202
rect 21586 71153 22318 71199
rect 21586 71150 21598 71153
rect 22306 71150 22318 71153
rect 22370 71150 22382 71202
rect 20302 71138 20354 71150
rect 14814 71090 14866 71102
rect 14814 71026 14866 71038
rect 15262 71090 15314 71102
rect 15262 71026 15314 71038
rect 16046 71090 16098 71102
rect 16046 71026 16098 71038
rect 22318 71090 22370 71102
rect 25666 71038 25678 71090
rect 25730 71038 25742 71090
rect 22318 71026 22370 71038
rect 19966 70978 20018 70990
rect 19282 70926 19294 70978
rect 19346 70926 19358 70978
rect 19966 70914 20018 70926
rect 21422 70978 21474 70990
rect 21422 70914 21474 70926
rect 24222 70978 24274 70990
rect 32398 70978 32450 70990
rect 25106 70926 25118 70978
rect 25170 70926 25182 70978
rect 24222 70914 24274 70926
rect 32398 70914 32450 70926
rect 32622 70978 32674 70990
rect 32622 70914 32674 70926
rect 33070 70978 33122 70990
rect 33506 70926 33518 70978
rect 33570 70926 33582 70978
rect 33070 70914 33122 70926
rect 2830 70866 2882 70878
rect 2830 70802 2882 70814
rect 3166 70866 3218 70878
rect 19394 70814 19406 70866
rect 19458 70814 19470 70866
rect 3166 70802 3218 70814
rect 1710 70754 1762 70766
rect 1710 70690 1762 70702
rect 2606 70754 2658 70766
rect 2606 70690 2658 70702
rect 11118 70754 11170 70766
rect 11118 70690 11170 70702
rect 21870 70754 21922 70766
rect 21870 70690 21922 70702
rect 31838 70754 31890 70766
rect 36542 70754 36594 70766
rect 32050 70702 32062 70754
rect 32114 70702 32126 70754
rect 35746 70702 35758 70754
rect 35810 70702 35822 70754
rect 31838 70690 31890 70702
rect 36542 70690 36594 70702
rect 1344 70586 38640 70620
rect 1344 70534 14024 70586
rect 14076 70534 14148 70586
rect 14200 70534 14272 70586
rect 14324 70534 14396 70586
rect 14448 70534 14520 70586
rect 14572 70534 14644 70586
rect 14696 70534 14768 70586
rect 14820 70534 14892 70586
rect 14944 70534 15016 70586
rect 15068 70534 15140 70586
rect 15192 70534 34024 70586
rect 34076 70534 34148 70586
rect 34200 70534 34272 70586
rect 34324 70534 34396 70586
rect 34448 70534 34520 70586
rect 34572 70534 34644 70586
rect 34696 70534 34768 70586
rect 34820 70534 34892 70586
rect 34944 70534 35016 70586
rect 35068 70534 35140 70586
rect 35192 70534 38640 70586
rect 1344 70500 38640 70534
rect 7982 70418 8034 70430
rect 15150 70418 15202 70430
rect 13570 70366 13582 70418
rect 13634 70366 13646 70418
rect 7982 70354 8034 70366
rect 15150 70354 15202 70366
rect 16606 70418 16658 70430
rect 16606 70354 16658 70366
rect 33182 70418 33234 70430
rect 33182 70354 33234 70366
rect 1710 70306 1762 70318
rect 1710 70242 1762 70254
rect 9662 70306 9714 70318
rect 9662 70242 9714 70254
rect 16046 70306 16098 70318
rect 33406 70306 33458 70318
rect 18162 70254 18174 70306
rect 18226 70254 18238 70306
rect 18610 70254 18622 70306
rect 18674 70254 18686 70306
rect 16046 70242 16098 70254
rect 33406 70242 33458 70254
rect 36654 70306 36706 70318
rect 36654 70242 36706 70254
rect 7758 70194 7810 70206
rect 7758 70130 7810 70142
rect 8430 70194 8482 70206
rect 8430 70130 8482 70142
rect 9438 70194 9490 70206
rect 9438 70130 9490 70142
rect 9774 70194 9826 70206
rect 9774 70130 9826 70142
rect 10782 70194 10834 70206
rect 15598 70194 15650 70206
rect 11218 70142 11230 70194
rect 11282 70142 11294 70194
rect 10782 70130 10834 70142
rect 15598 70130 15650 70142
rect 15934 70194 15986 70206
rect 15934 70130 15986 70142
rect 16270 70194 16322 70206
rect 16270 70130 16322 70142
rect 16718 70194 16770 70206
rect 25118 70194 25170 70206
rect 17490 70142 17502 70194
rect 17554 70142 17566 70194
rect 17714 70142 17726 70194
rect 17778 70142 17790 70194
rect 18498 70142 18510 70194
rect 18562 70142 18574 70194
rect 16718 70130 16770 70142
rect 25118 70130 25170 70142
rect 25566 70194 25618 70206
rect 25566 70130 25618 70142
rect 25790 70194 25842 70206
rect 25790 70130 25842 70142
rect 26350 70194 26402 70206
rect 26350 70130 26402 70142
rect 27134 70194 27186 70206
rect 31614 70194 31666 70206
rect 37550 70194 37602 70206
rect 27906 70142 27918 70194
rect 27970 70142 27982 70194
rect 32050 70142 32062 70194
rect 32114 70142 32126 70194
rect 33842 70142 33854 70194
rect 33906 70142 33918 70194
rect 34402 70142 34414 70194
rect 34466 70142 34478 70194
rect 27134 70130 27186 70142
rect 31614 70130 31666 70142
rect 37550 70130 37602 70142
rect 37886 70194 37938 70206
rect 37886 70130 37938 70142
rect 38110 70194 38162 70206
rect 38110 70130 38162 70142
rect 7422 70082 7474 70094
rect 7422 70018 7474 70030
rect 7870 70082 7922 70094
rect 7870 70018 7922 70030
rect 8990 70082 9042 70094
rect 8990 70018 9042 70030
rect 10334 70082 10386 70094
rect 10334 70018 10386 70030
rect 19406 70082 19458 70094
rect 19406 70018 19458 70030
rect 24670 70082 24722 70094
rect 24670 70018 24722 70030
rect 25342 70082 25394 70094
rect 25342 70018 25394 70030
rect 26462 70082 26514 70094
rect 26462 70018 26514 70030
rect 29822 70082 29874 70094
rect 29822 70018 29874 70030
rect 31166 70082 31218 70094
rect 31166 70018 31218 70030
rect 32510 70082 32562 70094
rect 37774 70082 37826 70094
rect 33058 70030 33070 70082
rect 33122 70030 33134 70082
rect 32510 70018 32562 70030
rect 37774 70018 37826 70030
rect 14254 69970 14306 69982
rect 14254 69906 14306 69918
rect 15486 69970 15538 69982
rect 15486 69906 15538 69918
rect 16830 69970 16882 69982
rect 16830 69906 16882 69918
rect 31502 69970 31554 69982
rect 31502 69906 31554 69918
rect 31838 69970 31890 69982
rect 31838 69906 31890 69918
rect 37438 69970 37490 69982
rect 37438 69906 37490 69918
rect 1344 69802 38640 69836
rect 1344 69750 4024 69802
rect 4076 69750 4148 69802
rect 4200 69750 4272 69802
rect 4324 69750 4396 69802
rect 4448 69750 4520 69802
rect 4572 69750 4644 69802
rect 4696 69750 4768 69802
rect 4820 69750 4892 69802
rect 4944 69750 5016 69802
rect 5068 69750 5140 69802
rect 5192 69750 24024 69802
rect 24076 69750 24148 69802
rect 24200 69750 24272 69802
rect 24324 69750 24396 69802
rect 24448 69750 24520 69802
rect 24572 69750 24644 69802
rect 24696 69750 24768 69802
rect 24820 69750 24892 69802
rect 24944 69750 25016 69802
rect 25068 69750 25140 69802
rect 25192 69750 38640 69802
rect 1344 69716 38640 69750
rect 11678 69634 11730 69646
rect 11678 69570 11730 69582
rect 12014 69634 12066 69646
rect 12014 69570 12066 69582
rect 27582 69634 27634 69646
rect 33742 69634 33794 69646
rect 29138 69582 29150 69634
rect 29202 69631 29214 69634
rect 29810 69631 29822 69634
rect 29202 69585 29822 69631
rect 29202 69582 29214 69585
rect 29810 69582 29822 69585
rect 29874 69582 29886 69634
rect 27582 69570 27634 69582
rect 33742 69570 33794 69582
rect 34638 69634 34690 69646
rect 34638 69570 34690 69582
rect 34974 69634 35026 69646
rect 35522 69582 35534 69634
rect 35586 69582 35598 69634
rect 34974 69570 35026 69582
rect 14926 69522 14978 69534
rect 29262 69522 29314 69534
rect 17490 69470 17502 69522
rect 17554 69470 17566 69522
rect 14926 69458 14978 69470
rect 29262 69458 29314 69470
rect 29822 69522 29874 69534
rect 29822 69458 29874 69470
rect 6974 69410 7026 69422
rect 10558 69410 10610 69422
rect 7410 69358 7422 69410
rect 7474 69358 7486 69410
rect 6974 69346 7026 69358
rect 10558 69346 10610 69358
rect 13358 69410 13410 69422
rect 13358 69346 13410 69358
rect 13806 69410 13858 69422
rect 18398 69410 18450 69422
rect 23886 69410 23938 69422
rect 34750 69410 34802 69422
rect 36094 69410 36146 69422
rect 16930 69358 16942 69410
rect 16994 69358 17006 69410
rect 17378 69358 17390 69410
rect 17442 69358 17454 69410
rect 18946 69358 18958 69410
rect 19010 69358 19022 69410
rect 24546 69358 24558 69410
rect 24610 69358 24622 69410
rect 30146 69358 30158 69410
rect 30210 69358 30222 69410
rect 30706 69358 30718 69410
rect 30770 69358 30782 69410
rect 35186 69358 35198 69410
rect 35250 69358 35262 69410
rect 36306 69358 36318 69410
rect 36370 69358 36382 69410
rect 13806 69346 13858 69358
rect 18398 69346 18450 69358
rect 23886 69346 23938 69358
rect 34750 69346 34802 69358
rect 36094 69346 36146 69358
rect 14030 69298 14082 69310
rect 12226 69246 12238 69298
rect 12290 69246 12302 69298
rect 12562 69246 12574 69298
rect 12626 69246 12638 69298
rect 14030 69234 14082 69246
rect 14814 69298 14866 69310
rect 14814 69234 14866 69246
rect 15038 69298 15090 69310
rect 15038 69234 15090 69246
rect 15598 69298 15650 69310
rect 15598 69234 15650 69246
rect 16046 69298 16098 69310
rect 18734 69298 18786 69310
rect 16370 69246 16382 69298
rect 16434 69246 16446 69298
rect 17938 69246 17950 69298
rect 18002 69246 18014 69298
rect 18498 69246 18510 69298
rect 18562 69246 18574 69298
rect 16046 69234 16098 69246
rect 18734 69234 18786 69246
rect 27918 69298 27970 69310
rect 27918 69234 27970 69246
rect 28366 69298 28418 69310
rect 28366 69234 28418 69246
rect 35982 69298 36034 69310
rect 35982 69234 36034 69246
rect 5742 69186 5794 69198
rect 5742 69122 5794 69134
rect 6190 69186 6242 69198
rect 11230 69186 11282 69198
rect 9874 69134 9886 69186
rect 9938 69134 9950 69186
rect 6190 69122 6242 69134
rect 11230 69122 11282 69134
rect 13582 69186 13634 69198
rect 13582 69122 13634 69134
rect 15486 69186 15538 69198
rect 15486 69122 15538 69134
rect 15822 69186 15874 69198
rect 15822 69122 15874 69134
rect 19406 69186 19458 69198
rect 19406 69122 19458 69134
rect 19742 69186 19794 69198
rect 27806 69186 27858 69198
rect 34302 69186 34354 69198
rect 27010 69134 27022 69186
rect 27074 69134 27086 69186
rect 33170 69134 33182 69186
rect 33234 69134 33246 69186
rect 19742 69122 19794 69134
rect 27806 69122 27858 69134
rect 34302 69122 34354 69134
rect 1344 69018 38640 69052
rect 1344 68966 14024 69018
rect 14076 68966 14148 69018
rect 14200 68966 14272 69018
rect 14324 68966 14396 69018
rect 14448 68966 14520 69018
rect 14572 68966 14644 69018
rect 14696 68966 14768 69018
rect 14820 68966 14892 69018
rect 14944 68966 15016 69018
rect 15068 68966 15140 69018
rect 15192 68966 34024 69018
rect 34076 68966 34148 69018
rect 34200 68966 34272 69018
rect 34324 68966 34396 69018
rect 34448 68966 34520 69018
rect 34572 68966 34644 69018
rect 34696 68966 34768 69018
rect 34820 68966 34892 69018
rect 34944 68966 35016 69018
rect 35068 68966 35140 69018
rect 35192 68966 38640 69018
rect 1344 68932 38640 68966
rect 7198 68850 7250 68862
rect 6178 68798 6190 68850
rect 6242 68798 6254 68850
rect 7198 68786 7250 68798
rect 10446 68850 10498 68862
rect 10446 68786 10498 68798
rect 11790 68850 11842 68862
rect 15934 68850 15986 68862
rect 15362 68798 15374 68850
rect 15426 68798 15438 68850
rect 11790 68786 11842 68798
rect 15934 68786 15986 68798
rect 18286 68850 18338 68862
rect 18286 68786 18338 68798
rect 19070 68850 19122 68862
rect 28814 68850 28866 68862
rect 28242 68798 28254 68850
rect 28306 68798 28318 68850
rect 19070 68786 19122 68798
rect 28814 68786 28866 68798
rect 29150 68850 29202 68862
rect 29150 68786 29202 68798
rect 30830 68850 30882 68862
rect 30830 68786 30882 68798
rect 35646 68850 35698 68862
rect 35646 68786 35698 68798
rect 35982 68850 36034 68862
rect 35982 68786 36034 68798
rect 1710 68738 1762 68750
rect 1710 68674 1762 68686
rect 11678 68738 11730 68750
rect 11678 68674 11730 68686
rect 11902 68738 11954 68750
rect 11902 68674 11954 68686
rect 19742 68738 19794 68750
rect 19742 68674 19794 68686
rect 19966 68738 20018 68750
rect 19966 68674 20018 68686
rect 12238 68626 12290 68638
rect 16494 68626 16546 68638
rect 3266 68574 3278 68626
rect 3330 68574 3342 68626
rect 3714 68574 3726 68626
rect 3778 68574 3790 68626
rect 12898 68574 12910 68626
rect 12962 68574 12974 68626
rect 12238 68562 12290 68574
rect 16494 68562 16546 68574
rect 17502 68626 17554 68638
rect 17502 68562 17554 68574
rect 17726 68626 17778 68638
rect 17726 68562 17778 68574
rect 18174 68626 18226 68638
rect 18174 68562 18226 68574
rect 18398 68626 18450 68638
rect 18398 68562 18450 68574
rect 18734 68626 18786 68638
rect 18734 68562 18786 68574
rect 19182 68626 19234 68638
rect 19182 68562 19234 68574
rect 19406 68626 19458 68638
rect 19406 68562 19458 68574
rect 20638 68626 20690 68638
rect 20638 68562 20690 68574
rect 23774 68626 23826 68638
rect 23774 68562 23826 68574
rect 23998 68626 24050 68638
rect 23998 68562 24050 68574
rect 24222 68626 24274 68638
rect 24222 68562 24274 68574
rect 24446 68626 24498 68638
rect 24446 68562 24498 68574
rect 24670 68626 24722 68638
rect 24670 68562 24722 68574
rect 25342 68626 25394 68638
rect 31390 68626 31442 68638
rect 25666 68574 25678 68626
rect 25730 68574 25742 68626
rect 31042 68574 31054 68626
rect 31106 68574 31118 68626
rect 25342 68562 25394 68574
rect 31390 68562 31442 68574
rect 35534 68626 35586 68638
rect 35534 68562 35586 68574
rect 35758 68626 35810 68638
rect 35758 68562 35810 68574
rect 7646 68514 7698 68526
rect 7646 68450 7698 68462
rect 9998 68514 10050 68526
rect 9998 68450 10050 68462
rect 10894 68514 10946 68526
rect 10894 68450 10946 68462
rect 11454 68514 11506 68526
rect 11454 68450 11506 68462
rect 16718 68514 16770 68526
rect 16718 68450 16770 68462
rect 17950 68514 18002 68526
rect 30382 68514 30434 68526
rect 20066 68462 20078 68514
rect 20130 68462 20142 68514
rect 17950 68450 18002 68462
rect 30382 68450 30434 68462
rect 6862 68402 6914 68414
rect 20750 68402 20802 68414
rect 16146 68350 16158 68402
rect 16210 68350 16222 68402
rect 6862 68338 6914 68350
rect 20750 68338 20802 68350
rect 30718 68402 30770 68414
rect 30718 68338 30770 68350
rect 1344 68234 38640 68268
rect 1344 68182 4024 68234
rect 4076 68182 4148 68234
rect 4200 68182 4272 68234
rect 4324 68182 4396 68234
rect 4448 68182 4520 68234
rect 4572 68182 4644 68234
rect 4696 68182 4768 68234
rect 4820 68182 4892 68234
rect 4944 68182 5016 68234
rect 5068 68182 5140 68234
rect 5192 68182 24024 68234
rect 24076 68182 24148 68234
rect 24200 68182 24272 68234
rect 24324 68182 24396 68234
rect 24448 68182 24520 68234
rect 24572 68182 24644 68234
rect 24696 68182 24768 68234
rect 24820 68182 24892 68234
rect 24944 68182 25016 68234
rect 25068 68182 25140 68234
rect 25192 68182 38640 68234
rect 1344 68148 38640 68182
rect 8318 68066 8370 68078
rect 21422 68066 21474 68078
rect 31838 68066 31890 68078
rect 8530 68014 8542 68066
rect 8594 68063 8606 68066
rect 8754 68063 8766 68066
rect 8594 68017 8766 68063
rect 8594 68014 8606 68017
rect 8754 68014 8766 68017
rect 8818 68014 8830 68066
rect 26674 68014 26686 68066
rect 26738 68014 26750 68066
rect 8318 68002 8370 68014
rect 21422 68002 21474 68014
rect 31838 68002 31890 68014
rect 8766 67954 8818 67966
rect 27582 67954 27634 67966
rect 34974 67954 35026 67966
rect 7970 67902 7982 67954
rect 8034 67902 8046 67954
rect 14802 67902 14814 67954
rect 14866 67902 14878 67954
rect 26786 67902 26798 67954
rect 26850 67902 26862 67954
rect 29810 67902 29822 67954
rect 29874 67902 29886 67954
rect 8766 67890 8818 67902
rect 27582 67890 27634 67902
rect 34974 67890 35026 67902
rect 35422 67954 35474 67966
rect 35422 67890 35474 67902
rect 3054 67842 3106 67854
rect 3054 67778 3106 67790
rect 4174 67842 4226 67854
rect 14478 67842 14530 67854
rect 17390 67842 17442 67854
rect 4946 67790 4958 67842
rect 5010 67790 5022 67842
rect 15250 67790 15262 67842
rect 15314 67790 15326 67842
rect 4174 67778 4226 67790
rect 14478 67778 14530 67790
rect 17390 67778 17442 67790
rect 20638 67842 20690 67854
rect 25118 67842 25170 67854
rect 31390 67842 31442 67854
rect 24434 67790 24446 67842
rect 24498 67790 24510 67842
rect 25554 67790 25566 67842
rect 25618 67790 25630 67842
rect 26002 67790 26014 67842
rect 26066 67790 26078 67842
rect 26450 67790 26462 67842
rect 26514 67790 26526 67842
rect 31154 67790 31166 67842
rect 31218 67790 31230 67842
rect 20638 67778 20690 67790
rect 25118 67778 25170 67790
rect 31390 67778 31442 67790
rect 32174 67842 32226 67854
rect 32174 67778 32226 67790
rect 35646 67842 35698 67854
rect 37102 67842 37154 67854
rect 35858 67790 35870 67842
rect 35922 67790 35934 67842
rect 37314 67790 37326 67842
rect 37378 67790 37390 67842
rect 35646 67778 35698 67790
rect 37102 67778 37154 67790
rect 5854 67730 5906 67742
rect 4722 67678 4734 67730
rect 4786 67678 4798 67730
rect 5854 67666 5906 67678
rect 5966 67730 6018 67742
rect 5966 67666 6018 67678
rect 6302 67730 6354 67742
rect 6302 67666 6354 67678
rect 14030 67730 14082 67742
rect 14030 67666 14082 67678
rect 14254 67730 14306 67742
rect 14254 67666 14306 67678
rect 16494 67730 16546 67742
rect 16494 67666 16546 67678
rect 17950 67730 18002 67742
rect 17950 67666 18002 67678
rect 22206 67730 22258 67742
rect 22206 67666 22258 67678
rect 29374 67730 29426 67742
rect 29374 67666 29426 67678
rect 30158 67730 30210 67742
rect 30158 67666 30210 67678
rect 30494 67730 30546 67742
rect 30494 67666 30546 67678
rect 32398 67730 32450 67742
rect 32398 67666 32450 67678
rect 35310 67730 35362 67742
rect 35310 67666 35362 67678
rect 36990 67730 37042 67742
rect 36990 67666 37042 67678
rect 1710 67618 1762 67630
rect 1710 67554 1762 67566
rect 3502 67618 3554 67630
rect 3502 67554 3554 67566
rect 3838 67618 3890 67630
rect 3838 67554 3890 67566
rect 5630 67618 5682 67630
rect 5630 67554 5682 67566
rect 6414 67618 6466 67630
rect 6414 67554 6466 67566
rect 6638 67618 6690 67630
rect 6638 67554 6690 67566
rect 6974 67618 7026 67630
rect 6974 67554 7026 67566
rect 7758 67618 7810 67630
rect 7758 67554 7810 67566
rect 8094 67618 8146 67630
rect 8094 67554 8146 67566
rect 9438 67618 9490 67630
rect 9438 67554 9490 67566
rect 9886 67618 9938 67630
rect 9886 67554 9938 67566
rect 11230 67618 11282 67630
rect 11230 67554 11282 67566
rect 14702 67618 14754 67630
rect 14702 67554 14754 67566
rect 14814 67618 14866 67630
rect 19630 67618 19682 67630
rect 17602 67566 17614 67618
rect 17666 67566 17678 67618
rect 14814 67554 14866 67566
rect 19630 67554 19682 67566
rect 19966 67618 20018 67630
rect 19966 67554 20018 67566
rect 20078 67618 20130 67630
rect 20078 67554 20130 67566
rect 20190 67618 20242 67630
rect 20190 67554 20242 67566
rect 29486 67618 29538 67630
rect 29486 67554 29538 67566
rect 29934 67618 29986 67630
rect 29934 67554 29986 67566
rect 32958 67618 33010 67630
rect 32958 67554 33010 67566
rect 1344 67450 38640 67484
rect 1344 67398 14024 67450
rect 14076 67398 14148 67450
rect 14200 67398 14272 67450
rect 14324 67398 14396 67450
rect 14448 67398 14520 67450
rect 14572 67398 14644 67450
rect 14696 67398 14768 67450
rect 14820 67398 14892 67450
rect 14944 67398 15016 67450
rect 15068 67398 15140 67450
rect 15192 67398 34024 67450
rect 34076 67398 34148 67450
rect 34200 67398 34272 67450
rect 34324 67398 34396 67450
rect 34448 67398 34520 67450
rect 34572 67398 34644 67450
rect 34696 67398 34768 67450
rect 34820 67398 34892 67450
rect 34944 67398 35016 67450
rect 35068 67398 35140 67450
rect 35192 67398 38640 67450
rect 1344 67364 38640 67398
rect 19854 67282 19906 67294
rect 26126 67282 26178 67294
rect 37662 67282 37714 67294
rect 6066 67230 6078 67282
rect 6130 67230 6142 67282
rect 12562 67230 12574 67282
rect 12626 67230 12638 67282
rect 15698 67230 15710 67282
rect 15762 67230 15774 67282
rect 18050 67230 18062 67282
rect 18114 67230 18126 67282
rect 23874 67230 23886 67282
rect 23938 67230 23950 67282
rect 31826 67230 31838 67282
rect 31890 67230 31902 67282
rect 19854 67218 19906 67230
rect 26126 67218 26178 67230
rect 37662 67218 37714 67230
rect 13470 67170 13522 67182
rect 3938 67118 3950 67170
rect 4002 67118 4014 67170
rect 4498 67118 4510 67170
rect 4562 67118 4574 67170
rect 13470 67106 13522 67118
rect 13918 67170 13970 67182
rect 25454 67170 25506 67182
rect 15474 67118 15486 67170
rect 15538 67118 15550 67170
rect 17602 67118 17614 67170
rect 17666 67118 17678 67170
rect 17938 67118 17950 67170
rect 18002 67118 18014 67170
rect 13918 67106 13970 67118
rect 25454 67106 25506 67118
rect 26014 67170 26066 67182
rect 26014 67106 26066 67118
rect 33182 67170 33234 67182
rect 33182 67106 33234 67118
rect 33294 67170 33346 67182
rect 33294 67106 33346 67118
rect 36878 67170 36930 67182
rect 36878 67106 36930 67118
rect 3726 67058 3778 67070
rect 9102 67058 9154 67070
rect 8418 67006 8430 67058
rect 8482 67006 8494 67058
rect 3726 66994 3778 67006
rect 9102 66994 9154 67006
rect 9662 67058 9714 67070
rect 18958 67058 19010 67070
rect 10098 67006 10110 67058
rect 10162 67006 10174 67058
rect 15250 67006 15262 67058
rect 15314 67006 15326 67058
rect 16258 67006 16270 67058
rect 16322 67006 16334 67058
rect 16706 67006 16718 67058
rect 16770 67006 16782 67058
rect 17378 67006 17390 67058
rect 17442 67006 17454 67058
rect 9662 66994 9714 67006
rect 18958 66994 19010 67006
rect 19070 67058 19122 67070
rect 19070 66994 19122 67006
rect 19182 67058 19234 67070
rect 19182 66994 19234 67006
rect 19630 67058 19682 67070
rect 19630 66994 19682 67006
rect 20974 67058 21026 67070
rect 28926 67058 28978 67070
rect 33966 67058 34018 67070
rect 21410 67006 21422 67058
rect 21474 67006 21486 67058
rect 29250 67006 29262 67058
rect 29314 67006 29326 67058
rect 34514 67006 34526 67058
rect 34578 67006 34590 67058
rect 20974 66994 21026 67006
rect 28926 66994 28978 67006
rect 33966 66994 34018 67006
rect 5406 66946 5458 66958
rect 5406 66882 5458 66894
rect 14926 66946 14978 66958
rect 14926 66882 14978 66894
rect 20190 66946 20242 66958
rect 20190 66882 20242 66894
rect 25230 66946 25282 66958
rect 26238 66946 26290 66958
rect 25554 66894 25566 66946
rect 25618 66894 25630 66946
rect 25230 66882 25282 66894
rect 26238 66882 26290 66894
rect 26686 66946 26738 66958
rect 26686 66882 26738 66894
rect 33742 66946 33794 66958
rect 33742 66882 33794 66894
rect 3390 66834 3442 66846
rect 3390 66770 3442 66782
rect 13134 66834 13186 66846
rect 13134 66770 13186 66782
rect 24446 66834 24498 66846
rect 24446 66770 24498 66782
rect 32398 66834 32450 66846
rect 32398 66770 32450 66782
rect 33182 66834 33234 66846
rect 33182 66770 33234 66782
rect 1344 66666 38640 66700
rect 1344 66614 4024 66666
rect 4076 66614 4148 66666
rect 4200 66614 4272 66666
rect 4324 66614 4396 66666
rect 4448 66614 4520 66666
rect 4572 66614 4644 66666
rect 4696 66614 4768 66666
rect 4820 66614 4892 66666
rect 4944 66614 5016 66666
rect 5068 66614 5140 66666
rect 5192 66614 24024 66666
rect 24076 66614 24148 66666
rect 24200 66614 24272 66666
rect 24324 66614 24396 66666
rect 24448 66614 24520 66666
rect 24572 66614 24644 66666
rect 24696 66614 24768 66666
rect 24820 66614 24892 66666
rect 24944 66614 25016 66666
rect 25068 66614 25140 66666
rect 25192 66614 38640 66666
rect 1344 66580 38640 66614
rect 6750 66498 6802 66510
rect 6750 66434 6802 66446
rect 7310 66498 7362 66510
rect 7310 66434 7362 66446
rect 7534 66498 7586 66510
rect 10670 66498 10722 66510
rect 8754 66446 8766 66498
rect 8818 66446 8830 66498
rect 7534 66434 7586 66446
rect 10670 66434 10722 66446
rect 11006 66498 11058 66510
rect 20638 66498 20690 66510
rect 19618 66446 19630 66498
rect 19682 66446 19694 66498
rect 11006 66434 11058 66446
rect 20638 66434 20690 66446
rect 21422 66498 21474 66510
rect 21422 66434 21474 66446
rect 21758 66498 21810 66510
rect 21758 66434 21810 66446
rect 37326 66498 37378 66510
rect 37326 66434 37378 66446
rect 8430 66386 8482 66398
rect 8430 66322 8482 66334
rect 9214 66386 9266 66398
rect 9214 66322 9266 66334
rect 10222 66386 10274 66398
rect 16270 66386 16322 66398
rect 25566 66386 25618 66398
rect 37550 66386 37602 66398
rect 15922 66334 15934 66386
rect 15986 66334 15998 66386
rect 19170 66334 19182 66386
rect 19234 66334 19246 66386
rect 36978 66334 36990 66386
rect 37042 66334 37054 66386
rect 10222 66322 10274 66334
rect 16270 66322 16322 66334
rect 25566 66322 25618 66334
rect 37550 66322 37602 66334
rect 6414 66274 6466 66286
rect 4946 66222 4958 66274
rect 5010 66222 5022 66274
rect 6414 66210 6466 66222
rect 6974 66274 7026 66286
rect 6974 66210 7026 66222
rect 8206 66274 8258 66286
rect 8206 66210 8258 66222
rect 17166 66274 17218 66286
rect 29038 66274 29090 66286
rect 19058 66222 19070 66274
rect 19122 66222 19134 66274
rect 29586 66222 29598 66274
rect 29650 66222 29662 66274
rect 17166 66210 17218 66222
rect 29038 66210 29090 66222
rect 2158 66162 2210 66174
rect 2158 66098 2210 66110
rect 4510 66162 4562 66174
rect 18510 66162 18562 66174
rect 11218 66110 11230 66162
rect 11282 66110 11294 66162
rect 11666 66110 11678 66162
rect 11730 66110 11742 66162
rect 4510 66098 4562 66110
rect 18510 66098 18562 66110
rect 20638 66162 20690 66174
rect 20638 66098 20690 66110
rect 20750 66162 20802 66174
rect 31950 66162 32002 66174
rect 21970 66110 21982 66162
rect 22034 66110 22046 66162
rect 22530 66110 22542 66162
rect 22594 66110 22606 66162
rect 20750 66098 20802 66110
rect 31950 66098 32002 66110
rect 36094 66162 36146 66174
rect 36094 66098 36146 66110
rect 1710 66050 1762 66062
rect 1710 65986 1762 65998
rect 4062 66050 4114 66062
rect 4062 65986 4114 65998
rect 4398 66050 4450 66062
rect 4398 65986 4450 65998
rect 4622 66050 4674 66062
rect 4622 65986 4674 65998
rect 5742 66050 5794 66062
rect 5742 65986 5794 65998
rect 7646 66050 7698 66062
rect 7646 65986 7698 65998
rect 9774 66050 9826 66062
rect 9774 65986 9826 65998
rect 17614 66050 17666 66062
rect 17614 65986 17666 65998
rect 18062 66050 18114 66062
rect 18062 65986 18114 65998
rect 24558 66050 24610 66062
rect 24558 65986 24610 65998
rect 25006 66050 25058 66062
rect 25006 65986 25058 65998
rect 25902 66050 25954 66062
rect 25902 65986 25954 65998
rect 26350 66050 26402 66062
rect 26350 65986 26402 65998
rect 28590 66050 28642 66062
rect 28590 65986 28642 65998
rect 32734 66050 32786 66062
rect 32734 65986 32786 65998
rect 36206 66050 36258 66062
rect 36206 65986 36258 65998
rect 36318 66050 36370 66062
rect 36318 65986 36370 65998
rect 1344 65882 38640 65916
rect 1344 65830 14024 65882
rect 14076 65830 14148 65882
rect 14200 65830 14272 65882
rect 14324 65830 14396 65882
rect 14448 65830 14520 65882
rect 14572 65830 14644 65882
rect 14696 65830 14768 65882
rect 14820 65830 14892 65882
rect 14944 65830 15016 65882
rect 15068 65830 15140 65882
rect 15192 65830 34024 65882
rect 34076 65830 34148 65882
rect 34200 65830 34272 65882
rect 34324 65830 34396 65882
rect 34448 65830 34520 65882
rect 34572 65830 34644 65882
rect 34696 65830 34768 65882
rect 34820 65830 34892 65882
rect 34944 65830 35016 65882
rect 35068 65830 35140 65882
rect 35192 65830 38640 65882
rect 1344 65796 38640 65830
rect 7870 65714 7922 65726
rect 4722 65662 4734 65714
rect 4786 65662 4798 65714
rect 7870 65650 7922 65662
rect 13246 65714 13298 65726
rect 13246 65650 13298 65662
rect 18734 65714 18786 65726
rect 33742 65714 33794 65726
rect 20962 65662 20974 65714
rect 21026 65662 21038 65714
rect 28354 65662 28366 65714
rect 28418 65662 28430 65714
rect 36866 65662 36878 65714
rect 36930 65662 36942 65714
rect 18734 65650 18786 65662
rect 33742 65650 33794 65662
rect 14030 65602 14082 65614
rect 14030 65538 14082 65550
rect 19070 65602 19122 65614
rect 19070 65538 19122 65550
rect 1822 65490 1874 65502
rect 5294 65490 5346 65502
rect 2258 65438 2270 65490
rect 2322 65438 2334 65490
rect 1822 65426 1874 65438
rect 5294 65426 5346 65438
rect 5630 65490 5682 65502
rect 5630 65426 5682 65438
rect 6190 65490 6242 65502
rect 6190 65426 6242 65438
rect 9998 65490 10050 65502
rect 9998 65426 10050 65438
rect 10670 65490 10722 65502
rect 19182 65490 19234 65502
rect 13570 65438 13582 65490
rect 13634 65438 13646 65490
rect 13794 65438 13806 65490
rect 13858 65438 13870 65490
rect 10670 65426 10722 65438
rect 19182 65426 19234 65438
rect 19630 65490 19682 65502
rect 19630 65426 19682 65438
rect 20526 65490 20578 65502
rect 21310 65490 21362 65502
rect 20850 65438 20862 65490
rect 20914 65438 20926 65490
rect 20526 65426 20578 65438
rect 21310 65426 21362 65438
rect 21534 65490 21586 65502
rect 21534 65426 21586 65438
rect 25342 65490 25394 65502
rect 29374 65490 29426 65502
rect 26002 65438 26014 65490
rect 26066 65438 26078 65490
rect 25342 65426 25394 65438
rect 29374 65426 29426 65438
rect 30830 65490 30882 65502
rect 31502 65490 31554 65502
rect 31266 65438 31278 65490
rect 31330 65438 31342 65490
rect 30830 65426 30882 65438
rect 31502 65426 31554 65438
rect 31614 65490 31666 65502
rect 31614 65426 31666 65438
rect 31838 65490 31890 65502
rect 31838 65426 31890 65438
rect 33966 65490 34018 65502
rect 37662 65490 37714 65502
rect 34626 65438 34638 65490
rect 34690 65438 34702 65490
rect 33966 65426 34018 65438
rect 37662 65426 37714 65438
rect 12798 65378 12850 65390
rect 12798 65314 12850 65326
rect 14478 65378 14530 65390
rect 14478 65314 14530 65326
rect 17838 65378 17890 65390
rect 17838 65314 17890 65326
rect 18286 65378 18338 65390
rect 18286 65314 18338 65326
rect 19742 65378 19794 65390
rect 19742 65314 19794 65326
rect 21982 65378 22034 65390
rect 21982 65314 22034 65326
rect 14142 65266 14194 65278
rect 14142 65202 14194 65214
rect 19966 65266 20018 65278
rect 19966 65202 20018 65214
rect 20190 65266 20242 65278
rect 20190 65202 20242 65214
rect 20302 65266 20354 65278
rect 20302 65202 20354 65214
rect 21086 65266 21138 65278
rect 21086 65202 21138 65214
rect 29038 65266 29090 65278
rect 29038 65202 29090 65214
rect 1344 65098 38640 65132
rect 1344 65046 4024 65098
rect 4076 65046 4148 65098
rect 4200 65046 4272 65098
rect 4324 65046 4396 65098
rect 4448 65046 4520 65098
rect 4572 65046 4644 65098
rect 4696 65046 4768 65098
rect 4820 65046 4892 65098
rect 4944 65046 5016 65098
rect 5068 65046 5140 65098
rect 5192 65046 24024 65098
rect 24076 65046 24148 65098
rect 24200 65046 24272 65098
rect 24324 65046 24396 65098
rect 24448 65046 24520 65098
rect 24572 65046 24644 65098
rect 24696 65046 24768 65098
rect 24820 65046 24892 65098
rect 24944 65046 25016 65098
rect 25068 65046 25140 65098
rect 25192 65046 38640 65098
rect 1344 65012 38640 65046
rect 3838 64930 3890 64942
rect 11342 64930 11394 64942
rect 35534 64930 35586 64942
rect 10098 64878 10110 64930
rect 10162 64878 10174 64930
rect 16146 64878 16158 64930
rect 16210 64878 16222 64930
rect 3838 64866 3890 64878
rect 11342 64866 11394 64878
rect 35534 64866 35586 64878
rect 35870 64930 35922 64942
rect 37326 64930 37378 64942
rect 36978 64878 36990 64930
rect 37042 64878 37054 64930
rect 35870 64866 35922 64878
rect 37326 64866 37378 64878
rect 10446 64818 10498 64830
rect 8530 64766 8542 64818
rect 8594 64766 8606 64818
rect 10446 64754 10498 64766
rect 10670 64818 10722 64830
rect 11790 64818 11842 64830
rect 17166 64818 17218 64830
rect 18734 64818 18786 64830
rect 10994 64766 11006 64818
rect 11058 64766 11070 64818
rect 15474 64766 15486 64818
rect 15538 64766 15550 64818
rect 18162 64766 18174 64818
rect 18226 64766 18238 64818
rect 10670 64754 10722 64766
rect 11790 64754 11842 64766
rect 17166 64754 17218 64766
rect 18734 64754 18786 64766
rect 20302 64818 20354 64830
rect 20302 64754 20354 64766
rect 29262 64818 29314 64830
rect 29262 64754 29314 64766
rect 35198 64818 35250 64830
rect 35198 64754 35250 64766
rect 37550 64818 37602 64830
rect 37550 64754 37602 64766
rect 13918 64706 13970 64718
rect 7746 64654 7758 64706
rect 7810 64654 7822 64706
rect 13918 64642 13970 64654
rect 14030 64706 14082 64718
rect 14030 64642 14082 64654
rect 14814 64706 14866 64718
rect 16046 64706 16098 64718
rect 18958 64706 19010 64718
rect 15586 64654 15598 64706
rect 15650 64654 15662 64706
rect 18274 64654 18286 64706
rect 18338 64654 18350 64706
rect 14814 64642 14866 64654
rect 16046 64642 16098 64654
rect 18958 64642 19010 64654
rect 35646 64706 35698 64718
rect 36082 64654 36094 64706
rect 36146 64654 36158 64706
rect 35646 64642 35698 64654
rect 2830 64594 2882 64606
rect 2830 64530 2882 64542
rect 3166 64594 3218 64606
rect 3166 64530 3218 64542
rect 3726 64594 3778 64606
rect 3726 64530 3778 64542
rect 11118 64594 11170 64606
rect 12910 64594 12962 64606
rect 12562 64542 12574 64594
rect 12626 64542 12638 64594
rect 11118 64530 11170 64542
rect 12910 64530 12962 64542
rect 13470 64594 13522 64606
rect 13470 64530 13522 64542
rect 14478 64594 14530 64606
rect 14478 64530 14530 64542
rect 14590 64594 14642 64606
rect 14590 64530 14642 64542
rect 19518 64594 19570 64606
rect 19518 64530 19570 64542
rect 1710 64482 1762 64494
rect 1710 64418 1762 64430
rect 2606 64482 2658 64494
rect 2606 64418 2658 64430
rect 5742 64482 5794 64494
rect 5742 64418 5794 64430
rect 12238 64482 12290 64494
rect 12238 64418 12290 64430
rect 13694 64482 13746 64494
rect 13694 64418 13746 64430
rect 13806 64482 13858 64494
rect 13806 64418 13858 64430
rect 16718 64482 16770 64494
rect 16718 64418 16770 64430
rect 17614 64482 17666 64494
rect 17614 64418 17666 64430
rect 19294 64482 19346 64494
rect 19294 64418 19346 64430
rect 19630 64482 19682 64494
rect 19630 64418 19682 64430
rect 29822 64482 29874 64494
rect 29822 64418 29874 64430
rect 1344 64314 38640 64348
rect 1344 64262 14024 64314
rect 14076 64262 14148 64314
rect 14200 64262 14272 64314
rect 14324 64262 14396 64314
rect 14448 64262 14520 64314
rect 14572 64262 14644 64314
rect 14696 64262 14768 64314
rect 14820 64262 14892 64314
rect 14944 64262 15016 64314
rect 15068 64262 15140 64314
rect 15192 64262 34024 64314
rect 34076 64262 34148 64314
rect 34200 64262 34272 64314
rect 34324 64262 34396 64314
rect 34448 64262 34520 64314
rect 34572 64262 34644 64314
rect 34696 64262 34768 64314
rect 34820 64262 34892 64314
rect 34944 64262 35016 64314
rect 35068 64262 35140 64314
rect 35192 64262 38640 64314
rect 1344 64228 38640 64262
rect 5742 64146 5794 64158
rect 4834 64094 4846 64146
rect 4898 64094 4910 64146
rect 5742 64082 5794 64094
rect 6190 64146 6242 64158
rect 6190 64082 6242 64094
rect 8990 64146 9042 64158
rect 17278 64146 17330 64158
rect 30270 64146 30322 64158
rect 12450 64094 12462 64146
rect 12514 64094 12526 64146
rect 16034 64094 16046 64146
rect 16098 64094 16110 64146
rect 28242 64094 28254 64146
rect 28306 64094 28318 64146
rect 8990 64082 9042 64094
rect 17278 64082 17330 64094
rect 30270 64082 30322 64094
rect 14690 63982 14702 64034
rect 14754 63982 14766 64034
rect 16146 63982 16158 64034
rect 16210 63982 16222 64034
rect 29138 63982 29150 64034
rect 29202 63982 29214 64034
rect 1934 63922 1986 63934
rect 5406 63922 5458 63934
rect 2370 63870 2382 63922
rect 2434 63870 2446 63922
rect 1934 63858 1986 63870
rect 5406 63858 5458 63870
rect 9662 63922 9714 63934
rect 13134 63922 13186 63934
rect 20414 63922 20466 63934
rect 9986 63870 9998 63922
rect 10050 63870 10062 63922
rect 15250 63870 15262 63922
rect 15314 63870 15326 63922
rect 15586 63870 15598 63922
rect 15650 63870 15662 63922
rect 17938 63870 17950 63922
rect 18002 63870 18014 63922
rect 18274 63870 18286 63922
rect 18338 63870 18350 63922
rect 19506 63870 19518 63922
rect 19570 63870 19582 63922
rect 9662 63858 9714 63870
rect 13134 63858 13186 63870
rect 20414 63858 20466 63870
rect 25342 63922 25394 63934
rect 28814 63922 28866 63934
rect 31838 63922 31890 63934
rect 25666 63870 25678 63922
rect 25730 63870 25742 63922
rect 29250 63870 29262 63922
rect 29314 63870 29326 63922
rect 25342 63858 25394 63870
rect 28814 63858 28866 63870
rect 31838 63858 31890 63870
rect 13694 63810 13746 63822
rect 13694 63746 13746 63758
rect 13918 63810 13970 63822
rect 19966 63810 20018 63822
rect 18050 63758 18062 63810
rect 18114 63758 18126 63810
rect 19618 63758 19630 63810
rect 19682 63758 19694 63810
rect 13918 63746 13970 63758
rect 19966 63746 20018 63758
rect 29934 63810 29986 63822
rect 29934 63746 29986 63758
rect 31278 63810 31330 63822
rect 31278 63746 31330 63758
rect 14242 63646 14254 63698
rect 14306 63646 14318 63698
rect 1344 63530 38640 63564
rect 1344 63478 4024 63530
rect 4076 63478 4148 63530
rect 4200 63478 4272 63530
rect 4324 63478 4396 63530
rect 4448 63478 4520 63530
rect 4572 63478 4644 63530
rect 4696 63478 4768 63530
rect 4820 63478 4892 63530
rect 4944 63478 5016 63530
rect 5068 63478 5140 63530
rect 5192 63478 24024 63530
rect 24076 63478 24148 63530
rect 24200 63478 24272 63530
rect 24324 63478 24396 63530
rect 24448 63478 24520 63530
rect 24572 63478 24644 63530
rect 24696 63478 24768 63530
rect 24820 63478 24892 63530
rect 24944 63478 25016 63530
rect 25068 63478 25140 63530
rect 25192 63478 38640 63530
rect 1344 63444 38640 63478
rect 3838 63362 3890 63374
rect 3838 63298 3890 63310
rect 7534 63362 7586 63374
rect 7534 63298 7586 63310
rect 18062 63362 18114 63374
rect 31714 63310 31726 63362
rect 31778 63310 31790 63362
rect 18062 63298 18114 63310
rect 4174 63250 4226 63262
rect 4174 63186 4226 63198
rect 5742 63250 5794 63262
rect 5742 63186 5794 63198
rect 6862 63250 6914 63262
rect 13582 63250 13634 63262
rect 24782 63250 24834 63262
rect 12338 63198 12350 63250
rect 12402 63198 12414 63250
rect 15474 63198 15486 63250
rect 15538 63198 15550 63250
rect 16818 63198 16830 63250
rect 16882 63198 16894 63250
rect 34738 63198 34750 63250
rect 34802 63198 34814 63250
rect 6862 63186 6914 63198
rect 13582 63186 13634 63198
rect 24782 63186 24834 63198
rect 6190 63138 6242 63150
rect 8542 63138 8594 63150
rect 4946 63086 4958 63138
rect 5010 63086 5022 63138
rect 7186 63086 7198 63138
rect 7250 63086 7262 63138
rect 8306 63086 8318 63138
rect 8370 63086 8382 63138
rect 6190 63074 6242 63086
rect 8542 63074 8594 63086
rect 8766 63138 8818 63150
rect 8766 63074 8818 63086
rect 9550 63138 9602 63150
rect 20302 63138 20354 63150
rect 10098 63086 10110 63138
rect 10162 63086 10174 63138
rect 14914 63086 14926 63138
rect 14978 63086 14990 63138
rect 15922 63086 15934 63138
rect 15986 63086 15998 63138
rect 16370 63086 16382 63138
rect 16434 63086 16446 63138
rect 17266 63086 17278 63138
rect 17330 63086 17342 63138
rect 20066 63086 20078 63138
rect 20130 63086 20142 63138
rect 9550 63074 9602 63086
rect 20302 63074 20354 63086
rect 20526 63138 20578 63150
rect 20526 63074 20578 63086
rect 23774 63138 23826 63150
rect 23774 63074 23826 63086
rect 24894 63138 24946 63150
rect 30494 63138 30546 63150
rect 25218 63086 25230 63138
rect 25282 63086 25294 63138
rect 24894 63074 24946 63086
rect 30494 63074 30546 63086
rect 31054 63138 31106 63150
rect 31266 63086 31278 63138
rect 31330 63086 31342 63138
rect 31054 63074 31106 63086
rect 8990 63026 9042 63038
rect 4722 62974 4734 63026
rect 4786 62974 4798 63026
rect 8990 62962 9042 62974
rect 14478 63026 14530 63038
rect 16830 63026 16882 63038
rect 15250 62974 15262 63026
rect 15314 62974 15326 63026
rect 14478 62962 14530 62974
rect 16830 62962 16882 62974
rect 18174 63026 18226 63038
rect 18174 62962 18226 62974
rect 19406 63026 19458 63038
rect 19406 62962 19458 62974
rect 19854 63026 19906 63038
rect 19854 62962 19906 62974
rect 20638 63026 20690 63038
rect 20638 62962 20690 62974
rect 20750 63026 20802 63038
rect 20750 62962 20802 62974
rect 24110 63026 24162 63038
rect 24110 62962 24162 62974
rect 24670 63026 24722 63038
rect 24670 62962 24722 62974
rect 26574 63026 26626 63038
rect 26574 62962 26626 62974
rect 27022 63026 27074 63038
rect 27022 62962 27074 62974
rect 27134 63026 27186 63038
rect 27134 62962 27186 62974
rect 30718 63026 30770 63038
rect 30718 62962 30770 62974
rect 34862 63026 34914 63038
rect 34862 62962 34914 62974
rect 35086 63026 35138 63038
rect 35086 62962 35138 62974
rect 35870 63026 35922 63038
rect 35870 62962 35922 62974
rect 1710 62914 1762 62926
rect 1710 62850 1762 62862
rect 7422 62914 7474 62926
rect 14030 62914 14082 62926
rect 7970 62862 7982 62914
rect 8034 62862 8046 62914
rect 7422 62850 7474 62862
rect 14030 62850 14082 62862
rect 17054 62914 17106 62926
rect 17054 62850 17106 62862
rect 19070 62914 19122 62926
rect 19070 62850 19122 62862
rect 19518 62914 19570 62926
rect 19518 62850 19570 62862
rect 25678 62914 25730 62926
rect 25678 62850 25730 62862
rect 26798 62914 26850 62926
rect 26798 62850 26850 62862
rect 28590 62914 28642 62926
rect 28590 62850 28642 62862
rect 29262 62914 29314 62926
rect 29262 62850 29314 62862
rect 30158 62914 30210 62926
rect 30158 62850 30210 62862
rect 33630 62914 33682 62926
rect 33630 62850 33682 62862
rect 35534 62914 35586 62926
rect 35534 62850 35586 62862
rect 35758 62914 35810 62926
rect 35758 62850 35810 62862
rect 35982 62914 36034 62926
rect 35982 62850 36034 62862
rect 1344 62746 38640 62780
rect 1344 62694 14024 62746
rect 14076 62694 14148 62746
rect 14200 62694 14272 62746
rect 14324 62694 14396 62746
rect 14448 62694 14520 62746
rect 14572 62694 14644 62746
rect 14696 62694 14768 62746
rect 14820 62694 14892 62746
rect 14944 62694 15016 62746
rect 15068 62694 15140 62746
rect 15192 62694 34024 62746
rect 34076 62694 34148 62746
rect 34200 62694 34272 62746
rect 34324 62694 34396 62746
rect 34448 62694 34520 62746
rect 34572 62694 34644 62746
rect 34696 62694 34768 62746
rect 34820 62694 34892 62746
rect 34944 62694 35016 62746
rect 35068 62694 35140 62746
rect 35192 62694 38640 62746
rect 1344 62660 38640 62694
rect 8878 62578 8930 62590
rect 8306 62526 8318 62578
rect 8370 62526 8382 62578
rect 8878 62514 8930 62526
rect 9998 62578 10050 62590
rect 14366 62578 14418 62590
rect 13570 62526 13582 62578
rect 13634 62526 13646 62578
rect 9998 62514 10050 62526
rect 14366 62514 14418 62526
rect 16270 62578 16322 62590
rect 16270 62514 16322 62526
rect 16718 62578 16770 62590
rect 16718 62514 16770 62526
rect 20190 62578 20242 62590
rect 29598 62578 29650 62590
rect 37550 62578 37602 62590
rect 24098 62526 24110 62578
rect 24162 62526 24174 62578
rect 28242 62526 28254 62578
rect 28306 62526 28318 62578
rect 36754 62526 36766 62578
rect 36818 62526 36830 62578
rect 20190 62514 20242 62526
rect 29598 62514 29650 62526
rect 37550 62514 37602 62526
rect 1710 62466 1762 62478
rect 1710 62402 1762 62414
rect 4846 62466 4898 62478
rect 4846 62402 4898 62414
rect 9886 62466 9938 62478
rect 9886 62402 9938 62414
rect 10446 62466 10498 62478
rect 10446 62402 10498 62414
rect 15822 62466 15874 62478
rect 15822 62402 15874 62414
rect 19294 62466 19346 62478
rect 19294 62402 19346 62414
rect 24670 62466 24722 62478
rect 24670 62402 24722 62414
rect 30942 62466 30994 62478
rect 30942 62402 30994 62414
rect 31054 62466 31106 62478
rect 31054 62402 31106 62414
rect 4398 62354 4450 62366
rect 4398 62290 4450 62302
rect 4734 62354 4786 62366
rect 10222 62354 10274 62366
rect 5282 62302 5294 62354
rect 5346 62302 5358 62354
rect 5730 62302 5742 62354
rect 5794 62302 5806 62354
rect 4734 62290 4786 62302
rect 10222 62290 10274 62302
rect 10894 62354 10946 62366
rect 14814 62354 14866 62366
rect 11218 62302 11230 62354
rect 11282 62302 11294 62354
rect 10894 62290 10946 62302
rect 14814 62290 14866 62302
rect 14926 62354 14978 62366
rect 14926 62290 14978 62302
rect 15374 62354 15426 62366
rect 19742 62354 19794 62366
rect 16034 62302 16046 62354
rect 16098 62302 16110 62354
rect 15374 62290 15426 62302
rect 19742 62290 19794 62302
rect 19854 62354 19906 62366
rect 19854 62290 19906 62302
rect 20078 62354 20130 62366
rect 20078 62290 20130 62302
rect 20302 62354 20354 62366
rect 20302 62290 20354 62302
rect 20974 62354 21026 62366
rect 25342 62354 25394 62366
rect 29150 62354 29202 62366
rect 21522 62302 21534 62354
rect 21586 62302 21598 62354
rect 25778 62302 25790 62354
rect 25842 62302 25854 62354
rect 20974 62290 21026 62302
rect 25342 62290 25394 62302
rect 29150 62290 29202 62302
rect 30046 62354 30098 62366
rect 30046 62290 30098 62302
rect 30718 62354 30770 62366
rect 30718 62290 30770 62302
rect 33406 62354 33458 62366
rect 33406 62290 33458 62302
rect 33854 62354 33906 62366
rect 34402 62302 34414 62354
rect 34466 62302 34478 62354
rect 33854 62290 33906 62302
rect 14590 62242 14642 62254
rect 14590 62178 14642 62190
rect 28814 62242 28866 62254
rect 28814 62178 28866 62190
rect 4846 62130 4898 62142
rect 4846 62066 4898 62078
rect 15598 62130 15650 62142
rect 15598 62066 15650 62078
rect 15934 62130 15986 62142
rect 15934 62066 15986 62078
rect 1344 61962 38640 61996
rect 1344 61910 4024 61962
rect 4076 61910 4148 61962
rect 4200 61910 4272 61962
rect 4324 61910 4396 61962
rect 4448 61910 4520 61962
rect 4572 61910 4644 61962
rect 4696 61910 4768 61962
rect 4820 61910 4892 61962
rect 4944 61910 5016 61962
rect 5068 61910 5140 61962
rect 5192 61910 24024 61962
rect 24076 61910 24148 61962
rect 24200 61910 24272 61962
rect 24324 61910 24396 61962
rect 24448 61910 24520 61962
rect 24572 61910 24644 61962
rect 24696 61910 24768 61962
rect 24820 61910 24892 61962
rect 24944 61910 25016 61962
rect 25068 61910 25140 61962
rect 25192 61910 38640 61962
rect 1344 61876 38640 61910
rect 12798 61794 12850 61806
rect 12798 61730 12850 61742
rect 15598 61794 15650 61806
rect 15598 61730 15650 61742
rect 15822 61794 15874 61806
rect 15822 61730 15874 61742
rect 17166 61794 17218 61806
rect 17166 61730 17218 61742
rect 21422 61794 21474 61806
rect 21422 61730 21474 61742
rect 26014 61794 26066 61806
rect 26014 61730 26066 61742
rect 26350 61794 26402 61806
rect 36978 61742 36990 61794
rect 37042 61742 37054 61794
rect 26350 61730 26402 61742
rect 15374 61682 15426 61694
rect 6738 61630 6750 61682
rect 6802 61630 6814 61682
rect 11442 61630 11454 61682
rect 11506 61630 11518 61682
rect 14914 61630 14926 61682
rect 14978 61630 14990 61682
rect 15374 61618 15426 61630
rect 16942 61682 16994 61694
rect 16942 61618 16994 61630
rect 24222 61682 24274 61694
rect 24222 61618 24274 61630
rect 35534 61682 35586 61694
rect 35534 61618 35586 61630
rect 35982 61682 36034 61694
rect 35982 61618 36034 61630
rect 37550 61682 37602 61694
rect 37550 61618 37602 61630
rect 4062 61570 4114 61582
rect 9214 61570 9266 61582
rect 4610 61518 4622 61570
rect 4674 61518 4686 61570
rect 8194 61518 8206 61570
rect 8258 61518 8270 61570
rect 4062 61506 4114 61518
rect 9214 61506 9266 61518
rect 10334 61570 10386 61582
rect 10334 61506 10386 61518
rect 11790 61570 11842 61582
rect 11790 61506 11842 61518
rect 12014 61570 12066 61582
rect 12014 61506 12066 61518
rect 12910 61570 12962 61582
rect 20862 61570 20914 61582
rect 13570 61518 13582 61570
rect 13634 61518 13646 61570
rect 13794 61518 13806 61570
rect 13858 61518 13870 61570
rect 15026 61518 15038 61570
rect 15090 61518 15102 61570
rect 20178 61518 20190 61570
rect 20242 61518 20254 61570
rect 12910 61506 12962 61518
rect 20862 61506 20914 61518
rect 21758 61570 21810 61582
rect 21758 61506 21810 61518
rect 29374 61570 29426 61582
rect 36206 61570 36258 61582
rect 29922 61518 29934 61570
rect 29986 61518 29998 61570
rect 29374 61506 29426 61518
rect 36206 61506 36258 61518
rect 36318 61570 36370 61582
rect 36318 61506 36370 61518
rect 37326 61570 37378 61582
rect 37326 61506 37378 61518
rect 11118 61458 11170 61470
rect 4834 61406 4846 61458
rect 4898 61406 4910 61458
rect 11118 61394 11170 61406
rect 12350 61458 12402 61470
rect 24558 61458 24610 61470
rect 28478 61458 28530 61470
rect 14914 61406 14926 61458
rect 14978 61406 14990 61458
rect 21970 61406 21982 61458
rect 22034 61406 22046 61458
rect 22306 61406 22318 61458
rect 22370 61406 22382 61458
rect 25218 61406 25230 61458
rect 25282 61406 25294 61458
rect 25778 61406 25790 61458
rect 25842 61406 25854 61458
rect 12350 61394 12402 61406
rect 24558 61394 24610 61406
rect 28478 61394 28530 61406
rect 35870 61458 35922 61470
rect 35870 61394 35922 61406
rect 1710 61346 1762 61358
rect 1710 61282 1762 61294
rect 3726 61346 3778 61358
rect 3726 61282 3778 61294
rect 5742 61346 5794 61358
rect 5742 61282 5794 61294
rect 8878 61346 8930 61358
rect 8878 61282 8930 61294
rect 9102 61346 9154 61358
rect 9102 61282 9154 61294
rect 9886 61346 9938 61358
rect 9886 61282 9938 61294
rect 10782 61346 10834 61358
rect 10782 61282 10834 61294
rect 11342 61346 11394 61358
rect 11342 61282 11394 61294
rect 12126 61346 12178 61358
rect 12126 61282 12178 61294
rect 16270 61346 16322 61358
rect 28590 61346 28642 61358
rect 33070 61346 33122 61358
rect 17714 61294 17726 61346
rect 17778 61294 17790 61346
rect 32498 61294 32510 61346
rect 32562 61294 32574 61346
rect 16270 61282 16322 61294
rect 28590 61282 28642 61294
rect 33070 61282 33122 61294
rect 33406 61346 33458 61358
rect 33406 61282 33458 61294
rect 33854 61346 33906 61358
rect 33854 61282 33906 61294
rect 34414 61346 34466 61358
rect 34414 61282 34466 61294
rect 1344 61178 38640 61212
rect 1344 61126 14024 61178
rect 14076 61126 14148 61178
rect 14200 61126 14272 61178
rect 14324 61126 14396 61178
rect 14448 61126 14520 61178
rect 14572 61126 14644 61178
rect 14696 61126 14768 61178
rect 14820 61126 14892 61178
rect 14944 61126 15016 61178
rect 15068 61126 15140 61178
rect 15192 61126 34024 61178
rect 34076 61126 34148 61178
rect 34200 61126 34272 61178
rect 34324 61126 34396 61178
rect 34448 61126 34520 61178
rect 34572 61126 34644 61178
rect 34696 61126 34768 61178
rect 34820 61126 34892 61178
rect 34944 61126 35016 61178
rect 35068 61126 35140 61178
rect 35192 61126 38640 61178
rect 1344 61092 38640 61126
rect 5294 61010 5346 61022
rect 4722 60958 4734 61010
rect 4786 60958 4798 61010
rect 5294 60946 5346 60958
rect 5630 61010 5682 61022
rect 5630 60946 5682 60958
rect 13582 61010 13634 61022
rect 13582 60946 13634 60958
rect 13694 61010 13746 61022
rect 13694 60946 13746 60958
rect 21422 61010 21474 61022
rect 21422 60946 21474 60958
rect 33182 61010 33234 61022
rect 33182 60946 33234 60958
rect 34190 61010 34242 61022
rect 37762 60958 37774 61010
rect 37826 60958 37838 61010
rect 34190 60946 34242 60958
rect 7198 60898 7250 60910
rect 6626 60846 6638 60898
rect 6690 60846 6702 60898
rect 7198 60834 7250 60846
rect 7534 60898 7586 60910
rect 7534 60834 7586 60846
rect 29934 60898 29986 60910
rect 29934 60834 29986 60846
rect 30046 60898 30098 60910
rect 30046 60834 30098 60846
rect 1822 60786 1874 60798
rect 5966 60786 6018 60798
rect 7422 60786 7474 60798
rect 2258 60734 2270 60786
rect 2322 60734 2334 60786
rect 6738 60734 6750 60786
rect 6802 60734 6814 60786
rect 1822 60722 1874 60734
rect 5966 60722 6018 60734
rect 7422 60722 7474 60734
rect 7982 60786 8034 60798
rect 7982 60722 8034 60734
rect 8542 60786 8594 60798
rect 16382 60786 16434 60798
rect 30606 60786 30658 60798
rect 31502 60786 31554 60798
rect 15922 60734 15934 60786
rect 15986 60734 15998 60786
rect 27010 60734 27022 60786
rect 27074 60734 27086 60786
rect 31042 60734 31054 60786
rect 31106 60734 31118 60786
rect 8542 60722 8594 60734
rect 16382 60722 16434 60734
rect 30606 60722 30658 60734
rect 31502 60722 31554 60734
rect 31726 60786 31778 60798
rect 31726 60722 31778 60734
rect 32062 60786 32114 60798
rect 32062 60722 32114 60734
rect 32398 60786 32450 60798
rect 32398 60722 32450 60734
rect 33294 60786 33346 60798
rect 33294 60722 33346 60734
rect 34638 60786 34690 60798
rect 35298 60734 35310 60786
rect 35362 60734 35374 60786
rect 34638 60722 34690 60734
rect 8990 60674 9042 60686
rect 8990 60610 9042 60622
rect 9662 60674 9714 60686
rect 9662 60610 9714 60622
rect 10110 60674 10162 60686
rect 10110 60610 10162 60622
rect 20974 60674 21026 60686
rect 20974 60610 21026 60622
rect 25342 60674 25394 60686
rect 25342 60610 25394 60622
rect 26686 60674 26738 60686
rect 31950 60674 32002 60686
rect 28690 60622 28702 60674
rect 28754 60622 28766 60674
rect 26686 60610 26738 60622
rect 31950 60610 32002 60622
rect 33742 60674 33794 60686
rect 33742 60610 33794 60622
rect 7758 60562 7810 60574
rect 7758 60498 7810 60510
rect 13470 60562 13522 60574
rect 13470 60498 13522 60510
rect 16158 60562 16210 60574
rect 16158 60498 16210 60510
rect 16494 60562 16546 60574
rect 30046 60562 30098 60574
rect 20850 60510 20862 60562
rect 20914 60559 20926 60562
rect 21522 60559 21534 60562
rect 20914 60513 21534 60559
rect 20914 60510 20926 60513
rect 21522 60510 21534 60513
rect 21586 60510 21598 60562
rect 16494 60498 16546 60510
rect 30046 60498 30098 60510
rect 33182 60562 33234 60574
rect 33182 60498 33234 60510
rect 38334 60562 38386 60574
rect 38334 60498 38386 60510
rect 1344 60394 38640 60428
rect 1344 60342 4024 60394
rect 4076 60342 4148 60394
rect 4200 60342 4272 60394
rect 4324 60342 4396 60394
rect 4448 60342 4520 60394
rect 4572 60342 4644 60394
rect 4696 60342 4768 60394
rect 4820 60342 4892 60394
rect 4944 60342 5016 60394
rect 5068 60342 5140 60394
rect 5192 60342 24024 60394
rect 24076 60342 24148 60394
rect 24200 60342 24272 60394
rect 24324 60342 24396 60394
rect 24448 60342 24520 60394
rect 24572 60342 24644 60394
rect 24696 60342 24768 60394
rect 24820 60342 24892 60394
rect 24944 60342 25016 60394
rect 25068 60342 25140 60394
rect 25192 60342 38640 60394
rect 1344 60308 38640 60342
rect 28590 60226 28642 60238
rect 5954 60174 5966 60226
rect 6018 60223 6030 60226
rect 6178 60223 6190 60226
rect 6018 60177 6190 60223
rect 6018 60174 6030 60177
rect 6178 60174 6190 60177
rect 6242 60174 6254 60226
rect 28590 60162 28642 60174
rect 33966 60226 34018 60238
rect 36978 60174 36990 60226
rect 37042 60174 37054 60226
rect 33966 60162 34018 60174
rect 5742 60114 5794 60126
rect 5742 60050 5794 60062
rect 6190 60114 6242 60126
rect 6190 60050 6242 60062
rect 12798 60114 12850 60126
rect 12798 60050 12850 60062
rect 19630 60114 19682 60126
rect 19630 60050 19682 60062
rect 20526 60114 20578 60126
rect 29934 60114 29986 60126
rect 26002 60062 26014 60114
rect 26066 60062 26078 60114
rect 20526 60050 20578 60062
rect 29934 60050 29986 60062
rect 36318 60114 36370 60126
rect 36318 60050 36370 60062
rect 37550 60114 37602 60126
rect 37550 60050 37602 60062
rect 7086 60002 7138 60014
rect 30270 60002 30322 60014
rect 36430 60002 36482 60014
rect 23762 59950 23774 60002
rect 23826 59950 23838 60002
rect 30930 59950 30942 60002
rect 30994 59950 31006 60002
rect 7086 59938 7138 59950
rect 30270 59938 30322 59950
rect 36430 59938 36482 59950
rect 37326 60002 37378 60014
rect 37326 59938 37378 59950
rect 29598 59890 29650 59902
rect 19282 59838 19294 59890
rect 19346 59838 19358 59890
rect 29598 59826 29650 59838
rect 29822 59890 29874 59902
rect 29822 59826 29874 59838
rect 30046 59890 30098 59902
rect 30046 59826 30098 59838
rect 36206 59890 36258 59902
rect 36206 59826 36258 59838
rect 1710 59778 1762 59790
rect 1710 59714 1762 59726
rect 19070 59778 19122 59790
rect 19070 59714 19122 59726
rect 20190 59778 20242 59790
rect 20190 59714 20242 59726
rect 21534 59778 21586 59790
rect 21534 59714 21586 59726
rect 23438 59778 23490 59790
rect 23438 59714 23490 59726
rect 28030 59778 28082 59790
rect 28030 59714 28082 59726
rect 28366 59778 28418 59790
rect 28366 59714 28418 59726
rect 28478 59778 28530 59790
rect 34302 59778 34354 59790
rect 33170 59726 33182 59778
rect 33234 59726 33246 59778
rect 28478 59714 28530 59726
rect 34302 59714 34354 59726
rect 1344 59610 38640 59644
rect 1344 59558 14024 59610
rect 14076 59558 14148 59610
rect 14200 59558 14272 59610
rect 14324 59558 14396 59610
rect 14448 59558 14520 59610
rect 14572 59558 14644 59610
rect 14696 59558 14768 59610
rect 14820 59558 14892 59610
rect 14944 59558 15016 59610
rect 15068 59558 15140 59610
rect 15192 59558 34024 59610
rect 34076 59558 34148 59610
rect 34200 59558 34272 59610
rect 34324 59558 34396 59610
rect 34448 59558 34520 59610
rect 34572 59558 34644 59610
rect 34696 59558 34768 59610
rect 34820 59558 34892 59610
rect 34944 59558 35016 59610
rect 35068 59558 35140 59610
rect 35192 59558 38640 59610
rect 1344 59524 38640 59558
rect 11678 59442 11730 59454
rect 11678 59378 11730 59390
rect 18398 59442 18450 59454
rect 18398 59378 18450 59390
rect 19742 59442 19794 59454
rect 19742 59378 19794 59390
rect 19854 59442 19906 59454
rect 19854 59378 19906 59390
rect 20638 59442 20690 59454
rect 20638 59378 20690 59390
rect 20750 59442 20802 59454
rect 20750 59378 20802 59390
rect 25342 59442 25394 59454
rect 25342 59378 25394 59390
rect 30494 59442 30546 59454
rect 30494 59378 30546 59390
rect 31614 59442 31666 59454
rect 31614 59378 31666 59390
rect 31726 59442 31778 59454
rect 31726 59378 31778 59390
rect 13022 59330 13074 59342
rect 18510 59330 18562 59342
rect 15026 59278 15038 59330
rect 15090 59278 15102 59330
rect 13022 59266 13074 59278
rect 18510 59266 18562 59278
rect 21646 59330 21698 59342
rect 21646 59266 21698 59278
rect 28926 59330 28978 59342
rect 28926 59266 28978 59278
rect 31838 59330 31890 59342
rect 31838 59266 31890 59278
rect 33070 59330 33122 59342
rect 33070 59266 33122 59278
rect 33294 59330 33346 59342
rect 33294 59266 33346 59278
rect 14478 59218 14530 59230
rect 14018 59166 14030 59218
rect 14082 59166 14094 59218
rect 14478 59154 14530 59166
rect 14814 59218 14866 59230
rect 19070 59218 19122 59230
rect 15362 59166 15374 59218
rect 15426 59166 15438 59218
rect 16034 59166 16046 59218
rect 16098 59166 16110 59218
rect 18722 59166 18734 59218
rect 18786 59166 18798 59218
rect 14814 59154 14866 59166
rect 19070 59154 19122 59166
rect 19966 59218 20018 59230
rect 19966 59154 20018 59166
rect 20414 59218 20466 59230
rect 20414 59154 20466 59166
rect 20862 59218 20914 59230
rect 20862 59154 20914 59166
rect 21310 59218 21362 59230
rect 21310 59154 21362 59166
rect 21534 59218 21586 59230
rect 21534 59154 21586 59166
rect 26014 59218 26066 59230
rect 32286 59218 32338 59230
rect 26674 59166 26686 59218
rect 26738 59166 26750 59218
rect 29922 59166 29934 59218
rect 29986 59166 29998 59218
rect 31938 59166 31950 59218
rect 32002 59166 32014 59218
rect 26014 59154 26066 59166
rect 32286 59154 32338 59166
rect 11342 59106 11394 59118
rect 11342 59042 11394 59054
rect 12462 59106 12514 59118
rect 18062 59106 18114 59118
rect 13570 59054 13582 59106
rect 13634 59054 13646 59106
rect 12462 59042 12514 59054
rect 18062 59042 18114 59054
rect 19518 59106 19570 59118
rect 19518 59042 19570 59054
rect 22206 59106 22258 59118
rect 22206 59042 22258 59054
rect 25790 59106 25842 59118
rect 25790 59042 25842 59054
rect 14702 58994 14754 59006
rect 14702 58930 14754 58942
rect 21646 58994 21698 59006
rect 21646 58930 21698 58942
rect 29710 58994 29762 59006
rect 29710 58930 29762 58942
rect 33406 58994 33458 59006
rect 33406 58930 33458 58942
rect 1344 58826 38640 58860
rect 1344 58774 4024 58826
rect 4076 58774 4148 58826
rect 4200 58774 4272 58826
rect 4324 58774 4396 58826
rect 4448 58774 4520 58826
rect 4572 58774 4644 58826
rect 4696 58774 4768 58826
rect 4820 58774 4892 58826
rect 4944 58774 5016 58826
rect 5068 58774 5140 58826
rect 5192 58774 24024 58826
rect 24076 58774 24148 58826
rect 24200 58774 24272 58826
rect 24324 58774 24396 58826
rect 24448 58774 24520 58826
rect 24572 58774 24644 58826
rect 24696 58774 24768 58826
rect 24820 58774 24892 58826
rect 24944 58774 25016 58826
rect 25068 58774 25140 58826
rect 25192 58774 38640 58826
rect 1344 58740 38640 58774
rect 31278 58658 31330 58670
rect 31278 58594 31330 58606
rect 32174 58658 32226 58670
rect 32174 58594 32226 58606
rect 13582 58546 13634 58558
rect 3938 58494 3950 58546
rect 4002 58494 4014 58546
rect 13582 58482 13634 58494
rect 15262 58546 15314 58558
rect 15262 58482 15314 58494
rect 32286 58546 32338 58558
rect 32286 58482 32338 58494
rect 7870 58434 7922 58446
rect 2930 58382 2942 58434
rect 2994 58382 3006 58434
rect 7522 58382 7534 58434
rect 7586 58382 7598 58434
rect 7870 58370 7922 58382
rect 9214 58434 9266 58446
rect 17166 58434 17218 58446
rect 18510 58434 18562 58446
rect 9538 58382 9550 58434
rect 9602 58382 9614 58434
rect 14802 58382 14814 58434
rect 14866 58382 14878 58434
rect 15026 58382 15038 58434
rect 15090 58382 15102 58434
rect 17490 58382 17502 58434
rect 17554 58382 17566 58434
rect 9214 58370 9266 58382
rect 17166 58370 17218 58382
rect 18510 58370 18562 58382
rect 19070 58434 19122 58446
rect 19070 58370 19122 58382
rect 19294 58434 19346 58446
rect 19854 58434 19906 58446
rect 19506 58382 19518 58434
rect 19570 58382 19582 58434
rect 19294 58370 19346 58382
rect 19854 58370 19906 58382
rect 20414 58434 20466 58446
rect 20414 58370 20466 58382
rect 20750 58434 20802 58446
rect 20750 58370 20802 58382
rect 21310 58434 21362 58446
rect 21310 58370 21362 58382
rect 21646 58434 21698 58446
rect 27358 58434 27410 58446
rect 26674 58382 26686 58434
rect 26738 58382 26750 58434
rect 21646 58370 21698 58382
rect 27358 58370 27410 58382
rect 28142 58434 28194 58446
rect 28142 58370 28194 58382
rect 29934 58434 29986 58446
rect 29934 58370 29986 58382
rect 30270 58434 30322 58446
rect 30270 58370 30322 58382
rect 30606 58434 30658 58446
rect 34974 58434 35026 58446
rect 31602 58382 31614 58434
rect 31666 58382 31678 58434
rect 31826 58382 31838 58434
rect 31890 58382 31902 58434
rect 30606 58370 30658 58382
rect 34974 58370 35026 58382
rect 35198 58434 35250 58446
rect 35198 58370 35250 58382
rect 36878 58434 36930 58446
rect 36878 58370 36930 58382
rect 2494 58322 2546 58334
rect 15710 58322 15762 58334
rect 2494 58258 2546 58270
rect 7310 58266 7362 58278
rect 7198 58210 7250 58222
rect 15710 58258 15762 58270
rect 16158 58322 16210 58334
rect 16158 58258 16210 58270
rect 16606 58322 16658 58334
rect 16606 58258 16658 58270
rect 18062 58322 18114 58334
rect 18062 58258 18114 58270
rect 18398 58322 18450 58334
rect 18398 58258 18450 58270
rect 18846 58322 18898 58334
rect 18846 58258 18898 58270
rect 20078 58322 20130 58334
rect 20078 58258 20130 58270
rect 20190 58322 20242 58334
rect 20190 58258 20242 58270
rect 21982 58322 22034 58334
rect 37326 58322 37378 58334
rect 35522 58270 35534 58322
rect 35586 58270 35598 58322
rect 21982 58258 22034 58270
rect 37326 58258 37378 58270
rect 37550 58322 37602 58334
rect 37550 58258 37602 58270
rect 7310 58202 7362 58214
rect 8206 58210 8258 58222
rect 7198 58146 7250 58158
rect 8206 58146 8258 58158
rect 8766 58210 8818 58222
rect 12686 58210 12738 58222
rect 12114 58158 12126 58210
rect 12178 58158 12190 58210
rect 8766 58146 8818 58158
rect 12686 58146 12738 58158
rect 18734 58210 18786 58222
rect 18734 58146 18786 58158
rect 20638 58210 20690 58222
rect 20638 58146 20690 58158
rect 21646 58210 21698 58222
rect 21646 58146 21698 58158
rect 22542 58210 22594 58222
rect 22542 58146 22594 58158
rect 23662 58210 23714 58222
rect 27694 58210 27746 58222
rect 24210 58158 24222 58210
rect 24274 58158 24286 58210
rect 23662 58146 23714 58158
rect 27694 58146 27746 58158
rect 29598 58210 29650 58222
rect 29598 58146 29650 58158
rect 30270 58210 30322 58222
rect 30270 58146 30322 58158
rect 30942 58210 30994 58222
rect 30942 58146 30994 58158
rect 31390 58210 31442 58222
rect 31390 58146 31442 58158
rect 32734 58210 32786 58222
rect 32734 58146 32786 58158
rect 34414 58210 34466 58222
rect 34414 58146 34466 58158
rect 37102 58210 37154 58222
rect 37102 58146 37154 58158
rect 1344 58042 38640 58076
rect 1344 57990 14024 58042
rect 14076 57990 14148 58042
rect 14200 57990 14272 58042
rect 14324 57990 14396 58042
rect 14448 57990 14520 58042
rect 14572 57990 14644 58042
rect 14696 57990 14768 58042
rect 14820 57990 14892 58042
rect 14944 57990 15016 58042
rect 15068 57990 15140 58042
rect 15192 57990 34024 58042
rect 34076 57990 34148 58042
rect 34200 57990 34272 58042
rect 34324 57990 34396 58042
rect 34448 57990 34520 58042
rect 34572 57990 34644 58042
rect 34696 57990 34768 58042
rect 34820 57990 34892 58042
rect 34944 57990 35016 58042
rect 35068 57990 35140 58042
rect 35192 57990 38640 58042
rect 1344 57956 38640 57990
rect 6526 57874 6578 57886
rect 6526 57810 6578 57822
rect 7086 57874 7138 57886
rect 7086 57810 7138 57822
rect 7310 57874 7362 57886
rect 19294 57874 19346 57886
rect 8530 57822 8542 57874
rect 8594 57822 8606 57874
rect 12562 57822 12574 57874
rect 12626 57822 12638 57874
rect 7310 57810 7362 57822
rect 19294 57810 19346 57822
rect 20638 57874 20690 57886
rect 25342 57874 25394 57886
rect 24210 57822 24222 57874
rect 24274 57822 24286 57874
rect 20638 57810 20690 57822
rect 25342 57810 25394 57822
rect 28142 57874 28194 57886
rect 28142 57810 28194 57822
rect 29934 57874 29986 57886
rect 29934 57810 29986 57822
rect 30494 57874 30546 57886
rect 30494 57810 30546 57822
rect 30942 57874 30994 57886
rect 30942 57810 30994 57822
rect 33742 57874 33794 57886
rect 33742 57810 33794 57822
rect 34302 57874 34354 57886
rect 38334 57874 38386 57886
rect 37650 57822 37662 57874
rect 37714 57822 37726 57874
rect 34302 57810 34354 57822
rect 38334 57810 38386 57822
rect 18846 57762 18898 57774
rect 10546 57710 10558 57762
rect 10610 57710 10622 57762
rect 11890 57710 11902 57762
rect 11954 57710 11966 57762
rect 12674 57710 12686 57762
rect 12738 57710 12750 57762
rect 14242 57710 14254 57762
rect 14306 57710 14318 57762
rect 18846 57698 18898 57710
rect 24782 57762 24834 57774
rect 25890 57710 25902 57762
rect 25954 57710 25966 57762
rect 26226 57710 26238 57762
rect 26290 57710 26302 57762
rect 27234 57710 27246 57762
rect 27298 57710 27310 57762
rect 24782 57698 24834 57710
rect 6862 57650 6914 57662
rect 18622 57650 18674 57662
rect 19406 57650 19458 57662
rect 2818 57598 2830 57650
rect 2882 57598 2894 57650
rect 10770 57598 10782 57650
rect 10834 57598 10846 57650
rect 11778 57598 11790 57650
rect 11842 57598 11854 57650
rect 12786 57598 12798 57650
rect 12850 57598 12862 57650
rect 13794 57598 13806 57650
rect 13858 57598 13870 57650
rect 14354 57598 14366 57650
rect 14418 57598 14430 57650
rect 15362 57598 15374 57650
rect 15426 57598 15438 57650
rect 15810 57598 15822 57650
rect 15874 57598 15886 57650
rect 16370 57598 16382 57650
rect 16434 57598 16446 57650
rect 19170 57598 19182 57650
rect 19234 57598 19246 57650
rect 6862 57586 6914 57598
rect 18622 57586 18674 57598
rect 19406 57586 19458 57598
rect 19742 57650 19794 57662
rect 20750 57650 20802 57662
rect 20066 57598 20078 57650
rect 20130 57598 20142 57650
rect 19742 57586 19794 57598
rect 20750 57586 20802 57598
rect 21086 57650 21138 57662
rect 25678 57650 25730 57662
rect 27806 57650 27858 57662
rect 21634 57598 21646 57650
rect 21698 57598 21710 57650
rect 27122 57598 27134 57650
rect 27186 57598 27198 57650
rect 21086 57586 21138 57598
rect 25678 57586 25730 57598
rect 27806 57586 27858 57598
rect 34078 57650 34130 57662
rect 34078 57586 34130 57598
rect 34638 57650 34690 57662
rect 35298 57598 35310 57650
rect 35362 57598 35374 57650
rect 34638 57586 34690 57598
rect 2606 57538 2658 57550
rect 6974 57538 7026 57550
rect 3490 57486 3502 57538
rect 3554 57486 3566 57538
rect 2606 57474 2658 57486
rect 6974 57474 7026 57486
rect 7982 57538 8034 57550
rect 7982 57474 8034 57486
rect 9102 57538 9154 57550
rect 16830 57538 16882 57550
rect 15250 57486 15262 57538
rect 15314 57486 15326 57538
rect 9102 57474 9154 57486
rect 16830 57474 16882 57486
rect 17726 57538 17778 57550
rect 17726 57474 17778 57486
rect 18174 57538 18226 57550
rect 18174 57474 18226 57486
rect 20526 57538 20578 57550
rect 30818 57486 30830 57538
rect 30882 57486 30894 57538
rect 20526 57474 20578 57486
rect 8206 57426 8258 57438
rect 8206 57362 8258 57374
rect 9662 57426 9714 57438
rect 9662 57362 9714 57374
rect 9998 57426 10050 57438
rect 18510 57426 18562 57438
rect 17826 57374 17838 57426
rect 17890 57423 17902 57426
rect 18274 57423 18286 57426
rect 17890 57377 18286 57423
rect 17890 57374 17902 57377
rect 18274 57374 18286 57377
rect 18338 57374 18350 57426
rect 9998 57362 10050 57374
rect 18510 57362 18562 57374
rect 20302 57426 20354 57438
rect 20302 57362 20354 57374
rect 31166 57426 31218 57438
rect 31166 57362 31218 57374
rect 34414 57426 34466 57438
rect 34414 57362 34466 57374
rect 1344 57258 38640 57292
rect 1344 57206 4024 57258
rect 4076 57206 4148 57258
rect 4200 57206 4272 57258
rect 4324 57206 4396 57258
rect 4448 57206 4520 57258
rect 4572 57206 4644 57258
rect 4696 57206 4768 57258
rect 4820 57206 4892 57258
rect 4944 57206 5016 57258
rect 5068 57206 5140 57258
rect 5192 57206 24024 57258
rect 24076 57206 24148 57258
rect 24200 57206 24272 57258
rect 24324 57206 24396 57258
rect 24448 57206 24520 57258
rect 24572 57206 24644 57258
rect 24696 57206 24768 57258
rect 24820 57206 24892 57258
rect 24944 57206 25016 57258
rect 25068 57206 25140 57258
rect 25192 57206 38640 57258
rect 1344 57172 38640 57206
rect 6078 57090 6130 57102
rect 6078 57026 6130 57038
rect 12798 57090 12850 57102
rect 12798 57026 12850 57038
rect 13582 57090 13634 57102
rect 34862 57090 34914 57102
rect 25890 57038 25902 57090
rect 25954 57087 25966 57090
rect 26562 57087 26574 57090
rect 25954 57041 26574 57087
rect 25954 57038 25966 57041
rect 26562 57038 26574 57041
rect 26626 57038 26638 57090
rect 13582 57026 13634 57038
rect 34862 57026 34914 57038
rect 35870 57090 35922 57102
rect 35870 57026 35922 57038
rect 36206 57090 36258 57102
rect 36978 57038 36990 57090
rect 37042 57038 37054 57090
rect 36206 57026 36258 57038
rect 7422 56978 7474 56990
rect 7422 56914 7474 56926
rect 11678 56978 11730 56990
rect 26574 56978 26626 56990
rect 12450 56926 12462 56978
rect 12514 56926 12526 56978
rect 17378 56926 17390 56978
rect 17442 56926 17454 56978
rect 11678 56914 11730 56926
rect 26574 56914 26626 56926
rect 27470 56978 27522 56990
rect 27470 56914 27522 56926
rect 3614 56866 3666 56878
rect 7646 56866 7698 56878
rect 11342 56866 11394 56878
rect 4274 56814 4286 56866
rect 4338 56814 4350 56866
rect 6514 56814 6526 56866
rect 6578 56814 6590 56866
rect 8194 56814 8206 56866
rect 8258 56814 8270 56866
rect 3614 56802 3666 56814
rect 7646 56802 7698 56814
rect 11342 56802 11394 56814
rect 11566 56866 11618 56878
rect 11566 56802 11618 56814
rect 11902 56866 11954 56878
rect 11902 56802 11954 56814
rect 12126 56866 12178 56878
rect 21646 56866 21698 56878
rect 25790 56866 25842 56878
rect 14242 56814 14254 56866
rect 14306 56814 14318 56866
rect 15362 56814 15374 56866
rect 15426 56814 15438 56866
rect 16370 56814 16382 56866
rect 16434 56814 16446 56866
rect 17602 56814 17614 56866
rect 17666 56814 17678 56866
rect 18610 56814 18622 56866
rect 18674 56814 18686 56866
rect 19506 56814 19518 56866
rect 19570 56814 19582 56866
rect 20402 56814 20414 56866
rect 20466 56814 20478 56866
rect 25106 56814 25118 56866
rect 25170 56814 25182 56866
rect 12126 56802 12178 56814
rect 21646 56802 21698 56814
rect 25790 56802 25842 56814
rect 28590 56866 28642 56878
rect 28590 56802 28642 56814
rect 29038 56866 29090 56878
rect 35086 56866 35138 56878
rect 29698 56814 29710 56866
rect 29762 56814 29774 56866
rect 34626 56814 34638 56866
rect 34690 56814 34702 56866
rect 29038 56802 29090 56814
rect 35086 56802 35138 56814
rect 35982 56866 36034 56878
rect 37550 56866 37602 56878
rect 36418 56814 36430 56866
rect 36482 56814 36494 56866
rect 37762 56814 37774 56866
rect 37826 56814 37838 56866
rect 35982 56802 36034 56814
rect 37550 56802 37602 56814
rect 13470 56754 13522 56766
rect 18174 56754 18226 56766
rect 21310 56754 21362 56766
rect 4386 56702 4398 56754
rect 4450 56702 4462 56754
rect 6626 56702 6638 56754
rect 6690 56702 6702 56754
rect 14354 56702 14366 56754
rect 14418 56702 14430 56754
rect 15250 56702 15262 56754
rect 15314 56702 15326 56754
rect 19730 56702 19742 56754
rect 19794 56702 19806 56754
rect 20290 56702 20302 56754
rect 20354 56702 20366 56754
rect 13470 56690 13522 56702
rect 18174 56690 18226 56702
rect 21310 56690 21362 56702
rect 21870 56754 21922 56766
rect 21870 56690 21922 56702
rect 22878 56754 22930 56766
rect 22878 56690 22930 56702
rect 37438 56754 37490 56766
rect 37438 56690 37490 56702
rect 3278 56642 3330 56654
rect 3278 56578 3330 56590
rect 4958 56642 5010 56654
rect 4958 56578 5010 56590
rect 5742 56642 5794 56654
rect 12574 56642 12626 56654
rect 16830 56642 16882 56654
rect 21534 56642 21586 56654
rect 10546 56590 10558 56642
rect 10610 56590 10622 56642
rect 15026 56590 15038 56642
rect 15090 56590 15102 56642
rect 19618 56590 19630 56642
rect 19682 56590 19694 56642
rect 5742 56578 5794 56590
rect 12574 56578 12626 56590
rect 16830 56578 16882 56590
rect 21534 56578 21586 56590
rect 22094 56642 22146 56654
rect 22094 56578 22146 56590
rect 26126 56642 26178 56654
rect 26126 56578 26178 56590
rect 27022 56642 27074 56654
rect 27022 56578 27074 56590
rect 28142 56642 28194 56654
rect 32734 56642 32786 56654
rect 32050 56590 32062 56642
rect 32114 56590 32126 56642
rect 28142 56578 28194 56590
rect 32734 56578 32786 56590
rect 33854 56642 33906 56654
rect 33854 56578 33906 56590
rect 34302 56642 34354 56654
rect 34302 56578 34354 56590
rect 34750 56642 34802 56654
rect 34750 56578 34802 56590
rect 1344 56474 38640 56508
rect 1344 56422 14024 56474
rect 14076 56422 14148 56474
rect 14200 56422 14272 56474
rect 14324 56422 14396 56474
rect 14448 56422 14520 56474
rect 14572 56422 14644 56474
rect 14696 56422 14768 56474
rect 14820 56422 14892 56474
rect 14944 56422 15016 56474
rect 15068 56422 15140 56474
rect 15192 56422 34024 56474
rect 34076 56422 34148 56474
rect 34200 56422 34272 56474
rect 34324 56422 34396 56474
rect 34448 56422 34520 56474
rect 34572 56422 34644 56474
rect 34696 56422 34768 56474
rect 34820 56422 34892 56474
rect 34944 56422 35016 56474
rect 35068 56422 35140 56474
rect 35192 56422 38640 56474
rect 1344 56388 38640 56422
rect 9662 56306 9714 56318
rect 6626 56254 6638 56306
rect 6690 56254 6702 56306
rect 9662 56242 9714 56254
rect 18510 56306 18562 56318
rect 18510 56242 18562 56254
rect 18958 56306 19010 56318
rect 18958 56242 19010 56254
rect 20638 56306 20690 56318
rect 20638 56242 20690 56254
rect 22766 56306 22818 56318
rect 22766 56242 22818 56254
rect 24670 56306 24722 56318
rect 24670 56242 24722 56254
rect 25342 56306 25394 56318
rect 36766 56306 36818 56318
rect 36194 56254 36206 56306
rect 36258 56254 36270 56306
rect 25342 56242 25394 56254
rect 36766 56242 36818 56254
rect 36990 56306 37042 56318
rect 36990 56242 37042 56254
rect 37214 56306 37266 56318
rect 37214 56242 37266 56254
rect 8318 56194 8370 56206
rect 8318 56130 8370 56142
rect 20750 56194 20802 56206
rect 20750 56130 20802 56142
rect 22094 56194 22146 56206
rect 22094 56130 22146 56142
rect 22990 56194 23042 56206
rect 22990 56130 23042 56142
rect 32062 56194 32114 56206
rect 32062 56130 32114 56142
rect 37438 56194 37490 56206
rect 37438 56130 37490 56142
rect 2382 56082 2434 56094
rect 3726 56082 3778 56094
rect 13134 56082 13186 56094
rect 17390 56082 17442 56094
rect 2818 56030 2830 56082
rect 2882 56030 2894 56082
rect 4162 56030 4174 56082
rect 4226 56030 4238 56082
rect 7746 56030 7758 56082
rect 7810 56030 7822 56082
rect 11442 56030 11454 56082
rect 11506 56030 11518 56082
rect 11666 56030 11678 56082
rect 11730 56030 11742 56082
rect 12562 56030 12574 56082
rect 12626 56030 12638 56082
rect 15026 56030 15038 56082
rect 15090 56030 15102 56082
rect 16370 56030 16382 56082
rect 16434 56030 16446 56082
rect 2382 56018 2434 56030
rect 3726 56018 3778 56030
rect 13134 56018 13186 56030
rect 17390 56018 17442 56030
rect 17614 56082 17666 56094
rect 17614 56018 17666 56030
rect 20302 56082 20354 56094
rect 20302 56018 20354 56030
rect 21422 56082 21474 56094
rect 21422 56018 21474 56030
rect 22318 56082 22370 56094
rect 22318 56018 22370 56030
rect 32510 56082 32562 56094
rect 32510 56018 32562 56030
rect 33294 56082 33346 56094
rect 33730 56030 33742 56082
rect 33794 56030 33806 56082
rect 33294 56018 33346 56030
rect 3278 55970 3330 55982
rect 8766 55970 8818 55982
rect 7858 55918 7870 55970
rect 7922 55918 7934 55970
rect 3278 55906 3330 55918
rect 8766 55906 8818 55918
rect 10110 55970 10162 55982
rect 10110 55906 10162 55918
rect 10670 55970 10722 55982
rect 10670 55906 10722 55918
rect 11902 55970 11954 55982
rect 11902 55906 11954 55918
rect 13246 55970 13298 55982
rect 13246 55906 13298 55918
rect 13694 55970 13746 55982
rect 13694 55906 13746 55918
rect 14254 55970 14306 55982
rect 15486 55970 15538 55982
rect 16830 55970 16882 55982
rect 14578 55918 14590 55970
rect 14642 55918 14654 55970
rect 15922 55918 15934 55970
rect 15986 55918 15998 55970
rect 14254 55906 14306 55918
rect 15486 55906 15538 55918
rect 16830 55906 16882 55918
rect 18846 55970 18898 55982
rect 25790 55970 25842 55982
rect 21970 55918 21982 55970
rect 22034 55918 22046 55970
rect 18846 55906 18898 55918
rect 25790 55906 25842 55918
rect 37102 55970 37154 55982
rect 37102 55906 37154 55918
rect 7198 55858 7250 55870
rect 17838 55858 17890 55870
rect 8530 55806 8542 55858
rect 8594 55855 8606 55858
rect 9090 55855 9102 55858
rect 8594 55809 9102 55855
rect 8594 55806 8606 55809
rect 9090 55806 9102 55809
rect 9154 55806 9166 55858
rect 7198 55794 7250 55806
rect 17838 55794 17890 55806
rect 18062 55858 18114 55870
rect 18062 55794 18114 55806
rect 22654 55858 22706 55870
rect 22654 55794 22706 55806
rect 1344 55690 38640 55724
rect 1344 55638 4024 55690
rect 4076 55638 4148 55690
rect 4200 55638 4272 55690
rect 4324 55638 4396 55690
rect 4448 55638 4520 55690
rect 4572 55638 4644 55690
rect 4696 55638 4768 55690
rect 4820 55638 4892 55690
rect 4944 55638 5016 55690
rect 5068 55638 5140 55690
rect 5192 55638 24024 55690
rect 24076 55638 24148 55690
rect 24200 55638 24272 55690
rect 24324 55638 24396 55690
rect 24448 55638 24520 55690
rect 24572 55638 24644 55690
rect 24696 55638 24768 55690
rect 24820 55638 24892 55690
rect 24944 55638 25016 55690
rect 25068 55638 25140 55690
rect 25192 55638 38640 55690
rect 1344 55604 38640 55638
rect 3838 55522 3890 55534
rect 3838 55458 3890 55470
rect 7198 55522 7250 55534
rect 14590 55522 14642 55534
rect 11778 55470 11790 55522
rect 11842 55519 11854 55522
rect 12898 55519 12910 55522
rect 11842 55473 12910 55519
rect 11842 55470 11854 55473
rect 12898 55470 12910 55473
rect 12962 55470 12974 55522
rect 21858 55470 21870 55522
rect 21922 55519 21934 55522
rect 22642 55519 22654 55522
rect 21922 55473 22654 55519
rect 21922 55470 21934 55473
rect 22642 55470 22654 55473
rect 22706 55470 22718 55522
rect 7198 55458 7250 55470
rect 14590 55458 14642 55470
rect 11118 55410 11170 55422
rect 3266 55358 3278 55410
rect 3330 55358 3342 55410
rect 8530 55358 8542 55410
rect 8594 55358 8606 55410
rect 11118 55346 11170 55358
rect 13022 55410 13074 55422
rect 13022 55346 13074 55358
rect 14030 55410 14082 55422
rect 16830 55410 16882 55422
rect 16034 55358 16046 55410
rect 16098 55358 16110 55410
rect 14030 55346 14082 55358
rect 16830 55346 16882 55358
rect 21646 55410 21698 55422
rect 21646 55346 21698 55358
rect 22094 55410 22146 55422
rect 22094 55346 22146 55358
rect 22542 55410 22594 55422
rect 22542 55346 22594 55358
rect 35758 55410 35810 55422
rect 35758 55346 35810 55358
rect 36430 55410 36482 55422
rect 36430 55346 36482 55358
rect 37438 55410 37490 55422
rect 37438 55346 37490 55358
rect 4174 55298 4226 55310
rect 6190 55298 6242 55310
rect 10110 55298 10162 55310
rect 4834 55246 4846 55298
rect 4898 55246 4910 55298
rect 7970 55246 7982 55298
rect 8034 55246 8046 55298
rect 4174 55234 4226 55246
rect 6190 55234 6242 55246
rect 10110 55234 10162 55246
rect 13918 55298 13970 55310
rect 18958 55298 19010 55310
rect 14242 55246 14254 55298
rect 14306 55246 14318 55298
rect 16370 55246 16382 55298
rect 16434 55246 16446 55298
rect 13918 55234 13970 55246
rect 18958 55234 19010 55246
rect 37102 55298 37154 55310
rect 37102 55234 37154 55246
rect 37214 55298 37266 55310
rect 37214 55234 37266 55246
rect 37550 55298 37602 55310
rect 37550 55234 37602 55246
rect 7310 55186 7362 55198
rect 12462 55186 12514 55198
rect 4946 55134 4958 55186
rect 5010 55134 5022 55186
rect 8418 55134 8430 55186
rect 8482 55134 8494 55186
rect 7310 55122 7362 55134
rect 12462 55122 12514 55134
rect 18398 55186 18450 55198
rect 18398 55122 18450 55134
rect 18734 55186 18786 55198
rect 18734 55122 18786 55134
rect 19294 55186 19346 55198
rect 19294 55122 19346 55134
rect 2606 55074 2658 55086
rect 2606 55010 2658 55022
rect 2830 55074 2882 55086
rect 2830 55010 2882 55022
rect 5742 55074 5794 55086
rect 5742 55010 5794 55022
rect 6862 55074 6914 55086
rect 6862 55010 6914 55022
rect 11566 55074 11618 55086
rect 11566 55010 11618 55022
rect 12014 55074 12066 55086
rect 12014 55010 12066 55022
rect 14142 55074 14194 55086
rect 14142 55010 14194 55022
rect 15038 55074 15090 55086
rect 15038 55010 15090 55022
rect 15486 55074 15538 55086
rect 15486 55010 15538 55022
rect 18846 55074 18898 55086
rect 18846 55010 18898 55022
rect 35646 55074 35698 55086
rect 35646 55010 35698 55022
rect 1344 54906 38640 54940
rect 1344 54854 14024 54906
rect 14076 54854 14148 54906
rect 14200 54854 14272 54906
rect 14324 54854 14396 54906
rect 14448 54854 14520 54906
rect 14572 54854 14644 54906
rect 14696 54854 14768 54906
rect 14820 54854 14892 54906
rect 14944 54854 15016 54906
rect 15068 54854 15140 54906
rect 15192 54854 34024 54906
rect 34076 54854 34148 54906
rect 34200 54854 34272 54906
rect 34324 54854 34396 54906
rect 34448 54854 34520 54906
rect 34572 54854 34644 54906
rect 34696 54854 34768 54906
rect 34820 54854 34892 54906
rect 34944 54854 35016 54906
rect 35068 54854 35140 54906
rect 35192 54854 38640 54906
rect 1344 54820 38640 54854
rect 5294 54738 5346 54750
rect 4722 54686 4734 54738
rect 4786 54686 4798 54738
rect 5294 54674 5346 54686
rect 5630 54738 5682 54750
rect 5630 54674 5682 54686
rect 8094 54738 8146 54750
rect 8094 54674 8146 54686
rect 11902 54738 11954 54750
rect 21758 54738 21810 54750
rect 21186 54686 21198 54738
rect 21250 54686 21262 54738
rect 11902 54674 11954 54686
rect 21758 54674 21810 54686
rect 22094 54738 22146 54750
rect 22094 54674 22146 54686
rect 26462 54738 26514 54750
rect 31166 54738 31218 54750
rect 30258 54686 30270 54738
rect 30322 54686 30334 54738
rect 26462 54674 26514 54686
rect 31166 54674 31218 54686
rect 34078 54738 34130 54750
rect 37538 54686 37550 54738
rect 37602 54686 37614 54738
rect 34078 54674 34130 54686
rect 6302 54626 6354 54638
rect 6302 54562 6354 54574
rect 8990 54626 9042 54638
rect 10770 54574 10782 54626
rect 10834 54574 10846 54626
rect 8990 54562 9042 54574
rect 1822 54514 1874 54526
rect 6190 54514 6242 54526
rect 2258 54462 2270 54514
rect 2322 54462 2334 54514
rect 1822 54450 1874 54462
rect 6190 54450 6242 54462
rect 6526 54514 6578 54526
rect 6526 54450 6578 54462
rect 6750 54514 6802 54526
rect 6750 54450 6802 54462
rect 7086 54514 7138 54526
rect 7086 54450 7138 54462
rect 7198 54514 7250 54526
rect 9998 54514 10050 54526
rect 13470 54514 13522 54526
rect 18286 54514 18338 54526
rect 27358 54514 27410 54526
rect 34526 54514 34578 54526
rect 38222 54514 38274 54526
rect 7634 54462 7646 54514
rect 7698 54462 7710 54514
rect 10658 54462 10670 54514
rect 10722 54462 10734 54514
rect 13010 54462 13022 54514
rect 13074 54462 13086 54514
rect 15026 54462 15038 54514
rect 15090 54462 15102 54514
rect 18722 54462 18734 54514
rect 18786 54462 18798 54514
rect 27682 54462 27694 54514
rect 27746 54462 27758 54514
rect 35186 54462 35198 54514
rect 35250 54462 35262 54514
rect 7198 54450 7250 54462
rect 9998 54450 10050 54462
rect 13470 54450 13522 54462
rect 18286 54450 18338 54462
rect 27358 54450 27410 54462
rect 34526 54450 34578 54462
rect 38222 54450 38274 54462
rect 7422 54402 7474 54414
rect 7422 54338 7474 54350
rect 11454 54402 11506 54414
rect 11454 54338 11506 54350
rect 12350 54402 12402 54414
rect 15598 54402 15650 54414
rect 15250 54350 15262 54402
rect 15314 54350 15326 54402
rect 12350 54338 12402 54350
rect 15598 54338 15650 54350
rect 22542 54402 22594 54414
rect 22542 54338 22594 54350
rect 27022 54402 27074 54414
rect 27022 54338 27074 54350
rect 33630 54402 33682 54414
rect 33630 54338 33682 54350
rect 9662 54290 9714 54302
rect 9662 54226 9714 54238
rect 13246 54290 13298 54302
rect 13246 54226 13298 54238
rect 13694 54290 13746 54302
rect 13694 54226 13746 54238
rect 13806 54290 13858 54302
rect 13806 54226 13858 54238
rect 30830 54290 30882 54302
rect 30830 54226 30882 54238
rect 1344 54122 38640 54156
rect 1344 54070 4024 54122
rect 4076 54070 4148 54122
rect 4200 54070 4272 54122
rect 4324 54070 4396 54122
rect 4448 54070 4520 54122
rect 4572 54070 4644 54122
rect 4696 54070 4768 54122
rect 4820 54070 4892 54122
rect 4944 54070 5016 54122
rect 5068 54070 5140 54122
rect 5192 54070 24024 54122
rect 24076 54070 24148 54122
rect 24200 54070 24272 54122
rect 24324 54070 24396 54122
rect 24448 54070 24520 54122
rect 24572 54070 24644 54122
rect 24696 54070 24768 54122
rect 24820 54070 24892 54122
rect 24944 54070 25016 54122
rect 25068 54070 25140 54122
rect 25192 54070 38640 54122
rect 1344 54036 38640 54070
rect 14814 53954 14866 53966
rect 14814 53890 14866 53902
rect 15374 53954 15426 53966
rect 19294 53954 19346 53966
rect 18610 53902 18622 53954
rect 18674 53902 18686 53954
rect 15374 53890 15426 53902
rect 19294 53890 19346 53902
rect 19630 53954 19682 53966
rect 19630 53890 19682 53902
rect 26462 53954 26514 53966
rect 26462 53890 26514 53902
rect 27694 53954 27746 53966
rect 30370 53902 30382 53954
rect 30434 53951 30446 53954
rect 31042 53951 31054 53954
rect 30434 53905 31054 53951
rect 30434 53902 30446 53905
rect 31042 53902 31054 53905
rect 31106 53902 31118 53954
rect 27694 53890 27746 53902
rect 6974 53842 7026 53854
rect 3266 53790 3278 53842
rect 3330 53790 3342 53842
rect 6974 53778 7026 53790
rect 12910 53842 12962 53854
rect 12910 53778 12962 53790
rect 13470 53842 13522 53854
rect 15598 53842 15650 53854
rect 20078 53842 20130 53854
rect 14354 53790 14366 53842
rect 14418 53790 14430 53842
rect 15026 53790 15038 53842
rect 15090 53790 15102 53842
rect 18162 53790 18174 53842
rect 18226 53790 18238 53842
rect 13470 53778 13522 53790
rect 15598 53778 15650 53790
rect 20078 53778 20130 53790
rect 30382 53842 30434 53854
rect 30382 53778 30434 53790
rect 2494 53730 2546 53742
rect 2494 53666 2546 53678
rect 2830 53730 2882 53742
rect 2830 53666 2882 53678
rect 5630 53730 5682 53742
rect 5630 53666 5682 53678
rect 7870 53730 7922 53742
rect 11566 53730 11618 53742
rect 12798 53730 12850 53742
rect 24670 53730 24722 53742
rect 26798 53730 26850 53742
rect 8530 53678 8542 53730
rect 8594 53678 8606 53730
rect 12226 53678 12238 53730
rect 12290 53678 12302 53730
rect 13906 53678 13918 53730
rect 13970 53678 13982 53730
rect 18274 53678 18286 53730
rect 18338 53678 18350 53730
rect 25890 53678 25902 53730
rect 25954 53678 25966 53730
rect 7870 53666 7922 53678
rect 11566 53666 11618 53678
rect 12798 53666 12850 53678
rect 24670 53666 24722 53678
rect 26798 53666 26850 53678
rect 5742 53618 5794 53630
rect 5742 53554 5794 53566
rect 15038 53618 15090 53630
rect 15038 53554 15090 53566
rect 19406 53618 19458 53630
rect 30830 53618 30882 53630
rect 25666 53566 25678 53618
rect 25730 53566 25742 53618
rect 28018 53566 28030 53618
rect 28082 53566 28094 53618
rect 28466 53566 28478 53618
rect 28530 53566 28542 53618
rect 19406 53554 19458 53566
rect 30830 53554 30882 53566
rect 31278 53618 31330 53630
rect 31278 53554 31330 53566
rect 31390 53618 31442 53630
rect 31390 53554 31442 53566
rect 31950 53618 32002 53630
rect 31950 53554 32002 53566
rect 25118 53506 25170 53518
rect 10882 53454 10894 53506
rect 10946 53454 10958 53506
rect 25118 53442 25170 53454
rect 27358 53506 27410 53518
rect 27358 53442 27410 53454
rect 29374 53506 29426 53518
rect 29374 53442 29426 53454
rect 31614 53506 31666 53518
rect 31614 53442 31666 53454
rect 1344 53338 38640 53372
rect 1344 53286 14024 53338
rect 14076 53286 14148 53338
rect 14200 53286 14272 53338
rect 14324 53286 14396 53338
rect 14448 53286 14520 53338
rect 14572 53286 14644 53338
rect 14696 53286 14768 53338
rect 14820 53286 14892 53338
rect 14944 53286 15016 53338
rect 15068 53286 15140 53338
rect 15192 53286 34024 53338
rect 34076 53286 34148 53338
rect 34200 53286 34272 53338
rect 34324 53286 34396 53338
rect 34448 53286 34520 53338
rect 34572 53286 34644 53338
rect 34696 53286 34768 53338
rect 34820 53286 34892 53338
rect 34944 53286 35016 53338
rect 35068 53286 35140 53338
rect 35192 53286 38640 53338
rect 1344 53252 38640 53286
rect 4062 53170 4114 53182
rect 4062 53106 4114 53118
rect 5182 53170 5234 53182
rect 5182 53106 5234 53118
rect 5854 53170 5906 53182
rect 5854 53106 5906 53118
rect 6526 53170 6578 53182
rect 13134 53170 13186 53182
rect 12562 53118 12574 53170
rect 12626 53118 12638 53170
rect 6526 53106 6578 53118
rect 13134 53106 13186 53118
rect 18958 53170 19010 53182
rect 18958 53106 19010 53118
rect 21646 53170 21698 53182
rect 21646 53106 21698 53118
rect 22094 53170 22146 53182
rect 22094 53106 22146 53118
rect 22654 53170 22706 53182
rect 22654 53106 22706 53118
rect 22878 53170 22930 53182
rect 22878 53106 22930 53118
rect 24222 53170 24274 53182
rect 24222 53106 24274 53118
rect 25342 53170 25394 53182
rect 25342 53106 25394 53118
rect 26350 53170 26402 53182
rect 30270 53170 30322 53182
rect 29698 53118 29710 53170
rect 29762 53118 29774 53170
rect 26350 53106 26402 53118
rect 30270 53106 30322 53118
rect 6078 53058 6130 53070
rect 6078 52994 6130 53006
rect 13358 53058 13410 53070
rect 13358 52994 13410 53006
rect 23438 53058 23490 53070
rect 23438 52994 23490 53006
rect 23662 53058 23714 53070
rect 23662 52994 23714 53006
rect 23774 53058 23826 53070
rect 23774 52994 23826 53006
rect 30942 53058 30994 53070
rect 30942 52994 30994 53006
rect 2494 52946 2546 52958
rect 2494 52882 2546 52894
rect 2830 52946 2882 52958
rect 2830 52882 2882 52894
rect 3726 52946 3778 52958
rect 3726 52882 3778 52894
rect 5406 52946 5458 52958
rect 5406 52882 5458 52894
rect 9438 52946 9490 52958
rect 13918 52946 13970 52958
rect 10098 52894 10110 52946
rect 10162 52894 10174 52946
rect 9438 52882 9490 52894
rect 13918 52882 13970 52894
rect 23326 52946 23378 52958
rect 23326 52882 23378 52894
rect 26574 52946 26626 52958
rect 30830 52946 30882 52958
rect 27234 52894 27246 52946
rect 27298 52894 27310 52946
rect 26574 52882 26626 52894
rect 30830 52882 30882 52894
rect 31166 52946 31218 52958
rect 31166 52882 31218 52894
rect 31502 52946 31554 52958
rect 31502 52882 31554 52894
rect 31950 52946 32002 52958
rect 31950 52882 32002 52894
rect 32174 52946 32226 52958
rect 32174 52882 32226 52894
rect 2046 52834 2098 52846
rect 4734 52834 4786 52846
rect 3266 52782 3278 52834
rect 3330 52782 3342 52834
rect 2046 52770 2098 52782
rect 4734 52770 4786 52782
rect 5966 52834 6018 52846
rect 5966 52770 6018 52782
rect 14702 52834 14754 52846
rect 14702 52770 14754 52782
rect 20974 52834 21026 52846
rect 20974 52770 21026 52782
rect 22766 52834 22818 52846
rect 22766 52770 22818 52782
rect 25790 52834 25842 52846
rect 25790 52770 25842 52782
rect 32062 52834 32114 52846
rect 32062 52770 32114 52782
rect 13470 52722 13522 52734
rect 13470 52658 13522 52670
rect 1344 52554 38640 52588
rect 1344 52502 4024 52554
rect 4076 52502 4148 52554
rect 4200 52502 4272 52554
rect 4324 52502 4396 52554
rect 4448 52502 4520 52554
rect 4572 52502 4644 52554
rect 4696 52502 4768 52554
rect 4820 52502 4892 52554
rect 4944 52502 5016 52554
rect 5068 52502 5140 52554
rect 5192 52502 24024 52554
rect 24076 52502 24148 52554
rect 24200 52502 24272 52554
rect 24324 52502 24396 52554
rect 24448 52502 24520 52554
rect 24572 52502 24644 52554
rect 24696 52502 24768 52554
rect 24820 52502 24892 52554
rect 24944 52502 25016 52554
rect 25068 52502 25140 52554
rect 25192 52502 38640 52554
rect 1344 52468 38640 52502
rect 26574 52386 26626 52398
rect 26574 52322 26626 52334
rect 9774 52274 9826 52286
rect 9774 52210 9826 52222
rect 10558 52274 10610 52286
rect 10558 52210 10610 52222
rect 11006 52274 11058 52286
rect 19854 52274 19906 52286
rect 11778 52222 11790 52274
rect 11842 52222 11854 52274
rect 11006 52210 11058 52222
rect 19854 52210 19906 52222
rect 25454 52274 25506 52286
rect 25454 52210 25506 52222
rect 30046 52274 30098 52286
rect 30046 52210 30098 52222
rect 3614 52162 3666 52174
rect 5182 52162 5234 52174
rect 4050 52110 4062 52162
rect 4114 52110 4126 52162
rect 3614 52098 3666 52110
rect 5182 52098 5234 52110
rect 5518 52162 5570 52174
rect 11230 52162 11282 52174
rect 6066 52110 6078 52162
rect 6130 52110 6142 52162
rect 5518 52098 5570 52110
rect 11230 52098 11282 52110
rect 11454 52162 11506 52174
rect 11454 52098 11506 52110
rect 12126 52162 12178 52174
rect 12126 52098 12178 52110
rect 12574 52162 12626 52174
rect 12574 52098 12626 52110
rect 20302 52162 20354 52174
rect 20302 52098 20354 52110
rect 20414 52162 20466 52174
rect 20414 52098 20466 52110
rect 20862 52162 20914 52174
rect 20862 52098 20914 52110
rect 21198 52162 21250 52174
rect 21198 52098 21250 52110
rect 21534 52162 21586 52174
rect 30270 52162 30322 52174
rect 21858 52110 21870 52162
rect 21922 52110 21934 52162
rect 22418 52110 22430 52162
rect 22482 52110 22494 52162
rect 25890 52110 25902 52162
rect 25954 52110 25966 52162
rect 21534 52098 21586 52110
rect 30270 52098 30322 52110
rect 31166 52162 31218 52174
rect 31826 52110 31838 52162
rect 31890 52110 31902 52162
rect 31166 52098 31218 52110
rect 4846 52050 4898 52062
rect 4386 51998 4398 52050
rect 4450 51998 4462 52050
rect 4846 51986 4898 51998
rect 4958 52050 5010 52062
rect 4958 51986 5010 51998
rect 10894 52050 10946 52062
rect 10894 51986 10946 51998
rect 11902 52050 11954 52062
rect 11902 51986 11954 51998
rect 19406 52050 19458 52062
rect 19406 51986 19458 51998
rect 20190 52050 20242 52062
rect 27582 52050 27634 52062
rect 25778 51998 25790 52050
rect 25842 51998 25854 52050
rect 20190 51986 20242 51998
rect 27582 51986 27634 51998
rect 30718 52050 30770 52062
rect 30718 51986 30770 51998
rect 3278 51938 3330 51950
rect 9214 51938 9266 51950
rect 8530 51886 8542 51938
rect 8594 51886 8606 51938
rect 3278 51874 3330 51886
rect 9214 51874 9266 51886
rect 13582 51938 13634 51950
rect 13582 51874 13634 51886
rect 21422 51938 21474 51950
rect 26910 51938 26962 51950
rect 24882 51886 24894 51938
rect 24946 51886 24958 51938
rect 21422 51874 21474 51886
rect 26910 51874 26962 51886
rect 30830 51938 30882 51950
rect 30830 51874 30882 51886
rect 30942 51938 30994 51950
rect 34862 51938 34914 51950
rect 34066 51886 34078 51938
rect 34130 51886 34142 51938
rect 30942 51874 30994 51886
rect 34862 51874 34914 51886
rect 1344 51770 38640 51804
rect 1344 51718 14024 51770
rect 14076 51718 14148 51770
rect 14200 51718 14272 51770
rect 14324 51718 14396 51770
rect 14448 51718 14520 51770
rect 14572 51718 14644 51770
rect 14696 51718 14768 51770
rect 14820 51718 14892 51770
rect 14944 51718 15016 51770
rect 15068 51718 15140 51770
rect 15192 51718 34024 51770
rect 34076 51718 34148 51770
rect 34200 51718 34272 51770
rect 34324 51718 34396 51770
rect 34448 51718 34520 51770
rect 34572 51718 34644 51770
rect 34696 51718 34768 51770
rect 34820 51718 34892 51770
rect 34944 51718 35016 51770
rect 35068 51718 35140 51770
rect 35192 51718 38640 51770
rect 1344 51684 38640 51718
rect 5294 51602 5346 51614
rect 4722 51550 4734 51602
rect 4786 51550 4798 51602
rect 5294 51538 5346 51550
rect 11678 51602 11730 51614
rect 11678 51538 11730 51550
rect 14254 51602 14306 51614
rect 23438 51602 23490 51614
rect 22866 51550 22878 51602
rect 22930 51550 22942 51602
rect 14254 51538 14306 51550
rect 23438 51538 23490 51550
rect 23774 51602 23826 51614
rect 23774 51538 23826 51550
rect 24222 51602 24274 51614
rect 24222 51538 24274 51550
rect 25790 51602 25842 51614
rect 25790 51538 25842 51550
rect 27022 51602 27074 51614
rect 27022 51538 27074 51550
rect 27470 51602 27522 51614
rect 27470 51538 27522 51550
rect 30942 51602 30994 51614
rect 30942 51538 30994 51550
rect 15598 51490 15650 51502
rect 32398 51490 32450 51502
rect 7298 51438 7310 51490
rect 7362 51438 7374 51490
rect 14802 51438 14814 51490
rect 14866 51438 14878 51490
rect 16258 51438 16270 51490
rect 16322 51438 16334 51490
rect 28018 51438 28030 51490
rect 28082 51438 28094 51490
rect 28466 51438 28478 51490
rect 28530 51438 28542 51490
rect 15598 51426 15650 51438
rect 32398 51426 32450 51438
rect 1822 51378 1874 51390
rect 2258 51338 2270 51390
rect 2322 51338 2334 51390
rect 8542 51378 8594 51390
rect 19966 51378 20018 51390
rect 27806 51378 27858 51390
rect 33182 51378 33234 51390
rect 6066 51326 6078 51378
rect 6130 51326 6142 51378
rect 15362 51326 15374 51378
rect 15426 51326 15438 51378
rect 15698 51326 15710 51378
rect 15762 51326 15774 51378
rect 18274 51326 18286 51378
rect 18338 51326 18350 51378
rect 20290 51326 20302 51378
rect 20354 51326 20366 51378
rect 31938 51326 31950 51378
rect 32002 51326 32014 51378
rect 1822 51314 1874 51326
rect 8542 51314 8594 51326
rect 19966 51314 20018 51326
rect 27806 51314 27858 51326
rect 33182 51314 33234 51326
rect 9662 51266 9714 51278
rect 9662 51202 9714 51214
rect 14366 51266 14418 51278
rect 14366 51202 14418 51214
rect 17614 51266 17666 51278
rect 17614 51202 17666 51214
rect 17838 51266 17890 51278
rect 25342 51266 25394 51278
rect 18162 51214 18174 51266
rect 18226 51214 18238 51266
rect 31602 51214 31614 51266
rect 31666 51214 31678 51266
rect 17838 51202 17890 51214
rect 25342 51202 25394 51214
rect 17266 51102 17278 51154
rect 17330 51151 17342 51154
rect 17602 51151 17614 51154
rect 17330 51105 17614 51151
rect 17330 51102 17342 51105
rect 17602 51102 17614 51105
rect 17666 51102 17678 51154
rect 25330 51102 25342 51154
rect 25394 51151 25406 51154
rect 25890 51151 25902 51154
rect 25394 51105 25902 51151
rect 25394 51102 25406 51105
rect 25890 51102 25902 51105
rect 25954 51102 25966 51154
rect 1344 50986 38640 51020
rect 1344 50934 4024 50986
rect 4076 50934 4148 50986
rect 4200 50934 4272 50986
rect 4324 50934 4396 50986
rect 4448 50934 4520 50986
rect 4572 50934 4644 50986
rect 4696 50934 4768 50986
rect 4820 50934 4892 50986
rect 4944 50934 5016 50986
rect 5068 50934 5140 50986
rect 5192 50934 24024 50986
rect 24076 50934 24148 50986
rect 24200 50934 24272 50986
rect 24324 50934 24396 50986
rect 24448 50934 24520 50986
rect 24572 50934 24644 50986
rect 24696 50934 24768 50986
rect 24820 50934 24892 50986
rect 24944 50934 25016 50986
rect 25068 50934 25140 50986
rect 25192 50934 38640 50986
rect 1344 50900 38640 50934
rect 5506 50766 5518 50818
rect 5570 50815 5582 50818
rect 5730 50815 5742 50818
rect 5570 50769 5742 50815
rect 5570 50766 5582 50769
rect 5730 50766 5742 50769
rect 5794 50815 5806 50818
rect 6626 50815 6638 50818
rect 5794 50769 6638 50815
rect 5794 50766 5806 50769
rect 6626 50766 6638 50769
rect 6690 50766 6702 50818
rect 5742 50706 5794 50718
rect 5742 50642 5794 50654
rect 6190 50706 6242 50718
rect 6190 50642 6242 50654
rect 8318 50706 8370 50718
rect 8318 50642 8370 50654
rect 9102 50706 9154 50718
rect 9102 50642 9154 50654
rect 15262 50706 15314 50718
rect 15262 50642 15314 50654
rect 16830 50706 16882 50718
rect 16830 50642 16882 50654
rect 18622 50706 18674 50718
rect 19854 50706 19906 50718
rect 19170 50654 19182 50706
rect 19234 50654 19246 50706
rect 18622 50642 18674 50654
rect 19854 50642 19906 50654
rect 23102 50706 23154 50718
rect 24894 50706 24946 50718
rect 24322 50654 24334 50706
rect 24386 50654 24398 50706
rect 23102 50642 23154 50654
rect 24894 50642 24946 50654
rect 30718 50706 30770 50718
rect 30718 50642 30770 50654
rect 31166 50706 31218 50718
rect 31166 50642 31218 50654
rect 3838 50594 3890 50606
rect 3838 50530 3890 50542
rect 4174 50594 4226 50606
rect 15150 50594 15202 50606
rect 14802 50542 14814 50594
rect 14866 50542 14878 50594
rect 4174 50530 4226 50542
rect 15150 50530 15202 50542
rect 15934 50594 15986 50606
rect 31614 50594 31666 50606
rect 16146 50542 16158 50594
rect 16210 50542 16222 50594
rect 18162 50542 18174 50594
rect 18226 50542 18238 50594
rect 19394 50542 19406 50594
rect 19458 50542 19470 50594
rect 23874 50542 23886 50594
rect 23938 50542 23950 50594
rect 32162 50542 32174 50594
rect 32226 50542 32238 50594
rect 15934 50530 15986 50542
rect 31614 50530 31666 50542
rect 6638 50482 6690 50494
rect 4498 50430 4510 50482
rect 4562 50430 4574 50482
rect 4946 50430 4958 50482
rect 5010 50430 5022 50482
rect 6638 50418 6690 50430
rect 17278 50482 17330 50494
rect 23438 50482 23490 50494
rect 19282 50430 19294 50482
rect 19346 50430 19358 50482
rect 17278 50418 17330 50430
rect 23438 50418 23490 50430
rect 34526 50482 34578 50494
rect 34526 50418 34578 50430
rect 13918 50370 13970 50382
rect 13918 50306 13970 50318
rect 35310 50370 35362 50382
rect 35310 50306 35362 50318
rect 1344 50202 38640 50236
rect 1344 50150 14024 50202
rect 14076 50150 14148 50202
rect 14200 50150 14272 50202
rect 14324 50150 14396 50202
rect 14448 50150 14520 50202
rect 14572 50150 14644 50202
rect 14696 50150 14768 50202
rect 14820 50150 14892 50202
rect 14944 50150 15016 50202
rect 15068 50150 15140 50202
rect 15192 50150 34024 50202
rect 34076 50150 34148 50202
rect 34200 50150 34272 50202
rect 34324 50150 34396 50202
rect 34448 50150 34520 50202
rect 34572 50150 34644 50202
rect 34696 50150 34768 50202
rect 34820 50150 34892 50202
rect 34944 50150 35016 50202
rect 35068 50150 35140 50202
rect 35192 50150 38640 50202
rect 1344 50116 38640 50150
rect 5518 50034 5570 50046
rect 5518 49970 5570 49982
rect 7310 50034 7362 50046
rect 7310 49970 7362 49982
rect 8654 50034 8706 50046
rect 8654 49970 8706 49982
rect 9662 50034 9714 50046
rect 9662 49970 9714 49982
rect 14590 50034 14642 50046
rect 18162 49982 18174 50034
rect 18226 49982 18238 50034
rect 23986 49982 23998 50034
rect 24050 49982 24062 50034
rect 14590 49970 14642 49982
rect 7758 49922 7810 49934
rect 7758 49858 7810 49870
rect 7870 49922 7922 49934
rect 7870 49858 7922 49870
rect 13470 49922 13522 49934
rect 13470 49858 13522 49870
rect 16606 49922 16658 49934
rect 26462 49922 26514 49934
rect 18050 49870 18062 49922
rect 18114 49870 18126 49922
rect 19506 49870 19518 49922
rect 19570 49870 19582 49922
rect 28130 49870 28142 49922
rect 28194 49870 28206 49922
rect 28690 49870 28702 49922
rect 28754 49870 28766 49922
rect 16606 49858 16658 49870
rect 26462 49858 26514 49870
rect 2830 49810 2882 49822
rect 2830 49746 2882 49758
rect 7534 49810 7586 49822
rect 7534 49746 7586 49758
rect 10782 49810 10834 49822
rect 15374 49810 15426 49822
rect 21982 49810 22034 49822
rect 11218 49758 11230 49810
rect 11282 49758 11294 49810
rect 15922 49758 15934 49810
rect 15986 49758 15998 49810
rect 17938 49758 17950 49810
rect 18002 49758 18014 49810
rect 18946 49758 18958 49810
rect 19010 49758 19022 49810
rect 22418 49758 22430 49810
rect 22482 49758 22494 49810
rect 23538 49758 23550 49810
rect 23602 49758 23614 49810
rect 23762 49758 23774 49810
rect 23826 49758 23838 49810
rect 10782 49746 10834 49758
rect 15374 49746 15426 49758
rect 21982 49746 22034 49758
rect 2494 49698 2546 49710
rect 10334 49698 10386 49710
rect 17502 49698 17554 49710
rect 3266 49646 3278 49698
rect 3330 49646 3342 49698
rect 15698 49646 15710 49698
rect 15762 49646 15774 49698
rect 2494 49634 2546 49646
rect 10334 49634 10386 49646
rect 17502 49634 17554 49646
rect 22878 49698 22930 49710
rect 27134 49698 27186 49710
rect 23426 49646 23438 49698
rect 23490 49646 23502 49698
rect 22878 49634 22930 49646
rect 27134 49634 27186 49646
rect 32174 49698 32226 49710
rect 32174 49634 32226 49646
rect 32510 49698 32562 49710
rect 32510 49634 32562 49646
rect 33182 49698 33234 49710
rect 33182 49634 33234 49646
rect 8542 49586 8594 49598
rect 8542 49522 8594 49534
rect 8878 49586 8930 49598
rect 8878 49522 8930 49534
rect 14254 49586 14306 49598
rect 14254 49522 14306 49534
rect 27582 49586 27634 49598
rect 27582 49522 27634 49534
rect 27918 49586 27970 49598
rect 31938 49534 31950 49586
rect 32002 49583 32014 49586
rect 32498 49583 32510 49586
rect 32002 49537 32510 49583
rect 32002 49534 32014 49537
rect 32498 49534 32510 49537
rect 32562 49534 32574 49586
rect 27918 49522 27970 49534
rect 1344 49418 38640 49452
rect 1344 49366 4024 49418
rect 4076 49366 4148 49418
rect 4200 49366 4272 49418
rect 4324 49366 4396 49418
rect 4448 49366 4520 49418
rect 4572 49366 4644 49418
rect 4696 49366 4768 49418
rect 4820 49366 4892 49418
rect 4944 49366 5016 49418
rect 5068 49366 5140 49418
rect 5192 49366 24024 49418
rect 24076 49366 24148 49418
rect 24200 49366 24272 49418
rect 24324 49366 24396 49418
rect 24448 49366 24520 49418
rect 24572 49366 24644 49418
rect 24696 49366 24768 49418
rect 24820 49366 24892 49418
rect 24944 49366 25016 49418
rect 25068 49366 25140 49418
rect 25192 49366 38640 49418
rect 1344 49332 38640 49366
rect 19294 49250 19346 49262
rect 19294 49186 19346 49198
rect 26238 49250 26290 49262
rect 26238 49186 26290 49198
rect 27694 49250 27746 49262
rect 27694 49186 27746 49198
rect 28030 49250 28082 49262
rect 28030 49186 28082 49198
rect 33518 49250 33570 49262
rect 33518 49186 33570 49198
rect 11230 49138 11282 49150
rect 11230 49074 11282 49086
rect 11678 49138 11730 49150
rect 11678 49074 11730 49086
rect 15150 49138 15202 49150
rect 15150 49074 15202 49086
rect 16494 49138 16546 49150
rect 16494 49074 16546 49086
rect 20078 49138 20130 49150
rect 20078 49074 20130 49086
rect 23550 49138 23602 49150
rect 32174 49138 32226 49150
rect 31602 49086 31614 49138
rect 31666 49086 31678 49138
rect 23550 49074 23602 49086
rect 32174 49074 32226 49086
rect 6862 49026 6914 49038
rect 11566 49026 11618 49038
rect 7298 48974 7310 49026
rect 7362 48974 7374 49026
rect 6862 48962 6914 48974
rect 11566 48962 11618 48974
rect 12238 49026 12290 49038
rect 12238 48962 12290 48974
rect 12574 49026 12626 49038
rect 12574 48962 12626 48974
rect 12910 49026 12962 49038
rect 12910 48962 12962 48974
rect 13918 49026 13970 49038
rect 13918 48962 13970 48974
rect 14254 49026 14306 49038
rect 15598 49026 15650 49038
rect 17726 49026 17778 49038
rect 14690 48974 14702 49026
rect 14754 48974 14766 49026
rect 15810 48974 15822 49026
rect 15874 48974 15886 49026
rect 17042 48974 17054 49026
rect 17106 48974 17118 49026
rect 14254 48962 14306 48974
rect 15598 48962 15650 48974
rect 17726 48962 17778 48974
rect 18398 49026 18450 49038
rect 18398 48962 18450 48974
rect 18510 49026 18562 49038
rect 31278 49026 31330 49038
rect 33070 49026 33122 49038
rect 18834 48974 18846 49026
rect 18898 48974 18910 49026
rect 22866 48974 22878 49026
rect 22930 48974 22942 49026
rect 23314 48974 23326 49026
rect 23378 48974 23390 49026
rect 24322 48974 24334 49026
rect 24386 48974 24398 49026
rect 27010 48974 27022 49026
rect 27074 48974 27086 49026
rect 32834 48974 32846 49026
rect 32898 48974 32910 49026
rect 18510 48962 18562 48974
rect 31278 48962 31330 48974
rect 33070 48962 33122 48974
rect 33630 49026 33682 49038
rect 33630 48962 33682 48974
rect 5630 48914 5682 48926
rect 5630 48850 5682 48862
rect 12798 48914 12850 48926
rect 12798 48850 12850 48862
rect 13582 48914 13634 48926
rect 13582 48850 13634 48862
rect 17950 48914 18002 48926
rect 17950 48850 18002 48862
rect 18622 48914 18674 48926
rect 31614 48914 31666 48926
rect 26898 48862 26910 48914
rect 26962 48862 26974 48914
rect 18622 48850 18674 48862
rect 31614 48850 31666 48862
rect 5742 48802 5794 48814
rect 10334 48802 10386 48814
rect 9762 48750 9774 48802
rect 9826 48750 9838 48802
rect 5742 48738 5794 48750
rect 10334 48738 10386 48750
rect 11790 48802 11842 48814
rect 11790 48738 11842 48750
rect 13694 48802 13746 48814
rect 13694 48738 13746 48750
rect 19630 48802 19682 48814
rect 19630 48738 19682 48750
rect 22318 48802 22370 48814
rect 22318 48738 22370 48750
rect 28590 48802 28642 48814
rect 28590 48738 28642 48750
rect 31838 48802 31890 48814
rect 31838 48738 31890 48750
rect 33742 48802 33794 48814
rect 33742 48738 33794 48750
rect 34302 48802 34354 48814
rect 34302 48738 34354 48750
rect 1344 48634 38640 48668
rect 1344 48582 14024 48634
rect 14076 48582 14148 48634
rect 14200 48582 14272 48634
rect 14324 48582 14396 48634
rect 14448 48582 14520 48634
rect 14572 48582 14644 48634
rect 14696 48582 14768 48634
rect 14820 48582 14892 48634
rect 14944 48582 15016 48634
rect 15068 48582 15140 48634
rect 15192 48582 34024 48634
rect 34076 48582 34148 48634
rect 34200 48582 34272 48634
rect 34324 48582 34396 48634
rect 34448 48582 34520 48634
rect 34572 48582 34644 48634
rect 34696 48582 34768 48634
rect 34820 48582 34892 48634
rect 34944 48582 35016 48634
rect 35068 48582 35140 48634
rect 35192 48582 38640 48634
rect 1344 48548 38640 48582
rect 7534 48466 7586 48478
rect 6402 48414 6414 48466
rect 6466 48414 6478 48466
rect 7534 48402 7586 48414
rect 7646 48466 7698 48478
rect 7646 48402 7698 48414
rect 8542 48466 8594 48478
rect 8542 48402 8594 48414
rect 11006 48466 11058 48478
rect 15150 48466 15202 48478
rect 14578 48414 14590 48466
rect 14642 48414 14654 48466
rect 11006 48402 11058 48414
rect 15150 48402 15202 48414
rect 15486 48466 15538 48478
rect 15486 48402 15538 48414
rect 24446 48466 24498 48478
rect 24446 48402 24498 48414
rect 25342 48466 25394 48478
rect 25342 48402 25394 48414
rect 26238 48466 26290 48478
rect 26238 48402 26290 48414
rect 26686 48466 26738 48478
rect 30830 48466 30882 48478
rect 30146 48414 30158 48466
rect 30210 48414 30222 48466
rect 26686 48402 26738 48414
rect 30830 48402 30882 48414
rect 32510 48466 32562 48478
rect 36418 48414 36430 48466
rect 36482 48414 36494 48466
rect 32510 48402 32562 48414
rect 7870 48354 7922 48366
rect 5730 48302 5742 48354
rect 5794 48302 5806 48354
rect 7870 48290 7922 48302
rect 19070 48354 19122 48366
rect 19070 48290 19122 48302
rect 23662 48354 23714 48366
rect 23662 48290 23714 48302
rect 2494 48242 2546 48254
rect 7422 48242 7474 48254
rect 2930 48190 2942 48242
rect 2994 48190 3006 48242
rect 6962 48190 6974 48242
rect 7026 48190 7038 48242
rect 2494 48178 2546 48190
rect 7422 48178 7474 48190
rect 9998 48242 10050 48254
rect 9998 48178 10050 48190
rect 11678 48242 11730 48254
rect 15934 48242 15986 48254
rect 20974 48242 21026 48254
rect 27358 48242 27410 48254
rect 31166 48242 31218 48254
rect 12114 48190 12126 48242
rect 12178 48190 12190 48242
rect 18498 48190 18510 48242
rect 18562 48190 18574 48242
rect 21410 48190 21422 48242
rect 21474 48190 21486 48242
rect 27682 48190 27694 48242
rect 27746 48190 27758 48242
rect 11678 48178 11730 48190
rect 15934 48178 15986 48190
rect 20974 48178 21026 48190
rect 27358 48178 27410 48190
rect 31166 48178 31218 48190
rect 31838 48242 31890 48254
rect 31838 48178 31890 48190
rect 33070 48242 33122 48254
rect 33070 48178 33122 48190
rect 33742 48242 33794 48254
rect 34066 48190 34078 48242
rect 34130 48190 34142 48242
rect 33742 48178 33794 48190
rect 4622 48130 4674 48142
rect 3266 48078 3278 48130
rect 3330 48078 3342 48130
rect 4622 48066 4674 48078
rect 8990 48130 9042 48142
rect 8990 48066 9042 48078
rect 9886 48130 9938 48142
rect 9886 48066 9938 48078
rect 16718 48130 16770 48142
rect 16718 48066 16770 48078
rect 17838 48130 17890 48142
rect 25790 48130 25842 48142
rect 18162 48078 18174 48130
rect 18226 48078 18238 48130
rect 17838 48066 17890 48078
rect 25790 48066 25842 48078
rect 31614 48018 31666 48030
rect 9762 47966 9774 48018
rect 9826 47966 9838 48018
rect 31614 47954 31666 47966
rect 32174 48018 32226 48030
rect 32174 47954 32226 47966
rect 32398 48018 32450 48030
rect 32398 47954 32450 47966
rect 33182 48018 33234 48030
rect 33182 47954 33234 47966
rect 37214 48018 37266 48030
rect 37214 47954 37266 47966
rect 1344 47850 38640 47884
rect 1344 47798 4024 47850
rect 4076 47798 4148 47850
rect 4200 47798 4272 47850
rect 4324 47798 4396 47850
rect 4448 47798 4520 47850
rect 4572 47798 4644 47850
rect 4696 47798 4768 47850
rect 4820 47798 4892 47850
rect 4944 47798 5016 47850
rect 5068 47798 5140 47850
rect 5192 47798 24024 47850
rect 24076 47798 24148 47850
rect 24200 47798 24272 47850
rect 24324 47798 24396 47850
rect 24448 47798 24520 47850
rect 24572 47798 24644 47850
rect 24696 47798 24768 47850
rect 24820 47798 24892 47850
rect 24944 47798 25016 47850
rect 25068 47798 25140 47850
rect 25192 47798 38640 47850
rect 1344 47764 38640 47798
rect 22990 47682 23042 47694
rect 9874 47630 9886 47682
rect 9938 47630 9950 47682
rect 22990 47618 23042 47630
rect 13582 47570 13634 47582
rect 3266 47518 3278 47570
rect 3330 47518 3342 47570
rect 6290 47518 6302 47570
rect 6354 47518 6366 47570
rect 13582 47506 13634 47518
rect 22094 47570 22146 47582
rect 22094 47506 22146 47518
rect 29262 47570 29314 47582
rect 31390 47570 31442 47582
rect 30706 47518 30718 47570
rect 30770 47518 30782 47570
rect 29262 47506 29314 47518
rect 31390 47506 31442 47518
rect 4622 47458 4674 47470
rect 4622 47394 4674 47406
rect 4846 47458 4898 47470
rect 4846 47394 4898 47406
rect 5182 47458 5234 47470
rect 7758 47458 7810 47470
rect 13694 47458 13746 47470
rect 17614 47458 17666 47470
rect 23214 47458 23266 47470
rect 7074 47406 7086 47458
rect 7138 47406 7150 47458
rect 10994 47406 11006 47458
rect 11058 47406 11070 47458
rect 14690 47406 14702 47458
rect 14754 47406 14766 47458
rect 22530 47406 22542 47458
rect 22594 47406 22606 47458
rect 5182 47394 5234 47406
rect 7758 47394 7810 47406
rect 13694 47394 13746 47406
rect 17614 47394 17666 47406
rect 23214 47394 23266 47406
rect 23326 47458 23378 47470
rect 23326 47394 23378 47406
rect 23662 47458 23714 47470
rect 23662 47394 23714 47406
rect 24446 47458 24498 47470
rect 31278 47458 31330 47470
rect 24770 47406 24782 47458
rect 24834 47406 24846 47458
rect 31042 47406 31054 47458
rect 31106 47406 31118 47458
rect 24446 47394 24498 47406
rect 31278 47394 31330 47406
rect 31502 47458 31554 47470
rect 36318 47458 36370 47470
rect 31714 47406 31726 47458
rect 31778 47406 31790 47458
rect 32610 47406 32622 47458
rect 32674 47406 32686 47458
rect 31502 47394 31554 47406
rect 36318 47394 36370 47406
rect 37550 47458 37602 47470
rect 37550 47394 37602 47406
rect 2606 47346 2658 47358
rect 2606 47282 2658 47294
rect 3726 47346 3778 47358
rect 3726 47282 3778 47294
rect 4062 47346 4114 47358
rect 7422 47346 7474 47358
rect 6066 47294 6078 47346
rect 6130 47294 6142 47346
rect 4062 47282 4114 47294
rect 7422 47282 7474 47294
rect 9102 47346 9154 47358
rect 13918 47346 13970 47358
rect 11218 47294 11230 47346
rect 11282 47294 11294 47346
rect 9102 47282 9154 47294
rect 13918 47282 13970 47294
rect 22878 47346 22930 47358
rect 22878 47282 22930 47294
rect 23886 47346 23938 47358
rect 23886 47282 23938 47294
rect 23998 47346 24050 47358
rect 23998 47282 24050 47294
rect 30382 47346 30434 47358
rect 30382 47282 30434 47294
rect 33182 47346 33234 47358
rect 33182 47282 33234 47294
rect 35758 47346 35810 47358
rect 35758 47282 35810 47294
rect 2158 47234 2210 47246
rect 2158 47170 2210 47182
rect 2830 47234 2882 47246
rect 2830 47170 2882 47182
rect 4958 47234 5010 47246
rect 4958 47170 5010 47182
rect 7534 47234 7586 47246
rect 7534 47170 7586 47182
rect 8094 47234 8146 47246
rect 8094 47170 8146 47182
rect 9438 47234 9490 47246
rect 9438 47170 9490 47182
rect 12350 47234 12402 47246
rect 12350 47170 12402 47182
rect 13470 47234 13522 47246
rect 13470 47170 13522 47182
rect 15598 47234 15650 47246
rect 15598 47170 15650 47182
rect 21646 47234 21698 47246
rect 21646 47170 21698 47182
rect 21982 47234 22034 47246
rect 21982 47170 22034 47182
rect 22206 47234 22258 47246
rect 27918 47234 27970 47246
rect 27122 47182 27134 47234
rect 27186 47182 27198 47234
rect 22206 47170 22258 47182
rect 27918 47170 27970 47182
rect 28366 47234 28418 47246
rect 28366 47170 28418 47182
rect 30158 47234 30210 47246
rect 30158 47170 30210 47182
rect 30606 47234 30658 47246
rect 30606 47170 30658 47182
rect 32174 47234 32226 47246
rect 37102 47234 37154 47246
rect 33618 47182 33630 47234
rect 33682 47182 33694 47234
rect 32174 47170 32226 47182
rect 37102 47170 37154 47182
rect 37998 47234 38050 47246
rect 37998 47170 38050 47182
rect 1344 47066 38640 47100
rect 1344 47014 14024 47066
rect 14076 47014 14148 47066
rect 14200 47014 14272 47066
rect 14324 47014 14396 47066
rect 14448 47014 14520 47066
rect 14572 47014 14644 47066
rect 14696 47014 14768 47066
rect 14820 47014 14892 47066
rect 14944 47014 15016 47066
rect 15068 47014 15140 47066
rect 15192 47014 34024 47066
rect 34076 47014 34148 47066
rect 34200 47014 34272 47066
rect 34324 47014 34396 47066
rect 34448 47014 34520 47066
rect 34572 47014 34644 47066
rect 34696 47014 34768 47066
rect 34820 47014 34892 47066
rect 34944 47014 35016 47066
rect 35068 47014 35140 47066
rect 35192 47014 38640 47066
rect 1344 46980 38640 47014
rect 5518 46898 5570 46910
rect 4834 46846 4846 46898
rect 4898 46846 4910 46898
rect 5518 46834 5570 46846
rect 6078 46898 6130 46910
rect 15374 46898 15426 46910
rect 10770 46846 10782 46898
rect 10834 46846 10846 46898
rect 6078 46834 6130 46846
rect 15374 46834 15426 46846
rect 18958 46898 19010 46910
rect 18958 46834 19010 46846
rect 25342 46898 25394 46910
rect 25342 46834 25394 46846
rect 26462 46898 26514 46910
rect 26462 46834 26514 46846
rect 27134 46898 27186 46910
rect 27134 46834 27186 46846
rect 29598 46898 29650 46910
rect 29598 46834 29650 46846
rect 30606 46898 30658 46910
rect 30606 46834 30658 46846
rect 31166 46898 31218 46910
rect 31166 46834 31218 46846
rect 31390 46898 31442 46910
rect 31390 46834 31442 46846
rect 32174 46898 32226 46910
rect 32174 46834 32226 46846
rect 34078 46898 34130 46910
rect 34078 46834 34130 46846
rect 36542 46898 36594 46910
rect 36542 46834 36594 46846
rect 5742 46786 5794 46798
rect 5742 46722 5794 46734
rect 5854 46786 5906 46798
rect 5854 46722 5906 46734
rect 6414 46786 6466 46798
rect 31614 46786 31666 46798
rect 11442 46734 11454 46786
rect 11506 46734 11518 46786
rect 28018 46734 28030 46786
rect 28082 46734 28094 46786
rect 6414 46722 6466 46734
rect 31614 46722 31666 46734
rect 34526 46786 34578 46798
rect 34526 46722 34578 46734
rect 1822 46674 1874 46686
rect 9998 46674 10050 46686
rect 17502 46674 17554 46686
rect 26238 46674 26290 46686
rect 2482 46622 2494 46674
rect 2546 46622 2558 46674
rect 11778 46622 11790 46674
rect 11842 46622 11854 46674
rect 19282 46622 19294 46674
rect 19346 46622 19358 46674
rect 1822 46610 1874 46622
rect 9998 46610 10050 46622
rect 17502 46610 17554 46622
rect 26238 46610 26290 46622
rect 26574 46674 26626 46686
rect 28702 46674 28754 46686
rect 32286 46674 32338 46686
rect 27906 46622 27918 46674
rect 27970 46622 27982 46674
rect 30930 46622 30942 46674
rect 30994 46622 31006 46674
rect 26574 46610 26626 46622
rect 28702 46610 28754 46622
rect 32286 46610 32338 46622
rect 34190 46674 34242 46686
rect 34190 46610 34242 46622
rect 34638 46674 34690 46686
rect 36206 46674 36258 46686
rect 35186 46622 35198 46674
rect 35250 46622 35262 46674
rect 35970 46622 35982 46674
rect 36034 46622 36046 46674
rect 34638 46610 34690 46622
rect 36206 46610 36258 46622
rect 37102 46674 37154 46686
rect 37102 46610 37154 46622
rect 6974 46562 7026 46574
rect 6974 46498 7026 46510
rect 7310 46562 7362 46574
rect 7310 46498 7362 46510
rect 7758 46562 7810 46574
rect 7758 46498 7810 46510
rect 8206 46562 8258 46574
rect 8206 46498 8258 46510
rect 9102 46562 9154 46574
rect 9102 46498 9154 46510
rect 13134 46562 13186 46574
rect 13134 46498 13186 46510
rect 13582 46562 13634 46574
rect 13582 46498 13634 46510
rect 14030 46562 14082 46574
rect 14030 46498 14082 46510
rect 14478 46562 14530 46574
rect 26014 46562 26066 46574
rect 23762 46510 23774 46562
rect 23826 46510 23838 46562
rect 14478 46498 14530 46510
rect 26014 46498 26066 46510
rect 27470 46562 27522 46574
rect 27470 46498 27522 46510
rect 30158 46562 30210 46574
rect 30158 46498 30210 46510
rect 31278 46562 31330 46574
rect 31278 46498 31330 46510
rect 33182 46562 33234 46574
rect 33182 46498 33234 46510
rect 33630 46562 33682 46574
rect 33630 46498 33682 46510
rect 37550 46562 37602 46574
rect 37550 46498 37602 46510
rect 37998 46562 38050 46574
rect 37998 46498 38050 46510
rect 29038 46450 29090 46462
rect 7746 46398 7758 46450
rect 7810 46447 7822 46450
rect 7970 46447 7982 46450
rect 7810 46401 7982 46447
rect 7810 46398 7822 46401
rect 7970 46398 7982 46401
rect 8034 46398 8046 46450
rect 13458 46398 13470 46450
rect 13522 46447 13534 46450
rect 14018 46447 14030 46450
rect 13522 46401 14030 46447
rect 13522 46398 13534 46401
rect 14018 46398 14030 46401
rect 14082 46447 14094 46450
rect 14466 46447 14478 46450
rect 14082 46401 14478 46447
rect 14082 46398 14094 46401
rect 14466 46398 14478 46401
rect 14530 46398 14542 46450
rect 29038 46386 29090 46398
rect 1344 46282 38640 46316
rect 1344 46230 4024 46282
rect 4076 46230 4148 46282
rect 4200 46230 4272 46282
rect 4324 46230 4396 46282
rect 4448 46230 4520 46282
rect 4572 46230 4644 46282
rect 4696 46230 4768 46282
rect 4820 46230 4892 46282
rect 4944 46230 5016 46282
rect 5068 46230 5140 46282
rect 5192 46230 24024 46282
rect 24076 46230 24148 46282
rect 24200 46230 24272 46282
rect 24324 46230 24396 46282
rect 24448 46230 24520 46282
rect 24572 46230 24644 46282
rect 24696 46230 24768 46282
rect 24820 46230 24892 46282
rect 24944 46230 25016 46282
rect 25068 46230 25140 46282
rect 25192 46230 38640 46282
rect 1344 46196 38640 46230
rect 3838 46114 3890 46126
rect 3838 46050 3890 46062
rect 17278 46114 17330 46126
rect 17278 46050 17330 46062
rect 22318 46114 22370 46126
rect 22318 46050 22370 46062
rect 30158 46114 30210 46126
rect 34738 46062 34750 46114
rect 34802 46062 34814 46114
rect 30158 46050 30210 46062
rect 2494 46002 2546 46014
rect 5742 46002 5794 46014
rect 3266 45950 3278 46002
rect 3330 45950 3342 46002
rect 2494 45938 2546 45950
rect 5742 45938 5794 45950
rect 6862 46002 6914 46014
rect 16046 46002 16098 46014
rect 18286 46002 18338 46014
rect 12338 45950 12350 46002
rect 12402 45950 12414 46002
rect 16818 45950 16830 46002
rect 16882 45950 16894 46002
rect 6862 45938 6914 45950
rect 16046 45938 16098 45950
rect 18286 45938 18338 45950
rect 20302 46002 20354 46014
rect 20302 45938 20354 45950
rect 20750 46002 20802 46014
rect 20750 45938 20802 45950
rect 22766 46002 22818 46014
rect 24222 46002 24274 46014
rect 23538 45950 23550 46002
rect 23602 45950 23614 46002
rect 22766 45938 22818 45950
rect 24222 45938 24274 45950
rect 35534 46002 35586 46014
rect 35534 45938 35586 45950
rect 37550 46002 37602 46014
rect 37550 45938 37602 45950
rect 37998 46002 38050 46014
rect 37998 45938 38050 45950
rect 2830 45890 2882 45902
rect 2830 45826 2882 45838
rect 4174 45890 4226 45902
rect 4174 45826 4226 45838
rect 7310 45890 7362 45902
rect 10894 45890 10946 45902
rect 17502 45890 17554 45902
rect 7634 45838 7646 45890
rect 7698 45838 7710 45890
rect 11778 45838 11790 45890
rect 11842 45838 11854 45890
rect 13794 45838 13806 45890
rect 13858 45838 13870 45890
rect 16594 45838 16606 45890
rect 16658 45838 16670 45890
rect 7310 45826 7362 45838
rect 10894 45826 10946 45838
rect 17502 45826 17554 45838
rect 21310 45890 21362 45902
rect 21310 45826 21362 45838
rect 21982 45890 22034 45902
rect 21982 45826 22034 45838
rect 22206 45890 22258 45902
rect 24782 45890 24834 45902
rect 37102 45890 37154 45902
rect 23426 45838 23438 45890
rect 23490 45838 23502 45890
rect 25106 45838 25118 45890
rect 25170 45838 25182 45890
rect 25666 45838 25678 45890
rect 25730 45838 25742 45890
rect 30370 45838 30382 45890
rect 30434 45838 30446 45890
rect 31042 45838 31054 45890
rect 31106 45838 31118 45890
rect 33170 45838 33182 45890
rect 33234 45838 33246 45890
rect 35746 45838 35758 45890
rect 35810 45838 35822 45890
rect 22206 45826 22258 45838
rect 24782 45826 24834 45838
rect 37102 45826 37154 45838
rect 18062 45778 18114 45790
rect 4386 45726 4398 45778
rect 4450 45726 4462 45778
rect 4946 45726 4958 45778
rect 5010 45726 5022 45778
rect 11442 45726 11454 45778
rect 11506 45726 11518 45778
rect 13682 45726 13694 45778
rect 13746 45726 13758 45778
rect 17826 45726 17838 45778
rect 17890 45726 17902 45778
rect 18062 45714 18114 45726
rect 28702 45778 28754 45790
rect 28702 45714 28754 45726
rect 30046 45778 30098 45790
rect 30046 45714 30098 45726
rect 36990 45778 37042 45790
rect 36990 45714 37042 45726
rect 6526 45666 6578 45678
rect 15374 45666 15426 45678
rect 9986 45614 9998 45666
rect 10050 45614 10062 45666
rect 13570 45614 13582 45666
rect 13634 45614 13646 45666
rect 6526 45602 6578 45614
rect 15374 45602 15426 45614
rect 18734 45666 18786 45678
rect 18734 45602 18786 45614
rect 19294 45666 19346 45678
rect 19294 45602 19346 45614
rect 21422 45666 21474 45678
rect 21422 45602 21474 45614
rect 21534 45666 21586 45678
rect 21534 45602 21586 45614
rect 22318 45666 22370 45678
rect 22318 45602 22370 45614
rect 24110 45666 24162 45678
rect 24110 45602 24162 45614
rect 24334 45666 24386 45678
rect 29262 45666 29314 45678
rect 28130 45614 28142 45666
rect 28194 45614 28206 45666
rect 24334 45602 24386 45614
rect 29262 45602 29314 45614
rect 29710 45666 29762 45678
rect 29710 45602 29762 45614
rect 35982 45666 36034 45678
rect 35982 45602 36034 45614
rect 1344 45498 38640 45532
rect 1344 45446 14024 45498
rect 14076 45446 14148 45498
rect 14200 45446 14272 45498
rect 14324 45446 14396 45498
rect 14448 45446 14520 45498
rect 14572 45446 14644 45498
rect 14696 45446 14768 45498
rect 14820 45446 14892 45498
rect 14944 45446 15016 45498
rect 15068 45446 15140 45498
rect 15192 45446 34024 45498
rect 34076 45446 34148 45498
rect 34200 45446 34272 45498
rect 34324 45446 34396 45498
rect 34448 45446 34520 45498
rect 34572 45446 34644 45498
rect 34696 45446 34768 45498
rect 34820 45446 34892 45498
rect 34944 45446 35016 45498
rect 35068 45446 35140 45498
rect 35192 45446 38640 45498
rect 1344 45412 38640 45446
rect 7646 45330 7698 45342
rect 7646 45266 7698 45278
rect 10894 45330 10946 45342
rect 10894 45266 10946 45278
rect 11342 45330 11394 45342
rect 11342 45266 11394 45278
rect 12686 45330 12738 45342
rect 12686 45266 12738 45278
rect 13134 45330 13186 45342
rect 13134 45266 13186 45278
rect 13694 45330 13746 45342
rect 13694 45266 13746 45278
rect 14926 45330 14978 45342
rect 14926 45266 14978 45278
rect 16382 45330 16434 45342
rect 16382 45266 16434 45278
rect 19630 45330 19682 45342
rect 23550 45330 23602 45342
rect 22978 45278 22990 45330
rect 23042 45278 23054 45330
rect 19630 45266 19682 45278
rect 23550 45266 23602 45278
rect 24334 45330 24386 45342
rect 24334 45266 24386 45278
rect 25902 45330 25954 45342
rect 25902 45266 25954 45278
rect 27806 45330 27858 45342
rect 31154 45278 31166 45330
rect 31218 45278 31230 45330
rect 27806 45266 27858 45278
rect 5630 45218 5682 45230
rect 11790 45218 11842 45230
rect 6514 45166 6526 45218
rect 6578 45166 6590 45218
rect 5630 45154 5682 45166
rect 11790 45154 11842 45166
rect 16718 45218 16770 45230
rect 16718 45154 16770 45166
rect 17390 45218 17442 45230
rect 17390 45154 17442 45166
rect 34190 45218 34242 45230
rect 34190 45154 34242 45166
rect 34414 45218 34466 45230
rect 34414 45154 34466 45166
rect 34862 45218 34914 45230
rect 36978 45166 36990 45218
rect 37042 45166 37054 45218
rect 34862 45154 34914 45166
rect 2830 45106 2882 45118
rect 8430 45106 8482 45118
rect 6402 45054 6414 45106
rect 6466 45054 6478 45106
rect 7634 45054 7646 45106
rect 7698 45054 7710 45106
rect 8194 45054 8206 45106
rect 8258 45054 8270 45106
rect 2830 45042 2882 45054
rect 8430 45042 8482 45054
rect 9662 45106 9714 45118
rect 9662 45042 9714 45054
rect 13806 45106 13858 45118
rect 13806 45042 13858 45054
rect 14142 45106 14194 45118
rect 14142 45042 14194 45054
rect 14478 45106 14530 45118
rect 14478 45042 14530 45054
rect 15150 45106 15202 45118
rect 15150 45042 15202 45054
rect 17726 45106 17778 45118
rect 17726 45042 17778 45054
rect 17950 45106 18002 45118
rect 20078 45106 20130 45118
rect 25790 45106 25842 45118
rect 18274 45054 18286 45106
rect 18338 45054 18350 45106
rect 20514 45054 20526 45106
rect 20578 45054 20590 45106
rect 17950 45042 18002 45054
rect 20078 45042 20130 45054
rect 25790 45042 25842 45054
rect 26126 45106 26178 45118
rect 26126 45042 26178 45054
rect 26350 45106 26402 45118
rect 26350 45042 26402 45054
rect 27694 45106 27746 45118
rect 27694 45042 27746 45054
rect 30830 45106 30882 45118
rect 30830 45042 30882 45054
rect 34638 45106 34690 45118
rect 34638 45042 34690 45054
rect 35422 45106 35474 45118
rect 36306 45054 36318 45106
rect 36370 45054 36382 45106
rect 35422 45042 35474 45054
rect 2494 44994 2546 45006
rect 5294 44994 5346 45006
rect 3266 44942 3278 44994
rect 3330 44942 3342 44994
rect 2494 44930 2546 44942
rect 5294 44930 5346 44942
rect 7310 44994 7362 45006
rect 7310 44930 7362 44942
rect 8878 44994 8930 45006
rect 8878 44930 8930 44942
rect 10446 44994 10498 45006
rect 10446 44930 10498 44942
rect 14030 44994 14082 45006
rect 15934 44994 15986 45006
rect 14802 44942 14814 44994
rect 14866 44942 14878 44994
rect 14030 44930 14082 44942
rect 15934 44930 15986 44942
rect 16830 44994 16882 45006
rect 16830 44930 16882 44942
rect 17502 44994 17554 45006
rect 17502 44930 17554 44942
rect 19294 44994 19346 45006
rect 19294 44930 19346 44942
rect 19518 44994 19570 45006
rect 19518 44930 19570 44942
rect 23886 44994 23938 45006
rect 23886 44930 23938 44942
rect 25454 44994 25506 45006
rect 25454 44930 25506 44942
rect 27246 44994 27298 45006
rect 27246 44930 27298 44942
rect 27582 44994 27634 45006
rect 27582 44930 27634 44942
rect 29934 44994 29986 45006
rect 29934 44930 29986 44942
rect 30606 44994 30658 45006
rect 30606 44930 30658 44942
rect 32510 44994 32562 45006
rect 32510 44930 32562 44942
rect 33854 44994 33906 45006
rect 33854 44930 33906 44942
rect 5966 44882 6018 44894
rect 5966 44818 6018 44830
rect 7982 44882 8034 44894
rect 18286 44882 18338 44894
rect 10434 44830 10446 44882
rect 10498 44879 10510 44882
rect 11442 44879 11454 44882
rect 10498 44833 11454 44879
rect 10498 44830 10510 44833
rect 11442 44830 11454 44833
rect 11506 44830 11518 44882
rect 7982 44818 8034 44830
rect 18286 44818 18338 44830
rect 18622 44882 18674 44894
rect 18622 44818 18674 44830
rect 34750 44882 34802 44894
rect 34750 44818 34802 44830
rect 37662 44882 37714 44894
rect 37662 44818 37714 44830
rect 1344 44714 38640 44748
rect 1344 44662 4024 44714
rect 4076 44662 4148 44714
rect 4200 44662 4272 44714
rect 4324 44662 4396 44714
rect 4448 44662 4520 44714
rect 4572 44662 4644 44714
rect 4696 44662 4768 44714
rect 4820 44662 4892 44714
rect 4944 44662 5016 44714
rect 5068 44662 5140 44714
rect 5192 44662 24024 44714
rect 24076 44662 24148 44714
rect 24200 44662 24272 44714
rect 24324 44662 24396 44714
rect 24448 44662 24520 44714
rect 24572 44662 24644 44714
rect 24696 44662 24768 44714
rect 24820 44662 24892 44714
rect 24944 44662 25016 44714
rect 25068 44662 25140 44714
rect 25192 44662 38640 44714
rect 1344 44628 38640 44662
rect 7646 44546 7698 44558
rect 7646 44482 7698 44494
rect 8206 44546 8258 44558
rect 8206 44482 8258 44494
rect 8542 44546 8594 44558
rect 8542 44482 8594 44494
rect 17054 44546 17106 44558
rect 17054 44482 17106 44494
rect 35982 44546 36034 44558
rect 35982 44482 36034 44494
rect 7534 44434 7586 44446
rect 6738 44382 6750 44434
rect 6802 44382 6814 44434
rect 7534 44370 7586 44382
rect 9662 44434 9714 44446
rect 9662 44370 9714 44382
rect 10558 44434 10610 44446
rect 10558 44370 10610 44382
rect 12238 44434 12290 44446
rect 12238 44370 12290 44382
rect 12910 44434 12962 44446
rect 18510 44434 18562 44446
rect 17602 44382 17614 44434
rect 17666 44382 17678 44434
rect 12910 44370 12962 44382
rect 18510 44370 18562 44382
rect 18622 44434 18674 44446
rect 18622 44370 18674 44382
rect 19070 44434 19122 44446
rect 19070 44370 19122 44382
rect 20302 44434 20354 44446
rect 20302 44370 20354 44382
rect 21758 44434 21810 44446
rect 21758 44370 21810 44382
rect 34190 44434 34242 44446
rect 34190 44370 34242 44382
rect 4174 44322 4226 44334
rect 8318 44322 8370 44334
rect 17726 44322 17778 44334
rect 7298 44270 7310 44322
rect 7362 44270 7374 44322
rect 8754 44270 8766 44322
rect 8818 44270 8830 44322
rect 13458 44270 13470 44322
rect 13522 44270 13534 44322
rect 14018 44270 14030 44322
rect 14082 44270 14094 44322
rect 4174 44258 4226 44270
rect 8318 44258 8370 44270
rect 17726 44258 17778 44270
rect 18062 44322 18114 44334
rect 18062 44258 18114 44270
rect 21310 44322 21362 44334
rect 21310 44258 21362 44270
rect 21982 44322 22034 44334
rect 21982 44258 22034 44270
rect 34526 44322 34578 44334
rect 37438 44322 37490 44334
rect 35298 44270 35310 44322
rect 35362 44270 35374 44322
rect 34526 44258 34578 44270
rect 37438 44258 37490 44270
rect 37550 44322 37602 44334
rect 37550 44258 37602 44270
rect 6414 44210 6466 44222
rect 4386 44158 4398 44210
rect 4450 44158 4462 44210
rect 4946 44158 4958 44210
rect 5010 44158 5022 44210
rect 6414 44146 6466 44158
rect 11342 44210 11394 44222
rect 11342 44146 11394 44158
rect 11454 44210 11506 44222
rect 11454 44146 11506 44158
rect 17614 44210 17666 44222
rect 17614 44146 17666 44158
rect 20414 44210 20466 44222
rect 20414 44146 20466 44158
rect 21534 44210 21586 44222
rect 21534 44146 21586 44158
rect 34638 44210 34690 44222
rect 34638 44146 34690 44158
rect 34862 44210 34914 44222
rect 37662 44210 37714 44222
rect 35186 44158 35198 44210
rect 35250 44158 35262 44210
rect 34862 44146 34914 44158
rect 37662 44146 37714 44158
rect 3838 44098 3890 44110
rect 3838 44034 3890 44046
rect 6638 44098 6690 44110
rect 6638 44034 6690 44046
rect 9214 44098 9266 44110
rect 9214 44034 9266 44046
rect 10110 44098 10162 44110
rect 10110 44034 10162 44046
rect 11006 44098 11058 44110
rect 11006 44034 11058 44046
rect 11678 44098 11730 44110
rect 17950 44098 18002 44110
rect 16258 44046 16270 44098
rect 16322 44046 16334 44098
rect 11678 44034 11730 44046
rect 17950 44034 18002 44046
rect 18958 44098 19010 44110
rect 18958 44034 19010 44046
rect 19742 44098 19794 44110
rect 19742 44034 19794 44046
rect 20190 44098 20242 44110
rect 20190 44034 20242 44046
rect 23662 44098 23714 44110
rect 23662 44034 23714 44046
rect 24110 44098 24162 44110
rect 24110 44034 24162 44046
rect 33854 44098 33906 44110
rect 33854 44034 33906 44046
rect 36318 44098 36370 44110
rect 36978 44046 36990 44098
rect 37042 44046 37054 44098
rect 36318 44034 36370 44046
rect 1344 43930 38640 43964
rect 1344 43878 14024 43930
rect 14076 43878 14148 43930
rect 14200 43878 14272 43930
rect 14324 43878 14396 43930
rect 14448 43878 14520 43930
rect 14572 43878 14644 43930
rect 14696 43878 14768 43930
rect 14820 43878 14892 43930
rect 14944 43878 15016 43930
rect 15068 43878 15140 43930
rect 15192 43878 34024 43930
rect 34076 43878 34148 43930
rect 34200 43878 34272 43930
rect 34324 43878 34396 43930
rect 34448 43878 34520 43930
rect 34572 43878 34644 43930
rect 34696 43878 34768 43930
rect 34820 43878 34892 43930
rect 34944 43878 35016 43930
rect 35068 43878 35140 43930
rect 35192 43878 38640 43930
rect 1344 43844 38640 43878
rect 5294 43762 5346 43774
rect 4722 43710 4734 43762
rect 4786 43710 4798 43762
rect 5294 43698 5346 43710
rect 6078 43762 6130 43774
rect 6078 43698 6130 43710
rect 8766 43762 8818 43774
rect 8766 43698 8818 43710
rect 10670 43762 10722 43774
rect 10670 43698 10722 43710
rect 15822 43762 15874 43774
rect 15822 43698 15874 43710
rect 16718 43762 16770 43774
rect 16718 43698 16770 43710
rect 17614 43762 17666 43774
rect 17614 43698 17666 43710
rect 17726 43762 17778 43774
rect 17726 43698 17778 43710
rect 18734 43762 18786 43774
rect 18734 43698 18786 43710
rect 18846 43762 18898 43774
rect 18846 43698 18898 43710
rect 19966 43762 20018 43774
rect 19966 43698 20018 43710
rect 20414 43762 20466 43774
rect 20414 43698 20466 43710
rect 20974 43762 21026 43774
rect 20974 43698 21026 43710
rect 30270 43762 30322 43774
rect 30270 43698 30322 43710
rect 35198 43762 35250 43774
rect 36530 43710 36542 43762
rect 36594 43710 36606 43762
rect 35198 43698 35250 43710
rect 5630 43650 5682 43662
rect 5630 43586 5682 43598
rect 12350 43650 12402 43662
rect 12350 43586 12402 43598
rect 12798 43650 12850 43662
rect 12798 43586 12850 43598
rect 13918 43650 13970 43662
rect 13918 43586 13970 43598
rect 14254 43650 14306 43662
rect 14254 43586 14306 43598
rect 15486 43650 15538 43662
rect 15486 43586 15538 43598
rect 16494 43650 16546 43662
rect 16494 43586 16546 43598
rect 19742 43650 19794 43662
rect 19742 43586 19794 43598
rect 29150 43650 29202 43662
rect 29150 43586 29202 43598
rect 29822 43650 29874 43662
rect 35858 43598 35870 43650
rect 35922 43598 35934 43650
rect 36418 43598 36430 43650
rect 36482 43598 36494 43650
rect 29822 43586 29874 43598
rect 1822 43538 1874 43550
rect 14142 43538 14194 43550
rect 2258 43486 2270 43538
rect 2322 43486 2334 43538
rect 8530 43486 8542 43538
rect 8594 43486 8606 43538
rect 11442 43486 11454 43538
rect 11506 43486 11518 43538
rect 12562 43486 12574 43538
rect 12626 43486 12638 43538
rect 1822 43474 1874 43486
rect 14142 43474 14194 43486
rect 14478 43538 14530 43550
rect 16382 43538 16434 43550
rect 16146 43486 16158 43538
rect 16210 43486 16222 43538
rect 14478 43474 14530 43486
rect 16382 43474 16434 43486
rect 16606 43538 16658 43550
rect 17838 43538 17890 43550
rect 18622 43538 18674 43550
rect 17378 43486 17390 43538
rect 17442 43486 17454 43538
rect 18050 43486 18062 43538
rect 18114 43486 18126 43538
rect 18386 43486 18398 43538
rect 18450 43486 18462 43538
rect 16606 43474 16658 43486
rect 17838 43474 17890 43486
rect 18622 43474 18674 43486
rect 18958 43538 19010 43550
rect 18958 43474 19010 43486
rect 19294 43538 19346 43550
rect 36766 43538 36818 43550
rect 30146 43486 30158 43538
rect 30210 43486 30222 43538
rect 30482 43486 30494 43538
rect 30546 43486 30558 43538
rect 19294 43474 19346 43486
rect 36766 43474 36818 43486
rect 6974 43426 7026 43438
rect 6974 43362 7026 43374
rect 8206 43426 8258 43438
rect 8206 43362 8258 43374
rect 9998 43426 10050 43438
rect 9998 43362 10050 43374
rect 11006 43426 11058 43438
rect 13358 43426 13410 43438
rect 11778 43374 11790 43426
rect 11842 43374 11854 43426
rect 11006 43362 11058 43374
rect 13358 43362 13410 43374
rect 19854 43426 19906 43438
rect 19854 43362 19906 43374
rect 21422 43426 21474 43438
rect 21422 43362 21474 43374
rect 26798 43426 26850 43438
rect 26798 43362 26850 43374
rect 30942 43426 30994 43438
rect 30942 43362 30994 43374
rect 31726 43426 31778 43438
rect 31726 43362 31778 43374
rect 33742 43426 33794 43438
rect 33742 43362 33794 43374
rect 34638 43426 34690 43438
rect 34638 43362 34690 43374
rect 37662 43426 37714 43438
rect 37662 43362 37714 43374
rect 8878 43314 8930 43326
rect 6738 43262 6750 43314
rect 6802 43311 6814 43314
rect 7074 43311 7086 43314
rect 6802 43265 7086 43311
rect 6802 43262 6814 43265
rect 7074 43262 7086 43265
rect 7138 43262 7150 43314
rect 8878 43250 8930 43262
rect 12238 43314 12290 43326
rect 12238 43250 12290 43262
rect 29486 43314 29538 43326
rect 29486 43250 29538 43262
rect 29598 43314 29650 43326
rect 29598 43250 29650 43262
rect 31950 43314 32002 43326
rect 37550 43314 37602 43326
rect 32274 43262 32286 43314
rect 32338 43262 32350 43314
rect 31950 43250 32002 43262
rect 37550 43250 37602 43262
rect 1344 43146 38640 43180
rect 1344 43094 4024 43146
rect 4076 43094 4148 43146
rect 4200 43094 4272 43146
rect 4324 43094 4396 43146
rect 4448 43094 4520 43146
rect 4572 43094 4644 43146
rect 4696 43094 4768 43146
rect 4820 43094 4892 43146
rect 4944 43094 5016 43146
rect 5068 43094 5140 43146
rect 5192 43094 24024 43146
rect 24076 43094 24148 43146
rect 24200 43094 24272 43146
rect 24324 43094 24396 43146
rect 24448 43094 24520 43146
rect 24572 43094 24644 43146
rect 24696 43094 24768 43146
rect 24820 43094 24892 43146
rect 24944 43094 25016 43146
rect 25068 43094 25140 43146
rect 25192 43094 38640 43146
rect 1344 43060 38640 43094
rect 5742 42978 5794 42990
rect 19854 42978 19906 42990
rect 13570 42926 13582 42978
rect 13634 42975 13646 42978
rect 14018 42975 14030 42978
rect 13634 42929 14030 42975
rect 13634 42926 13646 42929
rect 14018 42926 14030 42929
rect 14082 42926 14094 42978
rect 5742 42914 5794 42926
rect 19854 42914 19906 42926
rect 21758 42978 21810 42990
rect 21758 42914 21810 42926
rect 6078 42866 6130 42878
rect 6078 42802 6130 42814
rect 7422 42866 7474 42878
rect 7422 42802 7474 42814
rect 8206 42866 8258 42878
rect 8206 42802 8258 42814
rect 8542 42866 8594 42878
rect 8542 42802 8594 42814
rect 9102 42866 9154 42878
rect 9102 42802 9154 42814
rect 10110 42866 10162 42878
rect 10110 42802 10162 42814
rect 10670 42866 10722 42878
rect 10670 42802 10722 42814
rect 12686 42866 12738 42878
rect 12686 42802 12738 42814
rect 14030 42866 14082 42878
rect 14030 42802 14082 42814
rect 16046 42866 16098 42878
rect 16046 42802 16098 42814
rect 25006 42866 25058 42878
rect 25006 42802 25058 42814
rect 26238 42866 26290 42878
rect 26238 42802 26290 42814
rect 30270 42866 30322 42878
rect 35186 42814 35198 42866
rect 35250 42814 35262 42866
rect 30270 42802 30322 42814
rect 9214 42754 9266 42766
rect 9214 42690 9266 42702
rect 9662 42754 9714 42766
rect 9662 42690 9714 42702
rect 10334 42754 10386 42766
rect 12014 42754 12066 42766
rect 11666 42702 11678 42754
rect 11730 42702 11742 42754
rect 10334 42690 10386 42702
rect 12014 42690 12066 42702
rect 16382 42754 16434 42766
rect 20750 42754 20802 42766
rect 26574 42754 26626 42766
rect 16706 42702 16718 42754
rect 16770 42702 16782 42754
rect 22306 42702 22318 42754
rect 22370 42702 22382 42754
rect 16382 42690 16434 42702
rect 20750 42690 20802 42702
rect 26574 42690 26626 42702
rect 26798 42754 26850 42766
rect 26798 42690 26850 42702
rect 27022 42754 27074 42766
rect 27022 42690 27074 42702
rect 27582 42754 27634 42766
rect 31054 42754 31106 42766
rect 33182 42754 33234 42766
rect 30818 42702 30830 42754
rect 30882 42702 30894 42754
rect 31378 42702 31390 42754
rect 31442 42702 31454 42754
rect 27582 42690 27634 42702
rect 31054 42690 31106 42702
rect 33182 42690 33234 42702
rect 34302 42754 34354 42766
rect 34302 42690 34354 42702
rect 34414 42754 34466 42766
rect 36990 42754 37042 42766
rect 34962 42702 34974 42754
rect 35026 42702 35038 42754
rect 36194 42702 36206 42754
rect 36258 42702 36270 42754
rect 34414 42690 34466 42702
rect 36990 42690 37042 42702
rect 2830 42642 2882 42654
rect 2830 42578 2882 42590
rect 3166 42642 3218 42654
rect 12126 42642 12178 42654
rect 6290 42590 6302 42642
rect 6354 42590 6366 42642
rect 6738 42590 6750 42642
rect 6802 42590 6814 42642
rect 3166 42578 3218 42590
rect 12126 42578 12178 42590
rect 13582 42642 13634 42654
rect 24558 42642 24610 42654
rect 22530 42590 22542 42642
rect 22594 42590 22606 42642
rect 13582 42578 13634 42590
rect 24558 42578 24610 42590
rect 32398 42642 32450 42654
rect 36430 42642 36482 42654
rect 35074 42590 35086 42642
rect 35138 42590 35150 42642
rect 32398 42578 32450 42590
rect 36430 42578 36482 42590
rect 37998 42642 38050 42654
rect 37998 42578 38050 42590
rect 2606 42530 2658 42542
rect 2606 42466 2658 42478
rect 5070 42530 5122 42542
rect 5070 42466 5122 42478
rect 8654 42530 8706 42542
rect 8654 42466 8706 42478
rect 8990 42530 9042 42542
rect 20190 42530 20242 42542
rect 19282 42478 19294 42530
rect 19346 42478 19358 42530
rect 8990 42466 9042 42478
rect 20190 42466 20242 42478
rect 21422 42530 21474 42542
rect 21422 42466 21474 42478
rect 26686 42530 26738 42542
rect 26686 42466 26738 42478
rect 29934 42530 29986 42542
rect 29934 42466 29986 42478
rect 32846 42530 32898 42542
rect 32846 42466 32898 42478
rect 37102 42530 37154 42542
rect 37102 42466 37154 42478
rect 37326 42530 37378 42542
rect 37326 42466 37378 42478
rect 37662 42530 37714 42542
rect 37662 42466 37714 42478
rect 37886 42530 37938 42542
rect 37886 42466 37938 42478
rect 1344 42362 38640 42396
rect 1344 42310 14024 42362
rect 14076 42310 14148 42362
rect 14200 42310 14272 42362
rect 14324 42310 14396 42362
rect 14448 42310 14520 42362
rect 14572 42310 14644 42362
rect 14696 42310 14768 42362
rect 14820 42310 14892 42362
rect 14944 42310 15016 42362
rect 15068 42310 15140 42362
rect 15192 42310 34024 42362
rect 34076 42310 34148 42362
rect 34200 42310 34272 42362
rect 34324 42310 34396 42362
rect 34448 42310 34520 42362
rect 34572 42310 34644 42362
rect 34696 42310 34768 42362
rect 34820 42310 34892 42362
rect 34944 42310 35016 42362
rect 35068 42310 35140 42362
rect 35192 42310 38640 42362
rect 1344 42276 38640 42310
rect 7198 42194 7250 42206
rect 7198 42130 7250 42142
rect 8654 42194 8706 42206
rect 13806 42194 13858 42206
rect 10546 42142 10558 42194
rect 10610 42142 10622 42194
rect 8654 42130 8706 42142
rect 13806 42130 13858 42142
rect 17838 42194 17890 42206
rect 17838 42130 17890 42142
rect 19070 42194 19122 42206
rect 30494 42194 30546 42206
rect 23650 42142 23662 42194
rect 23714 42142 23726 42194
rect 29922 42142 29934 42194
rect 29986 42142 29998 42194
rect 19070 42130 19122 42142
rect 30494 42130 30546 42142
rect 8878 42082 8930 42094
rect 12686 42082 12738 42094
rect 9650 42030 9662 42082
rect 9714 42030 9726 42082
rect 8878 42018 8930 42030
rect 12686 42018 12738 42030
rect 17726 42082 17778 42094
rect 17726 42018 17778 42030
rect 26014 42082 26066 42094
rect 26014 42018 26066 42030
rect 26126 42082 26178 42094
rect 32050 42030 32062 42082
rect 32114 42030 32126 42082
rect 33506 42030 33518 42082
rect 33570 42030 33582 42082
rect 35410 42030 35422 42082
rect 35474 42030 35486 42082
rect 26126 42018 26178 42030
rect 8430 41970 8482 41982
rect 8430 41906 8482 41918
rect 8990 41970 9042 41982
rect 20974 41970 21026 41982
rect 24446 41970 24498 41982
rect 9538 41918 9550 41970
rect 9602 41918 9614 41970
rect 11554 41918 11566 41970
rect 11618 41918 11630 41970
rect 21410 41918 21422 41970
rect 21474 41918 21486 41970
rect 8990 41906 9042 41918
rect 20974 41906 21026 41918
rect 24446 41906 24498 41918
rect 25342 41970 25394 41982
rect 27022 41970 27074 41982
rect 33294 41970 33346 41982
rect 25778 41918 25790 41970
rect 25842 41918 25854 41970
rect 27346 41918 27358 41970
rect 27410 41918 27422 41970
rect 31042 41918 31054 41970
rect 31106 41918 31118 41970
rect 32162 41918 32174 41970
rect 32226 41918 32238 41970
rect 33842 41918 33854 41970
rect 33906 41918 33918 41970
rect 34738 41918 34750 41970
rect 34802 41918 34814 41970
rect 35074 41918 35086 41970
rect 35138 41918 35150 41970
rect 37314 41918 37326 41970
rect 37378 41918 37390 41970
rect 37762 41918 37774 41970
rect 37826 41918 37838 41970
rect 25342 41906 25394 41918
rect 27022 41906 27074 41918
rect 33294 41906 33346 41918
rect 18398 41858 18450 41870
rect 18398 41794 18450 41806
rect 19966 41858 20018 41870
rect 31714 41806 31726 41858
rect 31778 41806 31790 41858
rect 35522 41806 35534 41858
rect 35586 41806 35598 41858
rect 19966 41794 20018 41806
rect 25454 41746 25506 41758
rect 33182 41746 33234 41758
rect 26562 41694 26574 41746
rect 26626 41694 26638 41746
rect 25454 41682 25506 41694
rect 33182 41682 33234 41694
rect 37774 41746 37826 41758
rect 37774 41682 37826 41694
rect 38110 41746 38162 41758
rect 38110 41682 38162 41694
rect 1344 41578 38640 41612
rect 1344 41526 4024 41578
rect 4076 41526 4148 41578
rect 4200 41526 4272 41578
rect 4324 41526 4396 41578
rect 4448 41526 4520 41578
rect 4572 41526 4644 41578
rect 4696 41526 4768 41578
rect 4820 41526 4892 41578
rect 4944 41526 5016 41578
rect 5068 41526 5140 41578
rect 5192 41526 24024 41578
rect 24076 41526 24148 41578
rect 24200 41526 24272 41578
rect 24324 41526 24396 41578
rect 24448 41526 24520 41578
rect 24572 41526 24644 41578
rect 24696 41526 24768 41578
rect 24820 41526 24892 41578
rect 24944 41526 25016 41578
rect 25068 41526 25140 41578
rect 25192 41526 38640 41578
rect 1344 41492 38640 41526
rect 11118 41410 11170 41422
rect 11118 41346 11170 41358
rect 11342 41410 11394 41422
rect 11342 41346 11394 41358
rect 11902 41410 11954 41422
rect 11902 41346 11954 41358
rect 12350 41410 12402 41422
rect 12350 41346 12402 41358
rect 12574 41410 12626 41422
rect 12574 41346 12626 41358
rect 17502 41410 17554 41422
rect 17502 41346 17554 41358
rect 26462 41410 26514 41422
rect 26462 41346 26514 41358
rect 26686 41410 26738 41422
rect 26686 41346 26738 41358
rect 28142 41410 28194 41422
rect 31614 41410 31666 41422
rect 29026 41358 29038 41410
rect 29090 41407 29102 41410
rect 29810 41407 29822 41410
rect 29090 41361 29822 41407
rect 29090 41358 29102 41361
rect 29810 41358 29822 41361
rect 29874 41358 29886 41410
rect 28142 41346 28194 41358
rect 31614 41346 31666 41358
rect 32174 41410 32226 41422
rect 32174 41346 32226 41358
rect 18398 41298 18450 41310
rect 3266 41246 3278 41298
rect 3330 41246 3342 41298
rect 9538 41246 9550 41298
rect 9602 41246 9614 41298
rect 18398 41234 18450 41246
rect 18734 41298 18786 41310
rect 18734 41234 18786 41246
rect 20750 41298 20802 41310
rect 20750 41234 20802 41246
rect 21534 41298 21586 41310
rect 21534 41234 21586 41246
rect 22654 41298 22706 41310
rect 22654 41234 22706 41246
rect 26014 41298 26066 41310
rect 28590 41298 28642 41310
rect 27234 41246 27246 41298
rect 27298 41246 27310 41298
rect 27794 41246 27806 41298
rect 27858 41246 27870 41298
rect 26014 41234 26066 41246
rect 28590 41234 28642 41246
rect 29262 41298 29314 41310
rect 29262 41234 29314 41246
rect 29710 41298 29762 41310
rect 29710 41234 29762 41246
rect 30270 41298 30322 41310
rect 30270 41234 30322 41246
rect 30606 41298 30658 41310
rect 30606 41234 30658 41246
rect 8318 41186 8370 41198
rect 10670 41186 10722 41198
rect 8530 41134 8542 41186
rect 8594 41134 8606 41186
rect 9426 41134 9438 41186
rect 9490 41134 9502 41186
rect 9986 41134 9998 41186
rect 10050 41134 10062 41186
rect 8318 41122 8370 41134
rect 10670 41122 10722 41134
rect 12014 41186 12066 41198
rect 24670 41186 24722 41198
rect 21858 41134 21870 41186
rect 21922 41134 21934 41186
rect 12014 41122 12066 41134
rect 24670 41122 24722 41134
rect 24782 41186 24834 41198
rect 24782 41122 24834 41134
rect 25454 41186 25506 41198
rect 25454 41122 25506 41134
rect 25790 41186 25842 41198
rect 25790 41122 25842 41134
rect 26910 41186 26962 41198
rect 26910 41122 26962 41134
rect 27134 41186 27186 41198
rect 27134 41122 27186 41134
rect 27358 41186 27410 41198
rect 27358 41122 27410 41134
rect 28478 41186 28530 41198
rect 28478 41122 28530 41134
rect 30718 41186 30770 41198
rect 35758 41186 35810 41198
rect 31714 41134 31726 41186
rect 31778 41134 31790 41186
rect 32050 41134 32062 41186
rect 32114 41134 32126 41186
rect 35298 41134 35310 41186
rect 35362 41134 35374 41186
rect 30718 41122 30770 41134
rect 35758 41122 35810 41134
rect 36094 41186 36146 41198
rect 36094 41122 36146 41134
rect 37102 41186 37154 41198
rect 37102 41122 37154 41134
rect 8094 41074 8146 41086
rect 8094 41010 8146 41022
rect 8206 41074 8258 41086
rect 10558 41074 10610 41086
rect 8978 41022 8990 41074
rect 9042 41022 9054 41074
rect 8206 41010 8258 41022
rect 10558 41010 10610 41022
rect 11790 41074 11842 41086
rect 11790 41010 11842 41022
rect 17614 41074 17666 41086
rect 24558 41074 24610 41086
rect 22082 41022 22094 41074
rect 22146 41022 22158 41074
rect 17614 41010 17666 41022
rect 24558 41010 24610 41022
rect 25230 41074 25282 41086
rect 36318 41074 36370 41086
rect 31378 41022 31390 41074
rect 31442 41022 31454 41074
rect 32722 41022 32734 41074
rect 32786 41022 32798 41074
rect 33618 41022 33630 41074
rect 33682 41022 33694 41074
rect 37202 41022 37214 41074
rect 37266 41022 37278 41074
rect 37762 41022 37774 41074
rect 37826 41022 37838 41074
rect 25230 41010 25282 41022
rect 36318 41010 36370 41022
rect 2606 40962 2658 40974
rect 2606 40898 2658 40910
rect 2830 40962 2882 40974
rect 2830 40898 2882 40910
rect 5742 40962 5794 40974
rect 5742 40898 5794 40910
rect 6302 40962 6354 40974
rect 6302 40898 6354 40910
rect 7534 40962 7586 40974
rect 7534 40898 7586 40910
rect 7982 40962 8034 40974
rect 7982 40898 8034 40910
rect 11454 40962 11506 40974
rect 11454 40898 11506 40910
rect 22990 40962 23042 40974
rect 22990 40898 23042 40910
rect 23886 40962 23938 40974
rect 23886 40898 23938 40910
rect 24334 40962 24386 40974
rect 24334 40898 24386 40910
rect 24446 40962 24498 40974
rect 24446 40898 24498 40910
rect 26126 40962 26178 40974
rect 26126 40898 26178 40910
rect 27918 40962 27970 40974
rect 27918 40898 27970 40910
rect 35870 40962 35922 40974
rect 35870 40898 35922 40910
rect 35982 40962 36034 40974
rect 37314 40910 37326 40962
rect 37378 40910 37390 40962
rect 35982 40898 36034 40910
rect 1344 40794 38640 40828
rect 1344 40742 14024 40794
rect 14076 40742 14148 40794
rect 14200 40742 14272 40794
rect 14324 40742 14396 40794
rect 14448 40742 14520 40794
rect 14572 40742 14644 40794
rect 14696 40742 14768 40794
rect 14820 40742 14892 40794
rect 14944 40742 15016 40794
rect 15068 40742 15140 40794
rect 15192 40742 34024 40794
rect 34076 40742 34148 40794
rect 34200 40742 34272 40794
rect 34324 40742 34396 40794
rect 34448 40742 34520 40794
rect 34572 40742 34644 40794
rect 34696 40742 34768 40794
rect 34820 40742 34892 40794
rect 34944 40742 35016 40794
rect 35068 40742 35140 40794
rect 35192 40742 38640 40794
rect 1344 40708 38640 40742
rect 5294 40626 5346 40638
rect 4722 40574 4734 40626
rect 4786 40574 4798 40626
rect 5294 40562 5346 40574
rect 7422 40626 7474 40638
rect 7422 40562 7474 40574
rect 7982 40626 8034 40638
rect 7982 40562 8034 40574
rect 8878 40626 8930 40638
rect 8878 40562 8930 40574
rect 11118 40626 11170 40638
rect 22206 40626 22258 40638
rect 14130 40574 14142 40626
rect 14194 40574 14206 40626
rect 29026 40574 29038 40626
rect 29090 40574 29102 40626
rect 33618 40574 33630 40626
rect 33682 40574 33694 40626
rect 37650 40574 37662 40626
rect 37714 40574 37726 40626
rect 11118 40562 11170 40574
rect 22206 40562 22258 40574
rect 5742 40514 5794 40526
rect 8318 40514 8370 40526
rect 6626 40462 6638 40514
rect 6690 40462 6702 40514
rect 5742 40450 5794 40462
rect 8318 40450 8370 40462
rect 9550 40514 9602 40526
rect 34078 40514 34130 40526
rect 23202 40462 23214 40514
rect 23266 40462 23278 40514
rect 23650 40462 23662 40514
rect 23714 40462 23726 40514
rect 31042 40462 31054 40514
rect 31106 40462 31118 40514
rect 37874 40462 37886 40514
rect 37938 40462 37950 40514
rect 9550 40450 9602 40462
rect 34078 40450 34130 40462
rect 1822 40402 1874 40414
rect 9662 40402 9714 40414
rect 11230 40402 11282 40414
rect 15038 40402 15090 40414
rect 2258 40350 2270 40402
rect 2322 40350 2334 40402
rect 6738 40350 6750 40402
rect 6802 40350 6814 40402
rect 9986 40350 9998 40402
rect 10050 40350 10062 40402
rect 11778 40350 11790 40402
rect 11842 40350 11854 40402
rect 1822 40338 1874 40350
rect 9662 40338 9714 40350
rect 11230 40338 11282 40350
rect 15038 40338 15090 40350
rect 15934 40402 15986 40414
rect 15934 40338 15986 40350
rect 22990 40402 23042 40414
rect 22990 40338 23042 40350
rect 25902 40402 25954 40414
rect 30606 40402 30658 40414
rect 33070 40402 33122 40414
rect 26450 40350 26462 40402
rect 26514 40350 26526 40402
rect 32162 40350 32174 40402
rect 32226 40350 32238 40402
rect 25902 40338 25954 40350
rect 30606 40338 30658 40350
rect 33070 40338 33122 40350
rect 34190 40402 34242 40414
rect 35074 40350 35086 40402
rect 35138 40350 35150 40402
rect 36306 40350 36318 40402
rect 36370 40350 36382 40402
rect 37986 40350 37998 40402
rect 38050 40350 38062 40402
rect 34190 40338 34242 40350
rect 15486 40290 15538 40302
rect 15486 40226 15538 40238
rect 33294 40290 33346 40302
rect 33294 40226 33346 40238
rect 6078 40178 6130 40190
rect 22654 40178 22706 40190
rect 7298 40126 7310 40178
rect 7362 40175 7374 40178
rect 8194 40175 8206 40178
rect 7362 40129 8206 40175
rect 7362 40126 7374 40129
rect 8194 40126 8206 40129
rect 8258 40126 8270 40178
rect 6078 40114 6130 40126
rect 22654 40114 22706 40126
rect 30046 40178 30098 40190
rect 32386 40126 32398 40178
rect 32450 40126 32462 40178
rect 30046 40114 30098 40126
rect 1344 40010 38640 40044
rect 1344 39958 4024 40010
rect 4076 39958 4148 40010
rect 4200 39958 4272 40010
rect 4324 39958 4396 40010
rect 4448 39958 4520 40010
rect 4572 39958 4644 40010
rect 4696 39958 4768 40010
rect 4820 39958 4892 40010
rect 4944 39958 5016 40010
rect 5068 39958 5140 40010
rect 5192 39958 24024 40010
rect 24076 39958 24148 40010
rect 24200 39958 24272 40010
rect 24324 39958 24396 40010
rect 24448 39958 24520 40010
rect 24572 39958 24644 40010
rect 24696 39958 24768 40010
rect 24820 39958 24892 40010
rect 24944 39958 25016 40010
rect 25068 39958 25140 40010
rect 25192 39958 38640 40010
rect 1344 39924 38640 39958
rect 3726 39842 3778 39854
rect 3726 39778 3778 39790
rect 4062 39842 4114 39854
rect 4062 39778 4114 39790
rect 15150 39842 15202 39854
rect 38222 39842 38274 39854
rect 18946 39790 18958 39842
rect 19010 39839 19022 39842
rect 19618 39839 19630 39842
rect 19010 39793 19630 39839
rect 19010 39790 19022 39793
rect 19618 39790 19630 39793
rect 19682 39790 19694 39842
rect 15150 39778 15202 39790
rect 38222 39778 38274 39790
rect 5742 39730 5794 39742
rect 10782 39730 10834 39742
rect 9426 39678 9438 39730
rect 9490 39678 9502 39730
rect 5742 39666 5794 39678
rect 10782 39666 10834 39678
rect 11230 39730 11282 39742
rect 11230 39666 11282 39678
rect 14926 39730 14978 39742
rect 14926 39666 14978 39678
rect 19182 39730 19234 39742
rect 19182 39666 19234 39678
rect 19630 39730 19682 39742
rect 19630 39666 19682 39678
rect 26126 39730 26178 39742
rect 26126 39666 26178 39678
rect 29486 39730 29538 39742
rect 29486 39666 29538 39678
rect 29822 39730 29874 39742
rect 31054 39730 31106 39742
rect 30258 39678 30270 39730
rect 30322 39678 30334 39730
rect 29822 39666 29874 39678
rect 31054 39666 31106 39678
rect 31502 39730 31554 39742
rect 37102 39730 37154 39742
rect 31938 39678 31950 39730
rect 32002 39678 32014 39730
rect 34626 39678 34638 39730
rect 34690 39678 34702 39730
rect 31502 39666 31554 39678
rect 37102 39666 37154 39678
rect 3278 39618 3330 39630
rect 3278 39554 3330 39566
rect 6526 39618 6578 39630
rect 6526 39554 6578 39566
rect 7310 39618 7362 39630
rect 7310 39554 7362 39566
rect 9774 39618 9826 39630
rect 18622 39618 18674 39630
rect 25678 39618 25730 39630
rect 9986 39566 9998 39618
rect 10050 39566 10062 39618
rect 18162 39566 18174 39618
rect 18226 39566 18238 39618
rect 21746 39566 21758 39618
rect 21810 39566 21822 39618
rect 22306 39566 22318 39618
rect 22370 39566 22382 39618
rect 9774 39554 9826 39566
rect 18622 39554 18674 39566
rect 25678 39554 25730 39566
rect 30158 39618 30210 39630
rect 37214 39618 37266 39630
rect 32498 39566 32510 39618
rect 32562 39566 32574 39618
rect 34514 39566 34526 39618
rect 34578 39566 34590 39618
rect 30158 39554 30210 39566
rect 37214 39554 37266 39566
rect 37550 39618 37602 39630
rect 37550 39554 37602 39566
rect 24558 39506 24610 39518
rect 4274 39454 4286 39506
rect 4338 39454 4350 39506
rect 4834 39454 4846 39506
rect 4898 39454 4910 39506
rect 7522 39454 7534 39506
rect 7586 39454 7598 39506
rect 7858 39454 7870 39506
rect 7922 39454 7934 39506
rect 24558 39442 24610 39454
rect 25342 39506 25394 39518
rect 25342 39442 25394 39454
rect 32174 39506 32226 39518
rect 35646 39506 35698 39518
rect 32610 39454 32622 39506
rect 32674 39454 32686 39506
rect 32174 39442 32226 39454
rect 35646 39442 35698 39454
rect 36990 39506 37042 39518
rect 36990 39442 37042 39454
rect 37886 39506 37938 39518
rect 37886 39442 37938 39454
rect 2494 39394 2546 39406
rect 2494 39330 2546 39342
rect 2718 39394 2770 39406
rect 2718 39330 2770 39342
rect 6974 39394 7026 39406
rect 6974 39330 7026 39342
rect 8990 39394 9042 39406
rect 8990 39330 9042 39342
rect 9438 39394 9490 39406
rect 9438 39330 9490 39342
rect 9550 39394 9602 39406
rect 38110 39394 38162 39406
rect 15810 39342 15822 39394
rect 15874 39342 15886 39394
rect 9550 39330 9602 39342
rect 38110 39330 38162 39342
rect 1344 39226 38640 39260
rect 1344 39174 14024 39226
rect 14076 39174 14148 39226
rect 14200 39174 14272 39226
rect 14324 39174 14396 39226
rect 14448 39174 14520 39226
rect 14572 39174 14644 39226
rect 14696 39174 14768 39226
rect 14820 39174 14892 39226
rect 14944 39174 15016 39226
rect 15068 39174 15140 39226
rect 15192 39174 34024 39226
rect 34076 39174 34148 39226
rect 34200 39174 34272 39226
rect 34324 39174 34396 39226
rect 34448 39174 34520 39226
rect 34572 39174 34644 39226
rect 34696 39174 34768 39226
rect 34820 39174 34892 39226
rect 34944 39174 35016 39226
rect 35068 39174 35140 39226
rect 35192 39174 38640 39226
rect 1344 39140 38640 39174
rect 8094 39058 8146 39070
rect 3154 39006 3166 39058
rect 3218 39006 3230 39058
rect 7298 39006 7310 39058
rect 7362 39006 7374 39058
rect 8094 38994 8146 39006
rect 8654 39058 8706 39070
rect 14926 39058 14978 39070
rect 14130 39006 14142 39058
rect 14194 39006 14206 39058
rect 8654 38994 8706 39006
rect 14926 38994 14978 39006
rect 15486 39058 15538 39070
rect 15486 38994 15538 39006
rect 17838 39058 17890 39070
rect 17838 38994 17890 39006
rect 18398 39058 18450 39070
rect 18398 38994 18450 39006
rect 19070 39058 19122 39070
rect 19070 38994 19122 39006
rect 33294 39058 33346 39070
rect 33294 38994 33346 39006
rect 33742 39058 33794 39070
rect 33742 38994 33794 39006
rect 34302 39058 34354 39070
rect 34302 38994 34354 39006
rect 16718 38946 16770 38958
rect 16718 38882 16770 38894
rect 17614 38946 17666 38958
rect 17614 38882 17666 38894
rect 18286 38946 18338 38958
rect 18286 38882 18338 38894
rect 22766 38946 22818 38958
rect 22766 38882 22818 38894
rect 24110 38946 24162 38958
rect 24110 38882 24162 38894
rect 32286 38946 32338 38958
rect 32286 38882 32338 38894
rect 32398 38946 32450 38958
rect 32398 38882 32450 38894
rect 34190 38946 34242 38958
rect 35074 38894 35086 38946
rect 35138 38894 35150 38946
rect 34190 38882 34242 38894
rect 2830 38834 2882 38846
rect 2830 38770 2882 38782
rect 4622 38834 4674 38846
rect 16158 38834 16210 38846
rect 5058 38782 5070 38834
rect 5122 38782 5134 38834
rect 11330 38782 11342 38834
rect 11394 38782 11406 38834
rect 11890 38782 11902 38834
rect 11954 38782 11966 38834
rect 4622 38770 4674 38782
rect 16158 38770 16210 38782
rect 17390 38834 17442 38846
rect 17390 38770 17442 38782
rect 17950 38834 18002 38846
rect 17950 38770 18002 38782
rect 19518 38834 19570 38846
rect 32622 38834 32674 38846
rect 22306 38782 22318 38834
rect 22370 38782 22382 38834
rect 23538 38782 23550 38834
rect 23602 38782 23614 38834
rect 19518 38770 19570 38782
rect 32622 38770 32674 38782
rect 33518 38834 33570 38846
rect 33518 38770 33570 38782
rect 33966 38834 34018 38846
rect 34738 38782 34750 38834
rect 34802 38782 34814 38834
rect 37650 38782 37662 38834
rect 37714 38782 37726 38834
rect 38210 38782 38222 38834
rect 38274 38782 38286 38834
rect 33966 38770 34018 38782
rect 2494 38722 2546 38734
rect 2494 38658 2546 38670
rect 16494 38722 16546 38734
rect 16818 38670 16830 38722
rect 16882 38670 16894 38722
rect 21970 38670 21982 38722
rect 22034 38670 22046 38722
rect 23202 38670 23214 38722
rect 23266 38670 23278 38722
rect 35970 38670 35982 38722
rect 36034 38670 36046 38722
rect 16494 38658 16546 38670
rect 1344 38442 38640 38476
rect 1344 38390 4024 38442
rect 4076 38390 4148 38442
rect 4200 38390 4272 38442
rect 4324 38390 4396 38442
rect 4448 38390 4520 38442
rect 4572 38390 4644 38442
rect 4696 38390 4768 38442
rect 4820 38390 4892 38442
rect 4944 38390 5016 38442
rect 5068 38390 5140 38442
rect 5192 38390 24024 38442
rect 24076 38390 24148 38442
rect 24200 38390 24272 38442
rect 24324 38390 24396 38442
rect 24448 38390 24520 38442
rect 24572 38390 24644 38442
rect 24696 38390 24768 38442
rect 24820 38390 24892 38442
rect 24944 38390 25016 38442
rect 25068 38390 25140 38442
rect 25192 38390 38640 38442
rect 1344 38356 38640 38390
rect 5854 38274 5906 38286
rect 5854 38210 5906 38222
rect 6190 38274 6242 38286
rect 6190 38210 6242 38222
rect 18734 38274 18786 38286
rect 18734 38210 18786 38222
rect 33182 38274 33234 38286
rect 33618 38222 33630 38274
rect 33682 38222 33694 38274
rect 35746 38222 35758 38274
rect 35810 38222 35822 38274
rect 33182 38210 33234 38222
rect 24894 38162 24946 38174
rect 24894 38098 24946 38110
rect 33742 38162 33794 38174
rect 37998 38162 38050 38174
rect 35298 38110 35310 38162
rect 35362 38110 35374 38162
rect 36082 38110 36094 38162
rect 36146 38110 36158 38162
rect 37202 38110 37214 38162
rect 37266 38110 37278 38162
rect 33742 38098 33794 38110
rect 37998 38098 38050 38110
rect 15262 38050 15314 38062
rect 19630 38050 19682 38062
rect 15698 37998 15710 38050
rect 15762 37998 15774 38050
rect 15262 37986 15314 37998
rect 19630 37986 19682 37998
rect 31726 38050 31778 38062
rect 31726 37986 31778 37998
rect 32062 38050 32114 38062
rect 32062 37986 32114 37998
rect 33854 38050 33906 38062
rect 37774 38050 37826 38062
rect 35186 37998 35198 38050
rect 35250 37998 35262 38050
rect 36194 37998 36206 38050
rect 36258 37998 36270 38050
rect 37426 37998 37438 38050
rect 37490 37998 37502 38050
rect 33854 37986 33906 37998
rect 37774 37986 37826 37998
rect 9662 37938 9714 37950
rect 31390 37938 31442 37950
rect 6402 37886 6414 37938
rect 6466 37886 6478 37938
rect 6962 37886 6974 37938
rect 7026 37886 7038 37938
rect 19842 37886 19854 37938
rect 19906 37886 19918 37938
rect 20178 37886 20190 37938
rect 20242 37886 20254 37938
rect 9662 37874 9714 37886
rect 31390 37874 31442 37886
rect 32510 37938 32562 37950
rect 32510 37874 32562 37886
rect 32846 37938 32898 37950
rect 32846 37874 32898 37886
rect 8430 37826 8482 37838
rect 8430 37762 8482 37774
rect 8878 37826 8930 37838
rect 8878 37762 8930 37774
rect 9774 37826 9826 37838
rect 9774 37762 9826 37774
rect 9998 37826 10050 37838
rect 9998 37762 10050 37774
rect 11678 37826 11730 37838
rect 11678 37762 11730 37774
rect 13694 37826 13746 37838
rect 19294 37826 19346 37838
rect 17938 37774 17950 37826
rect 18002 37774 18014 37826
rect 13694 37762 13746 37774
rect 19294 37762 19346 37774
rect 26686 37826 26738 37838
rect 26686 37762 26738 37774
rect 27806 37826 27858 37838
rect 27806 37762 27858 37774
rect 28254 37826 28306 37838
rect 28254 37762 28306 37774
rect 31054 37826 31106 37838
rect 31054 37762 31106 37774
rect 31726 37826 31778 37838
rect 31726 37762 31778 37774
rect 32174 37826 32226 37838
rect 32174 37762 32226 37774
rect 32398 37826 32450 37838
rect 32398 37762 32450 37774
rect 33070 37826 33122 37838
rect 33070 37762 33122 37774
rect 37102 37826 37154 37838
rect 37102 37762 37154 37774
rect 37326 37826 37378 37838
rect 37326 37762 37378 37774
rect 1344 37658 38640 37692
rect 1344 37606 14024 37658
rect 14076 37606 14148 37658
rect 14200 37606 14272 37658
rect 14324 37606 14396 37658
rect 14448 37606 14520 37658
rect 14572 37606 14644 37658
rect 14696 37606 14768 37658
rect 14820 37606 14892 37658
rect 14944 37606 15016 37658
rect 15068 37606 15140 37658
rect 15192 37606 34024 37658
rect 34076 37606 34148 37658
rect 34200 37606 34272 37658
rect 34324 37606 34396 37658
rect 34448 37606 34520 37658
rect 34572 37606 34644 37658
rect 34696 37606 34768 37658
rect 34820 37606 34892 37658
rect 34944 37606 35016 37658
rect 35068 37606 35140 37658
rect 35192 37606 38640 37658
rect 1344 37572 38640 37606
rect 9102 37490 9154 37502
rect 9102 37426 9154 37438
rect 12350 37490 12402 37502
rect 16158 37490 16210 37502
rect 13346 37438 13358 37490
rect 13410 37438 13422 37490
rect 14802 37438 14814 37490
rect 14866 37438 14878 37490
rect 12350 37426 12402 37438
rect 16158 37426 16210 37438
rect 16718 37490 16770 37502
rect 16718 37426 16770 37438
rect 17838 37490 17890 37502
rect 22094 37490 22146 37502
rect 21522 37438 21534 37490
rect 21586 37438 21598 37490
rect 17838 37426 17890 37438
rect 22094 37426 22146 37438
rect 24670 37490 24722 37502
rect 31950 37490 32002 37502
rect 37774 37490 37826 37502
rect 31154 37438 31166 37490
rect 31218 37438 31230 37490
rect 35298 37438 35310 37490
rect 35362 37438 35374 37490
rect 24670 37426 24722 37438
rect 31950 37426 32002 37438
rect 37774 37426 37826 37438
rect 8766 37378 8818 37390
rect 3154 37326 3166 37378
rect 3218 37326 3230 37378
rect 8766 37314 8818 37326
rect 8878 37378 8930 37390
rect 8878 37314 8930 37326
rect 9998 37378 10050 37390
rect 9998 37314 10050 37326
rect 12574 37378 12626 37390
rect 22430 37378 22482 37390
rect 27022 37378 27074 37390
rect 12898 37326 12910 37378
rect 12962 37326 12974 37378
rect 14018 37326 14030 37378
rect 14082 37326 14094 37378
rect 25890 37326 25902 37378
rect 25954 37326 25966 37378
rect 26450 37326 26462 37378
rect 26514 37326 26526 37378
rect 12574 37314 12626 37326
rect 22430 37314 22482 37326
rect 27022 37314 27074 37326
rect 27582 37378 27634 37390
rect 27582 37314 27634 37326
rect 28030 37378 28082 37390
rect 28030 37314 28082 37326
rect 34190 37378 34242 37390
rect 34190 37314 34242 37326
rect 36206 37378 36258 37390
rect 36206 37314 36258 37326
rect 2830 37266 2882 37278
rect 2830 37202 2882 37214
rect 10222 37266 10274 37278
rect 10222 37202 10274 37214
rect 12238 37266 12290 37278
rect 16494 37266 16546 37278
rect 12786 37214 12798 37266
rect 12850 37214 12862 37266
rect 15026 37214 15038 37266
rect 15090 37214 15102 37266
rect 12238 37202 12290 37214
rect 16494 37202 16546 37214
rect 17502 37266 17554 37278
rect 17502 37202 17554 37214
rect 17726 37266 17778 37278
rect 17726 37202 17778 37214
rect 18062 37266 18114 37278
rect 18062 37202 18114 37214
rect 18622 37266 18674 37278
rect 25678 37266 25730 37278
rect 27806 37266 27858 37278
rect 19058 37214 19070 37266
rect 19122 37214 19134 37266
rect 27346 37214 27358 37266
rect 27410 37214 27422 37266
rect 18622 37202 18674 37214
rect 25678 37202 25730 37214
rect 27806 37202 27858 37214
rect 28254 37266 28306 37278
rect 35198 37266 35250 37278
rect 28914 37214 28926 37266
rect 28978 37214 28990 37266
rect 28254 37202 28306 37214
rect 35198 37202 35250 37214
rect 35646 37266 35698 37278
rect 37650 37214 37662 37266
rect 37714 37214 37726 37266
rect 35646 37202 35698 37214
rect 2494 37154 2546 37166
rect 2494 37090 2546 37102
rect 11454 37154 11506 37166
rect 11454 37090 11506 37102
rect 11902 37154 11954 37166
rect 22878 37154 22930 37166
rect 16818 37102 16830 37154
rect 16882 37102 16894 37154
rect 11902 37090 11954 37102
rect 22878 37090 22930 37102
rect 24110 37154 24162 37166
rect 24110 37090 24162 37102
rect 27694 37154 27746 37166
rect 27694 37090 27746 37102
rect 25342 37042 25394 37054
rect 10546 36990 10558 37042
rect 10610 36990 10622 37042
rect 25342 36978 25394 36990
rect 37886 37042 37938 37054
rect 37886 36978 37938 36990
rect 38110 37042 38162 37054
rect 38110 36978 38162 36990
rect 1344 36874 38640 36908
rect 1344 36822 4024 36874
rect 4076 36822 4148 36874
rect 4200 36822 4272 36874
rect 4324 36822 4396 36874
rect 4448 36822 4520 36874
rect 4572 36822 4644 36874
rect 4696 36822 4768 36874
rect 4820 36822 4892 36874
rect 4944 36822 5016 36874
rect 5068 36822 5140 36874
rect 5192 36822 24024 36874
rect 24076 36822 24148 36874
rect 24200 36822 24272 36874
rect 24324 36822 24396 36874
rect 24448 36822 24520 36874
rect 24572 36822 24644 36874
rect 24696 36822 24768 36874
rect 24820 36822 24892 36874
rect 24944 36822 25016 36874
rect 25068 36822 25140 36874
rect 25192 36822 38640 36874
rect 1344 36788 38640 36822
rect 11890 36654 11902 36706
rect 11954 36703 11966 36706
rect 12898 36703 12910 36706
rect 11954 36657 12910 36703
rect 11954 36654 11966 36657
rect 12898 36654 12910 36657
rect 12962 36654 12974 36706
rect 35410 36654 35422 36706
rect 35474 36654 35486 36706
rect 10894 36594 10946 36606
rect 29598 36594 29650 36606
rect 6402 36542 6414 36594
rect 6466 36542 6478 36594
rect 8754 36542 8766 36594
rect 8818 36542 8830 36594
rect 12114 36542 12126 36594
rect 12178 36591 12190 36594
rect 12338 36591 12350 36594
rect 12178 36545 12350 36591
rect 12178 36542 12190 36545
rect 12338 36542 12350 36545
rect 12402 36542 12414 36594
rect 14242 36542 14254 36594
rect 14306 36542 14318 36594
rect 23314 36542 23326 36594
rect 23378 36542 23390 36594
rect 26674 36542 26686 36594
rect 26738 36542 26750 36594
rect 33282 36542 33294 36594
rect 33346 36542 33358 36594
rect 35634 36542 35646 36594
rect 35698 36542 35710 36594
rect 10894 36530 10946 36542
rect 29598 36530 29650 36542
rect 8990 36482 9042 36494
rect 11902 36482 11954 36494
rect 27694 36482 27746 36494
rect 6178 36430 6190 36482
rect 6242 36430 6254 36482
rect 10322 36430 10334 36482
rect 10386 36430 10398 36482
rect 13570 36430 13582 36482
rect 13634 36430 13646 36482
rect 21522 36430 21534 36482
rect 21586 36430 21598 36482
rect 24322 36430 24334 36482
rect 24386 36430 24398 36482
rect 8990 36418 9042 36430
rect 11902 36418 11954 36430
rect 27694 36418 27746 36430
rect 29038 36482 29090 36494
rect 29038 36418 29090 36430
rect 29486 36482 29538 36494
rect 29486 36418 29538 36430
rect 30382 36482 30434 36494
rect 33630 36482 33682 36494
rect 34526 36482 34578 36494
rect 37550 36482 37602 36494
rect 31154 36430 31166 36482
rect 31218 36430 31230 36482
rect 31938 36430 31950 36482
rect 32002 36430 32014 36482
rect 33730 36430 33742 36482
rect 33794 36430 33806 36482
rect 35410 36430 35422 36482
rect 35474 36430 35486 36482
rect 36530 36430 36542 36482
rect 36594 36430 36606 36482
rect 30382 36418 30434 36430
rect 33630 36418 33682 36430
rect 34526 36418 34578 36430
rect 37550 36418 37602 36430
rect 4622 36370 4674 36382
rect 4622 36306 4674 36318
rect 4846 36370 4898 36382
rect 4846 36306 4898 36318
rect 5182 36370 5234 36382
rect 8766 36370 8818 36382
rect 11342 36370 11394 36382
rect 14814 36370 14866 36382
rect 31614 36370 31666 36382
rect 5842 36318 5854 36370
rect 5906 36318 5918 36370
rect 9538 36318 9550 36370
rect 9602 36318 9614 36370
rect 10098 36318 10110 36370
rect 10162 36318 10174 36370
rect 13682 36318 13694 36370
rect 13746 36318 13758 36370
rect 28018 36318 28030 36370
rect 28082 36318 28094 36370
rect 28466 36318 28478 36370
rect 28530 36318 28542 36370
rect 5182 36306 5234 36318
rect 8766 36306 8818 36318
rect 11342 36306 11394 36318
rect 14814 36306 14866 36318
rect 31614 36306 31666 36318
rect 31726 36370 31778 36382
rect 36990 36370 37042 36382
rect 32162 36318 32174 36370
rect 32226 36318 32238 36370
rect 32610 36318 32622 36370
rect 32674 36318 32686 36370
rect 31726 36306 31778 36318
rect 36990 36306 37042 36318
rect 37326 36370 37378 36382
rect 37326 36306 37378 36318
rect 37998 36370 38050 36382
rect 37998 36306 38050 36318
rect 38222 36370 38274 36382
rect 38222 36306 38274 36318
rect 2606 36258 2658 36270
rect 2606 36194 2658 36206
rect 2830 36258 2882 36270
rect 4062 36258 4114 36270
rect 3154 36206 3166 36258
rect 3218 36206 3230 36258
rect 2830 36194 2882 36206
rect 4062 36194 4114 36206
rect 4958 36258 5010 36270
rect 4958 36194 5010 36206
rect 7534 36258 7586 36270
rect 7534 36194 7586 36206
rect 8318 36258 8370 36270
rect 12462 36258 12514 36270
rect 9762 36206 9774 36258
rect 9826 36206 9838 36258
rect 8318 36194 8370 36206
rect 12462 36194 12514 36206
rect 12910 36258 12962 36270
rect 12910 36194 12962 36206
rect 18846 36258 18898 36270
rect 18846 36194 18898 36206
rect 27358 36258 27410 36270
rect 27358 36194 27410 36206
rect 29710 36258 29762 36270
rect 29710 36194 29762 36206
rect 30046 36258 30098 36270
rect 30046 36194 30098 36206
rect 30270 36258 30322 36270
rect 30270 36194 30322 36206
rect 30830 36258 30882 36270
rect 30830 36194 30882 36206
rect 31390 36258 31442 36270
rect 31390 36194 31442 36206
rect 37102 36258 37154 36270
rect 37102 36194 37154 36206
rect 38110 36258 38162 36270
rect 38110 36194 38162 36206
rect 1344 36090 38640 36124
rect 1344 36038 14024 36090
rect 14076 36038 14148 36090
rect 14200 36038 14272 36090
rect 14324 36038 14396 36090
rect 14448 36038 14520 36090
rect 14572 36038 14644 36090
rect 14696 36038 14768 36090
rect 14820 36038 14892 36090
rect 14944 36038 15016 36090
rect 15068 36038 15140 36090
rect 15192 36038 34024 36090
rect 34076 36038 34148 36090
rect 34200 36038 34272 36090
rect 34324 36038 34396 36090
rect 34448 36038 34520 36090
rect 34572 36038 34644 36090
rect 34696 36038 34768 36090
rect 34820 36038 34892 36090
rect 34944 36038 35016 36090
rect 35068 36038 35140 36090
rect 35192 36038 38640 36090
rect 1344 36004 38640 36038
rect 5854 35922 5906 35934
rect 4946 35870 4958 35922
rect 5010 35870 5022 35922
rect 5854 35858 5906 35870
rect 6302 35922 6354 35934
rect 6302 35858 6354 35870
rect 7086 35922 7138 35934
rect 7086 35858 7138 35870
rect 7870 35922 7922 35934
rect 22878 35922 22930 35934
rect 22306 35870 22318 35922
rect 22370 35870 22382 35922
rect 7870 35858 7922 35870
rect 22878 35858 22930 35870
rect 23214 35922 23266 35934
rect 35982 35922 36034 35934
rect 34962 35870 34974 35922
rect 35026 35870 35038 35922
rect 23214 35858 23266 35870
rect 35982 35858 36034 35870
rect 36094 35922 36146 35934
rect 36094 35858 36146 35870
rect 37326 35922 37378 35934
rect 37326 35858 37378 35870
rect 37438 35922 37490 35934
rect 37438 35858 37490 35870
rect 38334 35922 38386 35934
rect 38334 35858 38386 35870
rect 8654 35810 8706 35822
rect 8418 35758 8430 35810
rect 8482 35758 8494 35810
rect 8654 35746 8706 35758
rect 8766 35810 8818 35822
rect 8766 35746 8818 35758
rect 9662 35810 9714 35822
rect 9662 35746 9714 35758
rect 9774 35810 9826 35822
rect 9774 35746 9826 35758
rect 9886 35810 9938 35822
rect 38110 35810 38162 35822
rect 9986 35758 9998 35810
rect 10050 35758 10062 35810
rect 14914 35758 14926 35810
rect 14978 35758 14990 35810
rect 16370 35758 16382 35810
rect 16434 35758 16446 35810
rect 25890 35758 25902 35810
rect 25954 35758 25966 35810
rect 26450 35758 26462 35810
rect 26514 35758 26526 35810
rect 27794 35758 27806 35810
rect 27858 35758 27870 35810
rect 28354 35758 28366 35810
rect 28418 35758 28430 35810
rect 33058 35758 33070 35810
rect 33122 35758 33134 35810
rect 9886 35746 9938 35758
rect 38110 35746 38162 35758
rect 1822 35698 1874 35710
rect 8990 35698 9042 35710
rect 2370 35646 2382 35698
rect 2434 35646 2446 35698
rect 1822 35634 1874 35646
rect 8990 35634 9042 35646
rect 9550 35698 9602 35710
rect 19406 35698 19458 35710
rect 23998 35698 24050 35710
rect 11890 35646 11902 35698
rect 11954 35646 11966 35698
rect 14018 35646 14030 35698
rect 14082 35646 14094 35698
rect 14690 35646 14702 35698
rect 14754 35646 14766 35698
rect 15138 35646 15150 35698
rect 15202 35646 15214 35698
rect 19842 35646 19854 35698
rect 19906 35646 19918 35698
rect 9550 35634 9602 35646
rect 19406 35634 19458 35646
rect 23998 35634 24050 35646
rect 25678 35698 25730 35710
rect 25678 35634 25730 35646
rect 27582 35698 27634 35710
rect 34862 35698 34914 35710
rect 31826 35646 31838 35698
rect 31890 35646 31902 35698
rect 33618 35646 33630 35698
rect 33682 35646 33694 35698
rect 34626 35646 34638 35698
rect 34690 35646 34702 35698
rect 27582 35634 27634 35646
rect 34862 35634 34914 35646
rect 36206 35698 36258 35710
rect 36206 35634 36258 35646
rect 36430 35698 36482 35710
rect 36430 35634 36482 35646
rect 36654 35698 36706 35710
rect 37214 35698 37266 35710
rect 37998 35698 38050 35710
rect 36978 35646 36990 35698
rect 37042 35646 37054 35698
rect 37650 35646 37662 35698
rect 37714 35646 37726 35698
rect 36654 35634 36706 35646
rect 37214 35634 37266 35646
rect 37998 35634 38050 35646
rect 7758 35586 7810 35598
rect 24446 35586 24498 35598
rect 8642 35534 8654 35586
rect 8706 35534 8718 35586
rect 31938 35534 31950 35586
rect 32002 35534 32014 35586
rect 33730 35534 33742 35586
rect 33794 35534 33806 35586
rect 34290 35534 34302 35586
rect 34354 35534 34366 35586
rect 7758 35522 7810 35534
rect 24446 35522 24498 35534
rect 5518 35474 5570 35486
rect 25342 35474 25394 35486
rect 10882 35422 10894 35474
rect 10946 35422 10958 35474
rect 5518 35410 5570 35422
rect 25342 35410 25394 35422
rect 27246 35474 27298 35486
rect 34850 35422 34862 35474
rect 34914 35471 34926 35474
rect 35186 35471 35198 35474
rect 34914 35425 35198 35471
rect 34914 35422 34926 35425
rect 35186 35422 35198 35425
rect 35250 35422 35262 35474
rect 27246 35410 27298 35422
rect 1344 35306 38640 35340
rect 1344 35254 4024 35306
rect 4076 35254 4148 35306
rect 4200 35254 4272 35306
rect 4324 35254 4396 35306
rect 4448 35254 4520 35306
rect 4572 35254 4644 35306
rect 4696 35254 4768 35306
rect 4820 35254 4892 35306
rect 4944 35254 5016 35306
rect 5068 35254 5140 35306
rect 5192 35254 24024 35306
rect 24076 35254 24148 35306
rect 24200 35254 24272 35306
rect 24324 35254 24396 35306
rect 24448 35254 24520 35306
rect 24572 35254 24644 35306
rect 24696 35254 24768 35306
rect 24820 35254 24892 35306
rect 24944 35254 25016 35306
rect 25068 35254 25140 35306
rect 25192 35254 38640 35306
rect 1344 35220 38640 35254
rect 2158 35138 2210 35150
rect 2158 35074 2210 35086
rect 10334 35138 10386 35150
rect 10334 35074 10386 35086
rect 10894 35138 10946 35150
rect 10894 35074 10946 35086
rect 12462 35138 12514 35150
rect 12462 35074 12514 35086
rect 12798 35138 12850 35150
rect 12798 35074 12850 35086
rect 13582 35138 13634 35150
rect 13582 35074 13634 35086
rect 17166 35138 17218 35150
rect 17166 35074 17218 35086
rect 20302 35138 20354 35150
rect 20302 35074 20354 35086
rect 20638 35138 20690 35150
rect 20638 35074 20690 35086
rect 26574 35138 26626 35150
rect 26574 35074 26626 35086
rect 32510 35138 32562 35150
rect 32510 35074 32562 35086
rect 37326 35138 37378 35150
rect 37326 35074 37378 35086
rect 14590 35026 14642 35038
rect 14590 34962 14642 34974
rect 15038 35026 15090 35038
rect 27022 35026 27074 35038
rect 17938 34974 17950 35026
rect 18002 34974 18014 35026
rect 15038 34962 15090 34974
rect 27022 34962 27074 34974
rect 27358 35026 27410 35038
rect 35198 35026 35250 35038
rect 33282 34974 33294 35026
rect 33346 34974 33358 35026
rect 27358 34962 27410 34974
rect 35198 34962 35250 34974
rect 35870 35026 35922 35038
rect 35870 34962 35922 34974
rect 36206 35026 36258 35038
rect 36206 34962 36258 34974
rect 2494 34914 2546 34926
rect 4174 34914 4226 34926
rect 11118 34914 11170 34926
rect 23102 34914 23154 34926
rect 35646 34914 35698 34926
rect 3042 34862 3054 34914
rect 3106 34862 3118 34914
rect 4722 34862 4734 34914
rect 4786 34862 4798 34914
rect 6738 34862 6750 34914
rect 6802 34862 6814 34914
rect 7298 34862 7310 34914
rect 7362 34862 7374 34914
rect 11778 34862 11790 34914
rect 11842 34862 11854 34914
rect 19618 34862 19630 34914
rect 19682 34862 19694 34914
rect 23538 34862 23550 34914
rect 23602 34862 23614 34914
rect 33170 34862 33182 34914
rect 33234 34862 33246 34914
rect 33842 34862 33854 34914
rect 33906 34862 33918 34914
rect 2494 34850 2546 34862
rect 4174 34850 4226 34862
rect 11118 34850 11170 34862
rect 23102 34850 23154 34862
rect 35646 34850 35698 34862
rect 36094 34914 36146 34926
rect 36094 34850 36146 34862
rect 6078 34802 6130 34814
rect 13470 34802 13522 34814
rect 3266 34750 3278 34802
rect 3330 34750 3342 34802
rect 4946 34750 4958 34802
rect 5010 34750 5022 34802
rect 10546 34750 10558 34802
rect 10610 34750 10622 34802
rect 11666 34750 11678 34802
rect 11730 34750 11742 34802
rect 6078 34738 6130 34750
rect 13470 34738 13522 34750
rect 17278 34802 17330 34814
rect 17278 34738 17330 34750
rect 17614 34802 17666 34814
rect 17614 34738 17666 34750
rect 18062 34802 18114 34814
rect 18062 34738 18114 34750
rect 18510 34802 18562 34814
rect 18510 34738 18562 34750
rect 19070 34802 19122 34814
rect 25790 34802 25842 34814
rect 19506 34750 19518 34802
rect 19570 34750 19582 34802
rect 19070 34738 19122 34750
rect 25790 34738 25842 34750
rect 27806 34802 27858 34814
rect 27806 34738 27858 34750
rect 32398 34802 32450 34814
rect 35086 34802 35138 34814
rect 32834 34750 32846 34802
rect 32898 34750 32910 34802
rect 32398 34738 32450 34750
rect 35086 34738 35138 34750
rect 36318 34802 36370 34814
rect 36318 34738 36370 34750
rect 36990 34802 37042 34814
rect 36990 34738 37042 34750
rect 37214 34802 37266 34814
rect 37214 34738 37266 34750
rect 37774 34802 37826 34814
rect 37774 34738 37826 34750
rect 37886 34802 37938 34814
rect 37886 34738 37938 34750
rect 3838 34690 3890 34702
rect 3838 34626 3890 34638
rect 5742 34690 5794 34702
rect 5742 34626 5794 34638
rect 6190 34690 6242 34702
rect 6190 34626 6242 34638
rect 6414 34690 6466 34702
rect 13582 34690 13634 34702
rect 9538 34638 9550 34690
rect 9602 34638 9614 34690
rect 6414 34626 6466 34638
rect 13582 34626 13634 34638
rect 14142 34690 14194 34702
rect 14142 34626 14194 34638
rect 16718 34690 16770 34702
rect 16718 34626 16770 34638
rect 17166 34690 17218 34702
rect 17166 34626 17218 34638
rect 17838 34690 17890 34702
rect 17838 34626 17890 34638
rect 28254 34690 28306 34702
rect 28254 34626 28306 34638
rect 29822 34690 29874 34702
rect 29822 34626 29874 34638
rect 34862 34690 34914 34702
rect 34862 34626 34914 34638
rect 35310 34690 35362 34702
rect 35310 34626 35362 34638
rect 37550 34690 37602 34702
rect 37550 34626 37602 34638
rect 1344 34522 38640 34556
rect 1344 34470 14024 34522
rect 14076 34470 14148 34522
rect 14200 34470 14272 34522
rect 14324 34470 14396 34522
rect 14448 34470 14520 34522
rect 14572 34470 14644 34522
rect 14696 34470 14768 34522
rect 14820 34470 14892 34522
rect 14944 34470 15016 34522
rect 15068 34470 15140 34522
rect 15192 34470 34024 34522
rect 34076 34470 34148 34522
rect 34200 34470 34272 34522
rect 34324 34470 34396 34522
rect 34448 34470 34520 34522
rect 34572 34470 34644 34522
rect 34696 34470 34768 34522
rect 34820 34470 34892 34522
rect 34944 34470 35016 34522
rect 35068 34470 35140 34522
rect 35192 34470 38640 34522
rect 1344 34436 38640 34470
rect 5294 34354 5346 34366
rect 4610 34302 4622 34354
rect 4674 34302 4686 34354
rect 5294 34290 5346 34302
rect 5630 34354 5682 34366
rect 5630 34290 5682 34302
rect 7086 34354 7138 34366
rect 7086 34290 7138 34302
rect 7310 34354 7362 34366
rect 7310 34290 7362 34302
rect 9886 34354 9938 34366
rect 9886 34290 9938 34302
rect 11230 34354 11282 34366
rect 11230 34290 11282 34302
rect 12126 34354 12178 34366
rect 12126 34290 12178 34302
rect 15822 34354 15874 34366
rect 15822 34290 15874 34302
rect 16270 34354 16322 34366
rect 16270 34290 16322 34302
rect 16718 34354 16770 34366
rect 16718 34290 16770 34302
rect 16942 34354 16994 34366
rect 16942 34290 16994 34302
rect 25342 34354 25394 34366
rect 29710 34354 29762 34366
rect 29138 34302 29150 34354
rect 29202 34302 29214 34354
rect 25342 34290 25394 34302
rect 29710 34290 29762 34302
rect 35758 34354 35810 34366
rect 35758 34290 35810 34302
rect 37438 34354 37490 34366
rect 37438 34290 37490 34302
rect 7422 34242 7474 34254
rect 6626 34190 6638 34242
rect 6690 34190 6702 34242
rect 7422 34178 7474 34190
rect 10558 34242 10610 34254
rect 10558 34178 10610 34190
rect 16606 34242 16658 34254
rect 16606 34178 16658 34190
rect 30158 34242 30210 34254
rect 30158 34178 30210 34190
rect 30270 34242 30322 34254
rect 33070 34242 33122 34254
rect 32498 34190 32510 34242
rect 32562 34190 32574 34242
rect 30270 34178 30322 34190
rect 33070 34178 33122 34190
rect 33518 34242 33570 34254
rect 34066 34190 34078 34242
rect 34130 34190 34142 34242
rect 36642 34190 36654 34242
rect 36706 34190 36718 34242
rect 33518 34178 33570 34190
rect 1822 34130 1874 34142
rect 8094 34130 8146 34142
rect 2258 34078 2270 34130
rect 2322 34078 2334 34130
rect 6402 34078 6414 34130
rect 6466 34078 6478 34130
rect 1822 34066 1874 34078
rect 8094 34066 8146 34078
rect 8430 34130 8482 34142
rect 8430 34066 8482 34078
rect 8654 34130 8706 34142
rect 8654 34066 8706 34078
rect 9550 34130 9602 34142
rect 9550 34066 9602 34078
rect 9886 34130 9938 34142
rect 9886 34066 9938 34078
rect 10222 34130 10274 34142
rect 10222 34066 10274 34078
rect 10446 34130 10498 34142
rect 26014 34130 26066 34142
rect 30494 34130 30546 34142
rect 33854 34130 33906 34142
rect 17490 34078 17502 34130
rect 17554 34078 17566 34130
rect 17826 34078 17838 34130
rect 17890 34078 17902 34130
rect 20066 34078 20078 34130
rect 20130 34078 20142 34130
rect 26674 34078 26686 34130
rect 26738 34078 26750 34130
rect 31154 34078 31166 34130
rect 31218 34078 31230 34130
rect 31490 34078 31502 34130
rect 31554 34078 31566 34130
rect 32274 34078 32286 34130
rect 32338 34078 32350 34130
rect 33282 34078 33294 34130
rect 33346 34078 33358 34130
rect 34514 34078 34526 34130
rect 34578 34078 34590 34130
rect 35186 34078 35198 34130
rect 35250 34078 35262 34130
rect 36866 34078 36878 34130
rect 36930 34078 36942 34130
rect 10446 34066 10498 34078
rect 26014 34066 26066 34078
rect 30494 34066 30546 34078
rect 33854 34066 33906 34078
rect 7870 34018 7922 34030
rect 11678 34018 11730 34030
rect 8194 33966 8206 34018
rect 8258 33966 8270 34018
rect 7870 33954 7922 33966
rect 11678 33954 11730 33966
rect 12910 34018 12962 34030
rect 12910 33954 12962 33966
rect 21758 34018 21810 34030
rect 21758 33954 21810 33966
rect 22206 34018 22258 34030
rect 22206 33954 22258 33966
rect 31726 34018 31778 34030
rect 37886 34018 37938 34030
rect 33394 33966 33406 34018
rect 33458 33966 33470 34018
rect 31726 33954 31778 33966
rect 37886 33954 37938 33966
rect 5966 33906 6018 33918
rect 36094 33906 36146 33918
rect 21186 33854 21198 33906
rect 21250 33854 21262 33906
rect 34962 33854 34974 33906
rect 35026 33854 35038 33906
rect 5966 33842 6018 33854
rect 36094 33842 36146 33854
rect 1344 33738 38640 33772
rect 1344 33686 4024 33738
rect 4076 33686 4148 33738
rect 4200 33686 4272 33738
rect 4324 33686 4396 33738
rect 4448 33686 4520 33738
rect 4572 33686 4644 33738
rect 4696 33686 4768 33738
rect 4820 33686 4892 33738
rect 4944 33686 5016 33738
rect 5068 33686 5140 33738
rect 5192 33686 24024 33738
rect 24076 33686 24148 33738
rect 24200 33686 24272 33738
rect 24324 33686 24396 33738
rect 24448 33686 24520 33738
rect 24572 33686 24644 33738
rect 24696 33686 24768 33738
rect 24820 33686 24892 33738
rect 24944 33686 25016 33738
rect 25068 33686 25140 33738
rect 25192 33686 38640 33738
rect 1344 33652 38640 33686
rect 16382 33570 16434 33582
rect 4610 33518 4622 33570
rect 4674 33567 4686 33570
rect 5170 33567 5182 33570
rect 4674 33521 5182 33567
rect 4674 33518 4686 33521
rect 5170 33518 5182 33521
rect 5234 33518 5246 33570
rect 35858 33518 35870 33570
rect 35922 33518 35934 33570
rect 37538 33518 37550 33570
rect 37602 33518 37614 33570
rect 16382 33506 16434 33518
rect 4622 33458 4674 33470
rect 4622 33394 4674 33406
rect 5070 33458 5122 33470
rect 5070 33394 5122 33406
rect 11566 33458 11618 33470
rect 11566 33394 11618 33406
rect 12014 33458 12066 33470
rect 12014 33394 12066 33406
rect 16942 33458 16994 33470
rect 18958 33458 19010 33470
rect 17266 33406 17278 33458
rect 17330 33406 17342 33458
rect 16942 33394 16994 33406
rect 18958 33394 19010 33406
rect 22542 33458 22594 33470
rect 22542 33394 22594 33406
rect 23886 33458 23938 33470
rect 23886 33394 23938 33406
rect 26238 33458 26290 33470
rect 36990 33458 37042 33470
rect 33954 33406 33966 33458
rect 34018 33406 34030 33458
rect 35410 33406 35422 33458
rect 35474 33406 35486 33458
rect 26238 33394 26290 33406
rect 36990 33394 37042 33406
rect 37998 33458 38050 33470
rect 37998 33394 38050 33406
rect 6078 33346 6130 33358
rect 7534 33346 7586 33358
rect 11230 33346 11282 33358
rect 6850 33294 6862 33346
rect 6914 33294 6926 33346
rect 10546 33294 10558 33346
rect 10610 33294 10622 33346
rect 6078 33282 6130 33294
rect 7534 33282 7586 33294
rect 11230 33282 11282 33294
rect 13918 33346 13970 33358
rect 13918 33282 13970 33294
rect 16270 33346 16322 33358
rect 31166 33346 31218 33358
rect 24434 33294 24446 33346
rect 24498 33294 24510 33346
rect 16270 33282 16322 33294
rect 31166 33282 31218 33294
rect 31838 33346 31890 33358
rect 31838 33282 31890 33294
rect 33294 33346 33346 33358
rect 37214 33346 37266 33358
rect 33842 33294 33854 33346
rect 33906 33294 33918 33346
rect 34738 33294 34750 33346
rect 34802 33294 34814 33346
rect 35522 33294 35534 33346
rect 35586 33294 35598 33346
rect 33294 33282 33346 33294
rect 37214 33282 37266 33294
rect 2494 33234 2546 33246
rect 2494 33170 2546 33182
rect 2830 33234 2882 33246
rect 17726 33234 17778 33246
rect 3154 33182 3166 33234
rect 3218 33182 3230 33234
rect 6626 33182 6638 33234
rect 6690 33182 6702 33234
rect 14130 33182 14142 33234
rect 14194 33182 14206 33234
rect 14466 33182 14478 33234
rect 14530 33182 14542 33234
rect 17602 33182 17614 33234
rect 17666 33182 17678 33234
rect 2830 33170 2882 33182
rect 17726 33170 17778 33182
rect 17838 33234 17890 33246
rect 24658 33182 24670 33234
rect 24722 33182 24734 33234
rect 33730 33182 33742 33234
rect 33794 33182 33806 33234
rect 17838 33170 17890 33182
rect 4174 33122 4226 33134
rect 4174 33058 4226 33070
rect 5742 33122 5794 33134
rect 13582 33122 13634 33134
rect 8306 33070 8318 33122
rect 8370 33070 8382 33122
rect 5742 33058 5794 33070
rect 13582 33058 13634 33070
rect 15934 33122 15986 33134
rect 15934 33058 15986 33070
rect 16382 33122 16434 33134
rect 16382 33058 16434 33070
rect 18062 33122 18114 33134
rect 18062 33058 18114 33070
rect 18510 33122 18562 33134
rect 18510 33058 18562 33070
rect 22990 33122 23042 33134
rect 22990 33058 23042 33070
rect 23550 33122 23602 33134
rect 23550 33058 23602 33070
rect 25230 33122 25282 33134
rect 25230 33058 25282 33070
rect 29822 33122 29874 33134
rect 29822 33058 29874 33070
rect 30270 33122 30322 33134
rect 30270 33058 30322 33070
rect 30942 33122 30994 33134
rect 30942 33058 30994 33070
rect 31614 33122 31666 33134
rect 31614 33058 31666 33070
rect 31726 33122 31778 33134
rect 31726 33058 31778 33070
rect 32286 33122 32338 33134
rect 32286 33058 32338 33070
rect 32734 33122 32786 33134
rect 32734 33058 32786 33070
rect 1344 32954 38640 32988
rect 1344 32902 14024 32954
rect 14076 32902 14148 32954
rect 14200 32902 14272 32954
rect 14324 32902 14396 32954
rect 14448 32902 14520 32954
rect 14572 32902 14644 32954
rect 14696 32902 14768 32954
rect 14820 32902 14892 32954
rect 14944 32902 15016 32954
rect 15068 32902 15140 32954
rect 15192 32902 34024 32954
rect 34076 32902 34148 32954
rect 34200 32902 34272 32954
rect 34324 32902 34396 32954
rect 34448 32902 34520 32954
rect 34572 32902 34644 32954
rect 34696 32902 34768 32954
rect 34820 32902 34892 32954
rect 34944 32902 35016 32954
rect 35068 32902 35140 32954
rect 35192 32902 38640 32954
rect 1344 32868 38640 32902
rect 4734 32786 4786 32798
rect 4734 32722 4786 32734
rect 5630 32786 5682 32798
rect 5630 32722 5682 32734
rect 6862 32786 6914 32798
rect 6862 32722 6914 32734
rect 12014 32786 12066 32798
rect 15934 32786 15986 32798
rect 15362 32734 15374 32786
rect 15426 32734 15438 32786
rect 12014 32722 12066 32734
rect 15934 32722 15986 32734
rect 16270 32786 16322 32798
rect 16270 32722 16322 32734
rect 16718 32786 16770 32798
rect 16718 32722 16770 32734
rect 17614 32786 17666 32798
rect 17614 32722 17666 32734
rect 18062 32786 18114 32798
rect 25342 32786 25394 32798
rect 23986 32734 23998 32786
rect 24050 32734 24062 32786
rect 18062 32722 18114 32734
rect 25342 32722 25394 32734
rect 25790 32786 25842 32798
rect 25790 32722 25842 32734
rect 31166 32786 31218 32798
rect 31166 32722 31218 32734
rect 31390 32786 31442 32798
rect 31390 32722 31442 32734
rect 31838 32786 31890 32798
rect 31838 32722 31890 32734
rect 32398 32786 32450 32798
rect 32398 32722 32450 32734
rect 34078 32786 34130 32798
rect 34078 32722 34130 32734
rect 36878 32786 36930 32798
rect 36878 32722 36930 32734
rect 36990 32786 37042 32798
rect 36990 32722 37042 32734
rect 37102 32786 37154 32798
rect 37102 32722 37154 32734
rect 6526 32674 6578 32686
rect 6526 32610 6578 32622
rect 6638 32674 6690 32686
rect 6638 32610 6690 32622
rect 26238 32674 26290 32686
rect 30942 32674 30994 32686
rect 27234 32622 27246 32674
rect 27298 32622 27310 32674
rect 27794 32622 27806 32674
rect 27858 32622 27870 32674
rect 26238 32610 26290 32622
rect 30942 32610 30994 32622
rect 32174 32674 32226 32686
rect 32174 32610 32226 32622
rect 34526 32674 34578 32686
rect 37426 32622 37438 32674
rect 37490 32622 37502 32674
rect 34526 32610 34578 32622
rect 7982 32562 8034 32574
rect 7982 32498 8034 32510
rect 12238 32562 12290 32574
rect 21310 32562 21362 32574
rect 27022 32562 27074 32574
rect 12898 32510 12910 32562
rect 12962 32510 12974 32562
rect 21746 32510 21758 32562
rect 21810 32510 21822 32562
rect 12238 32498 12290 32510
rect 21310 32498 21362 32510
rect 27022 32498 27074 32510
rect 33182 32562 33234 32574
rect 33182 32498 33234 32510
rect 33518 32562 33570 32574
rect 33518 32498 33570 32510
rect 34078 32562 34130 32574
rect 37314 32510 37326 32562
rect 37378 32510 37390 32562
rect 34078 32498 34130 32510
rect 5182 32450 5234 32462
rect 5182 32386 5234 32398
rect 6190 32450 6242 32462
rect 6190 32386 6242 32398
rect 7534 32450 7586 32462
rect 7534 32386 7586 32398
rect 35758 32450 35810 32462
rect 35758 32386 35810 32398
rect 24782 32338 24834 32350
rect 5618 32286 5630 32338
rect 5682 32335 5694 32338
rect 6066 32335 6078 32338
rect 5682 32289 6078 32335
rect 5682 32286 5694 32289
rect 6066 32286 6078 32289
rect 6130 32286 6142 32338
rect 24782 32274 24834 32286
rect 26686 32338 26738 32350
rect 26686 32274 26738 32286
rect 31054 32338 31106 32350
rect 31054 32274 31106 32286
rect 32510 32338 32562 32350
rect 32510 32274 32562 32286
rect 33070 32338 33122 32350
rect 33070 32274 33122 32286
rect 33406 32338 33458 32350
rect 33406 32274 33458 32286
rect 1344 32170 38640 32204
rect 1344 32118 4024 32170
rect 4076 32118 4148 32170
rect 4200 32118 4272 32170
rect 4324 32118 4396 32170
rect 4448 32118 4520 32170
rect 4572 32118 4644 32170
rect 4696 32118 4768 32170
rect 4820 32118 4892 32170
rect 4944 32118 5016 32170
rect 5068 32118 5140 32170
rect 5192 32118 24024 32170
rect 24076 32118 24148 32170
rect 24200 32118 24272 32170
rect 24324 32118 24396 32170
rect 24448 32118 24520 32170
rect 24572 32118 24644 32170
rect 24696 32118 24768 32170
rect 24820 32118 24892 32170
rect 24944 32118 25016 32170
rect 25068 32118 25140 32170
rect 25192 32118 38640 32170
rect 1344 32084 38640 32118
rect 6190 32002 6242 32014
rect 14590 32002 14642 32014
rect 32734 32002 32786 32014
rect 13794 31999 13806 32002
rect 6190 31938 6242 31950
rect 13473 31953 13806 31999
rect 3614 31890 3666 31902
rect 3614 31826 3666 31838
rect 8878 31890 8930 31902
rect 12686 31890 12738 31902
rect 11890 31838 11902 31890
rect 11954 31838 11966 31890
rect 8878 31826 8930 31838
rect 12686 31826 12738 31838
rect 5058 31726 5070 31778
rect 5122 31726 5134 31778
rect 9986 31726 9998 31778
rect 10050 31726 10062 31778
rect 13473 31666 13519 31953
rect 13794 31950 13806 31953
rect 13858 31950 13870 32002
rect 16258 31950 16270 32002
rect 16322 31999 16334 32002
rect 16594 31999 16606 32002
rect 16322 31953 16606 31999
rect 16322 31950 16334 31953
rect 16594 31950 16606 31953
rect 16658 31950 16670 32002
rect 14590 31938 14642 31950
rect 32734 31938 32786 31950
rect 16270 31890 16322 31902
rect 16270 31826 16322 31838
rect 16718 31890 16770 31902
rect 16718 31826 16770 31838
rect 22990 31890 23042 31902
rect 22990 31826 23042 31838
rect 23326 31890 23378 31902
rect 23326 31826 23378 31838
rect 36206 31890 36258 31902
rect 36206 31826 36258 31838
rect 37214 31890 37266 31902
rect 37214 31826 37266 31838
rect 14926 31778 14978 31790
rect 17278 31778 17330 31790
rect 15698 31726 15710 31778
rect 15762 31726 15774 31778
rect 17042 31726 17054 31778
rect 17106 31726 17118 31778
rect 14926 31714 14978 31726
rect 17278 31714 17330 31726
rect 18174 31778 18226 31790
rect 18174 31714 18226 31726
rect 18398 31778 18450 31790
rect 18398 31714 18450 31726
rect 22542 31778 22594 31790
rect 26238 31778 26290 31790
rect 23986 31726 23998 31778
rect 24050 31726 24062 31778
rect 22542 31714 22594 31726
rect 26238 31714 26290 31726
rect 27694 31778 27746 31790
rect 27694 31714 27746 31726
rect 29934 31778 29986 31790
rect 29934 31714 29986 31726
rect 30158 31778 30210 31790
rect 30158 31714 30210 31726
rect 30606 31778 30658 31790
rect 30606 31714 30658 31726
rect 31054 31778 31106 31790
rect 32958 31778 33010 31790
rect 31602 31726 31614 31778
rect 31666 31726 31678 31778
rect 32610 31726 32622 31778
rect 32674 31726 32686 31778
rect 31054 31714 31106 31726
rect 32958 31714 33010 31726
rect 33966 31778 34018 31790
rect 34178 31726 34190 31778
rect 34242 31726 34254 31778
rect 33966 31714 34018 31726
rect 13694 31666 13746 31678
rect 17390 31666 17442 31678
rect 5618 31614 5630 31666
rect 5682 31614 5694 31666
rect 13458 31614 13470 31666
rect 13522 31614 13534 31666
rect 15586 31614 15598 31666
rect 15650 31614 15662 31666
rect 13694 31602 13746 31614
rect 17390 31602 17442 31614
rect 18734 31666 18786 31678
rect 25566 31666 25618 31678
rect 23874 31614 23886 31666
rect 23938 31614 23950 31666
rect 18734 31602 18786 31614
rect 25566 31602 25618 31614
rect 26910 31666 26962 31678
rect 30942 31666 30994 31678
rect 28018 31614 28030 31666
rect 28082 31614 28094 31666
rect 28466 31614 28478 31666
rect 28530 31614 28542 31666
rect 26910 31602 26962 31614
rect 30942 31602 30994 31614
rect 34750 31666 34802 31678
rect 34750 31602 34802 31614
rect 2606 31554 2658 31566
rect 2606 31490 2658 31502
rect 4510 31554 4562 31566
rect 4510 31490 4562 31502
rect 7310 31554 7362 31566
rect 7310 31490 7362 31502
rect 7982 31554 8034 31566
rect 7982 31490 8034 31502
rect 8542 31554 8594 31566
rect 8542 31490 8594 31502
rect 14142 31554 14194 31566
rect 18510 31554 18562 31566
rect 17826 31502 17838 31554
rect 17890 31502 17902 31554
rect 14142 31490 14194 31502
rect 18510 31490 18562 31502
rect 25902 31554 25954 31566
rect 25902 31490 25954 31502
rect 26350 31554 26402 31566
rect 26350 31490 26402 31502
rect 26574 31554 26626 31566
rect 26574 31490 26626 31502
rect 27358 31554 27410 31566
rect 27358 31490 27410 31502
rect 29822 31554 29874 31566
rect 29822 31490 29874 31502
rect 30382 31554 30434 31566
rect 30382 31490 30434 31502
rect 32398 31554 32450 31566
rect 33730 31502 33742 31554
rect 33794 31502 33806 31554
rect 32398 31490 32450 31502
rect 1344 31386 38640 31420
rect 1344 31334 14024 31386
rect 14076 31334 14148 31386
rect 14200 31334 14272 31386
rect 14324 31334 14396 31386
rect 14448 31334 14520 31386
rect 14572 31334 14644 31386
rect 14696 31334 14768 31386
rect 14820 31334 14892 31386
rect 14944 31334 15016 31386
rect 15068 31334 15140 31386
rect 15192 31334 34024 31386
rect 34076 31334 34148 31386
rect 34200 31334 34272 31386
rect 34324 31334 34396 31386
rect 34448 31334 34520 31386
rect 34572 31334 34644 31386
rect 34696 31334 34768 31386
rect 34820 31334 34892 31386
rect 34944 31334 35016 31386
rect 35068 31334 35140 31386
rect 35192 31334 38640 31386
rect 1344 31300 38640 31334
rect 2158 31218 2210 31230
rect 2158 31154 2210 31166
rect 9662 31218 9714 31230
rect 9662 31154 9714 31166
rect 15262 31218 15314 31230
rect 15262 31154 15314 31166
rect 16270 31218 16322 31230
rect 16270 31154 16322 31166
rect 16830 31218 16882 31230
rect 33182 31218 33234 31230
rect 28354 31166 28366 31218
rect 28418 31166 28430 31218
rect 16830 31154 16882 31166
rect 33182 31154 33234 31166
rect 2830 31106 2882 31118
rect 2830 31042 2882 31054
rect 3166 31106 3218 31118
rect 3166 31042 3218 31054
rect 15598 31106 15650 31118
rect 15598 31042 15650 31054
rect 29038 31106 29090 31118
rect 36878 31106 36930 31118
rect 30482 31054 30494 31106
rect 30546 31054 30558 31106
rect 34066 31054 34078 31106
rect 34130 31054 34142 31106
rect 35074 31054 35086 31106
rect 35138 31054 35150 31106
rect 29038 31042 29090 31054
rect 36878 31042 36930 31054
rect 15486 30994 15538 31006
rect 5506 30942 5518 30994
rect 5570 30942 5582 30994
rect 8978 30942 8990 30994
rect 9042 30942 9054 30994
rect 15486 30930 15538 30942
rect 17502 30994 17554 31006
rect 17502 30930 17554 30942
rect 17950 30994 18002 31006
rect 17950 30930 18002 30942
rect 25566 30994 25618 31006
rect 31166 30994 31218 31006
rect 26002 30942 26014 30994
rect 26066 30942 26078 30994
rect 30594 30942 30606 30994
rect 30658 30942 30670 30994
rect 32274 30942 32286 30994
rect 32338 30942 32350 30994
rect 33506 30942 33518 30994
rect 33570 30942 33582 30994
rect 35186 30942 35198 30994
rect 35250 30942 35262 30994
rect 25566 30930 25618 30942
rect 31166 30930 31218 30942
rect 2606 30882 2658 30894
rect 13358 30882 13410 30894
rect 3826 30830 3838 30882
rect 3890 30830 3902 30882
rect 6738 30830 6750 30882
rect 6802 30830 6814 30882
rect 2606 30818 2658 30830
rect 13358 30818 13410 30830
rect 14366 30882 14418 30894
rect 14366 30818 14418 30830
rect 14702 30882 14754 30894
rect 29374 30882 29426 30894
rect 17714 30830 17726 30882
rect 17778 30830 17790 30882
rect 14702 30818 14754 30830
rect 29374 30818 29426 30830
rect 29822 30882 29874 30894
rect 32386 30830 32398 30882
rect 32450 30830 32462 30882
rect 29822 30818 29874 30830
rect 15598 30770 15650 30782
rect 15598 30706 15650 30718
rect 17390 30770 17442 30782
rect 17390 30706 17442 30718
rect 18174 30770 18226 30782
rect 18174 30706 18226 30718
rect 31502 30770 31554 30782
rect 31502 30706 31554 30718
rect 1344 30602 38640 30636
rect 1344 30550 4024 30602
rect 4076 30550 4148 30602
rect 4200 30550 4272 30602
rect 4324 30550 4396 30602
rect 4448 30550 4520 30602
rect 4572 30550 4644 30602
rect 4696 30550 4768 30602
rect 4820 30550 4892 30602
rect 4944 30550 5016 30602
rect 5068 30550 5140 30602
rect 5192 30550 24024 30602
rect 24076 30550 24148 30602
rect 24200 30550 24272 30602
rect 24324 30550 24396 30602
rect 24448 30550 24520 30602
rect 24572 30550 24644 30602
rect 24696 30550 24768 30602
rect 24820 30550 24892 30602
rect 24944 30550 25016 30602
rect 25068 30550 25140 30602
rect 25192 30550 38640 30602
rect 1344 30516 38640 30550
rect 6414 30434 6466 30446
rect 26574 30434 26626 30446
rect 10770 30382 10782 30434
rect 10834 30382 10846 30434
rect 6414 30370 6466 30382
rect 26574 30370 26626 30382
rect 26910 30434 26962 30446
rect 26910 30370 26962 30382
rect 29598 30434 29650 30446
rect 30706 30382 30718 30434
rect 30770 30431 30782 30434
rect 31378 30431 31390 30434
rect 30770 30385 31390 30431
rect 30770 30382 30782 30385
rect 31378 30382 31390 30385
rect 31442 30382 31454 30434
rect 36194 30382 36206 30434
rect 36258 30382 36270 30434
rect 29598 30370 29650 30382
rect 6078 30322 6130 30334
rect 4834 30270 4846 30322
rect 4898 30270 4910 30322
rect 6078 30258 6130 30270
rect 7646 30322 7698 30334
rect 30942 30322 30994 30334
rect 16034 30270 16046 30322
rect 16098 30270 16110 30322
rect 7646 30258 7698 30270
rect 30942 30258 30994 30270
rect 2830 30210 2882 30222
rect 2830 30146 2882 30158
rect 3502 30210 3554 30222
rect 3502 30146 3554 30158
rect 4062 30210 4114 30222
rect 4062 30146 4114 30158
rect 5854 30210 5906 30222
rect 5854 30146 5906 30158
rect 7310 30210 7362 30222
rect 11678 30210 11730 30222
rect 16606 30210 16658 30222
rect 20414 30210 20466 30222
rect 8530 30158 8542 30210
rect 8594 30158 8606 30210
rect 10210 30158 10222 30210
rect 10274 30158 10286 30210
rect 12450 30158 12462 30210
rect 12514 30158 12526 30210
rect 14242 30158 14254 30210
rect 14306 30158 14318 30210
rect 19730 30158 19742 30210
rect 19794 30158 19806 30210
rect 7310 30146 7362 30158
rect 11678 30146 11730 30158
rect 16606 30146 16658 30158
rect 20414 30146 20466 30158
rect 20862 30210 20914 30222
rect 20862 30146 20914 30158
rect 21422 30210 21474 30222
rect 31502 30210 31554 30222
rect 27682 30158 27694 30210
rect 27746 30158 27758 30210
rect 31826 30158 31838 30210
rect 31890 30158 31902 30210
rect 32498 30158 32510 30210
rect 32562 30158 32574 30210
rect 34626 30158 34638 30210
rect 34690 30158 34702 30210
rect 21422 30146 21474 30158
rect 31502 30146 31554 30158
rect 3166 30098 3218 30110
rect 3166 30034 3218 30046
rect 3950 30098 4002 30110
rect 3950 30034 4002 30046
rect 4510 30098 4562 30110
rect 4510 30034 4562 30046
rect 7870 30098 7922 30110
rect 28590 30098 28642 30110
rect 8866 30046 8878 30098
rect 8930 30046 8942 30098
rect 12226 30046 12238 30098
rect 12290 30046 12302 30098
rect 27458 30046 27470 30098
rect 27522 30046 27534 30098
rect 29810 30046 29822 30098
rect 29874 30046 29886 30098
rect 30370 30046 30382 30098
rect 30434 30046 30446 30098
rect 7870 30034 7922 30046
rect 28590 30034 28642 30046
rect 2158 29986 2210 29998
rect 2158 29922 2210 29934
rect 2606 29986 2658 29998
rect 2606 29922 2658 29934
rect 3726 29986 3778 29998
rect 3726 29922 3778 29934
rect 4734 29986 4786 29998
rect 4734 29922 4786 29934
rect 7758 29986 7810 29998
rect 7758 29922 7810 29934
rect 11342 29986 11394 29998
rect 26126 29986 26178 29998
rect 17266 29934 17278 29986
rect 17330 29934 17342 29986
rect 11342 29922 11394 29934
rect 26126 29922 26178 29934
rect 29262 29986 29314 29998
rect 29262 29922 29314 29934
rect 1344 29818 38640 29852
rect 1344 29766 14024 29818
rect 14076 29766 14148 29818
rect 14200 29766 14272 29818
rect 14324 29766 14396 29818
rect 14448 29766 14520 29818
rect 14572 29766 14644 29818
rect 14696 29766 14768 29818
rect 14820 29766 14892 29818
rect 14944 29766 15016 29818
rect 15068 29766 15140 29818
rect 15192 29766 34024 29818
rect 34076 29766 34148 29818
rect 34200 29766 34272 29818
rect 34324 29766 34396 29818
rect 34448 29766 34520 29818
rect 34572 29766 34644 29818
rect 34696 29766 34768 29818
rect 34820 29766 34892 29818
rect 34944 29766 35016 29818
rect 35068 29766 35140 29818
rect 35192 29766 38640 29818
rect 1344 29732 38640 29766
rect 5294 29650 5346 29662
rect 4610 29598 4622 29650
rect 4674 29598 4686 29650
rect 5294 29586 5346 29598
rect 10782 29650 10834 29662
rect 17726 29650 17778 29662
rect 14466 29598 14478 29650
rect 14530 29598 14542 29650
rect 10782 29586 10834 29598
rect 17726 29586 17778 29598
rect 19294 29650 19346 29662
rect 19294 29586 19346 29598
rect 21310 29650 21362 29662
rect 21310 29586 21362 29598
rect 26686 29650 26738 29662
rect 26686 29586 26738 29598
rect 5630 29538 5682 29550
rect 5630 29474 5682 29486
rect 5854 29538 5906 29550
rect 10334 29538 10386 29550
rect 17950 29538 18002 29550
rect 8082 29486 8094 29538
rect 8146 29486 8158 29538
rect 15922 29486 15934 29538
rect 15986 29486 15998 29538
rect 16482 29486 16494 29538
rect 16546 29486 16558 29538
rect 5854 29474 5906 29486
rect 10334 29474 10386 29486
rect 17950 29474 18002 29486
rect 22318 29538 22370 29550
rect 29822 29538 29874 29550
rect 23314 29486 23326 29538
rect 23378 29486 23390 29538
rect 23874 29486 23886 29538
rect 23938 29486 23950 29538
rect 22318 29474 22370 29486
rect 29822 29474 29874 29486
rect 33854 29538 33906 29550
rect 33854 29474 33906 29486
rect 1822 29426 1874 29438
rect 11566 29426 11618 29438
rect 15710 29426 15762 29438
rect 2258 29374 2270 29426
rect 2322 29374 2334 29426
rect 7074 29374 7086 29426
rect 7138 29374 7150 29426
rect 8530 29374 8542 29426
rect 8594 29374 8606 29426
rect 9762 29374 9774 29426
rect 9826 29374 9838 29426
rect 11890 29374 11902 29426
rect 11954 29374 11966 29426
rect 1822 29362 1874 29374
rect 11566 29362 11618 29374
rect 15710 29362 15762 29374
rect 17390 29426 17442 29438
rect 17390 29362 17442 29374
rect 17614 29426 17666 29438
rect 23102 29426 23154 29438
rect 18722 29374 18734 29426
rect 18786 29374 18798 29426
rect 17614 29362 17666 29374
rect 23102 29362 23154 29374
rect 27134 29426 27186 29438
rect 30942 29426 30994 29438
rect 27570 29374 27582 29426
rect 27634 29374 27646 29426
rect 27134 29362 27186 29374
rect 30942 29362 30994 29374
rect 33070 29426 33122 29438
rect 33282 29374 33294 29426
rect 33346 29374 33358 29426
rect 33070 29362 33122 29374
rect 31614 29314 31666 29326
rect 8306 29262 8318 29314
rect 8370 29262 8382 29314
rect 9650 29262 9662 29314
rect 9714 29262 9726 29314
rect 31614 29250 31666 29262
rect 5518 29202 5570 29214
rect 5518 29138 5570 29150
rect 15038 29202 15090 29214
rect 15038 29138 15090 29150
rect 15374 29202 15426 29214
rect 15374 29138 15426 29150
rect 22766 29202 22818 29214
rect 22766 29138 22818 29150
rect 30606 29202 30658 29214
rect 30606 29138 30658 29150
rect 1344 29034 38640 29068
rect 1344 28982 4024 29034
rect 4076 28982 4148 29034
rect 4200 28982 4272 29034
rect 4324 28982 4396 29034
rect 4448 28982 4520 29034
rect 4572 28982 4644 29034
rect 4696 28982 4768 29034
rect 4820 28982 4892 29034
rect 4944 28982 5016 29034
rect 5068 28982 5140 29034
rect 5192 28982 24024 29034
rect 24076 28982 24148 29034
rect 24200 28982 24272 29034
rect 24324 28982 24396 29034
rect 24448 28982 24520 29034
rect 24572 28982 24644 29034
rect 24696 28982 24768 29034
rect 24820 28982 24892 29034
rect 24944 28982 25016 29034
rect 25068 28982 25140 29034
rect 25192 28982 38640 29034
rect 1344 28948 38640 28982
rect 3166 28866 3218 28878
rect 3166 28802 3218 28814
rect 3502 28866 3554 28878
rect 3502 28802 3554 28814
rect 4958 28866 5010 28878
rect 4958 28802 5010 28814
rect 13022 28866 13074 28878
rect 13022 28802 13074 28814
rect 13582 28866 13634 28878
rect 13582 28802 13634 28814
rect 13918 28866 13970 28878
rect 13918 28802 13970 28814
rect 22654 28866 22706 28878
rect 22654 28802 22706 28814
rect 22990 28866 23042 28878
rect 22990 28802 23042 28814
rect 19742 28754 19794 28766
rect 7858 28702 7870 28754
rect 7922 28702 7934 28754
rect 19742 28690 19794 28702
rect 21646 28754 21698 28766
rect 21646 28690 21698 28702
rect 21982 28754 22034 28766
rect 26674 28702 26686 28754
rect 26738 28702 26750 28754
rect 21982 28690 22034 28702
rect 2494 28642 2546 28654
rect 4174 28642 4226 28654
rect 3154 28590 3166 28642
rect 3218 28590 3230 28642
rect 2494 28578 2546 28590
rect 4174 28578 4226 28590
rect 4510 28642 4562 28654
rect 4510 28578 4562 28590
rect 5630 28642 5682 28654
rect 5630 28578 5682 28590
rect 5854 28642 5906 28654
rect 9550 28642 9602 28654
rect 18958 28642 19010 28654
rect 6962 28590 6974 28642
rect 7026 28590 7038 28642
rect 9986 28590 9998 28642
rect 10050 28590 10062 28642
rect 14354 28590 14366 28642
rect 14418 28590 14430 28642
rect 18274 28590 18286 28642
rect 18338 28590 18350 28642
rect 5854 28578 5906 28590
rect 9550 28578 9602 28590
rect 18958 28578 19010 28590
rect 19294 28642 19346 28654
rect 28142 28642 28194 28654
rect 23426 28590 23438 28642
rect 23490 28590 23502 28642
rect 25442 28590 25454 28642
rect 25506 28590 25518 28642
rect 19294 28578 19346 28590
rect 28142 28578 28194 28590
rect 2270 28530 2322 28542
rect 2270 28466 2322 28478
rect 2830 28530 2882 28542
rect 2830 28466 2882 28478
rect 3950 28530 4002 28542
rect 3950 28466 4002 28478
rect 4846 28530 4898 28542
rect 4846 28466 4898 28478
rect 4958 28530 5010 28542
rect 14690 28478 14702 28530
rect 14754 28478 14766 28530
rect 23538 28478 23550 28530
rect 23602 28478 23614 28530
rect 4958 28466 5010 28478
rect 4286 28418 4338 28430
rect 15262 28418 15314 28430
rect 6178 28366 6190 28418
rect 6242 28366 6254 28418
rect 12450 28366 12462 28418
rect 12514 28366 12526 28418
rect 15810 28366 15822 28418
rect 15874 28366 15886 28418
rect 4286 28354 4338 28366
rect 15262 28354 15314 28366
rect 1344 28250 38640 28284
rect 1344 28198 14024 28250
rect 14076 28198 14148 28250
rect 14200 28198 14272 28250
rect 14324 28198 14396 28250
rect 14448 28198 14520 28250
rect 14572 28198 14644 28250
rect 14696 28198 14768 28250
rect 14820 28198 14892 28250
rect 14944 28198 15016 28250
rect 15068 28198 15140 28250
rect 15192 28198 34024 28250
rect 34076 28198 34148 28250
rect 34200 28198 34272 28250
rect 34324 28198 34396 28250
rect 34448 28198 34520 28250
rect 34572 28198 34644 28250
rect 34696 28198 34768 28250
rect 34820 28198 34892 28250
rect 34944 28198 35016 28250
rect 35068 28198 35140 28250
rect 35192 28198 38640 28250
rect 1344 28164 38640 28198
rect 1598 28082 1650 28094
rect 12014 28082 12066 28094
rect 2258 28030 2270 28082
rect 2322 28030 2334 28082
rect 10098 28030 10110 28082
rect 10162 28030 10174 28082
rect 1598 28018 1650 28030
rect 12014 28018 12066 28030
rect 15486 28082 15538 28094
rect 15486 28018 15538 28030
rect 16830 28082 16882 28094
rect 16830 28018 16882 28030
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 17726 28082 17778 28094
rect 17726 28018 17778 28030
rect 17950 28082 18002 28094
rect 17950 28018 18002 28030
rect 18398 28082 18450 28094
rect 18398 28018 18450 28030
rect 18846 28082 18898 28094
rect 25342 28082 25394 28094
rect 23650 28030 23662 28082
rect 23714 28030 23726 28082
rect 18846 28018 18898 28030
rect 25342 28018 25394 28030
rect 29710 28082 29762 28094
rect 29710 28018 29762 28030
rect 9550 27970 9602 27982
rect 14254 27970 14306 27982
rect 6738 27918 6750 27970
rect 6802 27918 6814 27970
rect 12674 27918 12686 27970
rect 12738 27918 12750 27970
rect 13122 27918 13134 27970
rect 13186 27918 13198 27970
rect 9550 27906 9602 27918
rect 14254 27906 14306 27918
rect 14366 27970 14418 27982
rect 14366 27906 14418 27918
rect 14590 27970 14642 27982
rect 14590 27906 14642 27918
rect 15710 27970 15762 27982
rect 30046 27970 30098 27982
rect 31726 27970 31778 27982
rect 20290 27918 20302 27970
rect 20354 27918 20366 27970
rect 30818 27918 30830 27970
rect 30882 27918 30894 27970
rect 31378 27918 31390 27970
rect 31442 27918 31454 27970
rect 15710 27906 15762 27918
rect 30046 27906 30098 27918
rect 31726 27906 31778 27918
rect 5294 27858 5346 27870
rect 4722 27806 4734 27858
rect 4786 27806 4798 27858
rect 5294 27794 5346 27806
rect 5966 27858 6018 27870
rect 5966 27794 6018 27806
rect 6190 27858 6242 27870
rect 6190 27794 6242 27806
rect 6414 27858 6466 27870
rect 13918 27858 13970 27870
rect 7522 27806 7534 27858
rect 7586 27806 7598 27858
rect 6414 27794 6466 27806
rect 13918 27794 13970 27806
rect 15822 27858 15874 27870
rect 15822 27794 15874 27806
rect 17838 27858 17890 27870
rect 17838 27794 17890 27806
rect 19630 27858 19682 27870
rect 20974 27858 21026 27870
rect 20066 27806 20078 27858
rect 20130 27806 20142 27858
rect 21410 27806 21422 27858
rect 21474 27806 21486 27858
rect 30594 27806 30606 27858
rect 30658 27806 30670 27858
rect 19630 27794 19682 27806
rect 20974 27794 21026 27806
rect 5630 27746 5682 27758
rect 11566 27746 11618 27758
rect 7634 27694 7646 27746
rect 7698 27694 7710 27746
rect 8866 27694 8878 27746
rect 8930 27694 8942 27746
rect 5630 27682 5682 27694
rect 11566 27682 11618 27694
rect 12350 27746 12402 27758
rect 12350 27682 12402 27694
rect 15262 27746 15314 27758
rect 15262 27682 15314 27694
rect 16382 27746 16434 27758
rect 16382 27682 16434 27694
rect 24446 27746 24498 27758
rect 24446 27682 24498 27694
rect 25790 27746 25842 27758
rect 25790 27682 25842 27694
rect 5518 27634 5570 27646
rect 5518 27570 5570 27582
rect 9774 27634 9826 27646
rect 9774 27570 9826 27582
rect 19294 27634 19346 27646
rect 19294 27570 19346 27582
rect 30158 27634 30210 27646
rect 30158 27570 30210 27582
rect 1344 27466 38640 27500
rect 1344 27414 4024 27466
rect 4076 27414 4148 27466
rect 4200 27414 4272 27466
rect 4324 27414 4396 27466
rect 4448 27414 4520 27466
rect 4572 27414 4644 27466
rect 4696 27414 4768 27466
rect 4820 27414 4892 27466
rect 4944 27414 5016 27466
rect 5068 27414 5140 27466
rect 5192 27414 24024 27466
rect 24076 27414 24148 27466
rect 24200 27414 24272 27466
rect 24324 27414 24396 27466
rect 24448 27414 24520 27466
rect 24572 27414 24644 27466
rect 24696 27414 24768 27466
rect 24820 27414 24892 27466
rect 24944 27414 25016 27466
rect 25068 27414 25140 27466
rect 25192 27414 38640 27466
rect 1344 27380 38640 27414
rect 3614 27298 3666 27310
rect 3614 27234 3666 27246
rect 4734 27298 4786 27310
rect 7086 27298 7138 27310
rect 8318 27298 8370 27310
rect 19630 27298 19682 27310
rect 6402 27246 6414 27298
rect 6466 27246 6478 27298
rect 7410 27246 7422 27298
rect 7474 27246 7486 27298
rect 8642 27246 8654 27298
rect 8706 27246 8718 27298
rect 4734 27234 4786 27246
rect 7086 27234 7138 27246
rect 8318 27234 8370 27246
rect 19630 27234 19682 27246
rect 25678 27298 25730 27310
rect 25890 27246 25902 27298
rect 25954 27295 25966 27298
rect 26450 27295 26462 27298
rect 25954 27249 26462 27295
rect 25954 27246 25966 27249
rect 26450 27246 26462 27249
rect 26514 27246 26526 27298
rect 25678 27234 25730 27246
rect 3390 27186 3442 27198
rect 3390 27122 3442 27134
rect 5070 27186 5122 27198
rect 5070 27122 5122 27134
rect 6078 27186 6130 27198
rect 6078 27122 6130 27134
rect 9326 27186 9378 27198
rect 9326 27122 9378 27134
rect 9774 27186 9826 27198
rect 9774 27122 9826 27134
rect 13022 27186 13074 27198
rect 13022 27122 13074 27134
rect 13694 27186 13746 27198
rect 13694 27122 13746 27134
rect 14030 27186 14082 27198
rect 14030 27122 14082 27134
rect 15150 27186 15202 27198
rect 15150 27122 15202 27134
rect 16942 27186 16994 27198
rect 16942 27122 16994 27134
rect 17390 27186 17442 27198
rect 17390 27122 17442 27134
rect 26014 27186 26066 27198
rect 26014 27122 26066 27134
rect 26462 27186 26514 27198
rect 26462 27122 26514 27134
rect 2158 27074 2210 27086
rect 4958 27074 5010 27086
rect 6862 27074 6914 27086
rect 4162 27022 4174 27074
rect 4226 27022 4238 27074
rect 4498 27022 4510 27074
rect 4562 27022 4574 27074
rect 5618 27022 5630 27074
rect 5682 27022 5694 27074
rect 2158 27010 2210 27022
rect 4958 27010 5010 27022
rect 2942 26962 2994 26974
rect 2942 26898 2994 26910
rect 3950 26962 4002 26974
rect 3950 26898 4002 26910
rect 2606 26850 2658 26862
rect 2606 26786 2658 26798
rect 3726 26850 3778 26862
rect 5633 26850 5679 27022
rect 6862 27010 6914 27022
rect 8094 27074 8146 27086
rect 8094 27010 8146 27022
rect 18846 27074 18898 27086
rect 18846 27010 18898 27022
rect 22206 27074 22258 27086
rect 29710 27074 29762 27086
rect 22642 27022 22654 27074
rect 22706 27022 22718 27074
rect 22206 27010 22258 27022
rect 29710 27010 29762 27022
rect 29934 27074 29986 27086
rect 33966 27074 34018 27086
rect 30258 27022 30270 27074
rect 30322 27022 30334 27074
rect 30706 27022 30718 27074
rect 30770 27022 30782 27074
rect 29934 27010 29986 27022
rect 33966 27010 34018 27022
rect 5854 26962 5906 26974
rect 5854 26898 5906 26910
rect 14702 26962 14754 26974
rect 24894 26962 24946 26974
rect 19842 26910 19854 26962
rect 19906 26910 19918 26962
rect 20402 26910 20414 26962
rect 20466 26910 20478 26962
rect 14702 26898 14754 26910
rect 24894 26898 24946 26910
rect 29374 26962 29426 26974
rect 29374 26898 29426 26910
rect 33070 26962 33122 26974
rect 33070 26898 33122 26910
rect 19294 26850 19346 26862
rect 5618 26798 5630 26850
rect 5682 26798 5694 26850
rect 3726 26786 3778 26798
rect 19294 26786 19346 26798
rect 29822 26850 29874 26862
rect 29822 26786 29874 26798
rect 1344 26682 38640 26716
rect 1344 26630 14024 26682
rect 14076 26630 14148 26682
rect 14200 26630 14272 26682
rect 14324 26630 14396 26682
rect 14448 26630 14520 26682
rect 14572 26630 14644 26682
rect 14696 26630 14768 26682
rect 14820 26630 14892 26682
rect 14944 26630 15016 26682
rect 15068 26630 15140 26682
rect 15192 26630 34024 26682
rect 34076 26630 34148 26682
rect 34200 26630 34272 26682
rect 34324 26630 34396 26682
rect 34448 26630 34520 26682
rect 34572 26630 34644 26682
rect 34696 26630 34768 26682
rect 34820 26630 34892 26682
rect 34944 26630 35016 26682
rect 35068 26630 35140 26682
rect 35192 26630 38640 26682
rect 1344 26596 38640 26630
rect 3502 26514 3554 26526
rect 3502 26450 3554 26462
rect 3838 26514 3890 26526
rect 3838 26450 3890 26462
rect 4846 26514 4898 26526
rect 4846 26450 4898 26462
rect 7086 26514 7138 26526
rect 7086 26450 7138 26462
rect 7758 26514 7810 26526
rect 7758 26450 7810 26462
rect 8318 26514 8370 26526
rect 21758 26514 21810 26526
rect 21186 26462 21198 26514
rect 21250 26462 21262 26514
rect 8318 26450 8370 26462
rect 21758 26450 21810 26462
rect 23214 26514 23266 26526
rect 23214 26450 23266 26462
rect 6750 26402 6802 26414
rect 26350 26402 26402 26414
rect 22082 26350 22094 26402
rect 22146 26350 22158 26402
rect 22642 26350 22654 26402
rect 22706 26350 22718 26402
rect 6750 26338 6802 26350
rect 26350 26338 26402 26350
rect 26462 26402 26514 26414
rect 30370 26350 30382 26402
rect 30434 26350 30446 26402
rect 30594 26350 30606 26402
rect 30658 26350 30670 26402
rect 26462 26338 26514 26350
rect 5294 26290 5346 26302
rect 4610 26238 4622 26290
rect 4674 26238 4686 26290
rect 5294 26226 5346 26238
rect 6414 26290 6466 26302
rect 6414 26226 6466 26238
rect 6638 26290 6690 26302
rect 6638 26226 6690 26238
rect 7198 26290 7250 26302
rect 26686 26290 26738 26302
rect 18162 26238 18174 26290
rect 18226 26238 18238 26290
rect 18722 26238 18734 26290
rect 18786 26238 18798 26290
rect 7198 26226 7250 26238
rect 26686 26226 26738 26238
rect 30942 26290 30994 26302
rect 30942 26226 30994 26238
rect 4286 26178 4338 26190
rect 4286 26114 4338 26126
rect 23774 26178 23826 26190
rect 23774 26114 23826 26126
rect 26014 26178 26066 26190
rect 26014 26114 26066 26126
rect 29262 26178 29314 26190
rect 29262 26114 29314 26126
rect 29710 26178 29762 26190
rect 29710 26114 29762 26126
rect 4958 26066 5010 26078
rect 3714 26014 3726 26066
rect 3778 26063 3790 26066
rect 4274 26063 4286 26066
rect 3778 26017 4286 26063
rect 3778 26014 3790 26017
rect 4274 26014 4286 26017
rect 4338 26014 4350 26066
rect 4958 26002 5010 26014
rect 5518 26066 5570 26078
rect 6302 26066 6354 26078
rect 5842 26014 5854 26066
rect 5906 26014 5918 26066
rect 5518 26002 5570 26014
rect 6302 26002 6354 26014
rect 22878 26066 22930 26078
rect 31278 26066 31330 26078
rect 29362 26014 29374 26066
rect 29426 26063 29438 26066
rect 29810 26063 29822 26066
rect 29426 26017 29822 26063
rect 29426 26014 29438 26017
rect 29810 26014 29822 26017
rect 29874 26014 29886 26066
rect 22878 26002 22930 26014
rect 31278 26002 31330 26014
rect 1344 25898 38640 25932
rect 1344 25846 4024 25898
rect 4076 25846 4148 25898
rect 4200 25846 4272 25898
rect 4324 25846 4396 25898
rect 4448 25846 4520 25898
rect 4572 25846 4644 25898
rect 4696 25846 4768 25898
rect 4820 25846 4892 25898
rect 4944 25846 5016 25898
rect 5068 25846 5140 25898
rect 5192 25846 24024 25898
rect 24076 25846 24148 25898
rect 24200 25846 24272 25898
rect 24324 25846 24396 25898
rect 24448 25846 24520 25898
rect 24572 25846 24644 25898
rect 24696 25846 24768 25898
rect 24820 25846 24892 25898
rect 24944 25846 25016 25898
rect 25068 25846 25140 25898
rect 25192 25846 38640 25898
rect 1344 25812 38640 25846
rect 5630 25730 5682 25742
rect 5630 25666 5682 25678
rect 5742 25730 5794 25742
rect 5742 25666 5794 25678
rect 5966 25730 6018 25742
rect 5966 25666 6018 25678
rect 9998 25730 10050 25742
rect 9998 25666 10050 25678
rect 23774 25730 23826 25742
rect 23774 25666 23826 25678
rect 34190 25730 34242 25742
rect 34190 25666 34242 25678
rect 4174 25618 4226 25630
rect 4174 25554 4226 25566
rect 5070 25618 5122 25630
rect 5070 25554 5122 25566
rect 7646 25618 7698 25630
rect 7646 25554 7698 25566
rect 8094 25618 8146 25630
rect 8094 25554 8146 25566
rect 14030 25618 14082 25630
rect 14030 25554 14082 25566
rect 21982 25618 22034 25630
rect 30158 25618 30210 25630
rect 29586 25566 29598 25618
rect 29650 25566 29662 25618
rect 21982 25554 22034 25566
rect 30158 25554 30210 25566
rect 6078 25506 6130 25518
rect 6078 25442 6130 25454
rect 14702 25506 14754 25518
rect 27470 25506 27522 25518
rect 30718 25506 30770 25518
rect 26786 25454 26798 25506
rect 26850 25454 26862 25506
rect 29362 25454 29374 25506
rect 29426 25454 29438 25506
rect 31154 25454 31166 25506
rect 31218 25454 31230 25506
rect 14702 25442 14754 25454
rect 27470 25442 27522 25454
rect 30718 25442 30770 25454
rect 4734 25394 4786 25406
rect 14366 25394 14418 25406
rect 10210 25342 10222 25394
rect 10274 25342 10286 25394
rect 10546 25342 10558 25394
rect 10610 25342 10622 25394
rect 4734 25330 4786 25342
rect 14366 25330 14418 25342
rect 14478 25394 14530 25406
rect 14478 25330 14530 25342
rect 27918 25394 27970 25406
rect 27918 25330 27970 25342
rect 6862 25282 6914 25294
rect 6862 25218 6914 25230
rect 9214 25282 9266 25294
rect 9214 25218 9266 25230
rect 9662 25282 9714 25294
rect 9662 25218 9714 25230
rect 13582 25282 13634 25294
rect 13582 25218 13634 25230
rect 15038 25282 15090 25294
rect 15038 25218 15090 25230
rect 22318 25282 22370 25294
rect 28254 25282 28306 25294
rect 24546 25230 24558 25282
rect 24610 25230 24622 25282
rect 33394 25230 33406 25282
rect 33458 25230 33470 25282
rect 22318 25218 22370 25230
rect 28254 25218 28306 25230
rect 1344 25114 38640 25148
rect 1344 25062 14024 25114
rect 14076 25062 14148 25114
rect 14200 25062 14272 25114
rect 14324 25062 14396 25114
rect 14448 25062 14520 25114
rect 14572 25062 14644 25114
rect 14696 25062 14768 25114
rect 14820 25062 14892 25114
rect 14944 25062 15016 25114
rect 15068 25062 15140 25114
rect 15192 25062 34024 25114
rect 34076 25062 34148 25114
rect 34200 25062 34272 25114
rect 34324 25062 34396 25114
rect 34448 25062 34520 25114
rect 34572 25062 34644 25114
rect 34696 25062 34768 25114
rect 34820 25062 34892 25114
rect 34944 25062 35016 25114
rect 35068 25062 35140 25114
rect 35192 25062 38640 25114
rect 1344 25028 38640 25062
rect 1822 24946 1874 24958
rect 8542 24946 8594 24958
rect 3154 24894 3166 24946
rect 3218 24894 3230 24946
rect 1822 24882 1874 24894
rect 8542 24882 8594 24894
rect 12574 24946 12626 24958
rect 12574 24882 12626 24894
rect 13022 24946 13074 24958
rect 13022 24882 13074 24894
rect 18734 24946 18786 24958
rect 18734 24882 18786 24894
rect 26126 24946 26178 24958
rect 26126 24882 26178 24894
rect 26686 24946 26738 24958
rect 26686 24882 26738 24894
rect 28478 24946 28530 24958
rect 29922 24894 29934 24946
rect 29986 24894 29998 24946
rect 28478 24882 28530 24894
rect 24670 24834 24722 24846
rect 10770 24782 10782 24834
rect 10834 24782 10846 24834
rect 14018 24782 14030 24834
rect 14082 24782 14094 24834
rect 14354 24782 14366 24834
rect 14418 24782 14430 24834
rect 15362 24782 15374 24834
rect 15426 24782 15438 24834
rect 19730 24782 19742 24834
rect 19794 24782 19806 24834
rect 20290 24782 20302 24834
rect 20354 24782 20366 24834
rect 24670 24770 24722 24782
rect 25454 24834 25506 24846
rect 25454 24770 25506 24782
rect 27134 24834 27186 24846
rect 27134 24770 27186 24782
rect 27470 24834 27522 24846
rect 27470 24770 27522 24782
rect 2830 24722 2882 24734
rect 2830 24658 2882 24670
rect 3838 24722 3890 24734
rect 8990 24722 9042 24734
rect 8082 24670 8094 24722
rect 8146 24670 8158 24722
rect 3838 24658 3890 24670
rect 8990 24658 9042 24670
rect 9998 24722 10050 24734
rect 13806 24722 13858 24734
rect 19518 24722 19570 24734
rect 10546 24670 10558 24722
rect 10610 24670 10622 24722
rect 15474 24670 15486 24722
rect 15538 24670 15550 24722
rect 9998 24658 10050 24670
rect 13806 24658 13858 24670
rect 19518 24658 19570 24670
rect 26462 24722 26514 24734
rect 26462 24658 26514 24670
rect 26910 24722 26962 24734
rect 26910 24658 26962 24670
rect 27806 24722 27858 24734
rect 27806 24658 27858 24670
rect 28142 24722 28194 24734
rect 28142 24658 28194 24670
rect 28814 24722 28866 24734
rect 29598 24722 29650 24734
rect 29362 24670 29374 24722
rect 29426 24670 29438 24722
rect 30258 24670 30270 24722
rect 30322 24670 30334 24722
rect 28814 24658 28866 24670
rect 29598 24658 29650 24670
rect 2494 24610 2546 24622
rect 2494 24546 2546 24558
rect 5294 24610 5346 24622
rect 5294 24546 5346 24558
rect 11566 24610 11618 24622
rect 18286 24610 18338 24622
rect 16594 24558 16606 24610
rect 16658 24558 16670 24610
rect 11566 24546 11618 24558
rect 18286 24546 18338 24558
rect 25790 24610 25842 24622
rect 25790 24546 25842 24558
rect 27918 24610 27970 24622
rect 27918 24546 27970 24558
rect 30942 24610 30994 24622
rect 30942 24546 30994 24558
rect 31390 24610 31442 24622
rect 31390 24546 31442 24558
rect 31838 24610 31890 24622
rect 31838 24546 31890 24558
rect 9662 24498 9714 24510
rect 9662 24434 9714 24446
rect 13470 24498 13522 24510
rect 13470 24434 13522 24446
rect 19182 24498 19234 24510
rect 19182 24434 19234 24446
rect 25230 24498 25282 24510
rect 25230 24434 25282 24446
rect 26014 24498 26066 24510
rect 26014 24434 26066 24446
rect 27022 24498 27074 24510
rect 27022 24434 27074 24446
rect 1344 24330 38640 24364
rect 1344 24278 4024 24330
rect 4076 24278 4148 24330
rect 4200 24278 4272 24330
rect 4324 24278 4396 24330
rect 4448 24278 4520 24330
rect 4572 24278 4644 24330
rect 4696 24278 4768 24330
rect 4820 24278 4892 24330
rect 4944 24278 5016 24330
rect 5068 24278 5140 24330
rect 5192 24278 24024 24330
rect 24076 24278 24148 24330
rect 24200 24278 24272 24330
rect 24324 24278 24396 24330
rect 24448 24278 24520 24330
rect 24572 24278 24644 24330
rect 24696 24278 24768 24330
rect 24820 24278 24892 24330
rect 24944 24278 25016 24330
rect 25068 24278 25140 24330
rect 25192 24278 38640 24330
rect 1344 24244 38640 24278
rect 11342 24162 11394 24174
rect 11342 24098 11394 24110
rect 19630 24162 19682 24174
rect 19630 24098 19682 24110
rect 30494 24162 30546 24174
rect 30494 24098 30546 24110
rect 30606 24162 30658 24174
rect 30606 24098 30658 24110
rect 31054 24050 31106 24062
rect 6626 23998 6638 24050
rect 6690 23998 6702 24050
rect 24546 23998 24558 24050
rect 24610 23998 24622 24050
rect 27794 23998 27806 24050
rect 27858 23998 27870 24050
rect 31054 23986 31106 23998
rect 2158 23938 2210 23950
rect 7870 23938 7922 23950
rect 11566 23938 11618 23950
rect 23102 23938 23154 23950
rect 24894 23938 24946 23950
rect 7410 23886 7422 23938
rect 7474 23886 7486 23938
rect 8306 23886 8318 23938
rect 8370 23886 8382 23938
rect 13458 23886 13470 23938
rect 13522 23886 13534 23938
rect 13906 23886 13918 23938
rect 13970 23886 13982 23938
rect 24434 23886 24446 23938
rect 24498 23886 24510 23938
rect 2158 23874 2210 23886
rect 7870 23874 7922 23886
rect 11566 23874 11618 23886
rect 23102 23874 23154 23886
rect 24894 23874 24946 23886
rect 25006 23938 25058 23950
rect 29038 23938 29090 23950
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 25006 23874 25058 23886
rect 29038 23874 29090 23886
rect 29486 23938 29538 23950
rect 29486 23874 29538 23886
rect 30158 23938 30210 23950
rect 30158 23874 30210 23886
rect 30270 23938 30322 23950
rect 30270 23874 30322 23886
rect 4510 23826 4562 23838
rect 11678 23826 11730 23838
rect 2818 23774 2830 23826
rect 2882 23774 2894 23826
rect 6178 23774 6190 23826
rect 6242 23774 6254 23826
rect 4510 23762 4562 23774
rect 11678 23762 11730 23774
rect 18846 23826 18898 23838
rect 22766 23826 22818 23838
rect 19842 23774 19854 23826
rect 19906 23774 19918 23826
rect 20402 23774 20414 23826
rect 20466 23774 20478 23826
rect 18846 23762 18898 23774
rect 22766 23762 22818 23774
rect 1934 23714 1986 23726
rect 1934 23650 1986 23662
rect 2494 23714 2546 23726
rect 2494 23650 2546 23662
rect 3390 23714 3442 23726
rect 3390 23650 3442 23662
rect 4398 23714 4450 23726
rect 4398 23650 4450 23662
rect 5070 23714 5122 23726
rect 11902 23714 11954 23726
rect 10770 23662 10782 23714
rect 10834 23662 10846 23714
rect 5070 23650 5122 23662
rect 11902 23650 11954 23662
rect 12238 23714 12290 23726
rect 17054 23714 17106 23726
rect 16482 23662 16494 23714
rect 16546 23662 16558 23714
rect 12238 23650 12290 23662
rect 17054 23650 17106 23662
rect 17390 23714 17442 23726
rect 17390 23650 17442 23662
rect 17838 23714 17890 23726
rect 17838 23650 17890 23662
rect 19294 23714 19346 23726
rect 19294 23650 19346 23662
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 21870 23714 21922 23726
rect 21870 23650 21922 23662
rect 22430 23714 22482 23726
rect 22430 23650 22482 23662
rect 22878 23714 22930 23726
rect 22878 23650 22930 23662
rect 24110 23714 24162 23726
rect 24110 23650 24162 23662
rect 24670 23714 24722 23726
rect 24670 23650 24722 23662
rect 28478 23714 28530 23726
rect 28478 23650 28530 23662
rect 29598 23714 29650 23726
rect 29598 23650 29650 23662
rect 29710 23714 29762 23726
rect 29710 23650 29762 23662
rect 31502 23714 31554 23726
rect 31502 23650 31554 23662
rect 31950 23714 32002 23726
rect 31950 23650 32002 23662
rect 1344 23546 38640 23580
rect 1344 23494 14024 23546
rect 14076 23494 14148 23546
rect 14200 23494 14272 23546
rect 14324 23494 14396 23546
rect 14448 23494 14520 23546
rect 14572 23494 14644 23546
rect 14696 23494 14768 23546
rect 14820 23494 14892 23546
rect 14944 23494 15016 23546
rect 15068 23494 15140 23546
rect 15192 23494 34024 23546
rect 34076 23494 34148 23546
rect 34200 23494 34272 23546
rect 34324 23494 34396 23546
rect 34448 23494 34520 23546
rect 34572 23494 34644 23546
rect 34696 23494 34768 23546
rect 34820 23494 34892 23546
rect 34944 23494 35016 23546
rect 35068 23494 35140 23546
rect 35192 23494 38640 23546
rect 1344 23460 38640 23494
rect 3838 23378 3890 23390
rect 3838 23314 3890 23326
rect 4062 23378 4114 23390
rect 15150 23378 15202 23390
rect 5170 23326 5182 23378
rect 5234 23326 5246 23378
rect 4062 23314 4114 23326
rect 15150 23314 15202 23326
rect 21758 23378 21810 23390
rect 31614 23378 31666 23390
rect 28130 23326 28142 23378
rect 28194 23326 28206 23378
rect 21758 23314 21810 23326
rect 31614 23314 31666 23326
rect 1934 23266 1986 23278
rect 1934 23202 1986 23214
rect 2270 23266 2322 23278
rect 13806 23266 13858 23278
rect 20974 23266 21026 23278
rect 5394 23214 5406 23266
rect 5458 23214 5470 23266
rect 16258 23214 16270 23266
rect 16322 23214 16334 23266
rect 16482 23214 16494 23266
rect 16546 23214 16558 23266
rect 2270 23202 2322 23214
rect 13806 23202 13858 23214
rect 20974 23202 21026 23214
rect 25342 23266 25394 23278
rect 25342 23202 25394 23214
rect 27022 23266 27074 23278
rect 27022 23202 27074 23214
rect 2606 23154 2658 23166
rect 2606 23090 2658 23102
rect 4286 23154 4338 23166
rect 11118 23154 11170 23166
rect 14590 23154 14642 23166
rect 5282 23102 5294 23154
rect 5346 23102 5358 23154
rect 5954 23102 5966 23154
rect 6018 23102 6030 23154
rect 11554 23102 11566 23154
rect 11618 23102 11630 23154
rect 4286 23090 4338 23102
rect 11118 23090 11170 23102
rect 14590 23090 14642 23102
rect 15934 23154 15986 23166
rect 15934 23090 15986 23102
rect 18286 23154 18338 23166
rect 31054 23154 31106 23166
rect 18722 23102 18734 23154
rect 18786 23102 18798 23154
rect 21970 23102 21982 23154
rect 22034 23102 22046 23154
rect 26338 23102 26350 23154
rect 26402 23102 26414 23154
rect 30594 23102 30606 23154
rect 30658 23102 30670 23154
rect 18286 23090 18338 23102
rect 31054 23090 31106 23102
rect 3950 23042 4002 23054
rect 17502 23042 17554 23054
rect 3378 22990 3390 23042
rect 3442 22990 3454 23042
rect 8082 22990 8094 23042
rect 8146 22990 8158 23042
rect 23650 22990 23662 23042
rect 23714 22990 23726 23042
rect 26674 22990 26686 23042
rect 26738 22990 26750 23042
rect 3950 22978 4002 22990
rect 17502 22978 17554 22990
rect 4510 22930 4562 22942
rect 4510 22866 4562 22878
rect 15598 22930 15650 22942
rect 15598 22866 15650 22878
rect 27582 22930 27634 22942
rect 27582 22866 27634 22878
rect 1344 22762 38640 22796
rect 1344 22710 4024 22762
rect 4076 22710 4148 22762
rect 4200 22710 4272 22762
rect 4324 22710 4396 22762
rect 4448 22710 4520 22762
rect 4572 22710 4644 22762
rect 4696 22710 4768 22762
rect 4820 22710 4892 22762
rect 4944 22710 5016 22762
rect 5068 22710 5140 22762
rect 5192 22710 24024 22762
rect 24076 22710 24148 22762
rect 24200 22710 24272 22762
rect 24324 22710 24396 22762
rect 24448 22710 24520 22762
rect 24572 22710 24644 22762
rect 24696 22710 24768 22762
rect 24820 22710 24892 22762
rect 24944 22710 25016 22762
rect 25068 22710 25140 22762
rect 25192 22710 38640 22762
rect 1344 22676 38640 22710
rect 4174 22594 4226 22606
rect 4174 22530 4226 22542
rect 13582 22594 13634 22606
rect 13582 22530 13634 22542
rect 13918 22594 13970 22606
rect 29150 22594 29202 22606
rect 28130 22542 28142 22594
rect 28194 22542 28206 22594
rect 13918 22530 13970 22542
rect 29150 22530 29202 22542
rect 20862 22482 20914 22494
rect 3266 22430 3278 22482
rect 3330 22430 3342 22482
rect 11554 22430 11566 22482
rect 11618 22430 11630 22482
rect 20862 22418 20914 22430
rect 21758 22482 21810 22494
rect 29486 22482 29538 22494
rect 23874 22430 23886 22482
rect 23938 22430 23950 22482
rect 27234 22430 27246 22482
rect 27298 22430 27310 22482
rect 21758 22418 21810 22430
rect 29486 22418 29538 22430
rect 30942 22482 30994 22494
rect 30942 22418 30994 22430
rect 31390 22482 31442 22494
rect 31390 22418 31442 22430
rect 2158 22370 2210 22382
rect 12798 22370 12850 22382
rect 4834 22318 4846 22370
rect 4898 22318 4910 22370
rect 5618 22318 5630 22370
rect 5682 22318 5694 22370
rect 6066 22318 6078 22370
rect 6130 22318 6142 22370
rect 11218 22318 11230 22370
rect 11282 22318 11294 22370
rect 12450 22318 12462 22370
rect 12514 22318 12526 22370
rect 2158 22306 2210 22318
rect 12798 22306 12850 22318
rect 15374 22370 15426 22382
rect 23102 22370 23154 22382
rect 29934 22370 29986 22382
rect 15922 22318 15934 22370
rect 15986 22318 15998 22370
rect 23986 22318 23998 22370
rect 24050 22318 24062 22370
rect 24658 22318 24670 22370
rect 24722 22318 24734 22370
rect 25442 22318 25454 22370
rect 25506 22318 25518 22370
rect 27346 22318 27358 22370
rect 27410 22318 27422 22370
rect 15374 22306 15426 22318
rect 23102 22306 23154 22318
rect 29934 22306 29986 22318
rect 30606 22370 30658 22382
rect 30606 22306 30658 22318
rect 2494 22258 2546 22270
rect 11566 22258 11618 22270
rect 4946 22206 4958 22258
rect 5010 22206 5022 22258
rect 2494 22194 2546 22206
rect 11566 22194 11618 22206
rect 12126 22258 12178 22270
rect 24894 22258 24946 22270
rect 30046 22258 30098 22270
rect 14130 22206 14142 22258
rect 14194 22206 14206 22258
rect 14690 22206 14702 22258
rect 14754 22206 14766 22258
rect 21970 22206 21982 22258
rect 22034 22206 22046 22258
rect 22530 22206 22542 22258
rect 22594 22206 22606 22258
rect 25778 22206 25790 22258
rect 25842 22206 25854 22258
rect 12126 22194 12178 22206
rect 24894 22194 24946 22206
rect 30046 22194 30098 22206
rect 1822 22146 1874 22158
rect 1822 22082 1874 22094
rect 2830 22146 2882 22158
rect 2830 22082 2882 22094
rect 3838 22146 3890 22158
rect 9214 22146 9266 22158
rect 8530 22094 8542 22146
rect 8594 22094 8606 22146
rect 3838 22082 3890 22094
rect 9214 22082 9266 22094
rect 9550 22146 9602 22158
rect 9550 22082 9602 22094
rect 9998 22146 10050 22158
rect 9998 22082 10050 22094
rect 11678 22146 11730 22158
rect 11678 22082 11730 22094
rect 11902 22146 11954 22158
rect 11902 22082 11954 22094
rect 12238 22146 12290 22158
rect 19070 22146 19122 22158
rect 18498 22094 18510 22146
rect 18562 22094 18574 22146
rect 12238 22082 12290 22094
rect 19070 22082 19122 22094
rect 19406 22146 19458 22158
rect 19406 22082 19458 22094
rect 20302 22146 20354 22158
rect 20302 22082 20354 22094
rect 21422 22146 21474 22158
rect 21422 22082 21474 22094
rect 23214 22146 23266 22158
rect 23214 22082 23266 22094
rect 23438 22146 23490 22158
rect 23438 22082 23490 22094
rect 29262 22146 29314 22158
rect 29262 22082 29314 22094
rect 30158 22146 30210 22158
rect 30158 22082 30210 22094
rect 1344 21978 38640 22012
rect 1344 21926 14024 21978
rect 14076 21926 14148 21978
rect 14200 21926 14272 21978
rect 14324 21926 14396 21978
rect 14448 21926 14520 21978
rect 14572 21926 14644 21978
rect 14696 21926 14768 21978
rect 14820 21926 14892 21978
rect 14944 21926 15016 21978
rect 15068 21926 15140 21978
rect 15192 21926 34024 21978
rect 34076 21926 34148 21978
rect 34200 21926 34272 21978
rect 34324 21926 34396 21978
rect 34448 21926 34520 21978
rect 34572 21926 34644 21978
rect 34696 21926 34768 21978
rect 34820 21926 34892 21978
rect 34944 21926 35016 21978
rect 35068 21926 35140 21978
rect 35192 21926 38640 21978
rect 1344 21892 38640 21926
rect 5854 21810 5906 21822
rect 4834 21758 4846 21810
rect 4898 21758 4910 21810
rect 5854 21746 5906 21758
rect 8430 21810 8482 21822
rect 8430 21746 8482 21758
rect 8878 21810 8930 21822
rect 8878 21746 8930 21758
rect 13694 21810 13746 21822
rect 15598 21810 15650 21822
rect 25342 21810 25394 21822
rect 13694 21746 13746 21758
rect 15150 21754 15202 21766
rect 8766 21698 8818 21710
rect 6962 21646 6974 21698
rect 7026 21646 7038 21698
rect 8766 21634 8818 21646
rect 12350 21698 12402 21710
rect 12350 21634 12402 21646
rect 15038 21698 15090 21710
rect 23986 21758 23998 21810
rect 24050 21758 24062 21810
rect 15598 21746 15650 21758
rect 25342 21746 25394 21758
rect 31838 21810 31890 21822
rect 31838 21746 31890 21758
rect 15150 21690 15202 21702
rect 26238 21698 26290 21710
rect 16706 21646 16718 21698
rect 16770 21646 16782 21698
rect 28914 21646 28926 21698
rect 28978 21646 28990 21698
rect 29698 21646 29710 21698
rect 29762 21646 29774 21698
rect 15038 21634 15090 21646
rect 26238 21634 26290 21646
rect 1710 21586 1762 21598
rect 6190 21586 6242 21598
rect 7534 21586 7586 21598
rect 2370 21534 2382 21586
rect 2434 21534 2446 21586
rect 6850 21534 6862 21586
rect 6914 21534 6926 21586
rect 1710 21522 1762 21534
rect 6190 21522 6242 21534
rect 7534 21522 7586 21534
rect 9662 21586 9714 21598
rect 15934 21586 15986 21598
rect 17502 21586 17554 21598
rect 10098 21534 10110 21586
rect 10162 21534 10174 21586
rect 16594 21534 16606 21586
rect 16658 21534 16670 21586
rect 9662 21522 9714 21534
rect 15934 21522 15986 21534
rect 17502 21522 17554 21534
rect 21310 21586 21362 21598
rect 27022 21586 27074 21598
rect 21746 21534 21758 21586
rect 21810 21534 21822 21586
rect 25218 21534 25230 21586
rect 25282 21534 25294 21586
rect 28578 21534 28590 21586
rect 28642 21534 28654 21586
rect 29810 21534 29822 21586
rect 29874 21534 29886 21586
rect 21310 21522 21362 21534
rect 27022 21522 27074 21534
rect 14142 21474 14194 21486
rect 14142 21410 14194 21422
rect 14590 21474 14642 21486
rect 14590 21410 14642 21422
rect 5406 21362 5458 21374
rect 5406 21298 5458 21310
rect 8878 21362 8930 21374
rect 8878 21298 8930 21310
rect 13134 21362 13186 21374
rect 13134 21298 13186 21310
rect 15038 21362 15090 21374
rect 15038 21298 15090 21310
rect 24782 21362 24834 21374
rect 24782 21298 24834 21310
rect 28254 21362 28306 21374
rect 28254 21298 28306 21310
rect 1344 21194 38640 21228
rect 1344 21142 4024 21194
rect 4076 21142 4148 21194
rect 4200 21142 4272 21194
rect 4324 21142 4396 21194
rect 4448 21142 4520 21194
rect 4572 21142 4644 21194
rect 4696 21142 4768 21194
rect 4820 21142 4892 21194
rect 4944 21142 5016 21194
rect 5068 21142 5140 21194
rect 5192 21142 24024 21194
rect 24076 21142 24148 21194
rect 24200 21142 24272 21194
rect 24324 21142 24396 21194
rect 24448 21142 24520 21194
rect 24572 21142 24644 21194
rect 24696 21142 24768 21194
rect 24820 21142 24892 21194
rect 24944 21142 25016 21194
rect 25068 21142 25140 21194
rect 25192 21142 38640 21194
rect 1344 21108 38640 21142
rect 4510 21026 4562 21038
rect 4510 20962 4562 20974
rect 20414 21026 20466 21038
rect 20414 20962 20466 20974
rect 21870 21026 21922 21038
rect 21870 20962 21922 20974
rect 22206 21026 22258 21038
rect 22206 20962 22258 20974
rect 33518 21026 33570 21038
rect 33518 20962 33570 20974
rect 1934 20914 1986 20926
rect 1934 20850 1986 20862
rect 6750 20914 6802 20926
rect 12238 20914 12290 20926
rect 10546 20862 10558 20914
rect 10610 20862 10622 20914
rect 6750 20850 6802 20862
rect 12238 20850 12290 20862
rect 12910 20914 12962 20926
rect 12910 20850 12962 20862
rect 15150 20914 15202 20926
rect 15150 20850 15202 20862
rect 15598 20914 15650 20926
rect 25442 20862 25454 20914
rect 25506 20862 25518 20914
rect 27458 20862 27470 20914
rect 27522 20862 27534 20914
rect 15598 20850 15650 20862
rect 4622 20802 4674 20814
rect 4622 20738 4674 20750
rect 6078 20802 6130 20814
rect 6078 20738 6130 20750
rect 8430 20802 8482 20814
rect 12126 20802 12178 20814
rect 21422 20802 21474 20814
rect 9090 20750 9102 20802
rect 9154 20750 9166 20802
rect 10322 20750 10334 20802
rect 10386 20750 10398 20802
rect 11778 20750 11790 20802
rect 11842 20750 11854 20802
rect 20738 20750 20750 20802
rect 20802 20750 20814 20802
rect 8430 20738 8482 20750
rect 12126 20738 12178 20750
rect 21422 20738 21474 20750
rect 23998 20802 24050 20814
rect 23998 20738 24050 20750
rect 24558 20802 24610 20814
rect 24558 20738 24610 20750
rect 24670 20802 24722 20814
rect 27806 20802 27858 20814
rect 29150 20802 29202 20814
rect 25218 20750 25230 20802
rect 25282 20750 25294 20802
rect 28242 20750 28254 20802
rect 28306 20750 28318 20802
rect 24670 20738 24722 20750
rect 27806 20738 27858 20750
rect 29150 20738 29202 20750
rect 29486 20802 29538 20814
rect 29486 20738 29538 20750
rect 30046 20802 30098 20814
rect 30370 20750 30382 20802
rect 30434 20750 30446 20802
rect 30046 20738 30098 20750
rect 2830 20690 2882 20702
rect 2830 20626 2882 20638
rect 3166 20690 3218 20702
rect 3166 20626 3218 20638
rect 6190 20690 6242 20702
rect 6190 20626 6242 20638
rect 9326 20690 9378 20702
rect 9326 20626 9378 20638
rect 10894 20690 10946 20702
rect 29262 20690 29314 20702
rect 22418 20638 22430 20690
rect 22482 20638 22494 20690
rect 22978 20638 22990 20690
rect 23042 20638 23054 20690
rect 10894 20626 10946 20638
rect 29262 20626 29314 20638
rect 32734 20690 32786 20702
rect 32734 20626 32786 20638
rect 2494 20578 2546 20590
rect 2494 20514 2546 20526
rect 5070 20578 5122 20590
rect 5070 20514 5122 20526
rect 5742 20578 5794 20590
rect 5742 20514 5794 20526
rect 6414 20578 6466 20590
rect 6414 20514 6466 20526
rect 8766 20578 8818 20590
rect 8766 20514 8818 20526
rect 9550 20578 9602 20590
rect 9550 20514 9602 20526
rect 9662 20578 9714 20590
rect 9662 20514 9714 20526
rect 13694 20578 13746 20590
rect 13694 20514 13746 20526
rect 14142 20578 14194 20590
rect 14142 20514 14194 20526
rect 20526 20578 20578 20590
rect 20526 20514 20578 20526
rect 23662 20578 23714 20590
rect 23662 20514 23714 20526
rect 23886 20578 23938 20590
rect 23886 20514 23938 20526
rect 1344 20410 38640 20444
rect 1344 20358 14024 20410
rect 14076 20358 14148 20410
rect 14200 20358 14272 20410
rect 14324 20358 14396 20410
rect 14448 20358 14520 20410
rect 14572 20358 14644 20410
rect 14696 20358 14768 20410
rect 14820 20358 14892 20410
rect 14944 20358 15016 20410
rect 15068 20358 15140 20410
rect 15192 20358 34024 20410
rect 34076 20358 34148 20410
rect 34200 20358 34272 20410
rect 34324 20358 34396 20410
rect 34448 20358 34520 20410
rect 34572 20358 34644 20410
rect 34696 20358 34768 20410
rect 34820 20358 34892 20410
rect 34944 20358 35016 20410
rect 35068 20358 35140 20410
rect 35192 20358 38640 20410
rect 1344 20324 38640 20358
rect 6190 20242 6242 20254
rect 6190 20178 6242 20190
rect 10670 20242 10722 20254
rect 10670 20178 10722 20190
rect 11566 20242 11618 20254
rect 11566 20178 11618 20190
rect 11678 20242 11730 20254
rect 11678 20178 11730 20190
rect 1934 20130 1986 20142
rect 1934 20066 1986 20078
rect 10334 20130 10386 20142
rect 10334 20066 10386 20078
rect 10446 20130 10498 20142
rect 10446 20066 10498 20078
rect 12126 20130 12178 20142
rect 12126 20066 12178 20078
rect 12350 20130 12402 20142
rect 12350 20066 12402 20078
rect 12574 20130 12626 20142
rect 12574 20066 12626 20078
rect 13918 20130 13970 20142
rect 13918 20066 13970 20078
rect 14142 20130 14194 20142
rect 14142 20066 14194 20078
rect 18286 20130 18338 20142
rect 18286 20066 18338 20078
rect 18622 20130 18674 20142
rect 18622 20066 18674 20078
rect 18734 20130 18786 20142
rect 31950 20130 32002 20142
rect 25778 20078 25790 20130
rect 25842 20078 25854 20130
rect 26786 20078 26798 20130
rect 26850 20078 26862 20130
rect 18734 20066 18786 20078
rect 31950 20066 32002 20078
rect 12686 20018 12738 20030
rect 9874 19966 9886 20018
rect 9938 19966 9950 20018
rect 11890 19966 11902 20018
rect 11954 19966 11966 20018
rect 12686 19954 12738 19966
rect 14366 20018 14418 20030
rect 14366 19954 14418 19966
rect 14814 20018 14866 20030
rect 14814 19954 14866 19966
rect 18958 20018 19010 20030
rect 29710 20018 29762 20030
rect 23650 19966 23662 20018
rect 23714 19966 23726 20018
rect 24770 19966 24782 20018
rect 24834 19966 24846 20018
rect 25330 19966 25342 20018
rect 25394 19966 25406 20018
rect 28466 19966 28478 20018
rect 28530 19966 28542 20018
rect 29138 19966 29150 20018
rect 29202 19966 29214 20018
rect 18958 19954 19010 19966
rect 29710 19954 29762 19966
rect 30158 20018 30210 20030
rect 30158 19954 30210 19966
rect 30270 20018 30322 20030
rect 30270 19954 30322 19966
rect 30718 20018 30770 20030
rect 30718 19954 30770 19966
rect 2494 19906 2546 19918
rect 2494 19842 2546 19854
rect 5742 19906 5794 19918
rect 14254 19906 14306 19918
rect 10322 19854 10334 19906
rect 10386 19854 10398 19906
rect 5742 19842 5794 19854
rect 14254 19842 14306 19854
rect 23550 19906 23602 19918
rect 29822 19906 29874 19918
rect 27010 19854 27022 19906
rect 27074 19854 27086 19906
rect 23550 19842 23602 19854
rect 29822 19842 29874 19854
rect 30942 19906 30994 19918
rect 30942 19842 30994 19854
rect 31502 19906 31554 19918
rect 31502 19842 31554 19854
rect 24222 19794 24274 19806
rect 24222 19730 24274 19742
rect 30270 19794 30322 19806
rect 30270 19730 30322 19742
rect 1344 19626 38640 19660
rect 1344 19574 4024 19626
rect 4076 19574 4148 19626
rect 4200 19574 4272 19626
rect 4324 19574 4396 19626
rect 4448 19574 4520 19626
rect 4572 19574 4644 19626
rect 4696 19574 4768 19626
rect 4820 19574 4892 19626
rect 4944 19574 5016 19626
rect 5068 19574 5140 19626
rect 5192 19574 24024 19626
rect 24076 19574 24148 19626
rect 24200 19574 24272 19626
rect 24324 19574 24396 19626
rect 24448 19574 24520 19626
rect 24572 19574 24644 19626
rect 24696 19574 24768 19626
rect 24820 19574 24892 19626
rect 24944 19574 25016 19626
rect 25068 19574 25140 19626
rect 25192 19574 38640 19626
rect 1344 19540 38640 19574
rect 26910 19458 26962 19470
rect 2034 19406 2046 19458
rect 2098 19455 2110 19458
rect 2594 19455 2606 19458
rect 2098 19409 2606 19455
rect 2098 19406 2110 19409
rect 2594 19406 2606 19409
rect 2658 19406 2670 19458
rect 23874 19406 23886 19458
rect 23938 19455 23950 19458
rect 24658 19455 24670 19458
rect 23938 19409 24670 19455
rect 23938 19406 23950 19409
rect 24658 19406 24670 19409
rect 24722 19406 24734 19458
rect 26114 19406 26126 19458
rect 26178 19406 26190 19458
rect 26910 19394 26962 19406
rect 2046 19346 2098 19358
rect 24670 19346 24722 19358
rect 14578 19294 14590 19346
rect 14642 19294 14654 19346
rect 2046 19282 2098 19294
rect 24670 19282 24722 19294
rect 28030 19346 28082 19358
rect 28030 19282 28082 19294
rect 18846 19234 18898 19246
rect 2930 19182 2942 19234
rect 2994 19182 3006 19234
rect 3602 19182 3614 19234
rect 3666 19182 3678 19234
rect 14690 19182 14702 19234
rect 14754 19182 14766 19234
rect 15026 19182 15038 19234
rect 15090 19182 15102 19234
rect 18846 19170 18898 19182
rect 18958 19234 19010 19246
rect 18958 19170 19010 19182
rect 20526 19234 20578 19246
rect 27134 19234 27186 19246
rect 27918 19234 27970 19246
rect 29150 19234 29202 19246
rect 32734 19234 32786 19246
rect 25106 19182 25118 19234
rect 25170 19182 25182 19234
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 26338 19182 26350 19234
rect 26402 19182 26414 19234
rect 27346 19182 27358 19234
rect 27410 19182 27422 19234
rect 27682 19182 27694 19234
rect 27746 19182 27758 19234
rect 28354 19182 28366 19234
rect 28418 19182 28430 19234
rect 32274 19182 32286 19234
rect 32338 19182 32350 19234
rect 20526 19170 20578 19182
rect 27134 19170 27186 19182
rect 27918 19170 27970 19182
rect 29150 19170 29202 19182
rect 32734 19170 32786 19182
rect 19182 19122 19234 19134
rect 19742 19122 19794 19134
rect 19506 19070 19518 19122
rect 19570 19070 19582 19122
rect 19182 19058 19234 19070
rect 19742 19058 19794 19070
rect 20190 19122 20242 19134
rect 20190 19058 20242 19070
rect 20302 19122 20354 19134
rect 26798 19122 26850 19134
rect 26450 19070 26462 19122
rect 26514 19070 26526 19122
rect 20302 19058 20354 19070
rect 26798 19058 26850 19070
rect 2494 19010 2546 19022
rect 2494 18946 2546 18958
rect 3166 19010 3218 19022
rect 3166 18946 3218 18958
rect 3838 19010 3890 19022
rect 3838 18946 3890 18958
rect 14254 19010 14306 19022
rect 14254 18946 14306 18958
rect 14478 19010 14530 19022
rect 14478 18946 14530 18958
rect 17166 19010 17218 19022
rect 17166 18946 17218 18958
rect 19630 19010 19682 19022
rect 19630 18946 19682 18958
rect 24222 19010 24274 19022
rect 24222 18946 24274 18958
rect 28142 19010 28194 19022
rect 29810 18958 29822 19010
rect 29874 18958 29886 19010
rect 28142 18946 28194 18958
rect 1344 18842 38640 18876
rect 1344 18790 14024 18842
rect 14076 18790 14148 18842
rect 14200 18790 14272 18842
rect 14324 18790 14396 18842
rect 14448 18790 14520 18842
rect 14572 18790 14644 18842
rect 14696 18790 14768 18842
rect 14820 18790 14892 18842
rect 14944 18790 15016 18842
rect 15068 18790 15140 18842
rect 15192 18790 34024 18842
rect 34076 18790 34148 18842
rect 34200 18790 34272 18842
rect 34324 18790 34396 18842
rect 34448 18790 34520 18842
rect 34572 18790 34644 18842
rect 34696 18790 34768 18842
rect 34820 18790 34892 18842
rect 34944 18790 35016 18842
rect 35068 18790 35140 18842
rect 35192 18790 38640 18842
rect 1344 18756 38640 18790
rect 15374 18674 15426 18686
rect 27358 18674 27410 18686
rect 16594 18622 16606 18674
rect 16658 18622 16670 18674
rect 20514 18622 20526 18674
rect 20578 18622 20590 18674
rect 15374 18610 15426 18622
rect 27358 18610 27410 18622
rect 27918 18674 27970 18686
rect 29586 18622 29598 18674
rect 29650 18622 29662 18674
rect 27918 18610 27970 18622
rect 3166 18562 3218 18574
rect 3166 18498 3218 18510
rect 12014 18562 12066 18574
rect 12014 18498 12066 18510
rect 12238 18562 12290 18574
rect 26798 18562 26850 18574
rect 13122 18510 13134 18562
rect 13186 18510 13198 18562
rect 13794 18510 13806 18562
rect 13858 18510 13870 18562
rect 15698 18510 15710 18562
rect 15762 18510 15774 18562
rect 21522 18510 21534 18562
rect 21586 18510 21598 18562
rect 29026 18510 29038 18562
rect 29090 18510 29102 18562
rect 12238 18498 12290 18510
rect 26798 18498 26850 18510
rect 2606 18450 2658 18462
rect 2606 18386 2658 18398
rect 2830 18450 2882 18462
rect 17390 18450 17442 18462
rect 21198 18450 21250 18462
rect 23214 18450 23266 18462
rect 30718 18450 30770 18462
rect 13234 18398 13246 18450
rect 13298 18398 13310 18450
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 14802 18398 14814 18450
rect 14866 18398 14878 18450
rect 15586 18398 15598 18450
rect 15650 18398 15662 18450
rect 16706 18398 16718 18450
rect 16770 18398 16782 18450
rect 18050 18398 18062 18450
rect 18114 18398 18126 18450
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 21858 18398 21870 18450
rect 21922 18398 21934 18450
rect 22530 18398 22542 18450
rect 22594 18398 22606 18450
rect 28578 18398 28590 18450
rect 28642 18398 28654 18450
rect 29698 18398 29710 18450
rect 29762 18398 29774 18450
rect 2830 18386 2882 18398
rect 17390 18386 17442 18398
rect 21198 18386 21250 18398
rect 23214 18386 23266 18398
rect 30718 18386 30770 18398
rect 28254 18338 28306 18350
rect 28254 18274 28306 18286
rect 30158 18338 30210 18350
rect 30158 18274 30210 18286
rect 11902 18226 11954 18238
rect 11902 18162 11954 18174
rect 21086 18226 21138 18238
rect 21086 18162 21138 18174
rect 23102 18226 23154 18238
rect 23102 18162 23154 18174
rect 1344 18058 38640 18092
rect 1344 18006 4024 18058
rect 4076 18006 4148 18058
rect 4200 18006 4272 18058
rect 4324 18006 4396 18058
rect 4448 18006 4520 18058
rect 4572 18006 4644 18058
rect 4696 18006 4768 18058
rect 4820 18006 4892 18058
rect 4944 18006 5016 18058
rect 5068 18006 5140 18058
rect 5192 18006 24024 18058
rect 24076 18006 24148 18058
rect 24200 18006 24272 18058
rect 24324 18006 24396 18058
rect 24448 18006 24520 18058
rect 24572 18006 24644 18058
rect 24696 18006 24768 18058
rect 24820 18006 24892 18058
rect 24944 18006 25016 18058
rect 25068 18006 25140 18058
rect 25192 18006 38640 18058
rect 1344 17972 38640 18006
rect 4174 17890 4226 17902
rect 4174 17826 4226 17838
rect 10446 17890 10498 17902
rect 10446 17826 10498 17838
rect 13582 17890 13634 17902
rect 13582 17826 13634 17838
rect 9550 17778 9602 17790
rect 9550 17714 9602 17726
rect 17950 17778 18002 17790
rect 17950 17714 18002 17726
rect 19742 17778 19794 17790
rect 19742 17714 19794 17726
rect 29262 17778 29314 17790
rect 29262 17714 29314 17726
rect 9998 17666 10050 17678
rect 4610 17614 4622 17666
rect 4674 17614 4686 17666
rect 5618 17614 5630 17666
rect 5682 17614 5694 17666
rect 6066 17614 6078 17666
rect 6130 17614 6142 17666
rect 9998 17602 10050 17614
rect 11118 17666 11170 17678
rect 17054 17666 17106 17678
rect 11890 17614 11902 17666
rect 11954 17614 11966 17666
rect 16594 17614 16606 17666
rect 16658 17614 16670 17666
rect 11118 17602 11170 17614
rect 17054 17602 17106 17614
rect 19294 17666 19346 17678
rect 19294 17602 19346 17614
rect 19406 17666 19458 17678
rect 20638 17666 20690 17678
rect 20402 17614 20414 17666
rect 20466 17614 20478 17666
rect 19406 17602 19458 17614
rect 20638 17602 20690 17614
rect 21646 17666 21698 17678
rect 21646 17602 21698 17614
rect 22094 17666 22146 17678
rect 22094 17602 22146 17614
rect 22318 17666 22370 17678
rect 22318 17602 22370 17614
rect 22654 17666 22706 17678
rect 23314 17614 23326 17666
rect 23378 17614 23390 17666
rect 23538 17614 23550 17666
rect 23602 17614 23614 17666
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 22654 17602 22706 17614
rect 9214 17554 9266 17566
rect 22766 17554 22818 17566
rect 4946 17502 4958 17554
rect 5010 17502 5022 17554
rect 12002 17502 12014 17554
rect 12066 17502 12078 17554
rect 12562 17502 12574 17554
rect 12626 17502 12638 17554
rect 18162 17502 18174 17554
rect 18226 17502 18238 17554
rect 18610 17502 18622 17554
rect 18674 17502 18686 17554
rect 9214 17490 9266 17502
rect 22766 17490 22818 17502
rect 2606 17442 2658 17454
rect 2606 17378 2658 17390
rect 2830 17442 2882 17454
rect 3838 17442 3890 17454
rect 10558 17442 10610 17454
rect 3154 17390 3166 17442
rect 3218 17390 3230 17442
rect 8530 17390 8542 17442
rect 8594 17390 8606 17442
rect 2830 17378 2882 17390
rect 3838 17378 3890 17390
rect 10558 17378 10610 17390
rect 10782 17442 10834 17454
rect 10782 17378 10834 17390
rect 11454 17442 11506 17454
rect 17614 17442 17666 17454
rect 12338 17390 12350 17442
rect 12402 17390 12414 17442
rect 14354 17390 14366 17442
rect 14418 17390 14430 17442
rect 11454 17378 11506 17390
rect 17614 17378 17666 17390
rect 21422 17442 21474 17454
rect 21422 17378 21474 17390
rect 22206 17442 22258 17454
rect 22206 17378 22258 17390
rect 22990 17442 23042 17454
rect 24894 17442 24946 17454
rect 23650 17390 23662 17442
rect 23714 17390 23726 17442
rect 22990 17378 23042 17390
rect 24894 17378 24946 17390
rect 28254 17442 28306 17454
rect 28254 17378 28306 17390
rect 1344 17274 38640 17308
rect 1344 17222 14024 17274
rect 14076 17222 14148 17274
rect 14200 17222 14272 17274
rect 14324 17222 14396 17274
rect 14448 17222 14520 17274
rect 14572 17222 14644 17274
rect 14696 17222 14768 17274
rect 14820 17222 14892 17274
rect 14944 17222 15016 17274
rect 15068 17222 15140 17274
rect 15192 17222 34024 17274
rect 34076 17222 34148 17274
rect 34200 17222 34272 17274
rect 34324 17222 34396 17274
rect 34448 17222 34520 17274
rect 34572 17222 34644 17274
rect 34696 17222 34768 17274
rect 34820 17222 34892 17274
rect 34944 17222 35016 17274
rect 35068 17222 35140 17274
rect 35192 17222 38640 17274
rect 1344 17188 38640 17222
rect 2494 17106 2546 17118
rect 2494 17042 2546 17054
rect 7422 17106 7474 17118
rect 7422 17042 7474 17054
rect 8654 17106 8706 17118
rect 8654 17042 8706 17054
rect 10110 17106 10162 17118
rect 10110 17042 10162 17054
rect 18510 17106 18562 17118
rect 18510 17042 18562 17054
rect 20862 17106 20914 17118
rect 20862 17042 20914 17054
rect 22430 17106 22482 17118
rect 22430 17042 22482 17054
rect 23886 17106 23938 17118
rect 23886 17042 23938 17054
rect 24110 17106 24162 17118
rect 24110 17042 24162 17054
rect 25566 17106 25618 17118
rect 25566 17042 25618 17054
rect 26238 17106 26290 17118
rect 26238 17042 26290 17054
rect 26798 17106 26850 17118
rect 26798 17042 26850 17054
rect 1934 16994 1986 17006
rect 1934 16930 1986 16942
rect 3166 16994 3218 17006
rect 8430 16994 8482 17006
rect 4722 16942 4734 16994
rect 4786 16942 4798 16994
rect 3166 16930 3218 16942
rect 8430 16930 8482 16942
rect 9662 16994 9714 17006
rect 10894 16994 10946 17006
rect 10434 16942 10446 16994
rect 10498 16942 10510 16994
rect 9662 16930 9714 16942
rect 10894 16930 10946 16942
rect 11006 16994 11058 17006
rect 11006 16930 11058 16942
rect 11118 16994 11170 17006
rect 16494 16994 16546 17006
rect 13346 16942 13358 16994
rect 13410 16942 13422 16994
rect 15474 16942 15486 16994
rect 15538 16942 15550 16994
rect 11118 16930 11170 16942
rect 16494 16930 16546 16942
rect 16606 16994 16658 17006
rect 16606 16930 16658 16942
rect 19742 16994 19794 17006
rect 22654 16994 22706 17006
rect 20066 16942 20078 16994
rect 20130 16942 20142 16994
rect 19742 16930 19794 16942
rect 22654 16930 22706 16942
rect 23214 16994 23266 17006
rect 23214 16930 23266 16942
rect 23662 16994 23714 17006
rect 23662 16930 23714 16942
rect 25230 16994 25282 17006
rect 25230 16930 25282 16942
rect 26126 16994 26178 17006
rect 26126 16930 26178 16942
rect 2158 16882 2210 16894
rect 5294 16882 5346 16894
rect 2930 16830 2942 16882
rect 2994 16830 3006 16882
rect 4610 16830 4622 16882
rect 4674 16830 4686 16882
rect 2158 16818 2210 16830
rect 5294 16818 5346 16830
rect 5742 16882 5794 16894
rect 5742 16818 5794 16830
rect 6974 16882 7026 16894
rect 8206 16882 8258 16894
rect 7186 16830 7198 16882
rect 7250 16830 7262 16882
rect 6974 16818 7026 16830
rect 8206 16818 8258 16830
rect 8878 16882 8930 16894
rect 8878 16818 8930 16830
rect 9550 16882 9602 16894
rect 14926 16882 14978 16894
rect 17614 16882 17666 16894
rect 12114 16830 12126 16882
rect 12178 16830 12190 16882
rect 15698 16830 15710 16882
rect 15762 16830 15774 16882
rect 9550 16818 9602 16830
rect 14926 16818 14978 16830
rect 17614 16818 17666 16830
rect 20190 16882 20242 16894
rect 21422 16882 21474 16894
rect 20402 16830 20414 16882
rect 20466 16830 20478 16882
rect 21074 16830 21086 16882
rect 21138 16830 21150 16882
rect 20190 16818 20242 16830
rect 21422 16818 21474 16830
rect 22094 16882 22146 16894
rect 22094 16818 22146 16830
rect 23326 16882 23378 16894
rect 23326 16818 23378 16830
rect 24222 16882 24274 16894
rect 24222 16818 24274 16830
rect 25454 16882 25506 16894
rect 25454 16818 25506 16830
rect 25902 16882 25954 16894
rect 25902 16818 25954 16830
rect 3614 16770 3666 16782
rect 3614 16706 3666 16718
rect 3950 16770 4002 16782
rect 18062 16770 18114 16782
rect 6850 16718 6862 16770
rect 6914 16718 6926 16770
rect 3950 16706 4002 16718
rect 18062 16706 18114 16718
rect 19406 16770 19458 16782
rect 19406 16706 19458 16718
rect 22318 16770 22370 16782
rect 22318 16706 22370 16718
rect 7758 16658 7810 16670
rect 1698 16606 1710 16658
rect 1762 16655 1774 16658
rect 1922 16655 1934 16658
rect 1762 16609 1934 16655
rect 1762 16606 1774 16609
rect 1922 16606 1934 16609
rect 1986 16606 1998 16658
rect 7758 16594 7810 16606
rect 7870 16658 7922 16670
rect 7870 16594 7922 16606
rect 8318 16658 8370 16670
rect 8318 16594 8370 16606
rect 14590 16658 14642 16670
rect 14590 16594 14642 16606
rect 16606 16658 16658 16670
rect 16606 16594 16658 16606
rect 19518 16658 19570 16670
rect 19518 16594 19570 16606
rect 20750 16658 20802 16670
rect 20750 16594 20802 16606
rect 23774 16658 23826 16670
rect 23774 16594 23826 16606
rect 26238 16658 26290 16670
rect 26238 16594 26290 16606
rect 1344 16490 38640 16524
rect 1344 16438 4024 16490
rect 4076 16438 4148 16490
rect 4200 16438 4272 16490
rect 4324 16438 4396 16490
rect 4448 16438 4520 16490
rect 4572 16438 4644 16490
rect 4696 16438 4768 16490
rect 4820 16438 4892 16490
rect 4944 16438 5016 16490
rect 5068 16438 5140 16490
rect 5192 16438 24024 16490
rect 24076 16438 24148 16490
rect 24200 16438 24272 16490
rect 24324 16438 24396 16490
rect 24448 16438 24520 16490
rect 24572 16438 24644 16490
rect 24696 16438 24768 16490
rect 24820 16438 24892 16490
rect 24944 16438 25016 16490
rect 25068 16438 25140 16490
rect 25192 16438 38640 16490
rect 1344 16404 38640 16438
rect 3390 16322 3442 16334
rect 3390 16258 3442 16270
rect 6078 16322 6130 16334
rect 6078 16258 6130 16270
rect 13694 16322 13746 16334
rect 13694 16258 13746 16270
rect 21646 16322 21698 16334
rect 21646 16258 21698 16270
rect 26798 16322 26850 16334
rect 26798 16258 26850 16270
rect 30382 16322 30434 16334
rect 30382 16258 30434 16270
rect 4734 16210 4786 16222
rect 7758 16210 7810 16222
rect 11230 16210 11282 16222
rect 7410 16158 7422 16210
rect 7474 16158 7486 16210
rect 9426 16158 9438 16210
rect 9490 16158 9502 16210
rect 4734 16146 4786 16158
rect 7758 16146 7810 16158
rect 11230 16146 11282 16158
rect 13582 16210 13634 16222
rect 13582 16146 13634 16158
rect 14030 16210 14082 16222
rect 14030 16146 14082 16158
rect 14702 16210 14754 16222
rect 14702 16146 14754 16158
rect 15038 16210 15090 16222
rect 15038 16146 15090 16158
rect 23774 16210 23826 16222
rect 23774 16146 23826 16158
rect 29374 16210 29426 16222
rect 29374 16146 29426 16158
rect 6302 16098 6354 16110
rect 17614 16098 17666 16110
rect 3938 16046 3950 16098
rect 4002 16046 4014 16098
rect 5842 16046 5854 16098
rect 5906 16046 5918 16098
rect 7074 16046 7086 16098
rect 7138 16046 7150 16098
rect 8642 16046 8654 16098
rect 8706 16046 8718 16098
rect 12338 16046 12350 16098
rect 12402 16046 12414 16098
rect 12674 16046 12686 16098
rect 12738 16046 12750 16098
rect 6302 16034 6354 16046
rect 17614 16034 17666 16046
rect 24334 16098 24386 16110
rect 24334 16034 24386 16046
rect 24558 16098 24610 16110
rect 29934 16098 29986 16110
rect 24770 16046 24782 16098
rect 24834 16046 24846 16098
rect 25778 16046 25790 16098
rect 25842 16046 25854 16098
rect 30258 16046 30270 16098
rect 30322 16046 30334 16098
rect 24558 16034 24610 16046
rect 29934 16034 29986 16046
rect 12910 15986 12962 15998
rect 4162 15934 4174 15986
rect 4226 15934 4238 15986
rect 12910 15922 12962 15934
rect 21758 15986 21810 15998
rect 21758 15922 21810 15934
rect 25118 15986 25170 15998
rect 25118 15922 25170 15934
rect 1822 15874 1874 15886
rect 1822 15810 1874 15822
rect 3054 15874 3106 15886
rect 3054 15810 3106 15822
rect 5966 15874 6018 15886
rect 5966 15810 6018 15822
rect 14142 15874 14194 15886
rect 14142 15810 14194 15822
rect 17166 15874 17218 15886
rect 17166 15810 17218 15822
rect 22206 15874 22258 15886
rect 22206 15810 22258 15822
rect 22654 15874 22706 15886
rect 22654 15810 22706 15822
rect 24222 15874 24274 15886
rect 24222 15810 24274 15822
rect 24446 15874 24498 15886
rect 24446 15810 24498 15822
rect 25230 15874 25282 15886
rect 25230 15810 25282 15822
rect 25342 15874 25394 15886
rect 25342 15810 25394 15822
rect 1344 15706 38640 15740
rect 1344 15654 14024 15706
rect 14076 15654 14148 15706
rect 14200 15654 14272 15706
rect 14324 15654 14396 15706
rect 14448 15654 14520 15706
rect 14572 15654 14644 15706
rect 14696 15654 14768 15706
rect 14820 15654 14892 15706
rect 14944 15654 15016 15706
rect 15068 15654 15140 15706
rect 15192 15654 34024 15706
rect 34076 15654 34148 15706
rect 34200 15654 34272 15706
rect 34324 15654 34396 15706
rect 34448 15654 34520 15706
rect 34572 15654 34644 15706
rect 34696 15654 34768 15706
rect 34820 15654 34892 15706
rect 34944 15654 35016 15706
rect 35068 15654 35140 15706
rect 35192 15654 38640 15706
rect 1344 15620 38640 15654
rect 5294 15538 5346 15550
rect 4722 15486 4734 15538
rect 4786 15486 4798 15538
rect 5294 15474 5346 15486
rect 5854 15538 5906 15550
rect 5854 15474 5906 15486
rect 6414 15538 6466 15550
rect 6414 15474 6466 15486
rect 8430 15538 8482 15550
rect 8430 15474 8482 15486
rect 8654 15538 8706 15550
rect 8654 15474 8706 15486
rect 9662 15538 9714 15550
rect 9662 15474 9714 15486
rect 9774 15538 9826 15550
rect 9774 15474 9826 15486
rect 10558 15538 10610 15550
rect 10558 15474 10610 15486
rect 12910 15538 12962 15550
rect 29038 15538 29090 15550
rect 13346 15486 13358 15538
rect 13410 15486 13422 15538
rect 21634 15486 21646 15538
rect 21698 15486 21710 15538
rect 28466 15486 28478 15538
rect 28530 15486 28542 15538
rect 12910 15474 12962 15486
rect 29038 15474 29090 15486
rect 29598 15538 29650 15550
rect 29598 15474 29650 15486
rect 5742 15426 5794 15438
rect 5742 15362 5794 15374
rect 6078 15426 6130 15438
rect 6078 15362 6130 15374
rect 7198 15426 7250 15438
rect 9550 15426 9602 15438
rect 7522 15374 7534 15426
rect 7586 15374 7598 15426
rect 7198 15362 7250 15374
rect 9550 15362 9602 15374
rect 13918 15426 13970 15438
rect 30046 15426 30098 15438
rect 23202 15374 23214 15426
rect 23266 15374 23278 15426
rect 23538 15374 23550 15426
rect 23602 15374 23614 15426
rect 13918 15362 13970 15374
rect 30046 15362 30098 15374
rect 1822 15314 1874 15326
rect 6862 15314 6914 15326
rect 2258 15262 2270 15314
rect 2322 15262 2334 15314
rect 1822 15250 1874 15262
rect 6862 15250 6914 15262
rect 7758 15314 7810 15326
rect 7758 15250 7810 15262
rect 8206 15314 8258 15326
rect 8206 15250 8258 15262
rect 8878 15314 8930 15326
rect 8878 15250 8930 15262
rect 10222 15314 10274 15326
rect 10222 15250 10274 15262
rect 11566 15314 11618 15326
rect 11566 15250 11618 15262
rect 12238 15314 12290 15326
rect 12238 15250 12290 15262
rect 12798 15314 12850 15326
rect 12798 15250 12850 15262
rect 13134 15314 13186 15326
rect 13134 15250 13186 15262
rect 13358 15314 13410 15326
rect 13358 15250 13410 15262
rect 18734 15314 18786 15326
rect 22990 15314 23042 15326
rect 19170 15262 19182 15314
rect 19234 15262 19246 15314
rect 18734 15250 18786 15262
rect 22990 15250 23042 15262
rect 25566 15314 25618 15326
rect 25890 15262 25902 15314
rect 25954 15262 25966 15314
rect 25566 15250 25618 15262
rect 11006 15202 11058 15214
rect 14366 15202 14418 15214
rect 7858 15150 7870 15202
rect 7922 15150 7934 15202
rect 12002 15150 12014 15202
rect 12066 15150 12078 15202
rect 11006 15138 11058 15150
rect 14366 15138 14418 15150
rect 22206 15202 22258 15214
rect 22206 15138 22258 15150
rect 6974 15090 7026 15102
rect 6974 15026 7026 15038
rect 8766 15090 8818 15102
rect 8766 15026 8818 15038
rect 11790 15090 11842 15102
rect 11790 15026 11842 15038
rect 12350 15090 12402 15102
rect 12350 15026 12402 15038
rect 22654 15090 22706 15102
rect 22654 15026 22706 15038
rect 1344 14922 38640 14956
rect 1344 14870 4024 14922
rect 4076 14870 4148 14922
rect 4200 14870 4272 14922
rect 4324 14870 4396 14922
rect 4448 14870 4520 14922
rect 4572 14870 4644 14922
rect 4696 14870 4768 14922
rect 4820 14870 4892 14922
rect 4944 14870 5016 14922
rect 5068 14870 5140 14922
rect 5192 14870 24024 14922
rect 24076 14870 24148 14922
rect 24200 14870 24272 14922
rect 24324 14870 24396 14922
rect 24448 14870 24520 14922
rect 24572 14870 24644 14922
rect 24696 14870 24768 14922
rect 24820 14870 24892 14922
rect 24944 14870 25016 14922
rect 25068 14870 25140 14922
rect 25192 14870 38640 14922
rect 1344 14836 38640 14870
rect 4062 14754 4114 14766
rect 23886 14754 23938 14766
rect 21634 14702 21646 14754
rect 21698 14751 21710 14754
rect 22418 14751 22430 14754
rect 21698 14705 22430 14751
rect 21698 14702 21710 14705
rect 22418 14702 22430 14705
rect 22482 14702 22494 14754
rect 4062 14690 4114 14702
rect 23886 14690 23938 14702
rect 5742 14642 5794 14654
rect 7758 14642 7810 14654
rect 12798 14642 12850 14654
rect 6962 14590 6974 14642
rect 7026 14590 7038 14642
rect 11442 14590 11454 14642
rect 11506 14590 11518 14642
rect 5742 14578 5794 14590
rect 7758 14578 7810 14590
rect 12798 14578 12850 14590
rect 13582 14642 13634 14654
rect 13582 14578 13634 14590
rect 17614 14642 17666 14654
rect 17614 14578 17666 14590
rect 18062 14642 18114 14654
rect 18062 14578 18114 14590
rect 18622 14642 18674 14654
rect 18622 14578 18674 14590
rect 19854 14642 19906 14654
rect 19854 14578 19906 14590
rect 21982 14642 22034 14654
rect 21982 14578 22034 14590
rect 8430 14530 8482 14542
rect 4834 14478 4846 14530
rect 4898 14478 4910 14530
rect 7074 14478 7086 14530
rect 7138 14478 7150 14530
rect 8430 14466 8482 14478
rect 9214 14530 9266 14542
rect 9214 14466 9266 14478
rect 9774 14530 9826 14542
rect 9774 14466 9826 14478
rect 11118 14530 11170 14542
rect 11118 14466 11170 14478
rect 11902 14530 11954 14542
rect 11902 14466 11954 14478
rect 12350 14530 12402 14542
rect 12350 14466 12402 14478
rect 19182 14530 19234 14542
rect 27582 14530 27634 14542
rect 20626 14478 20638 14530
rect 20690 14478 20702 14530
rect 26898 14478 26910 14530
rect 26962 14478 26974 14530
rect 19182 14466 19234 14478
rect 27582 14466 27634 14478
rect 8206 14418 8258 14430
rect 9998 14418 10050 14430
rect 4722 14366 4734 14418
rect 4786 14366 4798 14418
rect 8754 14366 8766 14418
rect 8818 14366 8830 14418
rect 9090 14366 9102 14418
rect 9154 14366 9166 14418
rect 8206 14354 8258 14366
rect 9998 14354 10050 14366
rect 10110 14418 10162 14430
rect 15150 14418 15202 14430
rect 10322 14366 10334 14418
rect 10386 14366 10398 14418
rect 10110 14354 10162 14366
rect 15150 14354 15202 14366
rect 18846 14418 18898 14430
rect 18846 14354 18898 14366
rect 18958 14418 19010 14430
rect 20514 14366 20526 14418
rect 20578 14366 20590 14418
rect 18958 14354 19010 14366
rect 3726 14306 3778 14318
rect 3726 14242 3778 14254
rect 6190 14306 6242 14318
rect 6190 14242 6242 14254
rect 9886 14306 9938 14318
rect 9886 14242 9938 14254
rect 19518 14306 19570 14318
rect 19518 14242 19570 14254
rect 22430 14306 22482 14318
rect 27918 14306 27970 14318
rect 24658 14254 24670 14306
rect 24722 14254 24734 14306
rect 22430 14242 22482 14254
rect 27918 14242 27970 14254
rect 28366 14306 28418 14318
rect 28366 14242 28418 14254
rect 1344 14138 38640 14172
rect 1344 14086 14024 14138
rect 14076 14086 14148 14138
rect 14200 14086 14272 14138
rect 14324 14086 14396 14138
rect 14448 14086 14520 14138
rect 14572 14086 14644 14138
rect 14696 14086 14768 14138
rect 14820 14086 14892 14138
rect 14944 14086 15016 14138
rect 15068 14086 15140 14138
rect 15192 14086 34024 14138
rect 34076 14086 34148 14138
rect 34200 14086 34272 14138
rect 34324 14086 34396 14138
rect 34448 14086 34520 14138
rect 34572 14086 34644 14138
rect 34696 14086 34768 14138
rect 34820 14086 34892 14138
rect 34944 14086 35016 14138
rect 35068 14086 35140 14138
rect 35192 14086 38640 14138
rect 1344 14052 38640 14086
rect 5294 13970 5346 13982
rect 5294 13906 5346 13918
rect 8094 13970 8146 13982
rect 8094 13906 8146 13918
rect 10558 13970 10610 13982
rect 10558 13906 10610 13918
rect 11118 13970 11170 13982
rect 11118 13906 11170 13918
rect 12350 13970 12402 13982
rect 12350 13906 12402 13918
rect 15598 13970 15650 13982
rect 15598 13906 15650 13918
rect 16046 13970 16098 13982
rect 16046 13906 16098 13918
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 25790 13970 25842 13982
rect 25790 13906 25842 13918
rect 25902 13970 25954 13982
rect 25902 13906 25954 13918
rect 26798 13970 26850 13982
rect 26798 13906 26850 13918
rect 27358 13970 27410 13982
rect 27358 13906 27410 13918
rect 9550 13858 9602 13870
rect 9550 13794 9602 13806
rect 9886 13858 9938 13870
rect 9886 13794 9938 13806
rect 11230 13858 11282 13870
rect 20190 13858 20242 13870
rect 18050 13806 18062 13858
rect 18114 13806 18126 13858
rect 18610 13806 18622 13858
rect 18674 13806 18686 13858
rect 21186 13806 21198 13858
rect 21250 13806 21262 13858
rect 21746 13806 21758 13858
rect 21810 13806 21822 13858
rect 11230 13794 11282 13806
rect 20190 13794 20242 13806
rect 7758 13746 7810 13758
rect 7758 13682 7810 13694
rect 9102 13746 9154 13758
rect 9102 13682 9154 13694
rect 10110 13746 10162 13758
rect 10110 13682 10162 13694
rect 10782 13746 10834 13758
rect 10782 13682 10834 13694
rect 11454 13746 11506 13758
rect 14814 13746 14866 13758
rect 14242 13694 14254 13746
rect 14306 13694 14318 13746
rect 11454 13682 11506 13694
rect 14814 13682 14866 13694
rect 17838 13746 17890 13758
rect 17838 13682 17890 13694
rect 20974 13746 21026 13758
rect 20974 13682 21026 13694
rect 26014 13746 26066 13758
rect 26014 13682 26066 13694
rect 26462 13746 26514 13758
rect 26462 13682 26514 13694
rect 26686 13746 26738 13758
rect 26686 13682 26738 13694
rect 8206 13634 8258 13646
rect 8206 13570 8258 13582
rect 9662 13634 9714 13646
rect 9662 13570 9714 13582
rect 12014 13634 12066 13646
rect 12014 13570 12066 13582
rect 14926 13634 14978 13646
rect 14926 13570 14978 13582
rect 17502 13522 17554 13534
rect 17502 13458 17554 13470
rect 20638 13522 20690 13534
rect 20638 13458 20690 13470
rect 26798 13522 26850 13534
rect 26798 13458 26850 13470
rect 1344 13354 38640 13388
rect 1344 13302 4024 13354
rect 4076 13302 4148 13354
rect 4200 13302 4272 13354
rect 4324 13302 4396 13354
rect 4448 13302 4520 13354
rect 4572 13302 4644 13354
rect 4696 13302 4768 13354
rect 4820 13302 4892 13354
rect 4944 13302 5016 13354
rect 5068 13302 5140 13354
rect 5192 13302 24024 13354
rect 24076 13302 24148 13354
rect 24200 13302 24272 13354
rect 24324 13302 24396 13354
rect 24448 13302 24520 13354
rect 24572 13302 24644 13354
rect 24696 13302 24768 13354
rect 24820 13302 24892 13354
rect 24944 13302 25016 13354
rect 25068 13302 25140 13354
rect 25192 13302 38640 13354
rect 1344 13268 38640 13302
rect 3502 13186 3554 13198
rect 14030 13186 14082 13198
rect 7634 13134 7646 13186
rect 7698 13134 7710 13186
rect 9314 13134 9326 13186
rect 9378 13183 9390 13186
rect 9650 13183 9662 13186
rect 9378 13137 9662 13183
rect 9378 13134 9390 13137
rect 9650 13134 9662 13137
rect 9714 13134 9726 13186
rect 3502 13122 3554 13134
rect 14030 13122 14082 13134
rect 19966 13186 20018 13198
rect 19966 13122 20018 13134
rect 23214 13186 23266 13198
rect 23214 13122 23266 13134
rect 24558 13186 24610 13198
rect 24558 13122 24610 13134
rect 4846 13074 4898 13086
rect 4846 13010 4898 13022
rect 5742 13074 5794 13086
rect 9550 13074 9602 13086
rect 8754 13022 8766 13074
rect 8818 13022 8830 13074
rect 5742 13010 5794 13022
rect 9550 13010 9602 13022
rect 22430 13074 22482 13086
rect 26562 13022 26574 13074
rect 26626 13022 26638 13074
rect 22430 13010 22482 13022
rect 6974 12962 7026 12974
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 6974 12898 7026 12910
rect 7198 12962 7250 12974
rect 10782 12962 10834 12974
rect 8306 12910 8318 12962
rect 8370 12910 8382 12962
rect 7198 12898 7250 12910
rect 10782 12898 10834 12910
rect 11230 12962 11282 12974
rect 11230 12898 11282 12910
rect 11454 12962 11506 12974
rect 11454 12898 11506 12910
rect 15822 12962 15874 12974
rect 24446 12962 24498 12974
rect 16370 12910 16382 12962
rect 16434 12910 16446 12962
rect 16930 12910 16942 12962
rect 16994 12910 17006 12962
rect 27794 12910 27806 12962
rect 27858 12910 27870 12962
rect 15822 12898 15874 12910
rect 24446 12898 24498 12910
rect 7086 12850 7138 12862
rect 4050 12798 4062 12850
rect 4114 12798 4126 12850
rect 7086 12786 7138 12798
rect 8766 12850 8818 12862
rect 8766 12786 8818 12798
rect 8878 12850 8930 12862
rect 8878 12786 8930 12798
rect 10334 12850 10386 12862
rect 10334 12786 10386 12798
rect 12910 12850 12962 12862
rect 14354 12798 14366 12850
rect 14418 12798 14430 12850
rect 14578 12798 14590 12850
rect 14642 12798 14654 12850
rect 23426 12798 23438 12850
rect 23490 12798 23502 12850
rect 23986 12798 23998 12850
rect 24050 12798 24062 12850
rect 12910 12786 12962 12798
rect 3166 12738 3218 12750
rect 3166 12674 3218 12686
rect 9102 12738 9154 12750
rect 9102 12674 9154 12686
rect 11342 12738 11394 12750
rect 11342 12674 11394 12686
rect 13694 12738 13746 12750
rect 13694 12674 13746 12686
rect 15374 12738 15426 12750
rect 15374 12674 15426 12686
rect 15598 12738 15650 12750
rect 15598 12674 15650 12686
rect 15710 12738 15762 12750
rect 20302 12738 20354 12750
rect 19170 12686 19182 12738
rect 19234 12686 19246 12738
rect 15710 12674 15762 12686
rect 20302 12674 20354 12686
rect 22878 12738 22930 12750
rect 22878 12674 22930 12686
rect 1344 12570 38640 12604
rect 1344 12518 14024 12570
rect 14076 12518 14148 12570
rect 14200 12518 14272 12570
rect 14324 12518 14396 12570
rect 14448 12518 14520 12570
rect 14572 12518 14644 12570
rect 14696 12518 14768 12570
rect 14820 12518 14892 12570
rect 14944 12518 15016 12570
rect 15068 12518 15140 12570
rect 15192 12518 34024 12570
rect 34076 12518 34148 12570
rect 34200 12518 34272 12570
rect 34324 12518 34396 12570
rect 34448 12518 34520 12570
rect 34572 12518 34644 12570
rect 34696 12518 34768 12570
rect 34820 12518 34892 12570
rect 34944 12518 35016 12570
rect 35068 12518 35140 12570
rect 35192 12518 38640 12570
rect 1344 12484 38640 12518
rect 6078 12402 6130 12414
rect 4834 12350 4846 12402
rect 4898 12350 4910 12402
rect 6078 12338 6130 12350
rect 8206 12402 8258 12414
rect 8206 12338 8258 12350
rect 8542 12402 8594 12414
rect 8542 12338 8594 12350
rect 8990 12402 9042 12414
rect 8990 12338 9042 12350
rect 10334 12402 10386 12414
rect 10334 12338 10386 12350
rect 10558 12402 10610 12414
rect 10558 12338 10610 12350
rect 10894 12402 10946 12414
rect 10894 12338 10946 12350
rect 13246 12402 13298 12414
rect 17502 12402 17554 12414
rect 13906 12350 13918 12402
rect 13970 12350 13982 12402
rect 13246 12338 13298 12350
rect 17502 12338 17554 12350
rect 20414 12402 20466 12414
rect 20414 12338 20466 12350
rect 28254 12402 28306 12414
rect 28254 12338 28306 12350
rect 6862 12290 6914 12302
rect 6862 12226 6914 12238
rect 6526 12178 6578 12190
rect 1810 12126 1822 12178
rect 1874 12126 1886 12178
rect 2370 12126 2382 12178
rect 2434 12126 2446 12178
rect 6526 12114 6578 12126
rect 6750 12178 6802 12190
rect 6750 12114 6802 12126
rect 7086 12178 7138 12190
rect 7086 12114 7138 12126
rect 7534 12178 7586 12190
rect 7534 12114 7586 12126
rect 7758 12178 7810 12190
rect 7758 12114 7810 12126
rect 10222 12178 10274 12190
rect 16718 12178 16770 12190
rect 16258 12126 16270 12178
rect 16322 12126 16334 12178
rect 19842 12126 19854 12178
rect 19906 12126 19918 12178
rect 27346 12126 27358 12178
rect 27410 12126 27422 12178
rect 10222 12114 10274 12126
rect 16718 12114 16770 12126
rect 7310 12066 7362 12078
rect 7310 12002 7362 12014
rect 17950 12066 18002 12078
rect 17950 12002 18002 12014
rect 22430 12066 22482 12078
rect 22430 12002 22482 12014
rect 5406 11954 5458 11966
rect 5406 11890 5458 11902
rect 25454 11954 25506 11966
rect 25454 11890 25506 11902
rect 1344 11786 38640 11820
rect 1344 11734 4024 11786
rect 4076 11734 4148 11786
rect 4200 11734 4272 11786
rect 4324 11734 4396 11786
rect 4448 11734 4520 11786
rect 4572 11734 4644 11786
rect 4696 11734 4768 11786
rect 4820 11734 4892 11786
rect 4944 11734 5016 11786
rect 5068 11734 5140 11786
rect 5192 11734 24024 11786
rect 24076 11734 24148 11786
rect 24200 11734 24272 11786
rect 24324 11734 24396 11786
rect 24448 11734 24520 11786
rect 24572 11734 24644 11786
rect 24696 11734 24768 11786
rect 24820 11734 24892 11786
rect 24944 11734 25016 11786
rect 25068 11734 25140 11786
rect 25192 11734 38640 11786
rect 1344 11700 38640 11734
rect 3390 11618 3442 11630
rect 3390 11554 3442 11566
rect 3726 11618 3778 11630
rect 3726 11554 3778 11566
rect 6974 11618 7026 11630
rect 6974 11554 7026 11566
rect 11678 11618 11730 11630
rect 11678 11554 11730 11566
rect 25790 11618 25842 11630
rect 25790 11554 25842 11566
rect 5070 11506 5122 11518
rect 5070 11442 5122 11454
rect 7534 11506 7586 11518
rect 7534 11442 7586 11454
rect 17390 11506 17442 11518
rect 17390 11442 17442 11454
rect 26126 11506 26178 11518
rect 26126 11442 26178 11454
rect 6862 11394 6914 11406
rect 4386 11342 4398 11394
rect 4450 11342 4462 11394
rect 6862 11330 6914 11342
rect 7982 11394 8034 11406
rect 13582 11394 13634 11406
rect 22318 11394 22370 11406
rect 8642 11342 8654 11394
rect 8706 11342 8718 11394
rect 13906 11342 13918 11394
rect 13970 11342 13982 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 7982 11330 8034 11342
rect 13582 11330 13634 11342
rect 22318 11330 22370 11342
rect 6974 11282 7026 11294
rect 4498 11230 4510 11282
rect 4562 11230 4574 11282
rect 6974 11218 7026 11230
rect 17838 11282 17890 11294
rect 17838 11218 17890 11230
rect 5742 11170 5794 11182
rect 12014 11170 12066 11182
rect 10882 11118 10894 11170
rect 10946 11118 10958 11170
rect 5742 11106 5794 11118
rect 12014 11106 12066 11118
rect 12462 11170 12514 11182
rect 17054 11170 17106 11182
rect 26574 11170 26626 11182
rect 16370 11118 16382 11170
rect 16434 11118 16446 11170
rect 24994 11118 25006 11170
rect 25058 11118 25070 11170
rect 12462 11106 12514 11118
rect 17054 11106 17106 11118
rect 26574 11106 26626 11118
rect 1344 11002 38640 11036
rect 1344 10950 14024 11002
rect 14076 10950 14148 11002
rect 14200 10950 14272 11002
rect 14324 10950 14396 11002
rect 14448 10950 14520 11002
rect 14572 10950 14644 11002
rect 14696 10950 14768 11002
rect 14820 10950 14892 11002
rect 14944 10950 15016 11002
rect 15068 10950 15140 11002
rect 15192 10950 34024 11002
rect 34076 10950 34148 11002
rect 34200 10950 34272 11002
rect 34324 10950 34396 11002
rect 34448 10950 34520 11002
rect 34572 10950 34644 11002
rect 34696 10950 34768 11002
rect 34820 10950 34892 11002
rect 34944 10950 35016 11002
rect 35068 10950 35140 11002
rect 35192 10950 38640 11002
rect 1344 10916 38640 10950
rect 5294 10834 5346 10846
rect 4722 10782 4734 10834
rect 4786 10782 4798 10834
rect 5294 10770 5346 10782
rect 5406 10834 5458 10846
rect 9662 10834 9714 10846
rect 5954 10782 5966 10834
rect 6018 10782 6030 10834
rect 5406 10770 5458 10782
rect 9662 10770 9714 10782
rect 10110 10834 10162 10846
rect 14030 10834 14082 10846
rect 13234 10782 13246 10834
rect 13298 10782 13310 10834
rect 10110 10770 10162 10782
rect 14030 10770 14082 10782
rect 14590 10834 14642 10846
rect 14590 10770 14642 10782
rect 15486 10834 15538 10846
rect 15486 10770 15538 10782
rect 15934 10834 15986 10846
rect 23214 10834 23266 10846
rect 22530 10782 22542 10834
rect 22594 10782 22606 10834
rect 15934 10770 15986 10782
rect 23214 10770 23266 10782
rect 23662 10834 23714 10846
rect 23662 10770 23714 10782
rect 15150 10722 15202 10734
rect 15150 10658 15202 10670
rect 15262 10722 15314 10734
rect 15262 10658 15314 10670
rect 23998 10722 24050 10734
rect 23998 10658 24050 10670
rect 1822 10610 1874 10622
rect 8878 10610 8930 10622
rect 2258 10558 2270 10610
rect 2322 10558 2334 10610
rect 8418 10558 8430 10610
rect 8482 10558 8494 10610
rect 1822 10546 1874 10558
rect 8878 10546 8930 10558
rect 10334 10610 10386 10622
rect 19742 10610 19794 10622
rect 10994 10558 11006 10610
rect 11058 10558 11070 10610
rect 20178 10558 20190 10610
rect 20242 10558 20254 10610
rect 10334 10546 10386 10558
rect 19742 10546 19794 10558
rect 1344 10218 38640 10252
rect 1344 10166 4024 10218
rect 4076 10166 4148 10218
rect 4200 10166 4272 10218
rect 4324 10166 4396 10218
rect 4448 10166 4520 10218
rect 4572 10166 4644 10218
rect 4696 10166 4768 10218
rect 4820 10166 4892 10218
rect 4944 10166 5016 10218
rect 5068 10166 5140 10218
rect 5192 10166 24024 10218
rect 24076 10166 24148 10218
rect 24200 10166 24272 10218
rect 24324 10166 24396 10218
rect 24448 10166 24520 10218
rect 24572 10166 24644 10218
rect 24696 10166 24768 10218
rect 24820 10166 24892 10218
rect 24944 10166 25016 10218
rect 25068 10166 25140 10218
rect 25192 10166 38640 10218
rect 1344 10132 38640 10166
rect 6190 9938 6242 9950
rect 27010 9886 27022 9938
rect 27074 9886 27086 9938
rect 6190 9874 6242 9886
rect 28018 9662 28030 9714
rect 28082 9662 28094 9714
rect 5742 9602 5794 9614
rect 5742 9538 5794 9550
rect 9214 9602 9266 9614
rect 9214 9538 9266 9550
rect 1344 9434 38640 9468
rect 1344 9382 14024 9434
rect 14076 9382 14148 9434
rect 14200 9382 14272 9434
rect 14324 9382 14396 9434
rect 14448 9382 14520 9434
rect 14572 9382 14644 9434
rect 14696 9382 14768 9434
rect 14820 9382 14892 9434
rect 14944 9382 15016 9434
rect 15068 9382 15140 9434
rect 15192 9382 34024 9434
rect 34076 9382 34148 9434
rect 34200 9382 34272 9434
rect 34324 9382 34396 9434
rect 34448 9382 34520 9434
rect 34572 9382 34644 9434
rect 34696 9382 34768 9434
rect 34820 9382 34892 9434
rect 34944 9382 35016 9434
rect 35068 9382 35140 9434
rect 35192 9382 38640 9434
rect 1344 9348 38640 9382
rect 18958 9154 19010 9166
rect 18958 9090 19010 9102
rect 28030 9154 28082 9166
rect 28030 9090 28082 9102
rect 29038 9154 29090 9166
rect 29038 9090 29090 9102
rect 18734 9042 18786 9054
rect 18734 8978 18786 8990
rect 19070 9042 19122 9054
rect 19070 8978 19122 8990
rect 25342 9042 25394 9054
rect 29598 9042 29650 9054
rect 25778 8990 25790 9042
rect 25842 8990 25854 9042
rect 25342 8978 25394 8990
rect 29598 8978 29650 8990
rect 22990 8818 23042 8830
rect 22990 8754 23042 8766
rect 28814 8818 28866 8830
rect 28814 8754 28866 8766
rect 1344 8650 38640 8684
rect 1344 8598 4024 8650
rect 4076 8598 4148 8650
rect 4200 8598 4272 8650
rect 4324 8598 4396 8650
rect 4448 8598 4520 8650
rect 4572 8598 4644 8650
rect 4696 8598 4768 8650
rect 4820 8598 4892 8650
rect 4944 8598 5016 8650
rect 5068 8598 5140 8650
rect 5192 8598 24024 8650
rect 24076 8598 24148 8650
rect 24200 8598 24272 8650
rect 24324 8598 24396 8650
rect 24448 8598 24520 8650
rect 24572 8598 24644 8650
rect 24696 8598 24768 8650
rect 24820 8598 24892 8650
rect 24944 8598 25016 8650
rect 25068 8598 25140 8650
rect 25192 8598 38640 8650
rect 1344 8564 38640 8598
rect 19406 8482 19458 8494
rect 19406 8418 19458 8430
rect 27582 8482 27634 8494
rect 27582 8418 27634 8430
rect 7982 8370 8034 8382
rect 7982 8306 8034 8318
rect 25902 8370 25954 8382
rect 25902 8306 25954 8318
rect 26350 8370 26402 8382
rect 26350 8306 26402 8318
rect 27246 8370 27298 8382
rect 27246 8306 27298 8318
rect 17950 8258 18002 8270
rect 17950 8194 18002 8206
rect 18398 8258 18450 8270
rect 19282 8206 19294 8258
rect 19346 8206 19358 8258
rect 22306 8206 22318 8258
rect 22370 8206 22382 8258
rect 22866 8206 22878 8258
rect 22930 8206 22942 8258
rect 28242 8206 28254 8258
rect 28306 8206 28318 8258
rect 18398 8194 18450 8206
rect 17614 8146 17666 8158
rect 17614 8082 17666 8094
rect 18062 8146 18114 8158
rect 18062 8082 18114 8094
rect 18734 8146 18786 8158
rect 18734 8082 18786 8094
rect 18958 8146 19010 8158
rect 18958 8082 19010 8094
rect 19966 8146 20018 8158
rect 19966 8082 20018 8094
rect 20302 8146 20354 8158
rect 28354 8094 28366 8146
rect 28418 8094 28430 8146
rect 20302 8082 20354 8094
rect 5854 8034 5906 8046
rect 5854 7970 5906 7982
rect 17838 8034 17890 8046
rect 17838 7970 17890 7982
rect 18510 8034 18562 8046
rect 18510 7970 18562 7982
rect 19518 8034 19570 8046
rect 19518 7970 19570 7982
rect 19742 8034 19794 8046
rect 19742 7970 19794 7982
rect 20190 8034 20242 8046
rect 25330 7982 25342 8034
rect 25394 7982 25406 8034
rect 20190 7970 20242 7982
rect 1344 7866 38640 7900
rect 1344 7814 14024 7866
rect 14076 7814 14148 7866
rect 14200 7814 14272 7866
rect 14324 7814 14396 7866
rect 14448 7814 14520 7866
rect 14572 7814 14644 7866
rect 14696 7814 14768 7866
rect 14820 7814 14892 7866
rect 14944 7814 15016 7866
rect 15068 7814 15140 7866
rect 15192 7814 34024 7866
rect 34076 7814 34148 7866
rect 34200 7814 34272 7866
rect 34324 7814 34396 7866
rect 34448 7814 34520 7866
rect 34572 7814 34644 7866
rect 34696 7814 34768 7866
rect 34820 7814 34892 7866
rect 34944 7814 35016 7866
rect 35068 7814 35140 7866
rect 35192 7814 38640 7866
rect 1344 7780 38640 7814
rect 6078 7698 6130 7710
rect 4722 7646 4734 7698
rect 4786 7646 4798 7698
rect 6078 7634 6130 7646
rect 15598 7698 15650 7710
rect 15598 7634 15650 7646
rect 16830 7698 16882 7710
rect 21198 7698 21250 7710
rect 20626 7646 20638 7698
rect 20690 7646 20702 7698
rect 16830 7634 16882 7646
rect 21198 7634 21250 7646
rect 21422 7698 21474 7710
rect 21422 7634 21474 7646
rect 7982 7586 8034 7598
rect 7982 7522 8034 7534
rect 8542 7586 8594 7598
rect 8542 7522 8594 7534
rect 11902 7586 11954 7598
rect 11902 7522 11954 7534
rect 24670 7586 24722 7598
rect 24670 7522 24722 7534
rect 26014 7586 26066 7598
rect 27582 7586 27634 7598
rect 27010 7534 27022 7586
rect 27074 7534 27086 7586
rect 26014 7522 26066 7534
rect 27582 7522 27634 7534
rect 1822 7474 1874 7486
rect 7534 7474 7586 7486
rect 2146 7422 2158 7474
rect 2210 7422 2222 7474
rect 6850 7422 6862 7474
rect 6914 7422 6926 7474
rect 1822 7410 1874 7422
rect 7534 7410 7586 7422
rect 8094 7474 8146 7486
rect 8094 7410 8146 7422
rect 8430 7474 8482 7486
rect 8430 7410 8482 7422
rect 8766 7474 8818 7486
rect 14590 7474 14642 7486
rect 14242 7422 14254 7474
rect 14306 7422 14318 7474
rect 8766 7410 8818 7422
rect 14590 7410 14642 7422
rect 15150 7474 15202 7486
rect 15150 7410 15202 7422
rect 17502 7474 17554 7486
rect 26350 7474 26402 7486
rect 18162 7422 18174 7474
rect 18226 7422 18238 7474
rect 27122 7422 27134 7474
rect 27186 7422 27198 7474
rect 17502 7410 17554 7422
rect 26350 7410 26402 7422
rect 5630 7362 5682 7374
rect 5630 7298 5682 7310
rect 6638 7362 6690 7374
rect 6638 7298 6690 7310
rect 9662 7362 9714 7374
rect 9662 7298 9714 7310
rect 10110 7362 10162 7374
rect 10110 7298 10162 7310
rect 21534 7362 21586 7374
rect 21534 7298 21586 7310
rect 5294 7250 5346 7262
rect 5294 7186 5346 7198
rect 6526 7250 6578 7262
rect 6526 7186 6578 7198
rect 7982 7250 8034 7262
rect 7982 7186 8034 7198
rect 11118 7250 11170 7262
rect 11118 7186 11170 7198
rect 1344 7082 38640 7116
rect 1344 7030 4024 7082
rect 4076 7030 4148 7082
rect 4200 7030 4272 7082
rect 4324 7030 4396 7082
rect 4448 7030 4520 7082
rect 4572 7030 4644 7082
rect 4696 7030 4768 7082
rect 4820 7030 4892 7082
rect 4944 7030 5016 7082
rect 5068 7030 5140 7082
rect 5192 7030 24024 7082
rect 24076 7030 24148 7082
rect 24200 7030 24272 7082
rect 24324 7030 24396 7082
rect 24448 7030 24520 7082
rect 24572 7030 24644 7082
rect 24696 7030 24768 7082
rect 24820 7030 24892 7082
rect 24944 7030 25016 7082
rect 25068 7030 25140 7082
rect 25192 7030 38640 7082
rect 1344 6996 38640 7030
rect 5742 6914 5794 6926
rect 5742 6850 5794 6862
rect 6190 6914 6242 6926
rect 6190 6850 6242 6862
rect 6302 6914 6354 6926
rect 6302 6850 6354 6862
rect 6750 6914 6802 6926
rect 6750 6850 6802 6862
rect 6974 6914 7026 6926
rect 6974 6850 7026 6862
rect 8094 6914 8146 6926
rect 8094 6850 8146 6862
rect 21310 6914 21362 6926
rect 21310 6850 21362 6862
rect 21422 6802 21474 6814
rect 4498 6750 4510 6802
rect 4562 6750 4574 6802
rect 15026 6750 15038 6802
rect 15090 6750 15102 6802
rect 26786 6750 26798 6802
rect 26850 6750 26862 6802
rect 21422 6738 21474 6750
rect 2270 6690 2322 6702
rect 2270 6626 2322 6638
rect 2494 6690 2546 6702
rect 5854 6690 5906 6702
rect 8542 6690 8594 6702
rect 4050 6638 4062 6690
rect 4114 6638 4126 6690
rect 7746 6638 7758 6690
rect 7810 6638 7822 6690
rect 2494 6626 2546 6638
rect 5854 6626 5906 6638
rect 8542 6626 8594 6638
rect 9214 6690 9266 6702
rect 9214 6626 9266 6638
rect 9326 6690 9378 6702
rect 17054 6690 17106 6702
rect 22094 6690 22146 6702
rect 9986 6638 9998 6690
rect 10050 6638 10062 6690
rect 17714 6638 17726 6690
rect 17778 6638 17790 6690
rect 22418 6638 22430 6690
rect 22482 6638 22494 6690
rect 9326 6626 9378 6638
rect 17054 6626 17106 6638
rect 22094 6626 22146 6638
rect 2606 6578 2658 6590
rect 2606 6514 2658 6526
rect 2942 6578 2994 6590
rect 6414 6578 6466 6590
rect 3602 6526 3614 6578
rect 3666 6526 3678 6578
rect 2942 6514 2994 6526
rect 6414 6514 6466 6526
rect 7534 6578 7586 6590
rect 7534 6514 7586 6526
rect 7982 6578 8034 6590
rect 7982 6514 8034 6526
rect 12238 6578 12290 6590
rect 12238 6514 12290 6526
rect 13022 6578 13074 6590
rect 16718 6578 16770 6590
rect 13906 6526 13918 6578
rect 13970 6526 13982 6578
rect 13022 6514 13074 6526
rect 16718 6514 16770 6526
rect 16830 6578 16882 6590
rect 16830 6514 16882 6526
rect 25566 6578 25618 6590
rect 27794 6526 27806 6578
rect 27858 6526 27870 6578
rect 25566 6514 25618 6526
rect 3054 6466 3106 6478
rect 3054 6402 3106 6414
rect 3278 6466 3330 6478
rect 3278 6402 3330 6414
rect 5742 6466 5794 6478
rect 5742 6402 5794 6414
rect 8654 6466 8706 6478
rect 8654 6402 8706 6414
rect 8766 6466 8818 6478
rect 8766 6402 8818 6414
rect 16494 6466 16546 6478
rect 20750 6466 20802 6478
rect 26014 6466 26066 6478
rect 20066 6414 20078 6466
rect 20130 6414 20142 6466
rect 24994 6414 25006 6466
rect 25058 6414 25070 6466
rect 16494 6402 16546 6414
rect 20750 6402 20802 6414
rect 26014 6402 26066 6414
rect 1344 6298 38640 6332
rect 1344 6246 14024 6298
rect 14076 6246 14148 6298
rect 14200 6246 14272 6298
rect 14324 6246 14396 6298
rect 14448 6246 14520 6298
rect 14572 6246 14644 6298
rect 14696 6246 14768 6298
rect 14820 6246 14892 6298
rect 14944 6246 15016 6298
rect 15068 6246 15140 6298
rect 15192 6246 34024 6298
rect 34076 6246 34148 6298
rect 34200 6246 34272 6298
rect 34324 6246 34396 6298
rect 34448 6246 34520 6298
rect 34572 6246 34644 6298
rect 34696 6246 34768 6298
rect 34820 6246 34892 6298
rect 34944 6246 35016 6298
rect 35068 6246 35140 6298
rect 35192 6246 38640 6298
rect 1344 6212 38640 6246
rect 7870 6130 7922 6142
rect 13246 6130 13298 6142
rect 17502 6130 17554 6142
rect 7298 6078 7310 6130
rect 7362 6078 7374 6130
rect 8978 6078 8990 6130
rect 9042 6078 9054 6130
rect 12338 6078 12350 6130
rect 12402 6078 12414 6130
rect 13794 6078 13806 6130
rect 13858 6078 13870 6130
rect 7870 6066 7922 6078
rect 13246 6066 13298 6078
rect 17502 6066 17554 6078
rect 18286 6130 18338 6142
rect 18286 6066 18338 6078
rect 18398 6130 18450 6142
rect 18398 6066 18450 6078
rect 18622 6130 18674 6142
rect 28814 6130 28866 6142
rect 28130 6078 28142 6130
rect 28194 6078 28206 6130
rect 18622 6066 18674 6078
rect 28814 6066 28866 6078
rect 2494 6018 2546 6030
rect 2494 5954 2546 5966
rect 3166 6018 3218 6030
rect 3166 5954 3218 5966
rect 3502 6018 3554 6030
rect 3502 5954 3554 5966
rect 8318 6018 8370 6030
rect 8318 5954 8370 5966
rect 17614 6018 17666 6030
rect 17614 5954 17666 5966
rect 2830 5906 2882 5918
rect 2830 5842 2882 5854
rect 4174 5906 4226 5918
rect 8430 5906 8482 5918
rect 4722 5854 4734 5906
rect 4786 5854 4798 5906
rect 4174 5842 4226 5854
rect 8430 5842 8482 5854
rect 8542 5906 8594 5918
rect 8542 5842 8594 5854
rect 9438 5906 9490 5918
rect 17278 5906 17330 5918
rect 9986 5854 9998 5906
rect 10050 5854 10062 5906
rect 16370 5854 16382 5906
rect 16434 5854 16446 5906
rect 16818 5854 16830 5906
rect 16882 5854 16894 5906
rect 9438 5842 9490 5854
rect 17278 5842 17330 5854
rect 18174 5906 18226 5918
rect 25342 5906 25394 5918
rect 24322 5854 24334 5906
rect 24386 5854 24398 5906
rect 25778 5854 25790 5906
rect 25842 5854 25854 5906
rect 18174 5842 18226 5854
rect 25342 5842 25394 5854
rect 2046 5794 2098 5806
rect 2046 5730 2098 5742
rect 3614 5794 3666 5806
rect 22306 5742 22318 5794
rect 22370 5742 22382 5794
rect 3614 5730 3666 5742
rect 2382 5682 2434 5694
rect 2382 5618 2434 5630
rect 13134 5682 13186 5694
rect 13134 5618 13186 5630
rect 1344 5514 38640 5548
rect 1344 5462 4024 5514
rect 4076 5462 4148 5514
rect 4200 5462 4272 5514
rect 4324 5462 4396 5514
rect 4448 5462 4520 5514
rect 4572 5462 4644 5514
rect 4696 5462 4768 5514
rect 4820 5462 4892 5514
rect 4944 5462 5016 5514
rect 5068 5462 5140 5514
rect 5192 5462 24024 5514
rect 24076 5462 24148 5514
rect 24200 5462 24272 5514
rect 24324 5462 24396 5514
rect 24448 5462 24520 5514
rect 24572 5462 24644 5514
rect 24696 5462 24768 5514
rect 24820 5462 24892 5514
rect 24944 5462 25016 5514
rect 25068 5462 25140 5514
rect 25192 5462 38640 5514
rect 1344 5428 38640 5462
rect 6862 5346 6914 5358
rect 6862 5282 6914 5294
rect 22206 5346 22258 5358
rect 22206 5282 22258 5294
rect 5966 5234 6018 5246
rect 5966 5170 6018 5182
rect 11342 5234 11394 5246
rect 11342 5170 11394 5182
rect 13582 5234 13634 5246
rect 13582 5170 13634 5182
rect 14030 5234 14082 5246
rect 14030 5170 14082 5182
rect 21310 5234 21362 5246
rect 25330 5182 25342 5234
rect 25394 5182 25406 5234
rect 21310 5170 21362 5182
rect 5742 5122 5794 5134
rect 5742 5058 5794 5070
rect 5854 5122 5906 5134
rect 5854 5058 5906 5070
rect 6078 5122 6130 5134
rect 10334 5122 10386 5134
rect 6290 5070 6302 5122
rect 6354 5070 6366 5122
rect 9874 5070 9886 5122
rect 9938 5070 9950 5122
rect 6078 5058 6130 5070
rect 10334 5058 10386 5070
rect 10894 5122 10946 5134
rect 20402 5070 20414 5122
rect 20466 5070 20478 5122
rect 22530 5070 22542 5122
rect 22594 5070 22606 5122
rect 10894 5058 10946 5070
rect 15362 4958 15374 5010
rect 15426 4958 15438 5010
rect 7522 4846 7534 4898
rect 7586 4846 7598 4898
rect 1344 4730 38640 4764
rect 1344 4678 14024 4730
rect 14076 4678 14148 4730
rect 14200 4678 14272 4730
rect 14324 4678 14396 4730
rect 14448 4678 14520 4730
rect 14572 4678 14644 4730
rect 14696 4678 14768 4730
rect 14820 4678 14892 4730
rect 14944 4678 15016 4730
rect 15068 4678 15140 4730
rect 15192 4678 34024 4730
rect 34076 4678 34148 4730
rect 34200 4678 34272 4730
rect 34324 4678 34396 4730
rect 34448 4678 34520 4730
rect 34572 4678 34644 4730
rect 34696 4678 34768 4730
rect 34820 4678 34892 4730
rect 34944 4678 35016 4730
rect 35068 4678 35140 4730
rect 35192 4678 38640 4730
rect 1344 4644 38640 4678
rect 6078 4562 6130 4574
rect 4722 4510 4734 4562
rect 4786 4510 4798 4562
rect 6078 4498 6130 4510
rect 6302 4562 6354 4574
rect 6302 4498 6354 4510
rect 6414 4562 6466 4574
rect 6414 4498 6466 4510
rect 6526 4562 6578 4574
rect 6526 4498 6578 4510
rect 8318 4562 8370 4574
rect 8318 4498 8370 4510
rect 8878 4562 8930 4574
rect 8878 4498 8930 4510
rect 9102 4562 9154 4574
rect 26910 4562 26962 4574
rect 12562 4510 12574 4562
rect 12626 4510 12638 4562
rect 16370 4510 16382 4562
rect 16434 4510 16446 4562
rect 9102 4498 9154 4510
rect 26910 4498 26962 4510
rect 5406 4450 5458 4462
rect 5406 4386 5458 4398
rect 7422 4450 7474 4462
rect 7422 4386 7474 4398
rect 8430 4450 8482 4462
rect 8430 4386 8482 4398
rect 8766 4450 8818 4462
rect 8766 4386 8818 4398
rect 18062 4450 18114 4462
rect 18062 4386 18114 4398
rect 23998 4450 24050 4462
rect 23998 4386 24050 4398
rect 24782 4450 24834 4462
rect 25890 4398 25902 4450
rect 25954 4398 25966 4450
rect 24782 4386 24834 4398
rect 6974 4338 7026 4350
rect 9662 4338 9714 4350
rect 13246 4338 13298 4350
rect 20974 4338 21026 4350
rect 1698 4286 1710 4338
rect 1762 4286 1774 4338
rect 2258 4286 2270 4338
rect 2322 4286 2334 4338
rect 8082 4286 8094 4338
rect 8146 4286 8158 4338
rect 10098 4286 10110 4338
rect 10162 4286 10174 4338
rect 13906 4286 13918 4338
rect 13970 4286 13982 4338
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 6974 4274 7026 4286
rect 9662 4274 9714 4286
rect 13246 4274 13298 4286
rect 20974 4274 21026 4286
rect 21086 4338 21138 4350
rect 21746 4286 21758 4338
rect 21810 4286 21822 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 21086 4274 21138 4286
rect 7310 4226 7362 4238
rect 7310 4162 7362 4174
rect 25454 4226 25506 4238
rect 25454 4162 25506 4174
rect 13134 4114 13186 4126
rect 13134 4050 13186 4062
rect 16942 4114 16994 4126
rect 16942 4050 16994 4062
rect 17278 4114 17330 4126
rect 17278 4050 17330 4062
rect 26574 4114 26626 4126
rect 26574 4050 26626 4062
rect 1344 3946 38640 3980
rect 1344 3894 4024 3946
rect 4076 3894 4148 3946
rect 4200 3894 4272 3946
rect 4324 3894 4396 3946
rect 4448 3894 4520 3946
rect 4572 3894 4644 3946
rect 4696 3894 4768 3946
rect 4820 3894 4892 3946
rect 4944 3894 5016 3946
rect 5068 3894 5140 3946
rect 5192 3894 24024 3946
rect 24076 3894 24148 3946
rect 24200 3894 24272 3946
rect 24324 3894 24396 3946
rect 24448 3894 24520 3946
rect 24572 3894 24644 3946
rect 24696 3894 24768 3946
rect 24820 3894 24892 3946
rect 24944 3894 25016 3946
rect 25068 3894 25140 3946
rect 25192 3894 38640 3946
rect 1344 3860 38640 3894
rect 19742 3778 19794 3790
rect 19742 3714 19794 3726
rect 5966 3666 6018 3678
rect 5966 3602 6018 3614
rect 6414 3666 6466 3678
rect 6414 3602 6466 3614
rect 8318 3666 8370 3678
rect 19854 3666 19906 3678
rect 16930 3614 16942 3666
rect 16994 3614 17006 3666
rect 21970 3614 21982 3666
rect 22034 3614 22046 3666
rect 8318 3602 8370 3614
rect 19854 3602 19906 3614
rect 13246 3442 13298 3454
rect 16158 3442 16210 3454
rect 18734 3442 18786 3454
rect 13682 3390 13694 3442
rect 13746 3390 13758 3442
rect 17938 3390 17950 3442
rect 18002 3390 18014 3442
rect 13246 3378 13298 3390
rect 16158 3378 16210 3390
rect 18734 3378 18786 3390
rect 19070 3442 19122 3454
rect 20850 3390 20862 3442
rect 20914 3390 20926 3442
rect 19070 3378 19122 3390
rect 1344 3162 38640 3196
rect 1344 3110 14024 3162
rect 14076 3110 14148 3162
rect 14200 3110 14272 3162
rect 14324 3110 14396 3162
rect 14448 3110 14520 3162
rect 14572 3110 14644 3162
rect 14696 3110 14768 3162
rect 14820 3110 14892 3162
rect 14944 3110 15016 3162
rect 15068 3110 15140 3162
rect 15192 3110 34024 3162
rect 34076 3110 34148 3162
rect 34200 3110 34272 3162
rect 34324 3110 34396 3162
rect 34448 3110 34520 3162
rect 34572 3110 34644 3162
rect 34696 3110 34768 3162
rect 34820 3110 34892 3162
rect 34944 3110 35016 3162
rect 35068 3110 35140 3162
rect 35192 3110 38640 3162
rect 1344 3076 38640 3110
<< via1 >>
rect 4024 96406 4076 96458
rect 4148 96406 4200 96458
rect 4272 96406 4324 96458
rect 4396 96406 4448 96458
rect 4520 96406 4572 96458
rect 4644 96406 4696 96458
rect 4768 96406 4820 96458
rect 4892 96406 4944 96458
rect 5016 96406 5068 96458
rect 5140 96406 5192 96458
rect 24024 96406 24076 96458
rect 24148 96406 24200 96458
rect 24272 96406 24324 96458
rect 24396 96406 24448 96458
rect 24520 96406 24572 96458
rect 24644 96406 24696 96458
rect 24768 96406 24820 96458
rect 24892 96406 24944 96458
rect 25016 96406 25068 96458
rect 25140 96406 25192 96458
rect 30270 96014 30322 96066
rect 30046 95902 30098 95954
rect 1710 95790 1762 95842
rect 29822 95790 29874 95842
rect 14024 95622 14076 95674
rect 14148 95622 14200 95674
rect 14272 95622 14324 95674
rect 14396 95622 14448 95674
rect 14520 95622 14572 95674
rect 14644 95622 14696 95674
rect 14768 95622 14820 95674
rect 14892 95622 14944 95674
rect 15016 95622 15068 95674
rect 15140 95622 15192 95674
rect 34024 95622 34076 95674
rect 34148 95622 34200 95674
rect 34272 95622 34324 95674
rect 34396 95622 34448 95674
rect 34520 95622 34572 95674
rect 34644 95622 34696 95674
rect 34768 95622 34820 95674
rect 34892 95622 34944 95674
rect 35016 95622 35068 95674
rect 35140 95622 35192 95674
rect 4024 94838 4076 94890
rect 4148 94838 4200 94890
rect 4272 94838 4324 94890
rect 4396 94838 4448 94890
rect 4520 94838 4572 94890
rect 4644 94838 4696 94890
rect 4768 94838 4820 94890
rect 4892 94838 4944 94890
rect 5016 94838 5068 94890
rect 5140 94838 5192 94890
rect 24024 94838 24076 94890
rect 24148 94838 24200 94890
rect 24272 94838 24324 94890
rect 24396 94838 24448 94890
rect 24520 94838 24572 94890
rect 24644 94838 24696 94890
rect 24768 94838 24820 94890
rect 24892 94838 24944 94890
rect 25016 94838 25068 94890
rect 25140 94838 25192 94890
rect 1710 94222 1762 94274
rect 14024 94054 14076 94106
rect 14148 94054 14200 94106
rect 14272 94054 14324 94106
rect 14396 94054 14448 94106
rect 14520 94054 14572 94106
rect 14644 94054 14696 94106
rect 14768 94054 14820 94106
rect 14892 94054 14944 94106
rect 15016 94054 15068 94106
rect 15140 94054 15192 94106
rect 34024 94054 34076 94106
rect 34148 94054 34200 94106
rect 34272 94054 34324 94106
rect 34396 94054 34448 94106
rect 34520 94054 34572 94106
rect 34644 94054 34696 94106
rect 34768 94054 34820 94106
rect 34892 94054 34944 94106
rect 35016 94054 35068 94106
rect 35140 94054 35192 94106
rect 1710 93774 1762 93826
rect 4024 93270 4076 93322
rect 4148 93270 4200 93322
rect 4272 93270 4324 93322
rect 4396 93270 4448 93322
rect 4520 93270 4572 93322
rect 4644 93270 4696 93322
rect 4768 93270 4820 93322
rect 4892 93270 4944 93322
rect 5016 93270 5068 93322
rect 5140 93270 5192 93322
rect 24024 93270 24076 93322
rect 24148 93270 24200 93322
rect 24272 93270 24324 93322
rect 24396 93270 24448 93322
rect 24520 93270 24572 93322
rect 24644 93270 24696 93322
rect 24768 93270 24820 93322
rect 24892 93270 24944 93322
rect 25016 93270 25068 93322
rect 25140 93270 25192 93322
rect 14024 92486 14076 92538
rect 14148 92486 14200 92538
rect 14272 92486 14324 92538
rect 14396 92486 14448 92538
rect 14520 92486 14572 92538
rect 14644 92486 14696 92538
rect 14768 92486 14820 92538
rect 14892 92486 14944 92538
rect 15016 92486 15068 92538
rect 15140 92486 15192 92538
rect 34024 92486 34076 92538
rect 34148 92486 34200 92538
rect 34272 92486 34324 92538
rect 34396 92486 34448 92538
rect 34520 92486 34572 92538
rect 34644 92486 34696 92538
rect 34768 92486 34820 92538
rect 34892 92486 34944 92538
rect 35016 92486 35068 92538
rect 35140 92486 35192 92538
rect 1710 92206 1762 92258
rect 4024 91702 4076 91754
rect 4148 91702 4200 91754
rect 4272 91702 4324 91754
rect 4396 91702 4448 91754
rect 4520 91702 4572 91754
rect 4644 91702 4696 91754
rect 4768 91702 4820 91754
rect 4892 91702 4944 91754
rect 5016 91702 5068 91754
rect 5140 91702 5192 91754
rect 24024 91702 24076 91754
rect 24148 91702 24200 91754
rect 24272 91702 24324 91754
rect 24396 91702 24448 91754
rect 24520 91702 24572 91754
rect 24644 91702 24696 91754
rect 24768 91702 24820 91754
rect 24892 91702 24944 91754
rect 25016 91702 25068 91754
rect 25140 91702 25192 91754
rect 1710 91086 1762 91138
rect 14024 90918 14076 90970
rect 14148 90918 14200 90970
rect 14272 90918 14324 90970
rect 14396 90918 14448 90970
rect 14520 90918 14572 90970
rect 14644 90918 14696 90970
rect 14768 90918 14820 90970
rect 14892 90918 14944 90970
rect 15016 90918 15068 90970
rect 15140 90918 15192 90970
rect 34024 90918 34076 90970
rect 34148 90918 34200 90970
rect 34272 90918 34324 90970
rect 34396 90918 34448 90970
rect 34520 90918 34572 90970
rect 34644 90918 34696 90970
rect 34768 90918 34820 90970
rect 34892 90918 34944 90970
rect 35016 90918 35068 90970
rect 35140 90918 35192 90970
rect 4024 90134 4076 90186
rect 4148 90134 4200 90186
rect 4272 90134 4324 90186
rect 4396 90134 4448 90186
rect 4520 90134 4572 90186
rect 4644 90134 4696 90186
rect 4768 90134 4820 90186
rect 4892 90134 4944 90186
rect 5016 90134 5068 90186
rect 5140 90134 5192 90186
rect 24024 90134 24076 90186
rect 24148 90134 24200 90186
rect 24272 90134 24324 90186
rect 24396 90134 24448 90186
rect 24520 90134 24572 90186
rect 24644 90134 24696 90186
rect 24768 90134 24820 90186
rect 24892 90134 24944 90186
rect 25016 90134 25068 90186
rect 25140 90134 25192 90186
rect 1710 89630 1762 89682
rect 13694 89518 13746 89570
rect 14024 89350 14076 89402
rect 14148 89350 14200 89402
rect 14272 89350 14324 89402
rect 14396 89350 14448 89402
rect 14520 89350 14572 89402
rect 14644 89350 14696 89402
rect 14768 89350 14820 89402
rect 14892 89350 14944 89402
rect 15016 89350 15068 89402
rect 15140 89350 15192 89402
rect 34024 89350 34076 89402
rect 34148 89350 34200 89402
rect 34272 89350 34324 89402
rect 34396 89350 34448 89402
rect 34520 89350 34572 89402
rect 34644 89350 34696 89402
rect 34768 89350 34820 89402
rect 34892 89350 34944 89402
rect 35016 89350 35068 89402
rect 35140 89350 35192 89402
rect 1710 89070 1762 89122
rect 12350 89070 12402 89122
rect 9438 88958 9490 89010
rect 9998 88958 10050 89010
rect 8542 88846 8594 88898
rect 8990 88846 9042 88898
rect 13582 88846 13634 88898
rect 13918 88846 13970 88898
rect 13134 88734 13186 88786
rect 4024 88566 4076 88618
rect 4148 88566 4200 88618
rect 4272 88566 4324 88618
rect 4396 88566 4448 88618
rect 4520 88566 4572 88618
rect 4644 88566 4696 88618
rect 4768 88566 4820 88618
rect 4892 88566 4944 88618
rect 5016 88566 5068 88618
rect 5140 88566 5192 88618
rect 24024 88566 24076 88618
rect 24148 88566 24200 88618
rect 24272 88566 24324 88618
rect 24396 88566 24448 88618
rect 24520 88566 24572 88618
rect 24644 88566 24696 88618
rect 24768 88566 24820 88618
rect 24892 88566 24944 88618
rect 25016 88566 25068 88618
rect 25140 88566 25192 88618
rect 9102 88174 9154 88226
rect 9774 88174 9826 88226
rect 13918 88174 13970 88226
rect 14142 88062 14194 88114
rect 14702 88062 14754 88114
rect 1710 87950 1762 88002
rect 8430 87950 8482 88002
rect 8878 87950 8930 88002
rect 12014 87950 12066 88002
rect 12798 87950 12850 88002
rect 13582 87950 13634 88002
rect 14024 87782 14076 87834
rect 14148 87782 14200 87834
rect 14272 87782 14324 87834
rect 14396 87782 14448 87834
rect 14520 87782 14572 87834
rect 14644 87782 14696 87834
rect 14768 87782 14820 87834
rect 14892 87782 14944 87834
rect 15016 87782 15068 87834
rect 15140 87782 15192 87834
rect 34024 87782 34076 87834
rect 34148 87782 34200 87834
rect 34272 87782 34324 87834
rect 34396 87782 34448 87834
rect 34520 87782 34572 87834
rect 34644 87782 34696 87834
rect 34768 87782 34820 87834
rect 34892 87782 34944 87834
rect 35016 87782 35068 87834
rect 35140 87782 35192 87834
rect 8430 87614 8482 87666
rect 9886 87614 9938 87666
rect 10334 87614 10386 87666
rect 15038 87614 15090 87666
rect 16382 87614 16434 87666
rect 20414 87614 20466 87666
rect 10894 87502 10946 87554
rect 11454 87502 11506 87554
rect 5630 87390 5682 87442
rect 6078 87390 6130 87442
rect 9102 87390 9154 87442
rect 12126 87390 12178 87442
rect 12574 87390 12626 87442
rect 17390 87390 17442 87442
rect 17950 87390 18002 87442
rect 20974 87390 21026 87442
rect 21310 87390 21362 87442
rect 16046 87278 16098 87330
rect 16942 87278 16994 87330
rect 10670 87166 10722 87218
rect 15598 87166 15650 87218
rect 16046 87166 16098 87218
rect 16942 87166 16994 87218
rect 4024 86998 4076 87050
rect 4148 86998 4200 87050
rect 4272 86998 4324 87050
rect 4396 86998 4448 87050
rect 4520 86998 4572 87050
rect 4644 86998 4696 87050
rect 4768 86998 4820 87050
rect 4892 86998 4944 87050
rect 5016 86998 5068 87050
rect 5140 86998 5192 87050
rect 24024 86998 24076 87050
rect 24148 86998 24200 87050
rect 24272 86998 24324 87050
rect 24396 86998 24448 87050
rect 24520 86998 24572 87050
rect 24644 86998 24696 87050
rect 24768 86998 24820 87050
rect 24892 86998 24944 87050
rect 25016 86998 25068 87050
rect 25140 86998 25192 87050
rect 7646 86830 7698 86882
rect 12238 86830 12290 86882
rect 13022 86830 13074 86882
rect 18398 86830 18450 86882
rect 9998 86718 10050 86770
rect 12014 86718 12066 86770
rect 12910 86718 12962 86770
rect 7982 86606 8034 86658
rect 8766 86606 8818 86658
rect 9326 86606 9378 86658
rect 9886 86606 9938 86658
rect 10334 86606 10386 86658
rect 10894 86606 10946 86658
rect 12462 86606 12514 86658
rect 13582 86606 13634 86658
rect 14366 86606 14418 86658
rect 15038 86606 15090 86658
rect 18734 86606 18786 86658
rect 7310 86494 7362 86546
rect 8542 86494 8594 86546
rect 10222 86494 10274 86546
rect 11902 86494 11954 86546
rect 14030 86494 14082 86546
rect 18958 86494 19010 86546
rect 19406 86494 19458 86546
rect 1710 86382 1762 86434
rect 17278 86382 17330 86434
rect 18062 86382 18114 86434
rect 14024 86214 14076 86266
rect 14148 86214 14200 86266
rect 14272 86214 14324 86266
rect 14396 86214 14448 86266
rect 14520 86214 14572 86266
rect 14644 86214 14696 86266
rect 14768 86214 14820 86266
rect 14892 86214 14944 86266
rect 15016 86214 15068 86266
rect 15140 86214 15192 86266
rect 34024 86214 34076 86266
rect 34148 86214 34200 86266
rect 34272 86214 34324 86266
rect 34396 86214 34448 86266
rect 34520 86214 34572 86266
rect 34644 86214 34696 86266
rect 34768 86214 34820 86266
rect 34892 86214 34944 86266
rect 35016 86214 35068 86266
rect 35140 86214 35192 86266
rect 9662 86046 9714 86098
rect 10222 86046 10274 86098
rect 10782 86046 10834 86098
rect 13582 86046 13634 86098
rect 15374 86046 15426 86098
rect 23102 86046 23154 86098
rect 1710 85934 1762 85986
rect 9998 85934 10050 85986
rect 15710 85934 15762 85986
rect 16606 85934 16658 85986
rect 14142 85822 14194 85874
rect 15038 85822 15090 85874
rect 15374 85822 15426 85874
rect 20078 85822 20130 85874
rect 20638 85822 20690 85874
rect 24558 85822 24610 85874
rect 7422 85710 7474 85762
rect 10334 85710 10386 85762
rect 14814 85710 14866 85762
rect 16158 85710 16210 85762
rect 16494 85710 16546 85762
rect 16830 85710 16882 85762
rect 18174 85710 18226 85762
rect 18622 85710 18674 85762
rect 23662 85710 23714 85762
rect 23998 85710 24050 85762
rect 4024 85430 4076 85482
rect 4148 85430 4200 85482
rect 4272 85430 4324 85482
rect 4396 85430 4448 85482
rect 4520 85430 4572 85482
rect 4644 85430 4696 85482
rect 4768 85430 4820 85482
rect 4892 85430 4944 85482
rect 5016 85430 5068 85482
rect 5140 85430 5192 85482
rect 24024 85430 24076 85482
rect 24148 85430 24200 85482
rect 24272 85430 24324 85482
rect 24396 85430 24448 85482
rect 24520 85430 24572 85482
rect 24644 85430 24696 85482
rect 24768 85430 24820 85482
rect 24892 85430 24944 85482
rect 25016 85430 25068 85482
rect 25140 85430 25192 85482
rect 21422 85262 21474 85314
rect 4846 85150 4898 85202
rect 14366 85150 14418 85202
rect 6526 85038 6578 85090
rect 6974 85038 7026 85090
rect 10782 85038 10834 85090
rect 14254 85038 14306 85090
rect 21758 85038 21810 85090
rect 9214 84926 9266 84978
rect 13918 84926 13970 84978
rect 14478 84926 14530 84978
rect 20750 84926 20802 84978
rect 21982 84926 22034 84978
rect 22542 84926 22594 84978
rect 5854 84814 5906 84866
rect 9998 84814 10050 84866
rect 10334 84814 10386 84866
rect 12574 84814 12626 84866
rect 13022 84814 13074 84866
rect 13694 84814 13746 84866
rect 18174 84814 18226 84866
rect 14024 84646 14076 84698
rect 14148 84646 14200 84698
rect 14272 84646 14324 84698
rect 14396 84646 14448 84698
rect 14520 84646 14572 84698
rect 14644 84646 14696 84698
rect 14768 84646 14820 84698
rect 14892 84646 14944 84698
rect 15016 84646 15068 84698
rect 15140 84646 15192 84698
rect 34024 84646 34076 84698
rect 34148 84646 34200 84698
rect 34272 84646 34324 84698
rect 34396 84646 34448 84698
rect 34520 84646 34572 84698
rect 34644 84646 34696 84698
rect 34768 84646 34820 84698
rect 34892 84646 34944 84698
rect 35016 84646 35068 84698
rect 35140 84646 35192 84698
rect 6750 84478 6802 84530
rect 8318 84478 8370 84530
rect 9662 84478 9714 84530
rect 12238 84478 12290 84530
rect 12686 84478 12738 84530
rect 18734 84478 18786 84530
rect 22094 84478 22146 84530
rect 1710 84366 1762 84418
rect 8542 84366 8594 84418
rect 9774 84366 9826 84418
rect 13358 84366 13410 84418
rect 13582 84366 13634 84418
rect 14478 84366 14530 84418
rect 14590 84366 14642 84418
rect 15038 84366 15090 84418
rect 19294 84366 19346 84418
rect 19630 84366 19682 84418
rect 21086 84366 21138 84418
rect 3838 84254 3890 84306
rect 4174 84254 4226 84306
rect 8094 84254 8146 84306
rect 8766 84254 8818 84306
rect 12574 84254 12626 84306
rect 12798 84254 12850 84306
rect 13246 84254 13298 84306
rect 13694 84254 13746 84306
rect 20526 84254 20578 84306
rect 20974 84254 21026 84306
rect 7870 84142 7922 84194
rect 11790 84142 11842 84194
rect 17502 84142 17554 84194
rect 18286 84142 18338 84194
rect 7310 84030 7362 84082
rect 14478 84030 14530 84082
rect 19070 84030 19122 84082
rect 21758 84030 21810 84082
rect 4024 83862 4076 83914
rect 4148 83862 4200 83914
rect 4272 83862 4324 83914
rect 4396 83862 4448 83914
rect 4520 83862 4572 83914
rect 4644 83862 4696 83914
rect 4768 83862 4820 83914
rect 4892 83862 4944 83914
rect 5016 83862 5068 83914
rect 5140 83862 5192 83914
rect 24024 83862 24076 83914
rect 24148 83862 24200 83914
rect 24272 83862 24324 83914
rect 24396 83862 24448 83914
rect 24520 83862 24572 83914
rect 24644 83862 24696 83914
rect 24768 83862 24820 83914
rect 24892 83862 24944 83914
rect 25016 83862 25068 83914
rect 25140 83862 25192 83914
rect 5966 83694 6018 83746
rect 6302 83694 6354 83746
rect 8766 83694 8818 83746
rect 12126 83694 12178 83746
rect 12574 83582 12626 83634
rect 20302 83582 20354 83634
rect 3726 83470 3778 83522
rect 4286 83470 4338 83522
rect 7086 83470 7138 83522
rect 8766 83470 8818 83522
rect 12462 83470 12514 83522
rect 13470 83470 13522 83522
rect 14030 83470 14082 83522
rect 17614 83470 17666 83522
rect 17838 83470 17890 83522
rect 18286 83470 18338 83522
rect 18958 83470 19010 83522
rect 19182 83470 19234 83522
rect 19406 83470 19458 83522
rect 22990 83470 23042 83522
rect 4510 83358 4562 83410
rect 6862 83358 6914 83410
rect 8206 83358 8258 83410
rect 8430 83358 8482 83410
rect 18398 83358 18450 83410
rect 18734 83358 18786 83410
rect 19070 83358 19122 83410
rect 1710 83246 1762 83298
rect 3390 83246 3442 83298
rect 5070 83246 5122 83298
rect 7646 83246 7698 83298
rect 9214 83246 9266 83298
rect 16494 83246 16546 83298
rect 17054 83246 17106 83298
rect 17502 83246 17554 83298
rect 22542 83246 22594 83298
rect 22654 83246 22706 83298
rect 22878 83246 22930 83298
rect 14024 83078 14076 83130
rect 14148 83078 14200 83130
rect 14272 83078 14324 83130
rect 14396 83078 14448 83130
rect 14520 83078 14572 83130
rect 14644 83078 14696 83130
rect 14768 83078 14820 83130
rect 14892 83078 14944 83130
rect 15016 83078 15068 83130
rect 15140 83078 15192 83130
rect 34024 83078 34076 83130
rect 34148 83078 34200 83130
rect 34272 83078 34324 83130
rect 34396 83078 34448 83130
rect 34520 83078 34572 83130
rect 34644 83078 34696 83130
rect 34768 83078 34820 83130
rect 34892 83078 34944 83130
rect 35016 83078 35068 83130
rect 35140 83078 35192 83130
rect 4734 82910 4786 82962
rect 5294 82910 5346 82962
rect 5630 82910 5682 82962
rect 6190 82910 6242 82962
rect 11118 82910 11170 82962
rect 12910 82910 12962 82962
rect 15934 82910 15986 82962
rect 16718 82910 16770 82962
rect 25342 82910 25394 82962
rect 5518 82798 5570 82850
rect 13022 82798 13074 82850
rect 13582 82798 13634 82850
rect 14366 82798 14418 82850
rect 16270 82798 16322 82850
rect 17390 82798 17442 82850
rect 21870 82798 21922 82850
rect 1822 82686 1874 82738
rect 2270 82686 2322 82738
rect 6302 82686 6354 82738
rect 10670 82686 10722 82738
rect 10894 82686 10946 82738
rect 11342 82686 11394 82738
rect 14142 82686 14194 82738
rect 14478 82686 14530 82738
rect 16494 82686 16546 82738
rect 16830 82686 16882 82738
rect 17614 82686 17666 82738
rect 17838 82686 17890 82738
rect 24110 82686 24162 82738
rect 24558 82686 24610 82738
rect 25790 82686 25842 82738
rect 6750 82574 6802 82626
rect 7198 82574 7250 82626
rect 7646 82574 7698 82626
rect 11230 82574 11282 82626
rect 12574 82574 12626 82626
rect 13358 82574 13410 82626
rect 13694 82574 13746 82626
rect 15486 82574 15538 82626
rect 18846 82574 18898 82626
rect 5630 82462 5682 82514
rect 6190 82462 6242 82514
rect 15486 82462 15538 82514
rect 16046 82462 16098 82514
rect 21086 82462 21138 82514
rect 4024 82294 4076 82346
rect 4148 82294 4200 82346
rect 4272 82294 4324 82346
rect 4396 82294 4448 82346
rect 4520 82294 4572 82346
rect 4644 82294 4696 82346
rect 4768 82294 4820 82346
rect 4892 82294 4944 82346
rect 5016 82294 5068 82346
rect 5140 82294 5192 82346
rect 24024 82294 24076 82346
rect 24148 82294 24200 82346
rect 24272 82294 24324 82346
rect 24396 82294 24448 82346
rect 24520 82294 24572 82346
rect 24644 82294 24696 82346
rect 24768 82294 24820 82346
rect 24892 82294 24944 82346
rect 25016 82294 25068 82346
rect 25140 82294 25192 82346
rect 20638 82126 20690 82178
rect 4510 82014 4562 82066
rect 5966 82014 6018 82066
rect 6414 82014 6466 82066
rect 9438 82014 9490 82066
rect 10446 82014 10498 82066
rect 14478 82014 14530 82066
rect 21422 82014 21474 82066
rect 22430 82014 22482 82066
rect 10110 81902 10162 81954
rect 10334 81902 10386 81954
rect 10558 81902 10610 81954
rect 11118 81902 11170 81954
rect 11342 81902 11394 81954
rect 11454 81902 11506 81954
rect 11790 81902 11842 81954
rect 12126 81902 12178 81954
rect 15038 81902 15090 81954
rect 15262 81902 15314 81954
rect 16158 81902 16210 81954
rect 16270 81902 16322 81954
rect 16606 81902 16658 81954
rect 16942 81902 16994 81954
rect 17502 81902 17554 81954
rect 1710 81790 1762 81842
rect 4846 81790 4898 81842
rect 9886 81790 9938 81842
rect 10894 81790 10946 81842
rect 12350 81790 12402 81842
rect 13694 81790 13746 81842
rect 13806 81790 13858 81842
rect 14814 81790 14866 81842
rect 15486 81790 15538 81842
rect 22766 81790 22818 81842
rect 4398 81678 4450 81730
rect 4622 81678 4674 81730
rect 11230 81678 11282 81730
rect 12462 81678 12514 81730
rect 14702 81678 14754 81730
rect 16382 81678 16434 81730
rect 16494 81678 16546 81730
rect 20078 81678 20130 81730
rect 21982 81678 22034 81730
rect 22318 81678 22370 81730
rect 22542 81678 22594 81730
rect 14024 81510 14076 81562
rect 14148 81510 14200 81562
rect 14272 81510 14324 81562
rect 14396 81510 14448 81562
rect 14520 81510 14572 81562
rect 14644 81510 14696 81562
rect 14768 81510 14820 81562
rect 14892 81510 14944 81562
rect 15016 81510 15068 81562
rect 15140 81510 15192 81562
rect 34024 81510 34076 81562
rect 34148 81510 34200 81562
rect 34272 81510 34324 81562
rect 34396 81510 34448 81562
rect 34520 81510 34572 81562
rect 34644 81510 34696 81562
rect 34768 81510 34820 81562
rect 34892 81510 34944 81562
rect 35016 81510 35068 81562
rect 35140 81510 35192 81562
rect 15374 81342 15426 81394
rect 1710 81230 1762 81282
rect 8318 81230 8370 81282
rect 10894 81230 10946 81282
rect 15262 81230 15314 81282
rect 15934 81230 15986 81282
rect 5630 81118 5682 81170
rect 6078 81118 6130 81170
rect 9662 81118 9714 81170
rect 10334 81118 10386 81170
rect 10446 81118 10498 81170
rect 10558 81118 10610 81170
rect 11678 81118 11730 81170
rect 11902 81118 11954 81170
rect 12350 81118 12402 81170
rect 14814 81118 14866 81170
rect 15038 81118 15090 81170
rect 15486 81118 15538 81170
rect 16046 81118 16098 81170
rect 16494 81118 16546 81170
rect 16718 81118 16770 81170
rect 17390 81118 17442 81170
rect 18286 81118 18338 81170
rect 19294 81118 19346 81170
rect 22542 81118 22594 81170
rect 5182 81006 5234 81058
rect 9886 81006 9938 81058
rect 12126 81006 12178 81058
rect 13470 81006 13522 81058
rect 13918 81006 13970 81058
rect 14366 81006 14418 81058
rect 16270 81006 16322 81058
rect 18062 81006 18114 81058
rect 19182 81006 19234 81058
rect 20078 81006 20130 81058
rect 20526 81006 20578 81058
rect 22206 81006 22258 81058
rect 22318 81006 22370 81058
rect 23662 81006 23714 81058
rect 9102 80894 9154 80946
rect 11118 80894 11170 80946
rect 11230 80894 11282 80946
rect 12798 80894 12850 80946
rect 18958 80894 19010 80946
rect 4024 80726 4076 80778
rect 4148 80726 4200 80778
rect 4272 80726 4324 80778
rect 4396 80726 4448 80778
rect 4520 80726 4572 80778
rect 4644 80726 4696 80778
rect 4768 80726 4820 80778
rect 4892 80726 4944 80778
rect 5016 80726 5068 80778
rect 5140 80726 5192 80778
rect 24024 80726 24076 80778
rect 24148 80726 24200 80778
rect 24272 80726 24324 80778
rect 24396 80726 24448 80778
rect 24520 80726 24572 80778
rect 24644 80726 24696 80778
rect 24768 80726 24820 80778
rect 24892 80726 24944 80778
rect 25016 80726 25068 80778
rect 25140 80726 25192 80778
rect 5966 80558 6018 80610
rect 6078 80558 6130 80610
rect 6750 80558 6802 80610
rect 6974 80558 7026 80610
rect 7758 80558 7810 80610
rect 7982 80558 8034 80610
rect 10334 80558 10386 80610
rect 15150 80558 15202 80610
rect 19406 80558 19458 80610
rect 9774 80446 9826 80498
rect 10110 80446 10162 80498
rect 11678 80446 11730 80498
rect 19966 80446 20018 80498
rect 6078 80334 6130 80386
rect 6526 80334 6578 80386
rect 7310 80334 7362 80386
rect 9886 80334 9938 80386
rect 11902 80334 11954 80386
rect 14142 80334 14194 80386
rect 14478 80334 14530 80386
rect 14590 80334 14642 80386
rect 14702 80334 14754 80386
rect 15822 80334 15874 80386
rect 16270 80334 16322 80386
rect 8318 80222 8370 80274
rect 8654 80222 8706 80274
rect 8766 80222 8818 80274
rect 9214 80222 9266 80274
rect 11230 80222 11282 80274
rect 13806 80222 13858 80274
rect 1710 80110 1762 80162
rect 8094 80110 8146 80162
rect 9662 80110 9714 80162
rect 11454 80110 11506 80162
rect 11678 80110 11730 80162
rect 12910 80110 12962 80162
rect 13918 80110 13970 80162
rect 18846 80110 18898 80162
rect 14024 79942 14076 79994
rect 14148 79942 14200 79994
rect 14272 79942 14324 79994
rect 14396 79942 14448 79994
rect 14520 79942 14572 79994
rect 14644 79942 14696 79994
rect 14768 79942 14820 79994
rect 14892 79942 14944 79994
rect 15016 79942 15068 79994
rect 15140 79942 15192 79994
rect 34024 79942 34076 79994
rect 34148 79942 34200 79994
rect 34272 79942 34324 79994
rect 34396 79942 34448 79994
rect 34520 79942 34572 79994
rect 34644 79942 34696 79994
rect 34768 79942 34820 79994
rect 34892 79942 34944 79994
rect 35016 79942 35068 79994
rect 35140 79942 35192 79994
rect 4734 79774 4786 79826
rect 5854 79774 5906 79826
rect 6302 79774 6354 79826
rect 6750 79774 6802 79826
rect 17502 79774 17554 79826
rect 7422 79662 7474 79714
rect 7534 79662 7586 79714
rect 14142 79662 14194 79714
rect 15150 79662 15202 79714
rect 1822 79550 1874 79602
rect 2270 79550 2322 79602
rect 5406 79550 5458 79602
rect 8318 79550 8370 79602
rect 8654 79550 8706 79602
rect 11006 79550 11058 79602
rect 11566 79550 11618 79602
rect 12014 79550 12066 79602
rect 13022 79550 13074 79602
rect 13246 79550 13298 79602
rect 13694 79550 13746 79602
rect 15262 79550 15314 79602
rect 22094 79550 22146 79602
rect 13806 79438 13858 79490
rect 20638 79438 20690 79490
rect 20974 79438 21026 79490
rect 22206 79438 22258 79490
rect 22654 79438 22706 79490
rect 7982 79326 8034 79378
rect 12910 79326 12962 79378
rect 20638 79326 20690 79378
rect 21422 79326 21474 79378
rect 4024 79158 4076 79210
rect 4148 79158 4200 79210
rect 4272 79158 4324 79210
rect 4396 79158 4448 79210
rect 4520 79158 4572 79210
rect 4644 79158 4696 79210
rect 4768 79158 4820 79210
rect 4892 79158 4944 79210
rect 5016 79158 5068 79210
rect 5140 79158 5192 79210
rect 24024 79158 24076 79210
rect 24148 79158 24200 79210
rect 24272 79158 24324 79210
rect 24396 79158 24448 79210
rect 24520 79158 24572 79210
rect 24644 79158 24696 79210
rect 24768 79158 24820 79210
rect 24892 79158 24944 79210
rect 25016 79158 25068 79210
rect 25140 79158 25192 79210
rect 3278 78990 3330 79042
rect 13918 78990 13970 79042
rect 3390 78878 3442 78930
rect 4510 78878 4562 78930
rect 6526 78878 6578 78930
rect 12014 78878 12066 78930
rect 15934 78878 15986 78930
rect 19966 78878 20018 78930
rect 23326 78878 23378 78930
rect 4622 78766 4674 78818
rect 6078 78766 6130 78818
rect 7534 78766 7586 78818
rect 8206 78766 8258 78818
rect 11230 78766 11282 78818
rect 11566 78766 11618 78818
rect 13918 78766 13970 78818
rect 14254 78766 14306 78818
rect 15598 78766 15650 78818
rect 16046 78766 16098 78818
rect 20302 78766 20354 78818
rect 22206 78766 22258 78818
rect 5070 78654 5122 78706
rect 5630 78654 5682 78706
rect 13582 78654 13634 78706
rect 15486 78654 15538 78706
rect 16270 78654 16322 78706
rect 20750 78654 20802 78706
rect 21422 78654 21474 78706
rect 21870 78654 21922 78706
rect 22990 78654 23042 78706
rect 23214 78654 23266 78706
rect 1710 78542 1762 78594
rect 4174 78542 4226 78594
rect 4510 78542 4562 78594
rect 4846 78542 4898 78594
rect 7086 78542 7138 78594
rect 10670 78542 10722 78594
rect 11454 78542 11506 78594
rect 22542 78542 22594 78594
rect 14024 78374 14076 78426
rect 14148 78374 14200 78426
rect 14272 78374 14324 78426
rect 14396 78374 14448 78426
rect 14520 78374 14572 78426
rect 14644 78374 14696 78426
rect 14768 78374 14820 78426
rect 14892 78374 14944 78426
rect 15016 78374 15068 78426
rect 15140 78374 15192 78426
rect 34024 78374 34076 78426
rect 34148 78374 34200 78426
rect 34272 78374 34324 78426
rect 34396 78374 34448 78426
rect 34520 78374 34572 78426
rect 34644 78374 34696 78426
rect 34768 78374 34820 78426
rect 34892 78374 34944 78426
rect 35016 78374 35068 78426
rect 35140 78374 35192 78426
rect 4734 78206 4786 78258
rect 5294 78206 5346 78258
rect 9886 78206 9938 78258
rect 15262 78206 15314 78258
rect 20302 78206 20354 78258
rect 20974 78206 21026 78258
rect 24334 78206 24386 78258
rect 25342 78206 25394 78258
rect 6190 78094 6242 78146
rect 6750 78094 6802 78146
rect 7310 78094 7362 78146
rect 8878 78094 8930 78146
rect 1822 77982 1874 78034
rect 2270 77982 2322 78034
rect 5966 77982 6018 78034
rect 7198 77982 7250 78034
rect 7758 77982 7810 78034
rect 9550 77982 9602 78034
rect 9886 77982 9938 78034
rect 10110 77982 10162 78034
rect 10558 77982 10610 78034
rect 12462 77982 12514 78034
rect 15150 77982 15202 78034
rect 15374 77982 15426 78034
rect 15822 77982 15874 78034
rect 23326 77982 23378 78034
rect 23886 77982 23938 78034
rect 8318 77870 8370 77922
rect 8990 77870 9042 77922
rect 11342 77870 11394 77922
rect 13582 77870 13634 77922
rect 15598 77870 15650 77922
rect 16382 77870 16434 77922
rect 5630 77758 5682 77810
rect 7310 77758 7362 77810
rect 7870 77758 7922 77810
rect 8654 77758 8706 77810
rect 4024 77590 4076 77642
rect 4148 77590 4200 77642
rect 4272 77590 4324 77642
rect 4396 77590 4448 77642
rect 4520 77590 4572 77642
rect 4644 77590 4696 77642
rect 4768 77590 4820 77642
rect 4892 77590 4944 77642
rect 5016 77590 5068 77642
rect 5140 77590 5192 77642
rect 24024 77590 24076 77642
rect 24148 77590 24200 77642
rect 24272 77590 24324 77642
rect 24396 77590 24448 77642
rect 24520 77590 24572 77642
rect 24644 77590 24696 77642
rect 24768 77590 24820 77642
rect 24892 77590 24944 77642
rect 25016 77590 25068 77642
rect 25140 77590 25192 77642
rect 3278 77422 3330 77474
rect 3614 77422 3666 77474
rect 25678 77310 25730 77362
rect 5070 77198 5122 77250
rect 5742 77198 5794 77250
rect 6638 77198 6690 77250
rect 6974 77198 7026 77250
rect 9662 77198 9714 77250
rect 10110 77198 10162 77250
rect 13806 77198 13858 77250
rect 14590 77198 14642 77250
rect 15486 77198 15538 77250
rect 21198 77198 21250 77250
rect 24222 77198 24274 77250
rect 24782 77198 24834 77250
rect 25230 77198 25282 77250
rect 1710 77086 1762 77138
rect 3838 77086 3890 77138
rect 4286 77086 4338 77138
rect 5966 77086 6018 77138
rect 6302 77086 6354 77138
rect 6750 77086 6802 77138
rect 7982 77086 8034 77138
rect 10558 77086 10610 77138
rect 14702 77086 14754 77138
rect 15374 77086 15426 77138
rect 21982 77086 22034 77138
rect 6078 76974 6130 77026
rect 7534 76974 7586 77026
rect 8430 76974 8482 77026
rect 15150 76974 15202 77026
rect 14024 76806 14076 76858
rect 14148 76806 14200 76858
rect 14272 76806 14324 76858
rect 14396 76806 14448 76858
rect 14520 76806 14572 76858
rect 14644 76806 14696 76858
rect 14768 76806 14820 76858
rect 14892 76806 14944 76858
rect 15016 76806 15068 76858
rect 15140 76806 15192 76858
rect 34024 76806 34076 76858
rect 34148 76806 34200 76858
rect 34272 76806 34324 76858
rect 34396 76806 34448 76858
rect 34520 76806 34572 76858
rect 34644 76806 34696 76858
rect 34768 76806 34820 76858
rect 34892 76806 34944 76858
rect 35016 76806 35068 76858
rect 35140 76806 35192 76858
rect 4734 76638 4786 76690
rect 5406 76638 5458 76690
rect 9774 76638 9826 76690
rect 13806 76638 13858 76690
rect 16830 76638 16882 76690
rect 18734 76638 18786 76690
rect 20302 76638 20354 76690
rect 22318 76638 22370 76690
rect 1710 76526 1762 76578
rect 14590 76526 14642 76578
rect 15262 76526 15314 76578
rect 15822 76526 15874 76578
rect 17390 76526 17442 76578
rect 17726 76526 17778 76578
rect 21310 76526 21362 76578
rect 21758 76526 21810 76578
rect 11118 76414 11170 76466
rect 11566 76414 11618 76466
rect 15934 76414 15986 76466
rect 16382 76414 16434 76466
rect 17838 76414 17890 76466
rect 18398 76414 18450 76466
rect 18846 76414 18898 76466
rect 21982 76414 22034 76466
rect 6526 76302 6578 76354
rect 10222 76302 10274 76354
rect 10670 76302 10722 76354
rect 14702 76302 14754 76354
rect 17502 76302 17554 76354
rect 18286 76302 18338 76354
rect 20750 76302 20802 76354
rect 4024 76022 4076 76074
rect 4148 76022 4200 76074
rect 4272 76022 4324 76074
rect 4396 76022 4448 76074
rect 4520 76022 4572 76074
rect 4644 76022 4696 76074
rect 4768 76022 4820 76074
rect 4892 76022 4944 76074
rect 5016 76022 5068 76074
rect 5140 76022 5192 76074
rect 24024 76022 24076 76074
rect 24148 76022 24200 76074
rect 24272 76022 24324 76074
rect 24396 76022 24448 76074
rect 24520 76022 24572 76074
rect 24644 76022 24696 76074
rect 24768 76022 24820 76074
rect 24892 76022 24944 76074
rect 25016 76022 25068 76074
rect 25140 76022 25192 76074
rect 11006 75854 11058 75906
rect 11678 75854 11730 75906
rect 12014 75854 12066 75906
rect 20190 75854 20242 75906
rect 4398 75742 4450 75794
rect 5854 75742 5906 75794
rect 6750 75742 6802 75794
rect 9662 75742 9714 75794
rect 14478 75742 14530 75794
rect 14926 75742 14978 75794
rect 15374 75742 15426 75794
rect 5630 75630 5682 75682
rect 6078 75630 6130 75682
rect 6302 75630 6354 75682
rect 8542 75630 8594 75682
rect 10894 75630 10946 75682
rect 12798 75630 12850 75682
rect 15710 75630 15762 75682
rect 16046 75630 16098 75682
rect 16494 75630 16546 75682
rect 17166 75630 17218 75682
rect 5854 75518 5906 75570
rect 12574 75518 12626 75570
rect 16270 75518 16322 75570
rect 1710 75406 1762 75458
rect 4286 75406 4338 75458
rect 15934 75406 15986 75458
rect 19406 75406 19458 75458
rect 20526 75406 20578 75458
rect 14024 75238 14076 75290
rect 14148 75238 14200 75290
rect 14272 75238 14324 75290
rect 14396 75238 14448 75290
rect 14520 75238 14572 75290
rect 14644 75238 14696 75290
rect 14768 75238 14820 75290
rect 14892 75238 14944 75290
rect 15016 75238 15068 75290
rect 15140 75238 15192 75290
rect 34024 75238 34076 75290
rect 34148 75238 34200 75290
rect 34272 75238 34324 75290
rect 34396 75238 34448 75290
rect 34520 75238 34572 75290
rect 34644 75238 34696 75290
rect 34768 75238 34820 75290
rect 34892 75238 34944 75290
rect 35016 75238 35068 75290
rect 35140 75238 35192 75290
rect 6078 75070 6130 75122
rect 6974 75070 7026 75122
rect 8878 75070 8930 75122
rect 13358 75070 13410 75122
rect 14254 75070 14306 75122
rect 15710 75070 15762 75122
rect 16158 75070 16210 75122
rect 17838 75070 17890 75122
rect 9886 74958 9938 75010
rect 9998 74958 10050 75010
rect 11678 74958 11730 75010
rect 12686 74958 12738 75010
rect 16606 74958 16658 75010
rect 16830 74958 16882 75010
rect 17726 74958 17778 75010
rect 17950 74958 18002 75010
rect 3166 74846 3218 74898
rect 3614 74846 3666 74898
rect 7982 74846 8034 74898
rect 8990 74846 9042 74898
rect 10222 74846 10274 74898
rect 10782 74846 10834 74898
rect 12238 74846 12290 74898
rect 12910 74846 12962 74898
rect 14366 74846 14418 74898
rect 7422 74734 7474 74786
rect 8542 74734 8594 74786
rect 10894 74734 10946 74786
rect 12462 74734 12514 74786
rect 15262 74734 15314 74786
rect 16494 74734 16546 74786
rect 18510 74734 18562 74786
rect 6638 74622 6690 74674
rect 7422 74622 7474 74674
rect 8318 74622 8370 74674
rect 8878 74622 8930 74674
rect 15262 74622 15314 74674
rect 16158 74622 16210 74674
rect 4024 74454 4076 74506
rect 4148 74454 4200 74506
rect 4272 74454 4324 74506
rect 4396 74454 4448 74506
rect 4520 74454 4572 74506
rect 4644 74454 4696 74506
rect 4768 74454 4820 74506
rect 4892 74454 4944 74506
rect 5016 74454 5068 74506
rect 5140 74454 5192 74506
rect 24024 74454 24076 74506
rect 24148 74454 24200 74506
rect 24272 74454 24324 74506
rect 24396 74454 24448 74506
rect 24520 74454 24572 74506
rect 24644 74454 24696 74506
rect 24768 74454 24820 74506
rect 24892 74454 24944 74506
rect 25016 74454 25068 74506
rect 25140 74454 25192 74506
rect 10894 74286 10946 74338
rect 12574 74286 12626 74338
rect 12910 74286 12962 74338
rect 19518 74286 19570 74338
rect 5742 74174 5794 74226
rect 6190 74174 6242 74226
rect 6638 74174 6690 74226
rect 11230 74174 11282 74226
rect 11790 74174 11842 74226
rect 3838 74062 3890 74114
rect 7198 74062 7250 74114
rect 7870 74062 7922 74114
rect 12238 74062 12290 74114
rect 15822 74062 15874 74114
rect 16382 74062 16434 74114
rect 3502 73950 3554 74002
rect 4062 73950 4114 74002
rect 4622 73950 4674 74002
rect 12798 73950 12850 74002
rect 1710 73838 1762 73890
rect 2158 73838 2210 73890
rect 10110 73838 10162 73890
rect 15598 73838 15650 73890
rect 18734 73838 18786 73890
rect 19854 73838 19906 73890
rect 14024 73670 14076 73722
rect 14148 73670 14200 73722
rect 14272 73670 14324 73722
rect 14396 73670 14448 73722
rect 14520 73670 14572 73722
rect 14644 73670 14696 73722
rect 14768 73670 14820 73722
rect 14892 73670 14944 73722
rect 15016 73670 15068 73722
rect 15140 73670 15192 73722
rect 34024 73670 34076 73722
rect 34148 73670 34200 73722
rect 34272 73670 34324 73722
rect 34396 73670 34448 73722
rect 34520 73670 34572 73722
rect 34644 73670 34696 73722
rect 34768 73670 34820 73722
rect 34892 73670 34944 73722
rect 35016 73670 35068 73722
rect 35140 73670 35192 73722
rect 4734 73502 4786 73554
rect 5294 73502 5346 73554
rect 9102 73502 9154 73554
rect 9662 73502 9714 73554
rect 14366 73502 14418 73554
rect 15150 73502 15202 73554
rect 15934 73502 15986 73554
rect 8318 73390 8370 73442
rect 20638 73390 20690 73442
rect 1822 73278 1874 73330
rect 2270 73278 2322 73330
rect 5630 73278 5682 73330
rect 6078 73278 6130 73330
rect 9550 73278 9602 73330
rect 9774 73278 9826 73330
rect 10222 73278 10274 73330
rect 11006 73278 11058 73330
rect 11454 73278 11506 73330
rect 12126 73278 12178 73330
rect 22878 73278 22930 73330
rect 23438 73278 23490 73330
rect 10558 73166 10610 73218
rect 15486 73166 15538 73218
rect 23886 73166 23938 73218
rect 24334 73166 24386 73218
rect 10782 73054 10834 73106
rect 11342 73054 11394 73106
rect 19854 73054 19906 73106
rect 4024 72886 4076 72938
rect 4148 72886 4200 72938
rect 4272 72886 4324 72938
rect 4396 72886 4448 72938
rect 4520 72886 4572 72938
rect 4644 72886 4696 72938
rect 4768 72886 4820 72938
rect 4892 72886 4944 72938
rect 5016 72886 5068 72938
rect 5140 72886 5192 72938
rect 24024 72886 24076 72938
rect 24148 72886 24200 72938
rect 24272 72886 24324 72938
rect 24396 72886 24448 72938
rect 24520 72886 24572 72938
rect 24644 72886 24696 72938
rect 24768 72886 24820 72938
rect 24892 72886 24944 72938
rect 25016 72886 25068 72938
rect 25140 72886 25192 72938
rect 3838 72718 3890 72770
rect 21534 72718 21586 72770
rect 7758 72606 7810 72658
rect 9550 72606 9602 72658
rect 4174 72494 4226 72546
rect 4734 72494 4786 72546
rect 5966 72494 6018 72546
rect 6078 72494 6130 72546
rect 7870 72494 7922 72546
rect 23550 72494 23602 72546
rect 4958 72382 5010 72434
rect 8094 72382 8146 72434
rect 1710 72270 1762 72322
rect 7646 72270 7698 72322
rect 8654 72270 8706 72322
rect 9886 72270 9938 72322
rect 24334 72270 24386 72322
rect 14024 72102 14076 72154
rect 14148 72102 14200 72154
rect 14272 72102 14324 72154
rect 14396 72102 14448 72154
rect 14520 72102 14572 72154
rect 14644 72102 14696 72154
rect 14768 72102 14820 72154
rect 14892 72102 14944 72154
rect 15016 72102 15068 72154
rect 15140 72102 15192 72154
rect 34024 72102 34076 72154
rect 34148 72102 34200 72154
rect 34272 72102 34324 72154
rect 34396 72102 34448 72154
rect 34520 72102 34572 72154
rect 34644 72102 34696 72154
rect 34768 72102 34820 72154
rect 34892 72102 34944 72154
rect 35016 72102 35068 72154
rect 35140 72102 35192 72154
rect 18286 71934 18338 71986
rect 21758 71934 21810 71986
rect 35534 71934 35586 71986
rect 22318 71822 22370 71874
rect 22654 71822 22706 71874
rect 20750 71710 20802 71762
rect 21198 71710 21250 71762
rect 27806 71710 27858 71762
rect 35870 71710 35922 71762
rect 36094 71710 36146 71762
rect 36318 71710 36370 71762
rect 5294 71598 5346 71650
rect 23438 71598 23490 71650
rect 27470 71598 27522 71650
rect 30158 71598 30210 71650
rect 35086 71598 35138 71650
rect 35982 71598 36034 71650
rect 17726 71486 17778 71538
rect 22094 71486 22146 71538
rect 34974 71486 35026 71538
rect 4024 71318 4076 71370
rect 4148 71318 4200 71370
rect 4272 71318 4324 71370
rect 4396 71318 4448 71370
rect 4520 71318 4572 71370
rect 4644 71318 4696 71370
rect 4768 71318 4820 71370
rect 4892 71318 4944 71370
rect 5016 71318 5068 71370
rect 5140 71318 5192 71370
rect 24024 71318 24076 71370
rect 24148 71318 24200 71370
rect 24272 71318 24324 71370
rect 24396 71318 24448 71370
rect 24520 71318 24572 71370
rect 24644 71318 24696 71370
rect 24768 71318 24820 71370
rect 24892 71318 24944 71370
rect 25016 71318 25068 71370
rect 25140 71318 25192 71370
rect 20302 71150 20354 71202
rect 21534 71150 21586 71202
rect 22318 71150 22370 71202
rect 14814 71038 14866 71090
rect 15262 71038 15314 71090
rect 16046 71038 16098 71090
rect 22318 71038 22370 71090
rect 25678 71038 25730 71090
rect 19294 70926 19346 70978
rect 19966 70926 20018 70978
rect 21422 70926 21474 70978
rect 24222 70926 24274 70978
rect 25118 70926 25170 70978
rect 32398 70926 32450 70978
rect 32622 70926 32674 70978
rect 33070 70926 33122 70978
rect 33518 70926 33570 70978
rect 2830 70814 2882 70866
rect 3166 70814 3218 70866
rect 19406 70814 19458 70866
rect 1710 70702 1762 70754
rect 2606 70702 2658 70754
rect 11118 70702 11170 70754
rect 21870 70702 21922 70754
rect 31838 70702 31890 70754
rect 32062 70702 32114 70754
rect 35758 70702 35810 70754
rect 36542 70702 36594 70754
rect 14024 70534 14076 70586
rect 14148 70534 14200 70586
rect 14272 70534 14324 70586
rect 14396 70534 14448 70586
rect 14520 70534 14572 70586
rect 14644 70534 14696 70586
rect 14768 70534 14820 70586
rect 14892 70534 14944 70586
rect 15016 70534 15068 70586
rect 15140 70534 15192 70586
rect 34024 70534 34076 70586
rect 34148 70534 34200 70586
rect 34272 70534 34324 70586
rect 34396 70534 34448 70586
rect 34520 70534 34572 70586
rect 34644 70534 34696 70586
rect 34768 70534 34820 70586
rect 34892 70534 34944 70586
rect 35016 70534 35068 70586
rect 35140 70534 35192 70586
rect 7982 70366 8034 70418
rect 13582 70366 13634 70418
rect 15150 70366 15202 70418
rect 16606 70366 16658 70418
rect 33182 70366 33234 70418
rect 1710 70254 1762 70306
rect 9662 70254 9714 70306
rect 16046 70254 16098 70306
rect 18174 70254 18226 70306
rect 18622 70254 18674 70306
rect 33406 70254 33458 70306
rect 36654 70254 36706 70306
rect 7758 70142 7810 70194
rect 8430 70142 8482 70194
rect 9438 70142 9490 70194
rect 9774 70142 9826 70194
rect 10782 70142 10834 70194
rect 11230 70142 11282 70194
rect 15598 70142 15650 70194
rect 15934 70142 15986 70194
rect 16270 70142 16322 70194
rect 16718 70142 16770 70194
rect 17502 70142 17554 70194
rect 17726 70142 17778 70194
rect 18510 70142 18562 70194
rect 25118 70142 25170 70194
rect 25566 70142 25618 70194
rect 25790 70142 25842 70194
rect 26350 70142 26402 70194
rect 27134 70142 27186 70194
rect 27918 70142 27970 70194
rect 31614 70142 31666 70194
rect 32062 70142 32114 70194
rect 33854 70142 33906 70194
rect 34414 70142 34466 70194
rect 37550 70142 37602 70194
rect 37886 70142 37938 70194
rect 38110 70142 38162 70194
rect 7422 70030 7474 70082
rect 7870 70030 7922 70082
rect 8990 70030 9042 70082
rect 10334 70030 10386 70082
rect 19406 70030 19458 70082
rect 24670 70030 24722 70082
rect 25342 70030 25394 70082
rect 26462 70030 26514 70082
rect 29822 70030 29874 70082
rect 31166 70030 31218 70082
rect 32510 70030 32562 70082
rect 33070 70030 33122 70082
rect 37774 70030 37826 70082
rect 14254 69918 14306 69970
rect 15486 69918 15538 69970
rect 16830 69918 16882 69970
rect 31502 69918 31554 69970
rect 31838 69918 31890 69970
rect 37438 69918 37490 69970
rect 4024 69750 4076 69802
rect 4148 69750 4200 69802
rect 4272 69750 4324 69802
rect 4396 69750 4448 69802
rect 4520 69750 4572 69802
rect 4644 69750 4696 69802
rect 4768 69750 4820 69802
rect 4892 69750 4944 69802
rect 5016 69750 5068 69802
rect 5140 69750 5192 69802
rect 24024 69750 24076 69802
rect 24148 69750 24200 69802
rect 24272 69750 24324 69802
rect 24396 69750 24448 69802
rect 24520 69750 24572 69802
rect 24644 69750 24696 69802
rect 24768 69750 24820 69802
rect 24892 69750 24944 69802
rect 25016 69750 25068 69802
rect 25140 69750 25192 69802
rect 11678 69582 11730 69634
rect 12014 69582 12066 69634
rect 27582 69582 27634 69634
rect 29150 69582 29202 69634
rect 29822 69582 29874 69634
rect 33742 69582 33794 69634
rect 34638 69582 34690 69634
rect 34974 69582 35026 69634
rect 35534 69582 35586 69634
rect 14926 69470 14978 69522
rect 17502 69470 17554 69522
rect 29262 69470 29314 69522
rect 29822 69470 29874 69522
rect 6974 69358 7026 69410
rect 7422 69358 7474 69410
rect 10558 69358 10610 69410
rect 13358 69358 13410 69410
rect 13806 69358 13858 69410
rect 16942 69358 16994 69410
rect 17390 69358 17442 69410
rect 18398 69358 18450 69410
rect 18958 69358 19010 69410
rect 23886 69358 23938 69410
rect 24558 69358 24610 69410
rect 30158 69358 30210 69410
rect 30718 69358 30770 69410
rect 34750 69358 34802 69410
rect 35198 69358 35250 69410
rect 36094 69358 36146 69410
rect 36318 69358 36370 69410
rect 12238 69246 12290 69298
rect 12574 69246 12626 69298
rect 14030 69246 14082 69298
rect 14814 69246 14866 69298
rect 15038 69246 15090 69298
rect 15598 69246 15650 69298
rect 16046 69246 16098 69298
rect 16382 69246 16434 69298
rect 17950 69246 18002 69298
rect 18510 69246 18562 69298
rect 18734 69246 18786 69298
rect 27918 69246 27970 69298
rect 28366 69246 28418 69298
rect 35982 69246 36034 69298
rect 5742 69134 5794 69186
rect 6190 69134 6242 69186
rect 9886 69134 9938 69186
rect 11230 69134 11282 69186
rect 13582 69134 13634 69186
rect 15486 69134 15538 69186
rect 15822 69134 15874 69186
rect 19406 69134 19458 69186
rect 19742 69134 19794 69186
rect 27022 69134 27074 69186
rect 27806 69134 27858 69186
rect 33182 69134 33234 69186
rect 34302 69134 34354 69186
rect 14024 68966 14076 69018
rect 14148 68966 14200 69018
rect 14272 68966 14324 69018
rect 14396 68966 14448 69018
rect 14520 68966 14572 69018
rect 14644 68966 14696 69018
rect 14768 68966 14820 69018
rect 14892 68966 14944 69018
rect 15016 68966 15068 69018
rect 15140 68966 15192 69018
rect 34024 68966 34076 69018
rect 34148 68966 34200 69018
rect 34272 68966 34324 69018
rect 34396 68966 34448 69018
rect 34520 68966 34572 69018
rect 34644 68966 34696 69018
rect 34768 68966 34820 69018
rect 34892 68966 34944 69018
rect 35016 68966 35068 69018
rect 35140 68966 35192 69018
rect 6190 68798 6242 68850
rect 7198 68798 7250 68850
rect 10446 68798 10498 68850
rect 11790 68798 11842 68850
rect 15374 68798 15426 68850
rect 15934 68798 15986 68850
rect 18286 68798 18338 68850
rect 19070 68798 19122 68850
rect 28254 68798 28306 68850
rect 28814 68798 28866 68850
rect 29150 68798 29202 68850
rect 30830 68798 30882 68850
rect 35646 68798 35698 68850
rect 35982 68798 36034 68850
rect 1710 68686 1762 68738
rect 11678 68686 11730 68738
rect 11902 68686 11954 68738
rect 19742 68686 19794 68738
rect 19966 68686 20018 68738
rect 3278 68574 3330 68626
rect 3726 68574 3778 68626
rect 12238 68574 12290 68626
rect 12910 68574 12962 68626
rect 16494 68574 16546 68626
rect 17502 68574 17554 68626
rect 17726 68574 17778 68626
rect 18174 68574 18226 68626
rect 18398 68574 18450 68626
rect 18734 68574 18786 68626
rect 19182 68574 19234 68626
rect 19406 68574 19458 68626
rect 20638 68574 20690 68626
rect 23774 68574 23826 68626
rect 23998 68574 24050 68626
rect 24222 68574 24274 68626
rect 24446 68574 24498 68626
rect 24670 68574 24722 68626
rect 25342 68574 25394 68626
rect 25678 68574 25730 68626
rect 31054 68574 31106 68626
rect 31390 68574 31442 68626
rect 35534 68574 35586 68626
rect 35758 68574 35810 68626
rect 7646 68462 7698 68514
rect 9998 68462 10050 68514
rect 10894 68462 10946 68514
rect 11454 68462 11506 68514
rect 16718 68462 16770 68514
rect 17950 68462 18002 68514
rect 20078 68462 20130 68514
rect 30382 68462 30434 68514
rect 6862 68350 6914 68402
rect 16158 68350 16210 68402
rect 20750 68350 20802 68402
rect 30718 68350 30770 68402
rect 4024 68182 4076 68234
rect 4148 68182 4200 68234
rect 4272 68182 4324 68234
rect 4396 68182 4448 68234
rect 4520 68182 4572 68234
rect 4644 68182 4696 68234
rect 4768 68182 4820 68234
rect 4892 68182 4944 68234
rect 5016 68182 5068 68234
rect 5140 68182 5192 68234
rect 24024 68182 24076 68234
rect 24148 68182 24200 68234
rect 24272 68182 24324 68234
rect 24396 68182 24448 68234
rect 24520 68182 24572 68234
rect 24644 68182 24696 68234
rect 24768 68182 24820 68234
rect 24892 68182 24944 68234
rect 25016 68182 25068 68234
rect 25140 68182 25192 68234
rect 8318 68014 8370 68066
rect 8542 68014 8594 68066
rect 8766 68014 8818 68066
rect 21422 68014 21474 68066
rect 26686 68014 26738 68066
rect 31838 68014 31890 68066
rect 7982 67902 8034 67954
rect 8766 67902 8818 67954
rect 14814 67902 14866 67954
rect 26798 67902 26850 67954
rect 27582 67902 27634 67954
rect 29822 67902 29874 67954
rect 34974 67902 35026 67954
rect 35422 67902 35474 67954
rect 3054 67790 3106 67842
rect 4174 67790 4226 67842
rect 4958 67790 5010 67842
rect 14478 67790 14530 67842
rect 15262 67790 15314 67842
rect 17390 67790 17442 67842
rect 20638 67790 20690 67842
rect 24446 67790 24498 67842
rect 25118 67790 25170 67842
rect 25566 67790 25618 67842
rect 26014 67790 26066 67842
rect 26462 67790 26514 67842
rect 31166 67790 31218 67842
rect 31390 67790 31442 67842
rect 32174 67790 32226 67842
rect 35646 67790 35698 67842
rect 35870 67790 35922 67842
rect 37102 67790 37154 67842
rect 37326 67790 37378 67842
rect 4734 67678 4786 67730
rect 5854 67678 5906 67730
rect 5966 67678 6018 67730
rect 6302 67678 6354 67730
rect 14030 67678 14082 67730
rect 14254 67678 14306 67730
rect 16494 67678 16546 67730
rect 17950 67678 18002 67730
rect 22206 67678 22258 67730
rect 29374 67678 29426 67730
rect 30158 67678 30210 67730
rect 30494 67678 30546 67730
rect 32398 67678 32450 67730
rect 35310 67678 35362 67730
rect 36990 67678 37042 67730
rect 1710 67566 1762 67618
rect 3502 67566 3554 67618
rect 3838 67566 3890 67618
rect 5630 67566 5682 67618
rect 6414 67566 6466 67618
rect 6638 67566 6690 67618
rect 6974 67566 7026 67618
rect 7758 67566 7810 67618
rect 8094 67566 8146 67618
rect 9438 67566 9490 67618
rect 9886 67566 9938 67618
rect 11230 67566 11282 67618
rect 14702 67566 14754 67618
rect 14814 67566 14866 67618
rect 17614 67566 17666 67618
rect 19630 67566 19682 67618
rect 19966 67566 20018 67618
rect 20078 67566 20130 67618
rect 20190 67566 20242 67618
rect 29486 67566 29538 67618
rect 29934 67566 29986 67618
rect 32958 67566 33010 67618
rect 14024 67398 14076 67450
rect 14148 67398 14200 67450
rect 14272 67398 14324 67450
rect 14396 67398 14448 67450
rect 14520 67398 14572 67450
rect 14644 67398 14696 67450
rect 14768 67398 14820 67450
rect 14892 67398 14944 67450
rect 15016 67398 15068 67450
rect 15140 67398 15192 67450
rect 34024 67398 34076 67450
rect 34148 67398 34200 67450
rect 34272 67398 34324 67450
rect 34396 67398 34448 67450
rect 34520 67398 34572 67450
rect 34644 67398 34696 67450
rect 34768 67398 34820 67450
rect 34892 67398 34944 67450
rect 35016 67398 35068 67450
rect 35140 67398 35192 67450
rect 6078 67230 6130 67282
rect 12574 67230 12626 67282
rect 15710 67230 15762 67282
rect 18062 67230 18114 67282
rect 19854 67230 19906 67282
rect 23886 67230 23938 67282
rect 26126 67230 26178 67282
rect 31838 67230 31890 67282
rect 37662 67230 37714 67282
rect 3950 67118 4002 67170
rect 4510 67118 4562 67170
rect 13470 67118 13522 67170
rect 13918 67118 13970 67170
rect 15486 67118 15538 67170
rect 17614 67118 17666 67170
rect 17950 67118 18002 67170
rect 25454 67118 25506 67170
rect 26014 67118 26066 67170
rect 33182 67118 33234 67170
rect 33294 67118 33346 67170
rect 36878 67118 36930 67170
rect 3726 67006 3778 67058
rect 8430 67006 8482 67058
rect 9102 67006 9154 67058
rect 9662 67006 9714 67058
rect 10110 67006 10162 67058
rect 15262 67006 15314 67058
rect 16270 67006 16322 67058
rect 16718 67006 16770 67058
rect 17390 67006 17442 67058
rect 18958 67006 19010 67058
rect 19070 67006 19122 67058
rect 19182 67006 19234 67058
rect 19630 67006 19682 67058
rect 20974 67006 21026 67058
rect 21422 67006 21474 67058
rect 28926 67006 28978 67058
rect 29262 67006 29314 67058
rect 33966 67006 34018 67058
rect 34526 67006 34578 67058
rect 5406 66894 5458 66946
rect 14926 66894 14978 66946
rect 20190 66894 20242 66946
rect 25230 66894 25282 66946
rect 25566 66894 25618 66946
rect 26238 66894 26290 66946
rect 26686 66894 26738 66946
rect 33742 66894 33794 66946
rect 3390 66782 3442 66834
rect 13134 66782 13186 66834
rect 24446 66782 24498 66834
rect 32398 66782 32450 66834
rect 33182 66782 33234 66834
rect 4024 66614 4076 66666
rect 4148 66614 4200 66666
rect 4272 66614 4324 66666
rect 4396 66614 4448 66666
rect 4520 66614 4572 66666
rect 4644 66614 4696 66666
rect 4768 66614 4820 66666
rect 4892 66614 4944 66666
rect 5016 66614 5068 66666
rect 5140 66614 5192 66666
rect 24024 66614 24076 66666
rect 24148 66614 24200 66666
rect 24272 66614 24324 66666
rect 24396 66614 24448 66666
rect 24520 66614 24572 66666
rect 24644 66614 24696 66666
rect 24768 66614 24820 66666
rect 24892 66614 24944 66666
rect 25016 66614 25068 66666
rect 25140 66614 25192 66666
rect 6750 66446 6802 66498
rect 7310 66446 7362 66498
rect 7534 66446 7586 66498
rect 8766 66446 8818 66498
rect 10670 66446 10722 66498
rect 11006 66446 11058 66498
rect 19630 66446 19682 66498
rect 20638 66446 20690 66498
rect 21422 66446 21474 66498
rect 21758 66446 21810 66498
rect 37326 66446 37378 66498
rect 8430 66334 8482 66386
rect 9214 66334 9266 66386
rect 10222 66334 10274 66386
rect 15934 66334 15986 66386
rect 16270 66334 16322 66386
rect 19182 66334 19234 66386
rect 25566 66334 25618 66386
rect 36990 66334 37042 66386
rect 37550 66334 37602 66386
rect 4958 66222 5010 66274
rect 6414 66222 6466 66274
rect 6974 66222 7026 66274
rect 8206 66222 8258 66274
rect 17166 66222 17218 66274
rect 19070 66222 19122 66274
rect 29038 66222 29090 66274
rect 29598 66222 29650 66274
rect 2158 66110 2210 66162
rect 4510 66110 4562 66162
rect 11230 66110 11282 66162
rect 11678 66110 11730 66162
rect 18510 66110 18562 66162
rect 20638 66110 20690 66162
rect 20750 66110 20802 66162
rect 21982 66110 22034 66162
rect 22542 66110 22594 66162
rect 31950 66110 32002 66162
rect 36094 66110 36146 66162
rect 1710 65998 1762 66050
rect 4062 65998 4114 66050
rect 4398 65998 4450 66050
rect 4622 65998 4674 66050
rect 5742 65998 5794 66050
rect 7646 65998 7698 66050
rect 9774 65998 9826 66050
rect 17614 65998 17666 66050
rect 18062 65998 18114 66050
rect 24558 65998 24610 66050
rect 25006 65998 25058 66050
rect 25902 65998 25954 66050
rect 26350 65998 26402 66050
rect 28590 65998 28642 66050
rect 32734 65998 32786 66050
rect 36206 65998 36258 66050
rect 36318 65998 36370 66050
rect 14024 65830 14076 65882
rect 14148 65830 14200 65882
rect 14272 65830 14324 65882
rect 14396 65830 14448 65882
rect 14520 65830 14572 65882
rect 14644 65830 14696 65882
rect 14768 65830 14820 65882
rect 14892 65830 14944 65882
rect 15016 65830 15068 65882
rect 15140 65830 15192 65882
rect 34024 65830 34076 65882
rect 34148 65830 34200 65882
rect 34272 65830 34324 65882
rect 34396 65830 34448 65882
rect 34520 65830 34572 65882
rect 34644 65830 34696 65882
rect 34768 65830 34820 65882
rect 34892 65830 34944 65882
rect 35016 65830 35068 65882
rect 35140 65830 35192 65882
rect 4734 65662 4786 65714
rect 7870 65662 7922 65714
rect 13246 65662 13298 65714
rect 18734 65662 18786 65714
rect 20974 65662 21026 65714
rect 28366 65662 28418 65714
rect 33742 65662 33794 65714
rect 36878 65662 36930 65714
rect 14030 65550 14082 65602
rect 19070 65550 19122 65602
rect 1822 65438 1874 65490
rect 2270 65438 2322 65490
rect 5294 65438 5346 65490
rect 5630 65438 5682 65490
rect 6190 65438 6242 65490
rect 9998 65438 10050 65490
rect 10670 65438 10722 65490
rect 13582 65438 13634 65490
rect 13806 65438 13858 65490
rect 19182 65438 19234 65490
rect 19630 65438 19682 65490
rect 20526 65438 20578 65490
rect 20862 65438 20914 65490
rect 21310 65438 21362 65490
rect 21534 65438 21586 65490
rect 25342 65438 25394 65490
rect 26014 65438 26066 65490
rect 29374 65438 29426 65490
rect 30830 65438 30882 65490
rect 31278 65438 31330 65490
rect 31502 65438 31554 65490
rect 31614 65438 31666 65490
rect 31838 65438 31890 65490
rect 33966 65438 34018 65490
rect 34638 65438 34690 65490
rect 37662 65438 37714 65490
rect 12798 65326 12850 65378
rect 14478 65326 14530 65378
rect 17838 65326 17890 65378
rect 18286 65326 18338 65378
rect 19742 65326 19794 65378
rect 21982 65326 22034 65378
rect 14142 65214 14194 65266
rect 19966 65214 20018 65266
rect 20190 65214 20242 65266
rect 20302 65214 20354 65266
rect 21086 65214 21138 65266
rect 29038 65214 29090 65266
rect 4024 65046 4076 65098
rect 4148 65046 4200 65098
rect 4272 65046 4324 65098
rect 4396 65046 4448 65098
rect 4520 65046 4572 65098
rect 4644 65046 4696 65098
rect 4768 65046 4820 65098
rect 4892 65046 4944 65098
rect 5016 65046 5068 65098
rect 5140 65046 5192 65098
rect 24024 65046 24076 65098
rect 24148 65046 24200 65098
rect 24272 65046 24324 65098
rect 24396 65046 24448 65098
rect 24520 65046 24572 65098
rect 24644 65046 24696 65098
rect 24768 65046 24820 65098
rect 24892 65046 24944 65098
rect 25016 65046 25068 65098
rect 25140 65046 25192 65098
rect 3838 64878 3890 64930
rect 10110 64878 10162 64930
rect 11342 64878 11394 64930
rect 16158 64878 16210 64930
rect 35534 64878 35586 64930
rect 35870 64878 35922 64930
rect 36990 64878 37042 64930
rect 37326 64878 37378 64930
rect 8542 64766 8594 64818
rect 10446 64766 10498 64818
rect 10670 64766 10722 64818
rect 11006 64766 11058 64818
rect 11790 64766 11842 64818
rect 15486 64766 15538 64818
rect 17166 64766 17218 64818
rect 18174 64766 18226 64818
rect 18734 64766 18786 64818
rect 20302 64766 20354 64818
rect 29262 64766 29314 64818
rect 35198 64766 35250 64818
rect 37550 64766 37602 64818
rect 7758 64654 7810 64706
rect 13918 64654 13970 64706
rect 14030 64654 14082 64706
rect 14814 64654 14866 64706
rect 15598 64654 15650 64706
rect 16046 64654 16098 64706
rect 18286 64654 18338 64706
rect 18958 64654 19010 64706
rect 35646 64654 35698 64706
rect 36094 64654 36146 64706
rect 2830 64542 2882 64594
rect 3166 64542 3218 64594
rect 3726 64542 3778 64594
rect 11118 64542 11170 64594
rect 12574 64542 12626 64594
rect 12910 64542 12962 64594
rect 13470 64542 13522 64594
rect 14478 64542 14530 64594
rect 14590 64542 14642 64594
rect 19518 64542 19570 64594
rect 1710 64430 1762 64482
rect 2606 64430 2658 64482
rect 5742 64430 5794 64482
rect 12238 64430 12290 64482
rect 13694 64430 13746 64482
rect 13806 64430 13858 64482
rect 16718 64430 16770 64482
rect 17614 64430 17666 64482
rect 19294 64430 19346 64482
rect 19630 64430 19682 64482
rect 29822 64430 29874 64482
rect 14024 64262 14076 64314
rect 14148 64262 14200 64314
rect 14272 64262 14324 64314
rect 14396 64262 14448 64314
rect 14520 64262 14572 64314
rect 14644 64262 14696 64314
rect 14768 64262 14820 64314
rect 14892 64262 14944 64314
rect 15016 64262 15068 64314
rect 15140 64262 15192 64314
rect 34024 64262 34076 64314
rect 34148 64262 34200 64314
rect 34272 64262 34324 64314
rect 34396 64262 34448 64314
rect 34520 64262 34572 64314
rect 34644 64262 34696 64314
rect 34768 64262 34820 64314
rect 34892 64262 34944 64314
rect 35016 64262 35068 64314
rect 35140 64262 35192 64314
rect 4846 64094 4898 64146
rect 5742 64094 5794 64146
rect 6190 64094 6242 64146
rect 8990 64094 9042 64146
rect 12462 64094 12514 64146
rect 16046 64094 16098 64146
rect 17278 64094 17330 64146
rect 28254 64094 28306 64146
rect 30270 64094 30322 64146
rect 14702 63982 14754 64034
rect 16158 63982 16210 64034
rect 29150 63982 29202 64034
rect 1934 63870 1986 63922
rect 2382 63870 2434 63922
rect 5406 63870 5458 63922
rect 9662 63870 9714 63922
rect 9998 63870 10050 63922
rect 13134 63870 13186 63922
rect 15262 63870 15314 63922
rect 15598 63870 15650 63922
rect 17950 63870 18002 63922
rect 18286 63870 18338 63922
rect 19518 63870 19570 63922
rect 20414 63870 20466 63922
rect 25342 63870 25394 63922
rect 25678 63870 25730 63922
rect 28814 63870 28866 63922
rect 29262 63870 29314 63922
rect 31838 63870 31890 63922
rect 13694 63758 13746 63810
rect 13918 63758 13970 63810
rect 18062 63758 18114 63810
rect 19630 63758 19682 63810
rect 19966 63758 20018 63810
rect 29934 63758 29986 63810
rect 31278 63758 31330 63810
rect 14254 63646 14306 63698
rect 4024 63478 4076 63530
rect 4148 63478 4200 63530
rect 4272 63478 4324 63530
rect 4396 63478 4448 63530
rect 4520 63478 4572 63530
rect 4644 63478 4696 63530
rect 4768 63478 4820 63530
rect 4892 63478 4944 63530
rect 5016 63478 5068 63530
rect 5140 63478 5192 63530
rect 24024 63478 24076 63530
rect 24148 63478 24200 63530
rect 24272 63478 24324 63530
rect 24396 63478 24448 63530
rect 24520 63478 24572 63530
rect 24644 63478 24696 63530
rect 24768 63478 24820 63530
rect 24892 63478 24944 63530
rect 25016 63478 25068 63530
rect 25140 63478 25192 63530
rect 3838 63310 3890 63362
rect 7534 63310 7586 63362
rect 18062 63310 18114 63362
rect 31726 63310 31778 63362
rect 4174 63198 4226 63250
rect 5742 63198 5794 63250
rect 6862 63198 6914 63250
rect 12350 63198 12402 63250
rect 13582 63198 13634 63250
rect 15486 63198 15538 63250
rect 16830 63198 16882 63250
rect 24782 63198 24834 63250
rect 34750 63198 34802 63250
rect 4958 63086 5010 63138
rect 6190 63086 6242 63138
rect 7198 63086 7250 63138
rect 8318 63086 8370 63138
rect 8542 63086 8594 63138
rect 8766 63086 8818 63138
rect 9550 63086 9602 63138
rect 10110 63086 10162 63138
rect 14926 63086 14978 63138
rect 15934 63086 15986 63138
rect 16382 63086 16434 63138
rect 17278 63086 17330 63138
rect 20078 63086 20130 63138
rect 20302 63086 20354 63138
rect 20526 63086 20578 63138
rect 23774 63086 23826 63138
rect 24894 63086 24946 63138
rect 25230 63086 25282 63138
rect 30494 63086 30546 63138
rect 31054 63086 31106 63138
rect 31278 63086 31330 63138
rect 4734 62974 4786 63026
rect 8990 62974 9042 63026
rect 14478 62974 14530 63026
rect 15262 62974 15314 63026
rect 16830 62974 16882 63026
rect 18174 62974 18226 63026
rect 19406 62974 19458 63026
rect 19854 62974 19906 63026
rect 20638 62974 20690 63026
rect 20750 62974 20802 63026
rect 24110 62974 24162 63026
rect 24670 62974 24722 63026
rect 26574 62974 26626 63026
rect 27022 62974 27074 63026
rect 27134 62974 27186 63026
rect 30718 62974 30770 63026
rect 34862 62974 34914 63026
rect 35086 62974 35138 63026
rect 35870 62974 35922 63026
rect 1710 62862 1762 62914
rect 7422 62862 7474 62914
rect 7982 62862 8034 62914
rect 14030 62862 14082 62914
rect 17054 62862 17106 62914
rect 19070 62862 19122 62914
rect 19518 62862 19570 62914
rect 25678 62862 25730 62914
rect 26798 62862 26850 62914
rect 28590 62862 28642 62914
rect 29262 62862 29314 62914
rect 30158 62862 30210 62914
rect 33630 62862 33682 62914
rect 35534 62862 35586 62914
rect 35758 62862 35810 62914
rect 35982 62862 36034 62914
rect 14024 62694 14076 62746
rect 14148 62694 14200 62746
rect 14272 62694 14324 62746
rect 14396 62694 14448 62746
rect 14520 62694 14572 62746
rect 14644 62694 14696 62746
rect 14768 62694 14820 62746
rect 14892 62694 14944 62746
rect 15016 62694 15068 62746
rect 15140 62694 15192 62746
rect 34024 62694 34076 62746
rect 34148 62694 34200 62746
rect 34272 62694 34324 62746
rect 34396 62694 34448 62746
rect 34520 62694 34572 62746
rect 34644 62694 34696 62746
rect 34768 62694 34820 62746
rect 34892 62694 34944 62746
rect 35016 62694 35068 62746
rect 35140 62694 35192 62746
rect 8318 62526 8370 62578
rect 8878 62526 8930 62578
rect 9998 62526 10050 62578
rect 13582 62526 13634 62578
rect 14366 62526 14418 62578
rect 16270 62526 16322 62578
rect 16718 62526 16770 62578
rect 20190 62526 20242 62578
rect 24110 62526 24162 62578
rect 28254 62526 28306 62578
rect 29598 62526 29650 62578
rect 36766 62526 36818 62578
rect 37550 62526 37602 62578
rect 1710 62414 1762 62466
rect 4846 62414 4898 62466
rect 9886 62414 9938 62466
rect 10446 62414 10498 62466
rect 15822 62414 15874 62466
rect 19294 62414 19346 62466
rect 24670 62414 24722 62466
rect 30942 62414 30994 62466
rect 31054 62414 31106 62466
rect 4398 62302 4450 62354
rect 4734 62302 4786 62354
rect 5294 62302 5346 62354
rect 5742 62302 5794 62354
rect 10222 62302 10274 62354
rect 10894 62302 10946 62354
rect 11230 62302 11282 62354
rect 14814 62302 14866 62354
rect 14926 62302 14978 62354
rect 15374 62302 15426 62354
rect 16046 62302 16098 62354
rect 19742 62302 19794 62354
rect 19854 62302 19906 62354
rect 20078 62302 20130 62354
rect 20302 62302 20354 62354
rect 20974 62302 21026 62354
rect 21534 62302 21586 62354
rect 25342 62302 25394 62354
rect 25790 62302 25842 62354
rect 29150 62302 29202 62354
rect 30046 62302 30098 62354
rect 30718 62302 30770 62354
rect 33406 62302 33458 62354
rect 33854 62302 33906 62354
rect 34414 62302 34466 62354
rect 14590 62190 14642 62242
rect 28814 62190 28866 62242
rect 4846 62078 4898 62130
rect 15598 62078 15650 62130
rect 15934 62078 15986 62130
rect 4024 61910 4076 61962
rect 4148 61910 4200 61962
rect 4272 61910 4324 61962
rect 4396 61910 4448 61962
rect 4520 61910 4572 61962
rect 4644 61910 4696 61962
rect 4768 61910 4820 61962
rect 4892 61910 4944 61962
rect 5016 61910 5068 61962
rect 5140 61910 5192 61962
rect 24024 61910 24076 61962
rect 24148 61910 24200 61962
rect 24272 61910 24324 61962
rect 24396 61910 24448 61962
rect 24520 61910 24572 61962
rect 24644 61910 24696 61962
rect 24768 61910 24820 61962
rect 24892 61910 24944 61962
rect 25016 61910 25068 61962
rect 25140 61910 25192 61962
rect 12798 61742 12850 61794
rect 15598 61742 15650 61794
rect 15822 61742 15874 61794
rect 17166 61742 17218 61794
rect 21422 61742 21474 61794
rect 26014 61742 26066 61794
rect 26350 61742 26402 61794
rect 36990 61742 37042 61794
rect 6750 61630 6802 61682
rect 11454 61630 11506 61682
rect 14926 61630 14978 61682
rect 15374 61630 15426 61682
rect 16942 61630 16994 61682
rect 24222 61630 24274 61682
rect 35534 61630 35586 61682
rect 35982 61630 36034 61682
rect 37550 61630 37602 61682
rect 4062 61518 4114 61570
rect 4622 61518 4674 61570
rect 8206 61518 8258 61570
rect 9214 61518 9266 61570
rect 10334 61518 10386 61570
rect 11790 61518 11842 61570
rect 12014 61518 12066 61570
rect 12910 61518 12962 61570
rect 13582 61518 13634 61570
rect 13806 61518 13858 61570
rect 15038 61518 15090 61570
rect 20190 61518 20242 61570
rect 20862 61518 20914 61570
rect 21758 61518 21810 61570
rect 29374 61518 29426 61570
rect 29934 61518 29986 61570
rect 36206 61518 36258 61570
rect 36318 61518 36370 61570
rect 37326 61518 37378 61570
rect 4846 61406 4898 61458
rect 11118 61406 11170 61458
rect 12350 61406 12402 61458
rect 14926 61406 14978 61458
rect 21982 61406 22034 61458
rect 22318 61406 22370 61458
rect 24558 61406 24610 61458
rect 25230 61406 25282 61458
rect 25790 61406 25842 61458
rect 28478 61406 28530 61458
rect 35870 61406 35922 61458
rect 1710 61294 1762 61346
rect 3726 61294 3778 61346
rect 5742 61294 5794 61346
rect 8878 61294 8930 61346
rect 9102 61294 9154 61346
rect 9886 61294 9938 61346
rect 10782 61294 10834 61346
rect 11342 61294 11394 61346
rect 12126 61294 12178 61346
rect 16270 61294 16322 61346
rect 17726 61294 17778 61346
rect 28590 61294 28642 61346
rect 32510 61294 32562 61346
rect 33070 61294 33122 61346
rect 33406 61294 33458 61346
rect 33854 61294 33906 61346
rect 34414 61294 34466 61346
rect 14024 61126 14076 61178
rect 14148 61126 14200 61178
rect 14272 61126 14324 61178
rect 14396 61126 14448 61178
rect 14520 61126 14572 61178
rect 14644 61126 14696 61178
rect 14768 61126 14820 61178
rect 14892 61126 14944 61178
rect 15016 61126 15068 61178
rect 15140 61126 15192 61178
rect 34024 61126 34076 61178
rect 34148 61126 34200 61178
rect 34272 61126 34324 61178
rect 34396 61126 34448 61178
rect 34520 61126 34572 61178
rect 34644 61126 34696 61178
rect 34768 61126 34820 61178
rect 34892 61126 34944 61178
rect 35016 61126 35068 61178
rect 35140 61126 35192 61178
rect 4734 60958 4786 61010
rect 5294 60958 5346 61010
rect 5630 60958 5682 61010
rect 13582 60958 13634 61010
rect 13694 60958 13746 61010
rect 21422 60958 21474 61010
rect 33182 60958 33234 61010
rect 34190 60958 34242 61010
rect 37774 60958 37826 61010
rect 6638 60846 6690 60898
rect 7198 60846 7250 60898
rect 7534 60846 7586 60898
rect 29934 60846 29986 60898
rect 30046 60846 30098 60898
rect 1822 60734 1874 60786
rect 2270 60734 2322 60786
rect 5966 60734 6018 60786
rect 6750 60734 6802 60786
rect 7422 60734 7474 60786
rect 7982 60734 8034 60786
rect 8542 60734 8594 60786
rect 15934 60734 15986 60786
rect 16382 60734 16434 60786
rect 27022 60734 27074 60786
rect 30606 60734 30658 60786
rect 31054 60734 31106 60786
rect 31502 60734 31554 60786
rect 31726 60734 31778 60786
rect 32062 60734 32114 60786
rect 32398 60734 32450 60786
rect 33294 60734 33346 60786
rect 34638 60734 34690 60786
rect 35310 60734 35362 60786
rect 8990 60622 9042 60674
rect 9662 60622 9714 60674
rect 10110 60622 10162 60674
rect 20974 60622 21026 60674
rect 25342 60622 25394 60674
rect 26686 60622 26738 60674
rect 28702 60622 28754 60674
rect 31950 60622 32002 60674
rect 33742 60622 33794 60674
rect 7758 60510 7810 60562
rect 13470 60510 13522 60562
rect 16158 60510 16210 60562
rect 16494 60510 16546 60562
rect 20862 60510 20914 60562
rect 21534 60510 21586 60562
rect 30046 60510 30098 60562
rect 33182 60510 33234 60562
rect 38334 60510 38386 60562
rect 4024 60342 4076 60394
rect 4148 60342 4200 60394
rect 4272 60342 4324 60394
rect 4396 60342 4448 60394
rect 4520 60342 4572 60394
rect 4644 60342 4696 60394
rect 4768 60342 4820 60394
rect 4892 60342 4944 60394
rect 5016 60342 5068 60394
rect 5140 60342 5192 60394
rect 24024 60342 24076 60394
rect 24148 60342 24200 60394
rect 24272 60342 24324 60394
rect 24396 60342 24448 60394
rect 24520 60342 24572 60394
rect 24644 60342 24696 60394
rect 24768 60342 24820 60394
rect 24892 60342 24944 60394
rect 25016 60342 25068 60394
rect 25140 60342 25192 60394
rect 5966 60174 6018 60226
rect 6190 60174 6242 60226
rect 28590 60174 28642 60226
rect 33966 60174 34018 60226
rect 36990 60174 37042 60226
rect 5742 60062 5794 60114
rect 6190 60062 6242 60114
rect 12798 60062 12850 60114
rect 19630 60062 19682 60114
rect 20526 60062 20578 60114
rect 26014 60062 26066 60114
rect 29934 60062 29986 60114
rect 36318 60062 36370 60114
rect 37550 60062 37602 60114
rect 7086 59950 7138 60002
rect 23774 59950 23826 60002
rect 30270 59950 30322 60002
rect 30942 59950 30994 60002
rect 36430 59950 36482 60002
rect 37326 59950 37378 60002
rect 19294 59838 19346 59890
rect 29598 59838 29650 59890
rect 29822 59838 29874 59890
rect 30046 59838 30098 59890
rect 36206 59838 36258 59890
rect 1710 59726 1762 59778
rect 19070 59726 19122 59778
rect 20190 59726 20242 59778
rect 21534 59726 21586 59778
rect 23438 59726 23490 59778
rect 28030 59726 28082 59778
rect 28366 59726 28418 59778
rect 28478 59726 28530 59778
rect 33182 59726 33234 59778
rect 34302 59726 34354 59778
rect 14024 59558 14076 59610
rect 14148 59558 14200 59610
rect 14272 59558 14324 59610
rect 14396 59558 14448 59610
rect 14520 59558 14572 59610
rect 14644 59558 14696 59610
rect 14768 59558 14820 59610
rect 14892 59558 14944 59610
rect 15016 59558 15068 59610
rect 15140 59558 15192 59610
rect 34024 59558 34076 59610
rect 34148 59558 34200 59610
rect 34272 59558 34324 59610
rect 34396 59558 34448 59610
rect 34520 59558 34572 59610
rect 34644 59558 34696 59610
rect 34768 59558 34820 59610
rect 34892 59558 34944 59610
rect 35016 59558 35068 59610
rect 35140 59558 35192 59610
rect 11678 59390 11730 59442
rect 18398 59390 18450 59442
rect 19742 59390 19794 59442
rect 19854 59390 19906 59442
rect 20638 59390 20690 59442
rect 20750 59390 20802 59442
rect 25342 59390 25394 59442
rect 30494 59390 30546 59442
rect 31614 59390 31666 59442
rect 31726 59390 31778 59442
rect 13022 59278 13074 59330
rect 15038 59278 15090 59330
rect 18510 59278 18562 59330
rect 21646 59278 21698 59330
rect 28926 59278 28978 59330
rect 31838 59278 31890 59330
rect 33070 59278 33122 59330
rect 33294 59278 33346 59330
rect 14030 59166 14082 59218
rect 14478 59166 14530 59218
rect 14814 59166 14866 59218
rect 15374 59166 15426 59218
rect 16046 59166 16098 59218
rect 18734 59166 18786 59218
rect 19070 59166 19122 59218
rect 19966 59166 20018 59218
rect 20414 59166 20466 59218
rect 20862 59166 20914 59218
rect 21310 59166 21362 59218
rect 21534 59166 21586 59218
rect 26014 59166 26066 59218
rect 26686 59166 26738 59218
rect 29934 59166 29986 59218
rect 31950 59166 32002 59218
rect 32286 59166 32338 59218
rect 11342 59054 11394 59106
rect 12462 59054 12514 59106
rect 13582 59054 13634 59106
rect 18062 59054 18114 59106
rect 19518 59054 19570 59106
rect 22206 59054 22258 59106
rect 25790 59054 25842 59106
rect 14702 58942 14754 58994
rect 21646 58942 21698 58994
rect 29710 58942 29762 58994
rect 33406 58942 33458 58994
rect 4024 58774 4076 58826
rect 4148 58774 4200 58826
rect 4272 58774 4324 58826
rect 4396 58774 4448 58826
rect 4520 58774 4572 58826
rect 4644 58774 4696 58826
rect 4768 58774 4820 58826
rect 4892 58774 4944 58826
rect 5016 58774 5068 58826
rect 5140 58774 5192 58826
rect 24024 58774 24076 58826
rect 24148 58774 24200 58826
rect 24272 58774 24324 58826
rect 24396 58774 24448 58826
rect 24520 58774 24572 58826
rect 24644 58774 24696 58826
rect 24768 58774 24820 58826
rect 24892 58774 24944 58826
rect 25016 58774 25068 58826
rect 25140 58774 25192 58826
rect 31278 58606 31330 58658
rect 32174 58606 32226 58658
rect 3950 58494 4002 58546
rect 13582 58494 13634 58546
rect 15262 58494 15314 58546
rect 32286 58494 32338 58546
rect 2942 58382 2994 58434
rect 7534 58382 7586 58434
rect 7870 58382 7922 58434
rect 9214 58382 9266 58434
rect 9550 58382 9602 58434
rect 14814 58382 14866 58434
rect 15038 58382 15090 58434
rect 17166 58382 17218 58434
rect 17502 58382 17554 58434
rect 18510 58382 18562 58434
rect 19070 58382 19122 58434
rect 19294 58382 19346 58434
rect 19518 58382 19570 58434
rect 19854 58382 19906 58434
rect 20414 58382 20466 58434
rect 20750 58382 20802 58434
rect 21310 58382 21362 58434
rect 21646 58382 21698 58434
rect 26686 58382 26738 58434
rect 27358 58382 27410 58434
rect 28142 58382 28194 58434
rect 29934 58382 29986 58434
rect 30270 58382 30322 58434
rect 30606 58382 30658 58434
rect 31614 58382 31666 58434
rect 31838 58382 31890 58434
rect 34974 58382 35026 58434
rect 35198 58382 35250 58434
rect 36878 58382 36930 58434
rect 2494 58270 2546 58322
rect 7198 58158 7250 58210
rect 7310 58214 7362 58266
rect 15710 58270 15762 58322
rect 16158 58270 16210 58322
rect 16606 58270 16658 58322
rect 18062 58270 18114 58322
rect 18398 58270 18450 58322
rect 18846 58270 18898 58322
rect 20078 58270 20130 58322
rect 20190 58270 20242 58322
rect 21982 58270 22034 58322
rect 35534 58270 35586 58322
rect 37326 58270 37378 58322
rect 37550 58270 37602 58322
rect 8206 58158 8258 58210
rect 8766 58158 8818 58210
rect 12126 58158 12178 58210
rect 12686 58158 12738 58210
rect 18734 58158 18786 58210
rect 20638 58158 20690 58210
rect 21646 58158 21698 58210
rect 22542 58158 22594 58210
rect 23662 58158 23714 58210
rect 24222 58158 24274 58210
rect 27694 58158 27746 58210
rect 29598 58158 29650 58210
rect 30270 58158 30322 58210
rect 30942 58158 30994 58210
rect 31390 58158 31442 58210
rect 32734 58158 32786 58210
rect 34414 58158 34466 58210
rect 37102 58158 37154 58210
rect 14024 57990 14076 58042
rect 14148 57990 14200 58042
rect 14272 57990 14324 58042
rect 14396 57990 14448 58042
rect 14520 57990 14572 58042
rect 14644 57990 14696 58042
rect 14768 57990 14820 58042
rect 14892 57990 14944 58042
rect 15016 57990 15068 58042
rect 15140 57990 15192 58042
rect 34024 57990 34076 58042
rect 34148 57990 34200 58042
rect 34272 57990 34324 58042
rect 34396 57990 34448 58042
rect 34520 57990 34572 58042
rect 34644 57990 34696 58042
rect 34768 57990 34820 58042
rect 34892 57990 34944 58042
rect 35016 57990 35068 58042
rect 35140 57990 35192 58042
rect 6526 57822 6578 57874
rect 7086 57822 7138 57874
rect 7310 57822 7362 57874
rect 8542 57822 8594 57874
rect 12574 57822 12626 57874
rect 19294 57822 19346 57874
rect 20638 57822 20690 57874
rect 24222 57822 24274 57874
rect 25342 57822 25394 57874
rect 28142 57822 28194 57874
rect 29934 57822 29986 57874
rect 30494 57822 30546 57874
rect 30942 57822 30994 57874
rect 33742 57822 33794 57874
rect 34302 57822 34354 57874
rect 37662 57822 37714 57874
rect 38334 57822 38386 57874
rect 10558 57710 10610 57762
rect 11902 57710 11954 57762
rect 12686 57710 12738 57762
rect 14254 57710 14306 57762
rect 18846 57710 18898 57762
rect 24782 57710 24834 57762
rect 25902 57710 25954 57762
rect 26238 57710 26290 57762
rect 27246 57710 27298 57762
rect 2830 57598 2882 57650
rect 6862 57598 6914 57650
rect 10782 57598 10834 57650
rect 11790 57598 11842 57650
rect 12798 57598 12850 57650
rect 13806 57598 13858 57650
rect 14366 57598 14418 57650
rect 15374 57598 15426 57650
rect 15822 57598 15874 57650
rect 16382 57598 16434 57650
rect 18622 57598 18674 57650
rect 19182 57598 19234 57650
rect 19406 57598 19458 57650
rect 19742 57598 19794 57650
rect 20078 57598 20130 57650
rect 20750 57598 20802 57650
rect 21086 57598 21138 57650
rect 21646 57598 21698 57650
rect 25678 57598 25730 57650
rect 27134 57598 27186 57650
rect 27806 57598 27858 57650
rect 34078 57598 34130 57650
rect 34638 57598 34690 57650
rect 35310 57598 35362 57650
rect 2606 57486 2658 57538
rect 3502 57486 3554 57538
rect 6974 57486 7026 57538
rect 7982 57486 8034 57538
rect 9102 57486 9154 57538
rect 15262 57486 15314 57538
rect 16830 57486 16882 57538
rect 17726 57486 17778 57538
rect 18174 57486 18226 57538
rect 20526 57486 20578 57538
rect 30830 57486 30882 57538
rect 8206 57374 8258 57426
rect 9662 57374 9714 57426
rect 9998 57374 10050 57426
rect 17838 57374 17890 57426
rect 18286 57374 18338 57426
rect 18510 57374 18562 57426
rect 20302 57374 20354 57426
rect 31166 57374 31218 57426
rect 34414 57374 34466 57426
rect 4024 57206 4076 57258
rect 4148 57206 4200 57258
rect 4272 57206 4324 57258
rect 4396 57206 4448 57258
rect 4520 57206 4572 57258
rect 4644 57206 4696 57258
rect 4768 57206 4820 57258
rect 4892 57206 4944 57258
rect 5016 57206 5068 57258
rect 5140 57206 5192 57258
rect 24024 57206 24076 57258
rect 24148 57206 24200 57258
rect 24272 57206 24324 57258
rect 24396 57206 24448 57258
rect 24520 57206 24572 57258
rect 24644 57206 24696 57258
rect 24768 57206 24820 57258
rect 24892 57206 24944 57258
rect 25016 57206 25068 57258
rect 25140 57206 25192 57258
rect 6078 57038 6130 57090
rect 12798 57038 12850 57090
rect 13582 57038 13634 57090
rect 25902 57038 25954 57090
rect 26574 57038 26626 57090
rect 34862 57038 34914 57090
rect 35870 57038 35922 57090
rect 36206 57038 36258 57090
rect 36990 57038 37042 57090
rect 7422 56926 7474 56978
rect 11678 56926 11730 56978
rect 12462 56926 12514 56978
rect 17390 56926 17442 56978
rect 26574 56926 26626 56978
rect 27470 56926 27522 56978
rect 3614 56814 3666 56866
rect 4286 56814 4338 56866
rect 6526 56814 6578 56866
rect 7646 56814 7698 56866
rect 8206 56814 8258 56866
rect 11342 56814 11394 56866
rect 11566 56814 11618 56866
rect 11902 56814 11954 56866
rect 12126 56814 12178 56866
rect 14254 56814 14306 56866
rect 15374 56814 15426 56866
rect 16382 56814 16434 56866
rect 17614 56814 17666 56866
rect 18622 56814 18674 56866
rect 19518 56814 19570 56866
rect 20414 56814 20466 56866
rect 21646 56814 21698 56866
rect 25118 56814 25170 56866
rect 25790 56814 25842 56866
rect 28590 56814 28642 56866
rect 29038 56814 29090 56866
rect 29710 56814 29762 56866
rect 34638 56814 34690 56866
rect 35086 56814 35138 56866
rect 35982 56814 36034 56866
rect 36430 56814 36482 56866
rect 37550 56814 37602 56866
rect 37774 56814 37826 56866
rect 4398 56702 4450 56754
rect 6638 56702 6690 56754
rect 13470 56702 13522 56754
rect 14366 56702 14418 56754
rect 15262 56702 15314 56754
rect 18174 56702 18226 56754
rect 19742 56702 19794 56754
rect 20302 56702 20354 56754
rect 21310 56702 21362 56754
rect 21870 56702 21922 56754
rect 22878 56702 22930 56754
rect 37438 56702 37490 56754
rect 3278 56590 3330 56642
rect 4958 56590 5010 56642
rect 5742 56590 5794 56642
rect 10558 56590 10610 56642
rect 12574 56590 12626 56642
rect 15038 56590 15090 56642
rect 16830 56590 16882 56642
rect 19630 56590 19682 56642
rect 21534 56590 21586 56642
rect 22094 56590 22146 56642
rect 26126 56590 26178 56642
rect 27022 56590 27074 56642
rect 28142 56590 28194 56642
rect 32062 56590 32114 56642
rect 32734 56590 32786 56642
rect 33854 56590 33906 56642
rect 34302 56590 34354 56642
rect 34750 56590 34802 56642
rect 14024 56422 14076 56474
rect 14148 56422 14200 56474
rect 14272 56422 14324 56474
rect 14396 56422 14448 56474
rect 14520 56422 14572 56474
rect 14644 56422 14696 56474
rect 14768 56422 14820 56474
rect 14892 56422 14944 56474
rect 15016 56422 15068 56474
rect 15140 56422 15192 56474
rect 34024 56422 34076 56474
rect 34148 56422 34200 56474
rect 34272 56422 34324 56474
rect 34396 56422 34448 56474
rect 34520 56422 34572 56474
rect 34644 56422 34696 56474
rect 34768 56422 34820 56474
rect 34892 56422 34944 56474
rect 35016 56422 35068 56474
rect 35140 56422 35192 56474
rect 6638 56254 6690 56306
rect 9662 56254 9714 56306
rect 18510 56254 18562 56306
rect 18958 56254 19010 56306
rect 20638 56254 20690 56306
rect 22766 56254 22818 56306
rect 24670 56254 24722 56306
rect 25342 56254 25394 56306
rect 36206 56254 36258 56306
rect 36766 56254 36818 56306
rect 36990 56254 37042 56306
rect 37214 56254 37266 56306
rect 8318 56142 8370 56194
rect 20750 56142 20802 56194
rect 22094 56142 22146 56194
rect 22990 56142 23042 56194
rect 32062 56142 32114 56194
rect 37438 56142 37490 56194
rect 2382 56030 2434 56082
rect 2830 56030 2882 56082
rect 3726 56030 3778 56082
rect 4174 56030 4226 56082
rect 7758 56030 7810 56082
rect 11454 56030 11506 56082
rect 11678 56030 11730 56082
rect 12574 56030 12626 56082
rect 13134 56030 13186 56082
rect 15038 56030 15090 56082
rect 16382 56030 16434 56082
rect 17390 56030 17442 56082
rect 17614 56030 17666 56082
rect 20302 56030 20354 56082
rect 21422 56030 21474 56082
rect 22318 56030 22370 56082
rect 32510 56030 32562 56082
rect 33294 56030 33346 56082
rect 33742 56030 33794 56082
rect 3278 55918 3330 55970
rect 7870 55918 7922 55970
rect 8766 55918 8818 55970
rect 10110 55918 10162 55970
rect 10670 55918 10722 55970
rect 11902 55918 11954 55970
rect 13246 55918 13298 55970
rect 13694 55918 13746 55970
rect 14254 55918 14306 55970
rect 14590 55918 14642 55970
rect 15486 55918 15538 55970
rect 15934 55918 15986 55970
rect 16830 55918 16882 55970
rect 18846 55918 18898 55970
rect 21982 55918 22034 55970
rect 25790 55918 25842 55970
rect 37102 55918 37154 55970
rect 7198 55806 7250 55858
rect 8542 55806 8594 55858
rect 9102 55806 9154 55858
rect 17838 55806 17890 55858
rect 18062 55806 18114 55858
rect 22654 55806 22706 55858
rect 4024 55638 4076 55690
rect 4148 55638 4200 55690
rect 4272 55638 4324 55690
rect 4396 55638 4448 55690
rect 4520 55638 4572 55690
rect 4644 55638 4696 55690
rect 4768 55638 4820 55690
rect 4892 55638 4944 55690
rect 5016 55638 5068 55690
rect 5140 55638 5192 55690
rect 24024 55638 24076 55690
rect 24148 55638 24200 55690
rect 24272 55638 24324 55690
rect 24396 55638 24448 55690
rect 24520 55638 24572 55690
rect 24644 55638 24696 55690
rect 24768 55638 24820 55690
rect 24892 55638 24944 55690
rect 25016 55638 25068 55690
rect 25140 55638 25192 55690
rect 3838 55470 3890 55522
rect 7198 55470 7250 55522
rect 11790 55470 11842 55522
rect 12910 55470 12962 55522
rect 14590 55470 14642 55522
rect 21870 55470 21922 55522
rect 22654 55470 22706 55522
rect 3278 55358 3330 55410
rect 8542 55358 8594 55410
rect 11118 55358 11170 55410
rect 13022 55358 13074 55410
rect 14030 55358 14082 55410
rect 16046 55358 16098 55410
rect 16830 55358 16882 55410
rect 21646 55358 21698 55410
rect 22094 55358 22146 55410
rect 22542 55358 22594 55410
rect 35758 55358 35810 55410
rect 36430 55358 36482 55410
rect 37438 55358 37490 55410
rect 4174 55246 4226 55298
rect 4846 55246 4898 55298
rect 6190 55246 6242 55298
rect 7982 55246 8034 55298
rect 10110 55246 10162 55298
rect 13918 55246 13970 55298
rect 14254 55246 14306 55298
rect 16382 55246 16434 55298
rect 18958 55246 19010 55298
rect 37102 55246 37154 55298
rect 37214 55246 37266 55298
rect 37550 55246 37602 55298
rect 4958 55134 5010 55186
rect 7310 55134 7362 55186
rect 8430 55134 8482 55186
rect 12462 55134 12514 55186
rect 18398 55134 18450 55186
rect 18734 55134 18786 55186
rect 19294 55134 19346 55186
rect 2606 55022 2658 55074
rect 2830 55022 2882 55074
rect 5742 55022 5794 55074
rect 6862 55022 6914 55074
rect 11566 55022 11618 55074
rect 12014 55022 12066 55074
rect 14142 55022 14194 55074
rect 15038 55022 15090 55074
rect 15486 55022 15538 55074
rect 18846 55022 18898 55074
rect 35646 55022 35698 55074
rect 14024 54854 14076 54906
rect 14148 54854 14200 54906
rect 14272 54854 14324 54906
rect 14396 54854 14448 54906
rect 14520 54854 14572 54906
rect 14644 54854 14696 54906
rect 14768 54854 14820 54906
rect 14892 54854 14944 54906
rect 15016 54854 15068 54906
rect 15140 54854 15192 54906
rect 34024 54854 34076 54906
rect 34148 54854 34200 54906
rect 34272 54854 34324 54906
rect 34396 54854 34448 54906
rect 34520 54854 34572 54906
rect 34644 54854 34696 54906
rect 34768 54854 34820 54906
rect 34892 54854 34944 54906
rect 35016 54854 35068 54906
rect 35140 54854 35192 54906
rect 4734 54686 4786 54738
rect 5294 54686 5346 54738
rect 5630 54686 5682 54738
rect 8094 54686 8146 54738
rect 11902 54686 11954 54738
rect 21198 54686 21250 54738
rect 21758 54686 21810 54738
rect 22094 54686 22146 54738
rect 26462 54686 26514 54738
rect 30270 54686 30322 54738
rect 31166 54686 31218 54738
rect 34078 54686 34130 54738
rect 37550 54686 37602 54738
rect 6302 54574 6354 54626
rect 8990 54574 9042 54626
rect 10782 54574 10834 54626
rect 1822 54462 1874 54514
rect 2270 54462 2322 54514
rect 6190 54462 6242 54514
rect 6526 54462 6578 54514
rect 6750 54462 6802 54514
rect 7086 54462 7138 54514
rect 7198 54462 7250 54514
rect 7646 54462 7698 54514
rect 9998 54462 10050 54514
rect 10670 54462 10722 54514
rect 13022 54462 13074 54514
rect 13470 54462 13522 54514
rect 15038 54462 15090 54514
rect 18286 54462 18338 54514
rect 18734 54462 18786 54514
rect 27358 54462 27410 54514
rect 27694 54462 27746 54514
rect 34526 54462 34578 54514
rect 35198 54462 35250 54514
rect 38222 54462 38274 54514
rect 7422 54350 7474 54402
rect 11454 54350 11506 54402
rect 12350 54350 12402 54402
rect 15262 54350 15314 54402
rect 15598 54350 15650 54402
rect 22542 54350 22594 54402
rect 27022 54350 27074 54402
rect 33630 54350 33682 54402
rect 9662 54238 9714 54290
rect 13246 54238 13298 54290
rect 13694 54238 13746 54290
rect 13806 54238 13858 54290
rect 30830 54238 30882 54290
rect 4024 54070 4076 54122
rect 4148 54070 4200 54122
rect 4272 54070 4324 54122
rect 4396 54070 4448 54122
rect 4520 54070 4572 54122
rect 4644 54070 4696 54122
rect 4768 54070 4820 54122
rect 4892 54070 4944 54122
rect 5016 54070 5068 54122
rect 5140 54070 5192 54122
rect 24024 54070 24076 54122
rect 24148 54070 24200 54122
rect 24272 54070 24324 54122
rect 24396 54070 24448 54122
rect 24520 54070 24572 54122
rect 24644 54070 24696 54122
rect 24768 54070 24820 54122
rect 24892 54070 24944 54122
rect 25016 54070 25068 54122
rect 25140 54070 25192 54122
rect 14814 53902 14866 53954
rect 15374 53902 15426 53954
rect 18622 53902 18674 53954
rect 19294 53902 19346 53954
rect 19630 53902 19682 53954
rect 26462 53902 26514 53954
rect 27694 53902 27746 53954
rect 30382 53902 30434 53954
rect 31054 53902 31106 53954
rect 3278 53790 3330 53842
rect 6974 53790 7026 53842
rect 12910 53790 12962 53842
rect 13470 53790 13522 53842
rect 14366 53790 14418 53842
rect 15038 53790 15090 53842
rect 15598 53790 15650 53842
rect 18174 53790 18226 53842
rect 20078 53790 20130 53842
rect 30382 53790 30434 53842
rect 2494 53678 2546 53730
rect 2830 53678 2882 53730
rect 5630 53678 5682 53730
rect 7870 53678 7922 53730
rect 8542 53678 8594 53730
rect 11566 53678 11618 53730
rect 12238 53678 12290 53730
rect 12798 53678 12850 53730
rect 13918 53678 13970 53730
rect 18286 53678 18338 53730
rect 24670 53678 24722 53730
rect 25902 53678 25954 53730
rect 26798 53678 26850 53730
rect 5742 53566 5794 53618
rect 15038 53566 15090 53618
rect 19406 53566 19458 53618
rect 25678 53566 25730 53618
rect 28030 53566 28082 53618
rect 28478 53566 28530 53618
rect 30830 53566 30882 53618
rect 31278 53566 31330 53618
rect 31390 53566 31442 53618
rect 31950 53566 32002 53618
rect 10894 53454 10946 53506
rect 25118 53454 25170 53506
rect 27358 53454 27410 53506
rect 29374 53454 29426 53506
rect 31614 53454 31666 53506
rect 14024 53286 14076 53338
rect 14148 53286 14200 53338
rect 14272 53286 14324 53338
rect 14396 53286 14448 53338
rect 14520 53286 14572 53338
rect 14644 53286 14696 53338
rect 14768 53286 14820 53338
rect 14892 53286 14944 53338
rect 15016 53286 15068 53338
rect 15140 53286 15192 53338
rect 34024 53286 34076 53338
rect 34148 53286 34200 53338
rect 34272 53286 34324 53338
rect 34396 53286 34448 53338
rect 34520 53286 34572 53338
rect 34644 53286 34696 53338
rect 34768 53286 34820 53338
rect 34892 53286 34944 53338
rect 35016 53286 35068 53338
rect 35140 53286 35192 53338
rect 4062 53118 4114 53170
rect 5182 53118 5234 53170
rect 5854 53118 5906 53170
rect 6526 53118 6578 53170
rect 12574 53118 12626 53170
rect 13134 53118 13186 53170
rect 18958 53118 19010 53170
rect 21646 53118 21698 53170
rect 22094 53118 22146 53170
rect 22654 53118 22706 53170
rect 22878 53118 22930 53170
rect 24222 53118 24274 53170
rect 25342 53118 25394 53170
rect 26350 53118 26402 53170
rect 29710 53118 29762 53170
rect 30270 53118 30322 53170
rect 6078 53006 6130 53058
rect 13358 53006 13410 53058
rect 23438 53006 23490 53058
rect 23662 53006 23714 53058
rect 23774 53006 23826 53058
rect 30942 53006 30994 53058
rect 2494 52894 2546 52946
rect 2830 52894 2882 52946
rect 3726 52894 3778 52946
rect 5406 52894 5458 52946
rect 9438 52894 9490 52946
rect 10110 52894 10162 52946
rect 13918 52894 13970 52946
rect 23326 52894 23378 52946
rect 26574 52894 26626 52946
rect 27246 52894 27298 52946
rect 30830 52894 30882 52946
rect 31166 52894 31218 52946
rect 31502 52894 31554 52946
rect 31950 52894 32002 52946
rect 32174 52894 32226 52946
rect 2046 52782 2098 52834
rect 3278 52782 3330 52834
rect 4734 52782 4786 52834
rect 5966 52782 6018 52834
rect 14702 52782 14754 52834
rect 20974 52782 21026 52834
rect 22766 52782 22818 52834
rect 25790 52782 25842 52834
rect 32062 52782 32114 52834
rect 13470 52670 13522 52722
rect 4024 52502 4076 52554
rect 4148 52502 4200 52554
rect 4272 52502 4324 52554
rect 4396 52502 4448 52554
rect 4520 52502 4572 52554
rect 4644 52502 4696 52554
rect 4768 52502 4820 52554
rect 4892 52502 4944 52554
rect 5016 52502 5068 52554
rect 5140 52502 5192 52554
rect 24024 52502 24076 52554
rect 24148 52502 24200 52554
rect 24272 52502 24324 52554
rect 24396 52502 24448 52554
rect 24520 52502 24572 52554
rect 24644 52502 24696 52554
rect 24768 52502 24820 52554
rect 24892 52502 24944 52554
rect 25016 52502 25068 52554
rect 25140 52502 25192 52554
rect 26574 52334 26626 52386
rect 9774 52222 9826 52274
rect 10558 52222 10610 52274
rect 11006 52222 11058 52274
rect 11790 52222 11842 52274
rect 19854 52222 19906 52274
rect 25454 52222 25506 52274
rect 30046 52222 30098 52274
rect 3614 52110 3666 52162
rect 4062 52110 4114 52162
rect 5182 52110 5234 52162
rect 5518 52110 5570 52162
rect 6078 52110 6130 52162
rect 11230 52110 11282 52162
rect 11454 52110 11506 52162
rect 12126 52110 12178 52162
rect 12574 52110 12626 52162
rect 20302 52110 20354 52162
rect 20414 52110 20466 52162
rect 20862 52110 20914 52162
rect 21198 52110 21250 52162
rect 21534 52110 21586 52162
rect 21870 52110 21922 52162
rect 22430 52110 22482 52162
rect 25902 52110 25954 52162
rect 30270 52110 30322 52162
rect 31166 52110 31218 52162
rect 31838 52110 31890 52162
rect 4398 51998 4450 52050
rect 4846 51998 4898 52050
rect 4958 51998 5010 52050
rect 10894 51998 10946 52050
rect 11902 51998 11954 52050
rect 19406 51998 19458 52050
rect 20190 51998 20242 52050
rect 25790 51998 25842 52050
rect 27582 51998 27634 52050
rect 30718 51998 30770 52050
rect 3278 51886 3330 51938
rect 8542 51886 8594 51938
rect 9214 51886 9266 51938
rect 13582 51886 13634 51938
rect 21422 51886 21474 51938
rect 24894 51886 24946 51938
rect 26910 51886 26962 51938
rect 30830 51886 30882 51938
rect 30942 51886 30994 51938
rect 34078 51886 34130 51938
rect 34862 51886 34914 51938
rect 14024 51718 14076 51770
rect 14148 51718 14200 51770
rect 14272 51718 14324 51770
rect 14396 51718 14448 51770
rect 14520 51718 14572 51770
rect 14644 51718 14696 51770
rect 14768 51718 14820 51770
rect 14892 51718 14944 51770
rect 15016 51718 15068 51770
rect 15140 51718 15192 51770
rect 34024 51718 34076 51770
rect 34148 51718 34200 51770
rect 34272 51718 34324 51770
rect 34396 51718 34448 51770
rect 34520 51718 34572 51770
rect 34644 51718 34696 51770
rect 34768 51718 34820 51770
rect 34892 51718 34944 51770
rect 35016 51718 35068 51770
rect 35140 51718 35192 51770
rect 4734 51550 4786 51602
rect 5294 51550 5346 51602
rect 11678 51550 11730 51602
rect 14254 51550 14306 51602
rect 22878 51550 22930 51602
rect 23438 51550 23490 51602
rect 23774 51550 23826 51602
rect 24222 51550 24274 51602
rect 25790 51550 25842 51602
rect 27022 51550 27074 51602
rect 27470 51550 27522 51602
rect 30942 51550 30994 51602
rect 7310 51438 7362 51490
rect 14814 51438 14866 51490
rect 15598 51438 15650 51490
rect 16270 51438 16322 51490
rect 28030 51438 28082 51490
rect 28478 51438 28530 51490
rect 32398 51438 32450 51490
rect 1822 51326 1874 51378
rect 2270 51338 2322 51390
rect 6078 51326 6130 51378
rect 8542 51326 8594 51378
rect 15374 51326 15426 51378
rect 15710 51326 15762 51378
rect 18286 51326 18338 51378
rect 19966 51326 20018 51378
rect 20302 51326 20354 51378
rect 27806 51326 27858 51378
rect 31950 51326 32002 51378
rect 33182 51326 33234 51378
rect 9662 51214 9714 51266
rect 14366 51214 14418 51266
rect 17614 51214 17666 51266
rect 17838 51214 17890 51266
rect 18174 51214 18226 51266
rect 25342 51214 25394 51266
rect 31614 51214 31666 51266
rect 17278 51102 17330 51154
rect 17614 51102 17666 51154
rect 25342 51102 25394 51154
rect 25902 51102 25954 51154
rect 4024 50934 4076 50986
rect 4148 50934 4200 50986
rect 4272 50934 4324 50986
rect 4396 50934 4448 50986
rect 4520 50934 4572 50986
rect 4644 50934 4696 50986
rect 4768 50934 4820 50986
rect 4892 50934 4944 50986
rect 5016 50934 5068 50986
rect 5140 50934 5192 50986
rect 24024 50934 24076 50986
rect 24148 50934 24200 50986
rect 24272 50934 24324 50986
rect 24396 50934 24448 50986
rect 24520 50934 24572 50986
rect 24644 50934 24696 50986
rect 24768 50934 24820 50986
rect 24892 50934 24944 50986
rect 25016 50934 25068 50986
rect 25140 50934 25192 50986
rect 5518 50766 5570 50818
rect 5742 50766 5794 50818
rect 6638 50766 6690 50818
rect 5742 50654 5794 50706
rect 6190 50654 6242 50706
rect 8318 50654 8370 50706
rect 9102 50654 9154 50706
rect 15262 50654 15314 50706
rect 16830 50654 16882 50706
rect 18622 50654 18674 50706
rect 19182 50654 19234 50706
rect 19854 50654 19906 50706
rect 23102 50654 23154 50706
rect 24334 50654 24386 50706
rect 24894 50654 24946 50706
rect 30718 50654 30770 50706
rect 31166 50654 31218 50706
rect 3838 50542 3890 50594
rect 4174 50542 4226 50594
rect 14814 50542 14866 50594
rect 15150 50542 15202 50594
rect 15934 50542 15986 50594
rect 16158 50542 16210 50594
rect 18174 50542 18226 50594
rect 19406 50542 19458 50594
rect 23886 50542 23938 50594
rect 31614 50542 31666 50594
rect 32174 50542 32226 50594
rect 4510 50430 4562 50482
rect 4958 50430 5010 50482
rect 6638 50430 6690 50482
rect 17278 50430 17330 50482
rect 19294 50430 19346 50482
rect 23438 50430 23490 50482
rect 34526 50430 34578 50482
rect 13918 50318 13970 50370
rect 35310 50318 35362 50370
rect 14024 50150 14076 50202
rect 14148 50150 14200 50202
rect 14272 50150 14324 50202
rect 14396 50150 14448 50202
rect 14520 50150 14572 50202
rect 14644 50150 14696 50202
rect 14768 50150 14820 50202
rect 14892 50150 14944 50202
rect 15016 50150 15068 50202
rect 15140 50150 15192 50202
rect 34024 50150 34076 50202
rect 34148 50150 34200 50202
rect 34272 50150 34324 50202
rect 34396 50150 34448 50202
rect 34520 50150 34572 50202
rect 34644 50150 34696 50202
rect 34768 50150 34820 50202
rect 34892 50150 34944 50202
rect 35016 50150 35068 50202
rect 35140 50150 35192 50202
rect 5518 49982 5570 50034
rect 7310 49982 7362 50034
rect 8654 49982 8706 50034
rect 9662 49982 9714 50034
rect 14590 49982 14642 50034
rect 18174 49982 18226 50034
rect 23998 49982 24050 50034
rect 7758 49870 7810 49922
rect 7870 49870 7922 49922
rect 13470 49870 13522 49922
rect 16606 49870 16658 49922
rect 18062 49870 18114 49922
rect 19518 49870 19570 49922
rect 26462 49870 26514 49922
rect 28142 49870 28194 49922
rect 28702 49870 28754 49922
rect 2830 49758 2882 49810
rect 7534 49758 7586 49810
rect 10782 49758 10834 49810
rect 11230 49758 11282 49810
rect 15374 49758 15426 49810
rect 15934 49758 15986 49810
rect 17950 49758 18002 49810
rect 18958 49758 19010 49810
rect 21982 49758 22034 49810
rect 22430 49758 22482 49810
rect 23550 49758 23602 49810
rect 23774 49758 23826 49810
rect 2494 49646 2546 49698
rect 3278 49646 3330 49698
rect 10334 49646 10386 49698
rect 15710 49646 15762 49698
rect 17502 49646 17554 49698
rect 22878 49646 22930 49698
rect 23438 49646 23490 49698
rect 27134 49646 27186 49698
rect 32174 49646 32226 49698
rect 32510 49646 32562 49698
rect 33182 49646 33234 49698
rect 8542 49534 8594 49586
rect 8878 49534 8930 49586
rect 14254 49534 14306 49586
rect 27582 49534 27634 49586
rect 27918 49534 27970 49586
rect 31950 49534 32002 49586
rect 32510 49534 32562 49586
rect 4024 49366 4076 49418
rect 4148 49366 4200 49418
rect 4272 49366 4324 49418
rect 4396 49366 4448 49418
rect 4520 49366 4572 49418
rect 4644 49366 4696 49418
rect 4768 49366 4820 49418
rect 4892 49366 4944 49418
rect 5016 49366 5068 49418
rect 5140 49366 5192 49418
rect 24024 49366 24076 49418
rect 24148 49366 24200 49418
rect 24272 49366 24324 49418
rect 24396 49366 24448 49418
rect 24520 49366 24572 49418
rect 24644 49366 24696 49418
rect 24768 49366 24820 49418
rect 24892 49366 24944 49418
rect 25016 49366 25068 49418
rect 25140 49366 25192 49418
rect 19294 49198 19346 49250
rect 26238 49198 26290 49250
rect 27694 49198 27746 49250
rect 28030 49198 28082 49250
rect 33518 49198 33570 49250
rect 11230 49086 11282 49138
rect 11678 49086 11730 49138
rect 15150 49086 15202 49138
rect 16494 49086 16546 49138
rect 20078 49086 20130 49138
rect 23550 49086 23602 49138
rect 31614 49086 31666 49138
rect 32174 49086 32226 49138
rect 6862 48974 6914 49026
rect 7310 48974 7362 49026
rect 11566 48974 11618 49026
rect 12238 48974 12290 49026
rect 12574 48974 12626 49026
rect 12910 48974 12962 49026
rect 13918 48974 13970 49026
rect 14254 48974 14306 49026
rect 14702 48974 14754 49026
rect 15598 48974 15650 49026
rect 15822 48974 15874 49026
rect 17054 48974 17106 49026
rect 17726 48974 17778 49026
rect 18398 48974 18450 49026
rect 18510 48974 18562 49026
rect 18846 48974 18898 49026
rect 22878 48974 22930 49026
rect 23326 48974 23378 49026
rect 24334 48974 24386 49026
rect 27022 48974 27074 49026
rect 31278 48974 31330 49026
rect 32846 48974 32898 49026
rect 33070 48974 33122 49026
rect 33630 48974 33682 49026
rect 5630 48862 5682 48914
rect 12798 48862 12850 48914
rect 13582 48862 13634 48914
rect 17950 48862 18002 48914
rect 18622 48862 18674 48914
rect 26910 48862 26962 48914
rect 31614 48862 31666 48914
rect 5742 48750 5794 48802
rect 9774 48750 9826 48802
rect 10334 48750 10386 48802
rect 11790 48750 11842 48802
rect 13694 48750 13746 48802
rect 19630 48750 19682 48802
rect 22318 48750 22370 48802
rect 28590 48750 28642 48802
rect 31838 48750 31890 48802
rect 33742 48750 33794 48802
rect 34302 48750 34354 48802
rect 14024 48582 14076 48634
rect 14148 48582 14200 48634
rect 14272 48582 14324 48634
rect 14396 48582 14448 48634
rect 14520 48582 14572 48634
rect 14644 48582 14696 48634
rect 14768 48582 14820 48634
rect 14892 48582 14944 48634
rect 15016 48582 15068 48634
rect 15140 48582 15192 48634
rect 34024 48582 34076 48634
rect 34148 48582 34200 48634
rect 34272 48582 34324 48634
rect 34396 48582 34448 48634
rect 34520 48582 34572 48634
rect 34644 48582 34696 48634
rect 34768 48582 34820 48634
rect 34892 48582 34944 48634
rect 35016 48582 35068 48634
rect 35140 48582 35192 48634
rect 6414 48414 6466 48466
rect 7534 48414 7586 48466
rect 7646 48414 7698 48466
rect 8542 48414 8594 48466
rect 11006 48414 11058 48466
rect 14590 48414 14642 48466
rect 15150 48414 15202 48466
rect 15486 48414 15538 48466
rect 24446 48414 24498 48466
rect 25342 48414 25394 48466
rect 26238 48414 26290 48466
rect 26686 48414 26738 48466
rect 30158 48414 30210 48466
rect 30830 48414 30882 48466
rect 32510 48414 32562 48466
rect 36430 48414 36482 48466
rect 5742 48302 5794 48354
rect 7870 48302 7922 48354
rect 19070 48302 19122 48354
rect 23662 48302 23714 48354
rect 2494 48190 2546 48242
rect 2942 48190 2994 48242
rect 6974 48190 7026 48242
rect 7422 48190 7474 48242
rect 9998 48190 10050 48242
rect 11678 48190 11730 48242
rect 12126 48190 12178 48242
rect 15934 48190 15986 48242
rect 18510 48190 18562 48242
rect 20974 48190 21026 48242
rect 21422 48190 21474 48242
rect 27358 48190 27410 48242
rect 27694 48190 27746 48242
rect 31166 48190 31218 48242
rect 31838 48190 31890 48242
rect 33070 48190 33122 48242
rect 33742 48190 33794 48242
rect 34078 48190 34130 48242
rect 3278 48078 3330 48130
rect 4622 48078 4674 48130
rect 8990 48078 9042 48130
rect 9886 48078 9938 48130
rect 16718 48078 16770 48130
rect 17838 48078 17890 48130
rect 18174 48078 18226 48130
rect 25790 48078 25842 48130
rect 9774 47966 9826 48018
rect 31614 47966 31666 48018
rect 32174 47966 32226 48018
rect 32398 47966 32450 48018
rect 33182 47966 33234 48018
rect 37214 47966 37266 48018
rect 4024 47798 4076 47850
rect 4148 47798 4200 47850
rect 4272 47798 4324 47850
rect 4396 47798 4448 47850
rect 4520 47798 4572 47850
rect 4644 47798 4696 47850
rect 4768 47798 4820 47850
rect 4892 47798 4944 47850
rect 5016 47798 5068 47850
rect 5140 47798 5192 47850
rect 24024 47798 24076 47850
rect 24148 47798 24200 47850
rect 24272 47798 24324 47850
rect 24396 47798 24448 47850
rect 24520 47798 24572 47850
rect 24644 47798 24696 47850
rect 24768 47798 24820 47850
rect 24892 47798 24944 47850
rect 25016 47798 25068 47850
rect 25140 47798 25192 47850
rect 9886 47630 9938 47682
rect 22990 47630 23042 47682
rect 3278 47518 3330 47570
rect 6302 47518 6354 47570
rect 13582 47518 13634 47570
rect 22094 47518 22146 47570
rect 29262 47518 29314 47570
rect 30718 47518 30770 47570
rect 31390 47518 31442 47570
rect 4622 47406 4674 47458
rect 4846 47406 4898 47458
rect 5182 47406 5234 47458
rect 7086 47406 7138 47458
rect 7758 47406 7810 47458
rect 11006 47406 11058 47458
rect 13694 47406 13746 47458
rect 14702 47406 14754 47458
rect 17614 47406 17666 47458
rect 22542 47406 22594 47458
rect 23214 47406 23266 47458
rect 23326 47406 23378 47458
rect 23662 47406 23714 47458
rect 24446 47406 24498 47458
rect 24782 47406 24834 47458
rect 31054 47406 31106 47458
rect 31278 47406 31330 47458
rect 31502 47406 31554 47458
rect 31726 47406 31778 47458
rect 32622 47406 32674 47458
rect 36318 47406 36370 47458
rect 37550 47406 37602 47458
rect 2606 47294 2658 47346
rect 3726 47294 3778 47346
rect 4062 47294 4114 47346
rect 6078 47294 6130 47346
rect 7422 47294 7474 47346
rect 9102 47294 9154 47346
rect 11230 47294 11282 47346
rect 13918 47294 13970 47346
rect 22878 47294 22930 47346
rect 23886 47294 23938 47346
rect 23998 47294 24050 47346
rect 30382 47294 30434 47346
rect 33182 47294 33234 47346
rect 35758 47294 35810 47346
rect 2158 47182 2210 47234
rect 2830 47182 2882 47234
rect 4958 47182 5010 47234
rect 7534 47182 7586 47234
rect 8094 47182 8146 47234
rect 9438 47182 9490 47234
rect 12350 47182 12402 47234
rect 13470 47182 13522 47234
rect 15598 47182 15650 47234
rect 21646 47182 21698 47234
rect 21982 47182 22034 47234
rect 22206 47182 22258 47234
rect 27134 47182 27186 47234
rect 27918 47182 27970 47234
rect 28366 47182 28418 47234
rect 30158 47182 30210 47234
rect 30606 47182 30658 47234
rect 32174 47182 32226 47234
rect 33630 47182 33682 47234
rect 37102 47182 37154 47234
rect 37998 47182 38050 47234
rect 14024 47014 14076 47066
rect 14148 47014 14200 47066
rect 14272 47014 14324 47066
rect 14396 47014 14448 47066
rect 14520 47014 14572 47066
rect 14644 47014 14696 47066
rect 14768 47014 14820 47066
rect 14892 47014 14944 47066
rect 15016 47014 15068 47066
rect 15140 47014 15192 47066
rect 34024 47014 34076 47066
rect 34148 47014 34200 47066
rect 34272 47014 34324 47066
rect 34396 47014 34448 47066
rect 34520 47014 34572 47066
rect 34644 47014 34696 47066
rect 34768 47014 34820 47066
rect 34892 47014 34944 47066
rect 35016 47014 35068 47066
rect 35140 47014 35192 47066
rect 4846 46846 4898 46898
rect 5518 46846 5570 46898
rect 6078 46846 6130 46898
rect 10782 46846 10834 46898
rect 15374 46846 15426 46898
rect 18958 46846 19010 46898
rect 25342 46846 25394 46898
rect 26462 46846 26514 46898
rect 27134 46846 27186 46898
rect 29598 46846 29650 46898
rect 30606 46846 30658 46898
rect 31166 46846 31218 46898
rect 31390 46846 31442 46898
rect 32174 46846 32226 46898
rect 34078 46846 34130 46898
rect 36542 46846 36594 46898
rect 5742 46734 5794 46786
rect 5854 46734 5906 46786
rect 6414 46734 6466 46786
rect 11454 46734 11506 46786
rect 28030 46734 28082 46786
rect 31614 46734 31666 46786
rect 34526 46734 34578 46786
rect 1822 46622 1874 46674
rect 2494 46622 2546 46674
rect 9998 46622 10050 46674
rect 11790 46622 11842 46674
rect 17502 46622 17554 46674
rect 19294 46622 19346 46674
rect 26238 46622 26290 46674
rect 26574 46622 26626 46674
rect 27918 46622 27970 46674
rect 28702 46622 28754 46674
rect 30942 46622 30994 46674
rect 32286 46622 32338 46674
rect 34190 46622 34242 46674
rect 34638 46622 34690 46674
rect 35198 46622 35250 46674
rect 35982 46622 36034 46674
rect 36206 46622 36258 46674
rect 37102 46622 37154 46674
rect 6974 46510 7026 46562
rect 7310 46510 7362 46562
rect 7758 46510 7810 46562
rect 8206 46510 8258 46562
rect 9102 46510 9154 46562
rect 13134 46510 13186 46562
rect 13582 46510 13634 46562
rect 14030 46510 14082 46562
rect 14478 46510 14530 46562
rect 23774 46510 23826 46562
rect 26014 46510 26066 46562
rect 27470 46510 27522 46562
rect 30158 46510 30210 46562
rect 31278 46510 31330 46562
rect 33182 46510 33234 46562
rect 33630 46510 33682 46562
rect 37550 46510 37602 46562
rect 37998 46510 38050 46562
rect 7758 46398 7810 46450
rect 7982 46398 8034 46450
rect 13470 46398 13522 46450
rect 14030 46398 14082 46450
rect 14478 46398 14530 46450
rect 29038 46398 29090 46450
rect 4024 46230 4076 46282
rect 4148 46230 4200 46282
rect 4272 46230 4324 46282
rect 4396 46230 4448 46282
rect 4520 46230 4572 46282
rect 4644 46230 4696 46282
rect 4768 46230 4820 46282
rect 4892 46230 4944 46282
rect 5016 46230 5068 46282
rect 5140 46230 5192 46282
rect 24024 46230 24076 46282
rect 24148 46230 24200 46282
rect 24272 46230 24324 46282
rect 24396 46230 24448 46282
rect 24520 46230 24572 46282
rect 24644 46230 24696 46282
rect 24768 46230 24820 46282
rect 24892 46230 24944 46282
rect 25016 46230 25068 46282
rect 25140 46230 25192 46282
rect 3838 46062 3890 46114
rect 17278 46062 17330 46114
rect 22318 46062 22370 46114
rect 30158 46062 30210 46114
rect 34750 46062 34802 46114
rect 2494 45950 2546 46002
rect 3278 45950 3330 46002
rect 5742 45950 5794 46002
rect 6862 45950 6914 46002
rect 12350 45950 12402 46002
rect 16046 45950 16098 46002
rect 16830 45950 16882 46002
rect 18286 45950 18338 46002
rect 20302 45950 20354 46002
rect 20750 45950 20802 46002
rect 22766 45950 22818 46002
rect 23550 45950 23602 46002
rect 24222 45950 24274 46002
rect 35534 45950 35586 46002
rect 37550 45950 37602 46002
rect 37998 45950 38050 46002
rect 2830 45838 2882 45890
rect 4174 45838 4226 45890
rect 7310 45838 7362 45890
rect 7646 45838 7698 45890
rect 10894 45838 10946 45890
rect 11790 45838 11842 45890
rect 13806 45838 13858 45890
rect 16606 45838 16658 45890
rect 17502 45838 17554 45890
rect 21310 45838 21362 45890
rect 21982 45838 22034 45890
rect 22206 45838 22258 45890
rect 23438 45838 23490 45890
rect 24782 45838 24834 45890
rect 25118 45838 25170 45890
rect 25678 45838 25730 45890
rect 30382 45838 30434 45890
rect 31054 45838 31106 45890
rect 33182 45838 33234 45890
rect 35758 45838 35810 45890
rect 37102 45838 37154 45890
rect 4398 45726 4450 45778
rect 4958 45726 5010 45778
rect 11454 45726 11506 45778
rect 13694 45726 13746 45778
rect 17838 45726 17890 45778
rect 18062 45726 18114 45778
rect 28702 45726 28754 45778
rect 30046 45726 30098 45778
rect 36990 45726 37042 45778
rect 6526 45614 6578 45666
rect 9998 45614 10050 45666
rect 13582 45614 13634 45666
rect 15374 45614 15426 45666
rect 18734 45614 18786 45666
rect 19294 45614 19346 45666
rect 21422 45614 21474 45666
rect 21534 45614 21586 45666
rect 22318 45614 22370 45666
rect 24110 45614 24162 45666
rect 24334 45614 24386 45666
rect 28142 45614 28194 45666
rect 29262 45614 29314 45666
rect 29710 45614 29762 45666
rect 35982 45614 36034 45666
rect 14024 45446 14076 45498
rect 14148 45446 14200 45498
rect 14272 45446 14324 45498
rect 14396 45446 14448 45498
rect 14520 45446 14572 45498
rect 14644 45446 14696 45498
rect 14768 45446 14820 45498
rect 14892 45446 14944 45498
rect 15016 45446 15068 45498
rect 15140 45446 15192 45498
rect 34024 45446 34076 45498
rect 34148 45446 34200 45498
rect 34272 45446 34324 45498
rect 34396 45446 34448 45498
rect 34520 45446 34572 45498
rect 34644 45446 34696 45498
rect 34768 45446 34820 45498
rect 34892 45446 34944 45498
rect 35016 45446 35068 45498
rect 35140 45446 35192 45498
rect 7646 45278 7698 45330
rect 10894 45278 10946 45330
rect 11342 45278 11394 45330
rect 12686 45278 12738 45330
rect 13134 45278 13186 45330
rect 13694 45278 13746 45330
rect 14926 45278 14978 45330
rect 16382 45278 16434 45330
rect 19630 45278 19682 45330
rect 22990 45278 23042 45330
rect 23550 45278 23602 45330
rect 24334 45278 24386 45330
rect 25902 45278 25954 45330
rect 27806 45278 27858 45330
rect 31166 45278 31218 45330
rect 5630 45166 5682 45218
rect 6526 45166 6578 45218
rect 11790 45166 11842 45218
rect 16718 45166 16770 45218
rect 17390 45166 17442 45218
rect 34190 45166 34242 45218
rect 34414 45166 34466 45218
rect 34862 45166 34914 45218
rect 36990 45166 37042 45218
rect 2830 45054 2882 45106
rect 6414 45054 6466 45106
rect 7646 45054 7698 45106
rect 8206 45054 8258 45106
rect 8430 45054 8482 45106
rect 9662 45054 9714 45106
rect 13806 45054 13858 45106
rect 14142 45054 14194 45106
rect 14478 45054 14530 45106
rect 15150 45054 15202 45106
rect 17726 45054 17778 45106
rect 17950 45054 18002 45106
rect 18286 45054 18338 45106
rect 20078 45054 20130 45106
rect 20526 45054 20578 45106
rect 25790 45054 25842 45106
rect 26126 45054 26178 45106
rect 26350 45054 26402 45106
rect 27694 45054 27746 45106
rect 30830 45054 30882 45106
rect 34638 45054 34690 45106
rect 35422 45054 35474 45106
rect 36318 45054 36370 45106
rect 2494 44942 2546 44994
rect 3278 44942 3330 44994
rect 5294 44942 5346 44994
rect 7310 44942 7362 44994
rect 8878 44942 8930 44994
rect 10446 44942 10498 44994
rect 14030 44942 14082 44994
rect 14814 44942 14866 44994
rect 15934 44942 15986 44994
rect 16830 44942 16882 44994
rect 17502 44942 17554 44994
rect 19294 44942 19346 44994
rect 19518 44942 19570 44994
rect 23886 44942 23938 44994
rect 25454 44942 25506 44994
rect 27246 44942 27298 44994
rect 27582 44942 27634 44994
rect 29934 44942 29986 44994
rect 30606 44942 30658 44994
rect 32510 44942 32562 44994
rect 33854 44942 33906 44994
rect 5966 44830 6018 44882
rect 7982 44830 8034 44882
rect 10446 44830 10498 44882
rect 11454 44830 11506 44882
rect 18286 44830 18338 44882
rect 18622 44830 18674 44882
rect 34750 44830 34802 44882
rect 37662 44830 37714 44882
rect 4024 44662 4076 44714
rect 4148 44662 4200 44714
rect 4272 44662 4324 44714
rect 4396 44662 4448 44714
rect 4520 44662 4572 44714
rect 4644 44662 4696 44714
rect 4768 44662 4820 44714
rect 4892 44662 4944 44714
rect 5016 44662 5068 44714
rect 5140 44662 5192 44714
rect 24024 44662 24076 44714
rect 24148 44662 24200 44714
rect 24272 44662 24324 44714
rect 24396 44662 24448 44714
rect 24520 44662 24572 44714
rect 24644 44662 24696 44714
rect 24768 44662 24820 44714
rect 24892 44662 24944 44714
rect 25016 44662 25068 44714
rect 25140 44662 25192 44714
rect 7646 44494 7698 44546
rect 8206 44494 8258 44546
rect 8542 44494 8594 44546
rect 17054 44494 17106 44546
rect 35982 44494 36034 44546
rect 6750 44382 6802 44434
rect 7534 44382 7586 44434
rect 9662 44382 9714 44434
rect 10558 44382 10610 44434
rect 12238 44382 12290 44434
rect 12910 44382 12962 44434
rect 17614 44382 17666 44434
rect 18510 44382 18562 44434
rect 18622 44382 18674 44434
rect 19070 44382 19122 44434
rect 20302 44382 20354 44434
rect 21758 44382 21810 44434
rect 34190 44382 34242 44434
rect 4174 44270 4226 44322
rect 7310 44270 7362 44322
rect 8318 44270 8370 44322
rect 8766 44270 8818 44322
rect 13470 44270 13522 44322
rect 14030 44270 14082 44322
rect 17726 44270 17778 44322
rect 18062 44270 18114 44322
rect 21310 44270 21362 44322
rect 21982 44270 22034 44322
rect 34526 44270 34578 44322
rect 35310 44270 35362 44322
rect 37438 44270 37490 44322
rect 37550 44270 37602 44322
rect 4398 44158 4450 44210
rect 4958 44158 5010 44210
rect 6414 44158 6466 44210
rect 11342 44158 11394 44210
rect 11454 44158 11506 44210
rect 17614 44158 17666 44210
rect 20414 44158 20466 44210
rect 21534 44158 21586 44210
rect 34638 44158 34690 44210
rect 34862 44158 34914 44210
rect 35198 44158 35250 44210
rect 37662 44158 37714 44210
rect 3838 44046 3890 44098
rect 6638 44046 6690 44098
rect 9214 44046 9266 44098
rect 10110 44046 10162 44098
rect 11006 44046 11058 44098
rect 11678 44046 11730 44098
rect 16270 44046 16322 44098
rect 17950 44046 18002 44098
rect 18958 44046 19010 44098
rect 19742 44046 19794 44098
rect 20190 44046 20242 44098
rect 23662 44046 23714 44098
rect 24110 44046 24162 44098
rect 33854 44046 33906 44098
rect 36318 44046 36370 44098
rect 36990 44046 37042 44098
rect 14024 43878 14076 43930
rect 14148 43878 14200 43930
rect 14272 43878 14324 43930
rect 14396 43878 14448 43930
rect 14520 43878 14572 43930
rect 14644 43878 14696 43930
rect 14768 43878 14820 43930
rect 14892 43878 14944 43930
rect 15016 43878 15068 43930
rect 15140 43878 15192 43930
rect 34024 43878 34076 43930
rect 34148 43878 34200 43930
rect 34272 43878 34324 43930
rect 34396 43878 34448 43930
rect 34520 43878 34572 43930
rect 34644 43878 34696 43930
rect 34768 43878 34820 43930
rect 34892 43878 34944 43930
rect 35016 43878 35068 43930
rect 35140 43878 35192 43930
rect 4734 43710 4786 43762
rect 5294 43710 5346 43762
rect 6078 43710 6130 43762
rect 8766 43710 8818 43762
rect 10670 43710 10722 43762
rect 15822 43710 15874 43762
rect 16718 43710 16770 43762
rect 17614 43710 17666 43762
rect 17726 43710 17778 43762
rect 18734 43710 18786 43762
rect 18846 43710 18898 43762
rect 19966 43710 20018 43762
rect 20414 43710 20466 43762
rect 20974 43710 21026 43762
rect 30270 43710 30322 43762
rect 35198 43710 35250 43762
rect 36542 43710 36594 43762
rect 5630 43598 5682 43650
rect 12350 43598 12402 43650
rect 12798 43598 12850 43650
rect 13918 43598 13970 43650
rect 14254 43598 14306 43650
rect 15486 43598 15538 43650
rect 16494 43598 16546 43650
rect 19742 43598 19794 43650
rect 29150 43598 29202 43650
rect 29822 43598 29874 43650
rect 35870 43598 35922 43650
rect 36430 43598 36482 43650
rect 1822 43486 1874 43538
rect 2270 43486 2322 43538
rect 8542 43486 8594 43538
rect 11454 43486 11506 43538
rect 12574 43486 12626 43538
rect 14142 43486 14194 43538
rect 14478 43486 14530 43538
rect 16158 43486 16210 43538
rect 16382 43486 16434 43538
rect 16606 43486 16658 43538
rect 17390 43486 17442 43538
rect 17838 43486 17890 43538
rect 18062 43486 18114 43538
rect 18398 43486 18450 43538
rect 18622 43486 18674 43538
rect 18958 43486 19010 43538
rect 19294 43486 19346 43538
rect 30158 43486 30210 43538
rect 30494 43486 30546 43538
rect 36766 43486 36818 43538
rect 6974 43374 7026 43426
rect 8206 43374 8258 43426
rect 9998 43374 10050 43426
rect 11006 43374 11058 43426
rect 11790 43374 11842 43426
rect 13358 43374 13410 43426
rect 19854 43374 19906 43426
rect 21422 43374 21474 43426
rect 26798 43374 26850 43426
rect 30942 43374 30994 43426
rect 31726 43374 31778 43426
rect 33742 43374 33794 43426
rect 34638 43374 34690 43426
rect 37662 43374 37714 43426
rect 6750 43262 6802 43314
rect 7086 43262 7138 43314
rect 8878 43262 8930 43314
rect 12238 43262 12290 43314
rect 29486 43262 29538 43314
rect 29598 43262 29650 43314
rect 31950 43262 32002 43314
rect 32286 43262 32338 43314
rect 37550 43262 37602 43314
rect 4024 43094 4076 43146
rect 4148 43094 4200 43146
rect 4272 43094 4324 43146
rect 4396 43094 4448 43146
rect 4520 43094 4572 43146
rect 4644 43094 4696 43146
rect 4768 43094 4820 43146
rect 4892 43094 4944 43146
rect 5016 43094 5068 43146
rect 5140 43094 5192 43146
rect 24024 43094 24076 43146
rect 24148 43094 24200 43146
rect 24272 43094 24324 43146
rect 24396 43094 24448 43146
rect 24520 43094 24572 43146
rect 24644 43094 24696 43146
rect 24768 43094 24820 43146
rect 24892 43094 24944 43146
rect 25016 43094 25068 43146
rect 25140 43094 25192 43146
rect 5742 42926 5794 42978
rect 13582 42926 13634 42978
rect 14030 42926 14082 42978
rect 19854 42926 19906 42978
rect 21758 42926 21810 42978
rect 6078 42814 6130 42866
rect 7422 42814 7474 42866
rect 8206 42814 8258 42866
rect 8542 42814 8594 42866
rect 9102 42814 9154 42866
rect 10110 42814 10162 42866
rect 10670 42814 10722 42866
rect 12686 42814 12738 42866
rect 14030 42814 14082 42866
rect 16046 42814 16098 42866
rect 25006 42814 25058 42866
rect 26238 42814 26290 42866
rect 30270 42814 30322 42866
rect 35198 42814 35250 42866
rect 9214 42702 9266 42754
rect 9662 42702 9714 42754
rect 10334 42702 10386 42754
rect 11678 42702 11730 42754
rect 12014 42702 12066 42754
rect 16382 42702 16434 42754
rect 16718 42702 16770 42754
rect 20750 42702 20802 42754
rect 22318 42702 22370 42754
rect 26574 42702 26626 42754
rect 26798 42702 26850 42754
rect 27022 42702 27074 42754
rect 27582 42702 27634 42754
rect 30830 42702 30882 42754
rect 31054 42702 31106 42754
rect 31390 42702 31442 42754
rect 33182 42702 33234 42754
rect 34302 42702 34354 42754
rect 34414 42702 34466 42754
rect 34974 42702 35026 42754
rect 36206 42702 36258 42754
rect 36990 42702 37042 42754
rect 2830 42590 2882 42642
rect 3166 42590 3218 42642
rect 6302 42590 6354 42642
rect 6750 42590 6802 42642
rect 12126 42590 12178 42642
rect 13582 42590 13634 42642
rect 22542 42590 22594 42642
rect 24558 42590 24610 42642
rect 32398 42590 32450 42642
rect 35086 42590 35138 42642
rect 36430 42590 36482 42642
rect 37998 42590 38050 42642
rect 2606 42478 2658 42530
rect 5070 42478 5122 42530
rect 8654 42478 8706 42530
rect 8990 42478 9042 42530
rect 19294 42478 19346 42530
rect 20190 42478 20242 42530
rect 21422 42478 21474 42530
rect 26686 42478 26738 42530
rect 29934 42478 29986 42530
rect 32846 42478 32898 42530
rect 37102 42478 37154 42530
rect 37326 42478 37378 42530
rect 37662 42478 37714 42530
rect 37886 42478 37938 42530
rect 14024 42310 14076 42362
rect 14148 42310 14200 42362
rect 14272 42310 14324 42362
rect 14396 42310 14448 42362
rect 14520 42310 14572 42362
rect 14644 42310 14696 42362
rect 14768 42310 14820 42362
rect 14892 42310 14944 42362
rect 15016 42310 15068 42362
rect 15140 42310 15192 42362
rect 34024 42310 34076 42362
rect 34148 42310 34200 42362
rect 34272 42310 34324 42362
rect 34396 42310 34448 42362
rect 34520 42310 34572 42362
rect 34644 42310 34696 42362
rect 34768 42310 34820 42362
rect 34892 42310 34944 42362
rect 35016 42310 35068 42362
rect 35140 42310 35192 42362
rect 7198 42142 7250 42194
rect 8654 42142 8706 42194
rect 10558 42142 10610 42194
rect 13806 42142 13858 42194
rect 17838 42142 17890 42194
rect 19070 42142 19122 42194
rect 23662 42142 23714 42194
rect 29934 42142 29986 42194
rect 30494 42142 30546 42194
rect 8878 42030 8930 42082
rect 9662 42030 9714 42082
rect 12686 42030 12738 42082
rect 17726 42030 17778 42082
rect 26014 42030 26066 42082
rect 26126 42030 26178 42082
rect 32062 42030 32114 42082
rect 33518 42030 33570 42082
rect 35422 42030 35474 42082
rect 8430 41918 8482 41970
rect 8990 41918 9042 41970
rect 9550 41918 9602 41970
rect 11566 41918 11618 41970
rect 20974 41918 21026 41970
rect 21422 41918 21474 41970
rect 24446 41918 24498 41970
rect 25342 41918 25394 41970
rect 25790 41918 25842 41970
rect 27022 41918 27074 41970
rect 27358 41918 27410 41970
rect 31054 41918 31106 41970
rect 32174 41918 32226 41970
rect 33294 41918 33346 41970
rect 33854 41918 33906 41970
rect 34750 41918 34802 41970
rect 35086 41918 35138 41970
rect 37326 41918 37378 41970
rect 37774 41918 37826 41970
rect 18398 41806 18450 41858
rect 19966 41806 20018 41858
rect 31726 41806 31778 41858
rect 35534 41806 35586 41858
rect 25454 41694 25506 41746
rect 26574 41694 26626 41746
rect 33182 41694 33234 41746
rect 37774 41694 37826 41746
rect 38110 41694 38162 41746
rect 4024 41526 4076 41578
rect 4148 41526 4200 41578
rect 4272 41526 4324 41578
rect 4396 41526 4448 41578
rect 4520 41526 4572 41578
rect 4644 41526 4696 41578
rect 4768 41526 4820 41578
rect 4892 41526 4944 41578
rect 5016 41526 5068 41578
rect 5140 41526 5192 41578
rect 24024 41526 24076 41578
rect 24148 41526 24200 41578
rect 24272 41526 24324 41578
rect 24396 41526 24448 41578
rect 24520 41526 24572 41578
rect 24644 41526 24696 41578
rect 24768 41526 24820 41578
rect 24892 41526 24944 41578
rect 25016 41526 25068 41578
rect 25140 41526 25192 41578
rect 11118 41358 11170 41410
rect 11342 41358 11394 41410
rect 11902 41358 11954 41410
rect 12350 41358 12402 41410
rect 12574 41358 12626 41410
rect 17502 41358 17554 41410
rect 26462 41358 26514 41410
rect 26686 41358 26738 41410
rect 28142 41358 28194 41410
rect 29038 41358 29090 41410
rect 29822 41358 29874 41410
rect 31614 41358 31666 41410
rect 32174 41358 32226 41410
rect 3278 41246 3330 41298
rect 9550 41246 9602 41298
rect 18398 41246 18450 41298
rect 18734 41246 18786 41298
rect 20750 41246 20802 41298
rect 21534 41246 21586 41298
rect 22654 41246 22706 41298
rect 26014 41246 26066 41298
rect 27246 41246 27298 41298
rect 27806 41246 27858 41298
rect 28590 41246 28642 41298
rect 29262 41246 29314 41298
rect 29710 41246 29762 41298
rect 30270 41246 30322 41298
rect 30606 41246 30658 41298
rect 8318 41134 8370 41186
rect 8542 41134 8594 41186
rect 9438 41134 9490 41186
rect 9998 41134 10050 41186
rect 10670 41134 10722 41186
rect 12014 41134 12066 41186
rect 21870 41134 21922 41186
rect 24670 41134 24722 41186
rect 24782 41134 24834 41186
rect 25454 41134 25506 41186
rect 25790 41134 25842 41186
rect 26910 41134 26962 41186
rect 27134 41134 27186 41186
rect 27358 41134 27410 41186
rect 28478 41134 28530 41186
rect 30718 41134 30770 41186
rect 31726 41134 31778 41186
rect 32062 41134 32114 41186
rect 35310 41134 35362 41186
rect 35758 41134 35810 41186
rect 36094 41134 36146 41186
rect 37102 41134 37154 41186
rect 8094 41022 8146 41074
rect 8206 41022 8258 41074
rect 8990 41022 9042 41074
rect 10558 41022 10610 41074
rect 11790 41022 11842 41074
rect 17614 41022 17666 41074
rect 22094 41022 22146 41074
rect 24558 41022 24610 41074
rect 25230 41022 25282 41074
rect 31390 41022 31442 41074
rect 32734 41022 32786 41074
rect 33630 41022 33682 41074
rect 36318 41022 36370 41074
rect 37214 41022 37266 41074
rect 37774 41022 37826 41074
rect 2606 40910 2658 40962
rect 2830 40910 2882 40962
rect 5742 40910 5794 40962
rect 6302 40910 6354 40962
rect 7534 40910 7586 40962
rect 7982 40910 8034 40962
rect 11454 40910 11506 40962
rect 22990 40910 23042 40962
rect 23886 40910 23938 40962
rect 24334 40910 24386 40962
rect 24446 40910 24498 40962
rect 26126 40910 26178 40962
rect 27918 40910 27970 40962
rect 35870 40910 35922 40962
rect 35982 40910 36034 40962
rect 37326 40910 37378 40962
rect 14024 40742 14076 40794
rect 14148 40742 14200 40794
rect 14272 40742 14324 40794
rect 14396 40742 14448 40794
rect 14520 40742 14572 40794
rect 14644 40742 14696 40794
rect 14768 40742 14820 40794
rect 14892 40742 14944 40794
rect 15016 40742 15068 40794
rect 15140 40742 15192 40794
rect 34024 40742 34076 40794
rect 34148 40742 34200 40794
rect 34272 40742 34324 40794
rect 34396 40742 34448 40794
rect 34520 40742 34572 40794
rect 34644 40742 34696 40794
rect 34768 40742 34820 40794
rect 34892 40742 34944 40794
rect 35016 40742 35068 40794
rect 35140 40742 35192 40794
rect 4734 40574 4786 40626
rect 5294 40574 5346 40626
rect 7422 40574 7474 40626
rect 7982 40574 8034 40626
rect 8878 40574 8930 40626
rect 11118 40574 11170 40626
rect 14142 40574 14194 40626
rect 22206 40574 22258 40626
rect 29038 40574 29090 40626
rect 33630 40574 33682 40626
rect 37662 40574 37714 40626
rect 5742 40462 5794 40514
rect 6638 40462 6690 40514
rect 8318 40462 8370 40514
rect 9550 40462 9602 40514
rect 23214 40462 23266 40514
rect 23662 40462 23714 40514
rect 31054 40462 31106 40514
rect 34078 40462 34130 40514
rect 37886 40462 37938 40514
rect 1822 40350 1874 40402
rect 2270 40350 2322 40402
rect 6750 40350 6802 40402
rect 9662 40350 9714 40402
rect 9998 40350 10050 40402
rect 11230 40350 11282 40402
rect 11790 40350 11842 40402
rect 15038 40350 15090 40402
rect 15934 40350 15986 40402
rect 22990 40350 23042 40402
rect 25902 40350 25954 40402
rect 26462 40350 26514 40402
rect 30606 40350 30658 40402
rect 32174 40350 32226 40402
rect 33070 40350 33122 40402
rect 34190 40350 34242 40402
rect 35086 40350 35138 40402
rect 36318 40350 36370 40402
rect 37998 40350 38050 40402
rect 15486 40238 15538 40290
rect 33294 40238 33346 40290
rect 6078 40126 6130 40178
rect 7310 40126 7362 40178
rect 8206 40126 8258 40178
rect 22654 40126 22706 40178
rect 30046 40126 30098 40178
rect 32398 40126 32450 40178
rect 4024 39958 4076 40010
rect 4148 39958 4200 40010
rect 4272 39958 4324 40010
rect 4396 39958 4448 40010
rect 4520 39958 4572 40010
rect 4644 39958 4696 40010
rect 4768 39958 4820 40010
rect 4892 39958 4944 40010
rect 5016 39958 5068 40010
rect 5140 39958 5192 40010
rect 24024 39958 24076 40010
rect 24148 39958 24200 40010
rect 24272 39958 24324 40010
rect 24396 39958 24448 40010
rect 24520 39958 24572 40010
rect 24644 39958 24696 40010
rect 24768 39958 24820 40010
rect 24892 39958 24944 40010
rect 25016 39958 25068 40010
rect 25140 39958 25192 40010
rect 3726 39790 3778 39842
rect 4062 39790 4114 39842
rect 15150 39790 15202 39842
rect 18958 39790 19010 39842
rect 19630 39790 19682 39842
rect 38222 39790 38274 39842
rect 5742 39678 5794 39730
rect 9438 39678 9490 39730
rect 10782 39678 10834 39730
rect 11230 39678 11282 39730
rect 14926 39678 14978 39730
rect 19182 39678 19234 39730
rect 19630 39678 19682 39730
rect 26126 39678 26178 39730
rect 29486 39678 29538 39730
rect 29822 39678 29874 39730
rect 30270 39678 30322 39730
rect 31054 39678 31106 39730
rect 31502 39678 31554 39730
rect 31950 39678 32002 39730
rect 34638 39678 34690 39730
rect 37102 39678 37154 39730
rect 3278 39566 3330 39618
rect 6526 39566 6578 39618
rect 7310 39566 7362 39618
rect 9774 39566 9826 39618
rect 9998 39566 10050 39618
rect 18174 39566 18226 39618
rect 18622 39566 18674 39618
rect 21758 39566 21810 39618
rect 22318 39566 22370 39618
rect 25678 39566 25730 39618
rect 30158 39566 30210 39618
rect 32510 39566 32562 39618
rect 34526 39566 34578 39618
rect 37214 39566 37266 39618
rect 37550 39566 37602 39618
rect 4286 39454 4338 39506
rect 4846 39454 4898 39506
rect 7534 39454 7586 39506
rect 7870 39454 7922 39506
rect 24558 39454 24610 39506
rect 25342 39454 25394 39506
rect 32174 39454 32226 39506
rect 32622 39454 32674 39506
rect 35646 39454 35698 39506
rect 36990 39454 37042 39506
rect 37886 39454 37938 39506
rect 2494 39342 2546 39394
rect 2718 39342 2770 39394
rect 6974 39342 7026 39394
rect 8990 39342 9042 39394
rect 9438 39342 9490 39394
rect 9550 39342 9602 39394
rect 15822 39342 15874 39394
rect 38110 39342 38162 39394
rect 14024 39174 14076 39226
rect 14148 39174 14200 39226
rect 14272 39174 14324 39226
rect 14396 39174 14448 39226
rect 14520 39174 14572 39226
rect 14644 39174 14696 39226
rect 14768 39174 14820 39226
rect 14892 39174 14944 39226
rect 15016 39174 15068 39226
rect 15140 39174 15192 39226
rect 34024 39174 34076 39226
rect 34148 39174 34200 39226
rect 34272 39174 34324 39226
rect 34396 39174 34448 39226
rect 34520 39174 34572 39226
rect 34644 39174 34696 39226
rect 34768 39174 34820 39226
rect 34892 39174 34944 39226
rect 35016 39174 35068 39226
rect 35140 39174 35192 39226
rect 3166 39006 3218 39058
rect 7310 39006 7362 39058
rect 8094 39006 8146 39058
rect 8654 39006 8706 39058
rect 14142 39006 14194 39058
rect 14926 39006 14978 39058
rect 15486 39006 15538 39058
rect 17838 39006 17890 39058
rect 18398 39006 18450 39058
rect 19070 39006 19122 39058
rect 33294 39006 33346 39058
rect 33742 39006 33794 39058
rect 34302 39006 34354 39058
rect 16718 38894 16770 38946
rect 17614 38894 17666 38946
rect 18286 38894 18338 38946
rect 22766 38894 22818 38946
rect 24110 38894 24162 38946
rect 32286 38894 32338 38946
rect 32398 38894 32450 38946
rect 34190 38894 34242 38946
rect 35086 38894 35138 38946
rect 2830 38782 2882 38834
rect 4622 38782 4674 38834
rect 5070 38782 5122 38834
rect 11342 38782 11394 38834
rect 11902 38782 11954 38834
rect 16158 38782 16210 38834
rect 17390 38782 17442 38834
rect 17950 38782 18002 38834
rect 19518 38782 19570 38834
rect 22318 38782 22370 38834
rect 23550 38782 23602 38834
rect 32622 38782 32674 38834
rect 33518 38782 33570 38834
rect 33966 38782 34018 38834
rect 34750 38782 34802 38834
rect 37662 38782 37714 38834
rect 38222 38782 38274 38834
rect 2494 38670 2546 38722
rect 16494 38670 16546 38722
rect 16830 38670 16882 38722
rect 21982 38670 22034 38722
rect 23214 38670 23266 38722
rect 35982 38670 36034 38722
rect 4024 38390 4076 38442
rect 4148 38390 4200 38442
rect 4272 38390 4324 38442
rect 4396 38390 4448 38442
rect 4520 38390 4572 38442
rect 4644 38390 4696 38442
rect 4768 38390 4820 38442
rect 4892 38390 4944 38442
rect 5016 38390 5068 38442
rect 5140 38390 5192 38442
rect 24024 38390 24076 38442
rect 24148 38390 24200 38442
rect 24272 38390 24324 38442
rect 24396 38390 24448 38442
rect 24520 38390 24572 38442
rect 24644 38390 24696 38442
rect 24768 38390 24820 38442
rect 24892 38390 24944 38442
rect 25016 38390 25068 38442
rect 25140 38390 25192 38442
rect 5854 38222 5906 38274
rect 6190 38222 6242 38274
rect 18734 38222 18786 38274
rect 33182 38222 33234 38274
rect 33630 38222 33682 38274
rect 35758 38222 35810 38274
rect 24894 38110 24946 38162
rect 33742 38110 33794 38162
rect 35310 38110 35362 38162
rect 36094 38110 36146 38162
rect 37214 38110 37266 38162
rect 37998 38110 38050 38162
rect 15262 37998 15314 38050
rect 15710 37998 15762 38050
rect 19630 37998 19682 38050
rect 31726 37998 31778 38050
rect 32062 37998 32114 38050
rect 33854 37998 33906 38050
rect 35198 37998 35250 38050
rect 36206 37998 36258 38050
rect 37438 37998 37490 38050
rect 37774 37998 37826 38050
rect 6414 37886 6466 37938
rect 6974 37886 7026 37938
rect 9662 37886 9714 37938
rect 19854 37886 19906 37938
rect 20190 37886 20242 37938
rect 31390 37886 31442 37938
rect 32510 37886 32562 37938
rect 32846 37886 32898 37938
rect 8430 37774 8482 37826
rect 8878 37774 8930 37826
rect 9774 37774 9826 37826
rect 9998 37774 10050 37826
rect 11678 37774 11730 37826
rect 13694 37774 13746 37826
rect 17950 37774 18002 37826
rect 19294 37774 19346 37826
rect 26686 37774 26738 37826
rect 27806 37774 27858 37826
rect 28254 37774 28306 37826
rect 31054 37774 31106 37826
rect 31726 37774 31778 37826
rect 32174 37774 32226 37826
rect 32398 37774 32450 37826
rect 33070 37774 33122 37826
rect 37102 37774 37154 37826
rect 37326 37774 37378 37826
rect 14024 37606 14076 37658
rect 14148 37606 14200 37658
rect 14272 37606 14324 37658
rect 14396 37606 14448 37658
rect 14520 37606 14572 37658
rect 14644 37606 14696 37658
rect 14768 37606 14820 37658
rect 14892 37606 14944 37658
rect 15016 37606 15068 37658
rect 15140 37606 15192 37658
rect 34024 37606 34076 37658
rect 34148 37606 34200 37658
rect 34272 37606 34324 37658
rect 34396 37606 34448 37658
rect 34520 37606 34572 37658
rect 34644 37606 34696 37658
rect 34768 37606 34820 37658
rect 34892 37606 34944 37658
rect 35016 37606 35068 37658
rect 35140 37606 35192 37658
rect 9102 37438 9154 37490
rect 12350 37438 12402 37490
rect 13358 37438 13410 37490
rect 14814 37438 14866 37490
rect 16158 37438 16210 37490
rect 16718 37438 16770 37490
rect 17838 37438 17890 37490
rect 21534 37438 21586 37490
rect 22094 37438 22146 37490
rect 24670 37438 24722 37490
rect 31166 37438 31218 37490
rect 31950 37438 32002 37490
rect 35310 37438 35362 37490
rect 37774 37438 37826 37490
rect 3166 37326 3218 37378
rect 8766 37326 8818 37378
rect 8878 37326 8930 37378
rect 9998 37326 10050 37378
rect 12574 37326 12626 37378
rect 12910 37326 12962 37378
rect 14030 37326 14082 37378
rect 22430 37326 22482 37378
rect 25902 37326 25954 37378
rect 26462 37326 26514 37378
rect 27022 37326 27074 37378
rect 27582 37326 27634 37378
rect 28030 37326 28082 37378
rect 34190 37326 34242 37378
rect 36206 37326 36258 37378
rect 2830 37214 2882 37266
rect 10222 37214 10274 37266
rect 12238 37214 12290 37266
rect 12798 37214 12850 37266
rect 15038 37214 15090 37266
rect 16494 37214 16546 37266
rect 17502 37214 17554 37266
rect 17726 37214 17778 37266
rect 18062 37214 18114 37266
rect 18622 37214 18674 37266
rect 19070 37214 19122 37266
rect 25678 37214 25730 37266
rect 27358 37214 27410 37266
rect 27806 37214 27858 37266
rect 28254 37214 28306 37266
rect 28926 37214 28978 37266
rect 35198 37214 35250 37266
rect 35646 37214 35698 37266
rect 37662 37214 37714 37266
rect 2494 37102 2546 37154
rect 11454 37102 11506 37154
rect 11902 37102 11954 37154
rect 16830 37102 16882 37154
rect 22878 37102 22930 37154
rect 24110 37102 24162 37154
rect 27694 37102 27746 37154
rect 10558 36990 10610 37042
rect 25342 36990 25394 37042
rect 37886 36990 37938 37042
rect 38110 36990 38162 37042
rect 4024 36822 4076 36874
rect 4148 36822 4200 36874
rect 4272 36822 4324 36874
rect 4396 36822 4448 36874
rect 4520 36822 4572 36874
rect 4644 36822 4696 36874
rect 4768 36822 4820 36874
rect 4892 36822 4944 36874
rect 5016 36822 5068 36874
rect 5140 36822 5192 36874
rect 24024 36822 24076 36874
rect 24148 36822 24200 36874
rect 24272 36822 24324 36874
rect 24396 36822 24448 36874
rect 24520 36822 24572 36874
rect 24644 36822 24696 36874
rect 24768 36822 24820 36874
rect 24892 36822 24944 36874
rect 25016 36822 25068 36874
rect 25140 36822 25192 36874
rect 11902 36654 11954 36706
rect 12910 36654 12962 36706
rect 35422 36654 35474 36706
rect 6414 36542 6466 36594
rect 8766 36542 8818 36594
rect 10894 36542 10946 36594
rect 12126 36542 12178 36594
rect 12350 36542 12402 36594
rect 14254 36542 14306 36594
rect 23326 36542 23378 36594
rect 26686 36542 26738 36594
rect 29598 36542 29650 36594
rect 33294 36542 33346 36594
rect 35646 36542 35698 36594
rect 6190 36430 6242 36482
rect 8990 36430 9042 36482
rect 10334 36430 10386 36482
rect 11902 36430 11954 36482
rect 13582 36430 13634 36482
rect 21534 36430 21586 36482
rect 24334 36430 24386 36482
rect 27694 36430 27746 36482
rect 29038 36430 29090 36482
rect 29486 36430 29538 36482
rect 30382 36430 30434 36482
rect 31166 36430 31218 36482
rect 31950 36430 32002 36482
rect 33630 36430 33682 36482
rect 33742 36430 33794 36482
rect 34526 36430 34578 36482
rect 35422 36430 35474 36482
rect 36542 36430 36594 36482
rect 37550 36430 37602 36482
rect 4622 36318 4674 36370
rect 4846 36318 4898 36370
rect 5182 36318 5234 36370
rect 5854 36318 5906 36370
rect 8766 36318 8818 36370
rect 9550 36318 9602 36370
rect 10110 36318 10162 36370
rect 11342 36318 11394 36370
rect 13694 36318 13746 36370
rect 14814 36318 14866 36370
rect 28030 36318 28082 36370
rect 28478 36318 28530 36370
rect 31614 36318 31666 36370
rect 31726 36318 31778 36370
rect 32174 36318 32226 36370
rect 32622 36318 32674 36370
rect 36990 36318 37042 36370
rect 37326 36318 37378 36370
rect 37998 36318 38050 36370
rect 38222 36318 38274 36370
rect 2606 36206 2658 36258
rect 2830 36206 2882 36258
rect 3166 36206 3218 36258
rect 4062 36206 4114 36258
rect 4958 36206 5010 36258
rect 7534 36206 7586 36258
rect 8318 36206 8370 36258
rect 9774 36206 9826 36258
rect 12462 36206 12514 36258
rect 12910 36206 12962 36258
rect 18846 36206 18898 36258
rect 27358 36206 27410 36258
rect 29710 36206 29762 36258
rect 30046 36206 30098 36258
rect 30270 36206 30322 36258
rect 30830 36206 30882 36258
rect 31390 36206 31442 36258
rect 37102 36206 37154 36258
rect 38110 36206 38162 36258
rect 14024 36038 14076 36090
rect 14148 36038 14200 36090
rect 14272 36038 14324 36090
rect 14396 36038 14448 36090
rect 14520 36038 14572 36090
rect 14644 36038 14696 36090
rect 14768 36038 14820 36090
rect 14892 36038 14944 36090
rect 15016 36038 15068 36090
rect 15140 36038 15192 36090
rect 34024 36038 34076 36090
rect 34148 36038 34200 36090
rect 34272 36038 34324 36090
rect 34396 36038 34448 36090
rect 34520 36038 34572 36090
rect 34644 36038 34696 36090
rect 34768 36038 34820 36090
rect 34892 36038 34944 36090
rect 35016 36038 35068 36090
rect 35140 36038 35192 36090
rect 4958 35870 5010 35922
rect 5854 35870 5906 35922
rect 6302 35870 6354 35922
rect 7086 35870 7138 35922
rect 7870 35870 7922 35922
rect 22318 35870 22370 35922
rect 22878 35870 22930 35922
rect 23214 35870 23266 35922
rect 34974 35870 35026 35922
rect 35982 35870 36034 35922
rect 36094 35870 36146 35922
rect 37326 35870 37378 35922
rect 37438 35870 37490 35922
rect 38334 35870 38386 35922
rect 8430 35758 8482 35810
rect 8654 35758 8706 35810
rect 8766 35758 8818 35810
rect 9662 35758 9714 35810
rect 9774 35758 9826 35810
rect 9886 35758 9938 35810
rect 9998 35758 10050 35810
rect 14926 35758 14978 35810
rect 16382 35758 16434 35810
rect 25902 35758 25954 35810
rect 26462 35758 26514 35810
rect 27806 35758 27858 35810
rect 28366 35758 28418 35810
rect 33070 35758 33122 35810
rect 38110 35758 38162 35810
rect 1822 35646 1874 35698
rect 2382 35646 2434 35698
rect 8990 35646 9042 35698
rect 9550 35646 9602 35698
rect 11902 35646 11954 35698
rect 14030 35646 14082 35698
rect 14702 35646 14754 35698
rect 15150 35646 15202 35698
rect 19406 35646 19458 35698
rect 19854 35646 19906 35698
rect 23998 35646 24050 35698
rect 25678 35646 25730 35698
rect 27582 35646 27634 35698
rect 31838 35646 31890 35698
rect 33630 35646 33682 35698
rect 34638 35646 34690 35698
rect 34862 35646 34914 35698
rect 36206 35646 36258 35698
rect 36430 35646 36482 35698
rect 36654 35646 36706 35698
rect 36990 35646 37042 35698
rect 37214 35646 37266 35698
rect 37662 35646 37714 35698
rect 37998 35646 38050 35698
rect 7758 35534 7810 35586
rect 8654 35534 8706 35586
rect 24446 35534 24498 35586
rect 31950 35534 32002 35586
rect 33742 35534 33794 35586
rect 34302 35534 34354 35586
rect 5518 35422 5570 35474
rect 10894 35422 10946 35474
rect 25342 35422 25394 35474
rect 27246 35422 27298 35474
rect 34862 35422 34914 35474
rect 35198 35422 35250 35474
rect 4024 35254 4076 35306
rect 4148 35254 4200 35306
rect 4272 35254 4324 35306
rect 4396 35254 4448 35306
rect 4520 35254 4572 35306
rect 4644 35254 4696 35306
rect 4768 35254 4820 35306
rect 4892 35254 4944 35306
rect 5016 35254 5068 35306
rect 5140 35254 5192 35306
rect 24024 35254 24076 35306
rect 24148 35254 24200 35306
rect 24272 35254 24324 35306
rect 24396 35254 24448 35306
rect 24520 35254 24572 35306
rect 24644 35254 24696 35306
rect 24768 35254 24820 35306
rect 24892 35254 24944 35306
rect 25016 35254 25068 35306
rect 25140 35254 25192 35306
rect 2158 35086 2210 35138
rect 10334 35086 10386 35138
rect 10894 35086 10946 35138
rect 12462 35086 12514 35138
rect 12798 35086 12850 35138
rect 13582 35086 13634 35138
rect 17166 35086 17218 35138
rect 20302 35086 20354 35138
rect 20638 35086 20690 35138
rect 26574 35086 26626 35138
rect 32510 35086 32562 35138
rect 37326 35086 37378 35138
rect 14590 34974 14642 35026
rect 15038 34974 15090 35026
rect 17950 34974 18002 35026
rect 27022 34974 27074 35026
rect 27358 34974 27410 35026
rect 33294 34974 33346 35026
rect 35198 34974 35250 35026
rect 35870 34974 35922 35026
rect 36206 34974 36258 35026
rect 2494 34862 2546 34914
rect 3054 34862 3106 34914
rect 4174 34862 4226 34914
rect 4734 34862 4786 34914
rect 6750 34862 6802 34914
rect 7310 34862 7362 34914
rect 11118 34862 11170 34914
rect 11790 34862 11842 34914
rect 19630 34862 19682 34914
rect 23102 34862 23154 34914
rect 23550 34862 23602 34914
rect 33182 34862 33234 34914
rect 33854 34862 33906 34914
rect 35646 34862 35698 34914
rect 36094 34862 36146 34914
rect 3278 34750 3330 34802
rect 4958 34750 5010 34802
rect 6078 34750 6130 34802
rect 10558 34750 10610 34802
rect 11678 34750 11730 34802
rect 13470 34750 13522 34802
rect 17278 34750 17330 34802
rect 17614 34750 17666 34802
rect 18062 34750 18114 34802
rect 18510 34750 18562 34802
rect 19070 34750 19122 34802
rect 19518 34750 19570 34802
rect 25790 34750 25842 34802
rect 27806 34750 27858 34802
rect 32398 34750 32450 34802
rect 32846 34750 32898 34802
rect 35086 34750 35138 34802
rect 36318 34750 36370 34802
rect 36990 34750 37042 34802
rect 37214 34750 37266 34802
rect 37774 34750 37826 34802
rect 37886 34750 37938 34802
rect 3838 34638 3890 34690
rect 5742 34638 5794 34690
rect 6190 34638 6242 34690
rect 6414 34638 6466 34690
rect 9550 34638 9602 34690
rect 13582 34638 13634 34690
rect 14142 34638 14194 34690
rect 16718 34638 16770 34690
rect 17166 34638 17218 34690
rect 17838 34638 17890 34690
rect 28254 34638 28306 34690
rect 29822 34638 29874 34690
rect 34862 34638 34914 34690
rect 35310 34638 35362 34690
rect 37550 34638 37602 34690
rect 14024 34470 14076 34522
rect 14148 34470 14200 34522
rect 14272 34470 14324 34522
rect 14396 34470 14448 34522
rect 14520 34470 14572 34522
rect 14644 34470 14696 34522
rect 14768 34470 14820 34522
rect 14892 34470 14944 34522
rect 15016 34470 15068 34522
rect 15140 34470 15192 34522
rect 34024 34470 34076 34522
rect 34148 34470 34200 34522
rect 34272 34470 34324 34522
rect 34396 34470 34448 34522
rect 34520 34470 34572 34522
rect 34644 34470 34696 34522
rect 34768 34470 34820 34522
rect 34892 34470 34944 34522
rect 35016 34470 35068 34522
rect 35140 34470 35192 34522
rect 4622 34302 4674 34354
rect 5294 34302 5346 34354
rect 5630 34302 5682 34354
rect 7086 34302 7138 34354
rect 7310 34302 7362 34354
rect 9886 34302 9938 34354
rect 11230 34302 11282 34354
rect 12126 34302 12178 34354
rect 15822 34302 15874 34354
rect 16270 34302 16322 34354
rect 16718 34302 16770 34354
rect 16942 34302 16994 34354
rect 25342 34302 25394 34354
rect 29150 34302 29202 34354
rect 29710 34302 29762 34354
rect 35758 34302 35810 34354
rect 37438 34302 37490 34354
rect 6638 34190 6690 34242
rect 7422 34190 7474 34242
rect 10558 34190 10610 34242
rect 16606 34190 16658 34242
rect 30158 34190 30210 34242
rect 30270 34190 30322 34242
rect 32510 34190 32562 34242
rect 33070 34190 33122 34242
rect 33518 34190 33570 34242
rect 34078 34190 34130 34242
rect 36654 34190 36706 34242
rect 1822 34078 1874 34130
rect 2270 34078 2322 34130
rect 6414 34078 6466 34130
rect 8094 34078 8146 34130
rect 8430 34078 8482 34130
rect 8654 34078 8706 34130
rect 9550 34078 9602 34130
rect 9886 34078 9938 34130
rect 10222 34078 10274 34130
rect 10446 34078 10498 34130
rect 17502 34078 17554 34130
rect 17838 34078 17890 34130
rect 20078 34078 20130 34130
rect 26014 34078 26066 34130
rect 26686 34078 26738 34130
rect 30494 34078 30546 34130
rect 31166 34078 31218 34130
rect 31502 34078 31554 34130
rect 32286 34078 32338 34130
rect 33294 34078 33346 34130
rect 33854 34078 33906 34130
rect 34526 34078 34578 34130
rect 35198 34078 35250 34130
rect 36878 34078 36930 34130
rect 7870 33966 7922 34018
rect 8206 33966 8258 34018
rect 11678 33966 11730 34018
rect 12910 33966 12962 34018
rect 21758 33966 21810 34018
rect 22206 33966 22258 34018
rect 31726 33966 31778 34018
rect 33406 33966 33458 34018
rect 37886 33966 37938 34018
rect 5966 33854 6018 33906
rect 21198 33854 21250 33906
rect 34974 33854 35026 33906
rect 36094 33854 36146 33906
rect 4024 33686 4076 33738
rect 4148 33686 4200 33738
rect 4272 33686 4324 33738
rect 4396 33686 4448 33738
rect 4520 33686 4572 33738
rect 4644 33686 4696 33738
rect 4768 33686 4820 33738
rect 4892 33686 4944 33738
rect 5016 33686 5068 33738
rect 5140 33686 5192 33738
rect 24024 33686 24076 33738
rect 24148 33686 24200 33738
rect 24272 33686 24324 33738
rect 24396 33686 24448 33738
rect 24520 33686 24572 33738
rect 24644 33686 24696 33738
rect 24768 33686 24820 33738
rect 24892 33686 24944 33738
rect 25016 33686 25068 33738
rect 25140 33686 25192 33738
rect 4622 33518 4674 33570
rect 5182 33518 5234 33570
rect 16382 33518 16434 33570
rect 35870 33518 35922 33570
rect 37550 33518 37602 33570
rect 4622 33406 4674 33458
rect 5070 33406 5122 33458
rect 11566 33406 11618 33458
rect 12014 33406 12066 33458
rect 16942 33406 16994 33458
rect 17278 33406 17330 33458
rect 18958 33406 19010 33458
rect 22542 33406 22594 33458
rect 23886 33406 23938 33458
rect 26238 33406 26290 33458
rect 33966 33406 34018 33458
rect 35422 33406 35474 33458
rect 36990 33406 37042 33458
rect 37998 33406 38050 33458
rect 6078 33294 6130 33346
rect 6862 33294 6914 33346
rect 7534 33294 7586 33346
rect 10558 33294 10610 33346
rect 11230 33294 11282 33346
rect 13918 33294 13970 33346
rect 16270 33294 16322 33346
rect 24446 33294 24498 33346
rect 31166 33294 31218 33346
rect 31838 33294 31890 33346
rect 33294 33294 33346 33346
rect 33854 33294 33906 33346
rect 34750 33294 34802 33346
rect 35534 33294 35586 33346
rect 37214 33294 37266 33346
rect 2494 33182 2546 33234
rect 2830 33182 2882 33234
rect 3166 33182 3218 33234
rect 6638 33182 6690 33234
rect 14142 33182 14194 33234
rect 14478 33182 14530 33234
rect 17614 33182 17666 33234
rect 17726 33182 17778 33234
rect 17838 33182 17890 33234
rect 24670 33182 24722 33234
rect 33742 33182 33794 33234
rect 4174 33070 4226 33122
rect 5742 33070 5794 33122
rect 8318 33070 8370 33122
rect 13582 33070 13634 33122
rect 15934 33070 15986 33122
rect 16382 33070 16434 33122
rect 18062 33070 18114 33122
rect 18510 33070 18562 33122
rect 22990 33070 23042 33122
rect 23550 33070 23602 33122
rect 25230 33070 25282 33122
rect 29822 33070 29874 33122
rect 30270 33070 30322 33122
rect 30942 33070 30994 33122
rect 31614 33070 31666 33122
rect 31726 33070 31778 33122
rect 32286 33070 32338 33122
rect 32734 33070 32786 33122
rect 14024 32902 14076 32954
rect 14148 32902 14200 32954
rect 14272 32902 14324 32954
rect 14396 32902 14448 32954
rect 14520 32902 14572 32954
rect 14644 32902 14696 32954
rect 14768 32902 14820 32954
rect 14892 32902 14944 32954
rect 15016 32902 15068 32954
rect 15140 32902 15192 32954
rect 34024 32902 34076 32954
rect 34148 32902 34200 32954
rect 34272 32902 34324 32954
rect 34396 32902 34448 32954
rect 34520 32902 34572 32954
rect 34644 32902 34696 32954
rect 34768 32902 34820 32954
rect 34892 32902 34944 32954
rect 35016 32902 35068 32954
rect 35140 32902 35192 32954
rect 4734 32734 4786 32786
rect 5630 32734 5682 32786
rect 6862 32734 6914 32786
rect 12014 32734 12066 32786
rect 15374 32734 15426 32786
rect 15934 32734 15986 32786
rect 16270 32734 16322 32786
rect 16718 32734 16770 32786
rect 17614 32734 17666 32786
rect 18062 32734 18114 32786
rect 23998 32734 24050 32786
rect 25342 32734 25394 32786
rect 25790 32734 25842 32786
rect 31166 32734 31218 32786
rect 31390 32734 31442 32786
rect 31838 32734 31890 32786
rect 32398 32734 32450 32786
rect 34078 32734 34130 32786
rect 36878 32734 36930 32786
rect 36990 32734 37042 32786
rect 37102 32734 37154 32786
rect 6526 32622 6578 32674
rect 6638 32622 6690 32674
rect 26238 32622 26290 32674
rect 27246 32622 27298 32674
rect 27806 32622 27858 32674
rect 30942 32622 30994 32674
rect 32174 32622 32226 32674
rect 34526 32622 34578 32674
rect 37438 32622 37490 32674
rect 7982 32510 8034 32562
rect 12238 32510 12290 32562
rect 12910 32510 12962 32562
rect 21310 32510 21362 32562
rect 21758 32510 21810 32562
rect 27022 32510 27074 32562
rect 33182 32510 33234 32562
rect 33518 32510 33570 32562
rect 34078 32510 34130 32562
rect 37326 32510 37378 32562
rect 5182 32398 5234 32450
rect 6190 32398 6242 32450
rect 7534 32398 7586 32450
rect 35758 32398 35810 32450
rect 5630 32286 5682 32338
rect 6078 32286 6130 32338
rect 24782 32286 24834 32338
rect 26686 32286 26738 32338
rect 31054 32286 31106 32338
rect 32510 32286 32562 32338
rect 33070 32286 33122 32338
rect 33406 32286 33458 32338
rect 4024 32118 4076 32170
rect 4148 32118 4200 32170
rect 4272 32118 4324 32170
rect 4396 32118 4448 32170
rect 4520 32118 4572 32170
rect 4644 32118 4696 32170
rect 4768 32118 4820 32170
rect 4892 32118 4944 32170
rect 5016 32118 5068 32170
rect 5140 32118 5192 32170
rect 24024 32118 24076 32170
rect 24148 32118 24200 32170
rect 24272 32118 24324 32170
rect 24396 32118 24448 32170
rect 24520 32118 24572 32170
rect 24644 32118 24696 32170
rect 24768 32118 24820 32170
rect 24892 32118 24944 32170
rect 25016 32118 25068 32170
rect 25140 32118 25192 32170
rect 6190 31950 6242 32002
rect 3614 31838 3666 31890
rect 8878 31838 8930 31890
rect 11902 31838 11954 31890
rect 12686 31838 12738 31890
rect 5070 31726 5122 31778
rect 9998 31726 10050 31778
rect 13806 31950 13858 32002
rect 14590 31950 14642 32002
rect 16270 31950 16322 32002
rect 16606 31950 16658 32002
rect 32734 31950 32786 32002
rect 16270 31838 16322 31890
rect 16718 31838 16770 31890
rect 22990 31838 23042 31890
rect 23326 31838 23378 31890
rect 36206 31838 36258 31890
rect 37214 31838 37266 31890
rect 14926 31726 14978 31778
rect 15710 31726 15762 31778
rect 17054 31726 17106 31778
rect 17278 31726 17330 31778
rect 18174 31726 18226 31778
rect 18398 31726 18450 31778
rect 22542 31726 22594 31778
rect 23998 31726 24050 31778
rect 26238 31726 26290 31778
rect 27694 31726 27746 31778
rect 29934 31726 29986 31778
rect 30158 31726 30210 31778
rect 30606 31726 30658 31778
rect 31054 31726 31106 31778
rect 31614 31726 31666 31778
rect 32622 31726 32674 31778
rect 32958 31726 33010 31778
rect 33966 31726 34018 31778
rect 34190 31726 34242 31778
rect 5630 31614 5682 31666
rect 13470 31614 13522 31666
rect 13694 31614 13746 31666
rect 15598 31614 15650 31666
rect 17390 31614 17442 31666
rect 18734 31614 18786 31666
rect 23886 31614 23938 31666
rect 25566 31614 25618 31666
rect 26910 31614 26962 31666
rect 28030 31614 28082 31666
rect 28478 31614 28530 31666
rect 30942 31614 30994 31666
rect 34750 31614 34802 31666
rect 2606 31502 2658 31554
rect 4510 31502 4562 31554
rect 7310 31502 7362 31554
rect 7982 31502 8034 31554
rect 8542 31502 8594 31554
rect 14142 31502 14194 31554
rect 17838 31502 17890 31554
rect 18510 31502 18562 31554
rect 25902 31502 25954 31554
rect 26350 31502 26402 31554
rect 26574 31502 26626 31554
rect 27358 31502 27410 31554
rect 29822 31502 29874 31554
rect 30382 31502 30434 31554
rect 32398 31502 32450 31554
rect 33742 31502 33794 31554
rect 14024 31334 14076 31386
rect 14148 31334 14200 31386
rect 14272 31334 14324 31386
rect 14396 31334 14448 31386
rect 14520 31334 14572 31386
rect 14644 31334 14696 31386
rect 14768 31334 14820 31386
rect 14892 31334 14944 31386
rect 15016 31334 15068 31386
rect 15140 31334 15192 31386
rect 34024 31334 34076 31386
rect 34148 31334 34200 31386
rect 34272 31334 34324 31386
rect 34396 31334 34448 31386
rect 34520 31334 34572 31386
rect 34644 31334 34696 31386
rect 34768 31334 34820 31386
rect 34892 31334 34944 31386
rect 35016 31334 35068 31386
rect 35140 31334 35192 31386
rect 2158 31166 2210 31218
rect 9662 31166 9714 31218
rect 15262 31166 15314 31218
rect 16270 31166 16322 31218
rect 16830 31166 16882 31218
rect 28366 31166 28418 31218
rect 33182 31166 33234 31218
rect 2830 31054 2882 31106
rect 3166 31054 3218 31106
rect 15598 31054 15650 31106
rect 29038 31054 29090 31106
rect 30494 31054 30546 31106
rect 34078 31054 34130 31106
rect 35086 31054 35138 31106
rect 36878 31054 36930 31106
rect 5518 30942 5570 30994
rect 8990 30942 9042 30994
rect 15486 30942 15538 30994
rect 17502 30942 17554 30994
rect 17950 30942 18002 30994
rect 25566 30942 25618 30994
rect 26014 30942 26066 30994
rect 30606 30942 30658 30994
rect 31166 30942 31218 30994
rect 32286 30942 32338 30994
rect 33518 30942 33570 30994
rect 35198 30942 35250 30994
rect 2606 30830 2658 30882
rect 3838 30830 3890 30882
rect 6750 30830 6802 30882
rect 13358 30830 13410 30882
rect 14366 30830 14418 30882
rect 14702 30830 14754 30882
rect 17726 30830 17778 30882
rect 29374 30830 29426 30882
rect 29822 30830 29874 30882
rect 32398 30830 32450 30882
rect 15598 30718 15650 30770
rect 17390 30718 17442 30770
rect 18174 30718 18226 30770
rect 31502 30718 31554 30770
rect 4024 30550 4076 30602
rect 4148 30550 4200 30602
rect 4272 30550 4324 30602
rect 4396 30550 4448 30602
rect 4520 30550 4572 30602
rect 4644 30550 4696 30602
rect 4768 30550 4820 30602
rect 4892 30550 4944 30602
rect 5016 30550 5068 30602
rect 5140 30550 5192 30602
rect 24024 30550 24076 30602
rect 24148 30550 24200 30602
rect 24272 30550 24324 30602
rect 24396 30550 24448 30602
rect 24520 30550 24572 30602
rect 24644 30550 24696 30602
rect 24768 30550 24820 30602
rect 24892 30550 24944 30602
rect 25016 30550 25068 30602
rect 25140 30550 25192 30602
rect 6414 30382 6466 30434
rect 10782 30382 10834 30434
rect 26574 30382 26626 30434
rect 26910 30382 26962 30434
rect 29598 30382 29650 30434
rect 30718 30382 30770 30434
rect 31390 30382 31442 30434
rect 36206 30382 36258 30434
rect 4846 30270 4898 30322
rect 6078 30270 6130 30322
rect 7646 30270 7698 30322
rect 16046 30270 16098 30322
rect 30942 30270 30994 30322
rect 2830 30158 2882 30210
rect 3502 30158 3554 30210
rect 4062 30158 4114 30210
rect 5854 30158 5906 30210
rect 7310 30158 7362 30210
rect 8542 30158 8594 30210
rect 10222 30158 10274 30210
rect 11678 30158 11730 30210
rect 12462 30158 12514 30210
rect 14254 30158 14306 30210
rect 16606 30158 16658 30210
rect 19742 30158 19794 30210
rect 20414 30158 20466 30210
rect 20862 30158 20914 30210
rect 21422 30158 21474 30210
rect 27694 30158 27746 30210
rect 31502 30158 31554 30210
rect 31838 30158 31890 30210
rect 32510 30158 32562 30210
rect 34638 30158 34690 30210
rect 3166 30046 3218 30098
rect 3950 30046 4002 30098
rect 4510 30046 4562 30098
rect 7870 30046 7922 30098
rect 8878 30046 8930 30098
rect 12238 30046 12290 30098
rect 27470 30046 27522 30098
rect 28590 30046 28642 30098
rect 29822 30046 29874 30098
rect 30382 30046 30434 30098
rect 2158 29934 2210 29986
rect 2606 29934 2658 29986
rect 3726 29934 3778 29986
rect 4734 29934 4786 29986
rect 7758 29934 7810 29986
rect 11342 29934 11394 29986
rect 17278 29934 17330 29986
rect 26126 29934 26178 29986
rect 29262 29934 29314 29986
rect 14024 29766 14076 29818
rect 14148 29766 14200 29818
rect 14272 29766 14324 29818
rect 14396 29766 14448 29818
rect 14520 29766 14572 29818
rect 14644 29766 14696 29818
rect 14768 29766 14820 29818
rect 14892 29766 14944 29818
rect 15016 29766 15068 29818
rect 15140 29766 15192 29818
rect 34024 29766 34076 29818
rect 34148 29766 34200 29818
rect 34272 29766 34324 29818
rect 34396 29766 34448 29818
rect 34520 29766 34572 29818
rect 34644 29766 34696 29818
rect 34768 29766 34820 29818
rect 34892 29766 34944 29818
rect 35016 29766 35068 29818
rect 35140 29766 35192 29818
rect 4622 29598 4674 29650
rect 5294 29598 5346 29650
rect 10782 29598 10834 29650
rect 14478 29598 14530 29650
rect 17726 29598 17778 29650
rect 19294 29598 19346 29650
rect 21310 29598 21362 29650
rect 26686 29598 26738 29650
rect 5630 29486 5682 29538
rect 5854 29486 5906 29538
rect 8094 29486 8146 29538
rect 10334 29486 10386 29538
rect 15934 29486 15986 29538
rect 16494 29486 16546 29538
rect 17950 29486 18002 29538
rect 22318 29486 22370 29538
rect 23326 29486 23378 29538
rect 23886 29486 23938 29538
rect 29822 29486 29874 29538
rect 33854 29486 33906 29538
rect 1822 29374 1874 29426
rect 2270 29374 2322 29426
rect 7086 29374 7138 29426
rect 8542 29374 8594 29426
rect 9774 29374 9826 29426
rect 11566 29374 11618 29426
rect 11902 29374 11954 29426
rect 15710 29374 15762 29426
rect 17390 29374 17442 29426
rect 17614 29374 17666 29426
rect 18734 29374 18786 29426
rect 23102 29374 23154 29426
rect 27134 29374 27186 29426
rect 27582 29374 27634 29426
rect 30942 29374 30994 29426
rect 33070 29374 33122 29426
rect 33294 29374 33346 29426
rect 8318 29262 8370 29314
rect 9662 29262 9714 29314
rect 31614 29262 31666 29314
rect 5518 29150 5570 29202
rect 15038 29150 15090 29202
rect 15374 29150 15426 29202
rect 22766 29150 22818 29202
rect 30606 29150 30658 29202
rect 4024 28982 4076 29034
rect 4148 28982 4200 29034
rect 4272 28982 4324 29034
rect 4396 28982 4448 29034
rect 4520 28982 4572 29034
rect 4644 28982 4696 29034
rect 4768 28982 4820 29034
rect 4892 28982 4944 29034
rect 5016 28982 5068 29034
rect 5140 28982 5192 29034
rect 24024 28982 24076 29034
rect 24148 28982 24200 29034
rect 24272 28982 24324 29034
rect 24396 28982 24448 29034
rect 24520 28982 24572 29034
rect 24644 28982 24696 29034
rect 24768 28982 24820 29034
rect 24892 28982 24944 29034
rect 25016 28982 25068 29034
rect 25140 28982 25192 29034
rect 3166 28814 3218 28866
rect 3502 28814 3554 28866
rect 4958 28814 5010 28866
rect 13022 28814 13074 28866
rect 13582 28814 13634 28866
rect 13918 28814 13970 28866
rect 22654 28814 22706 28866
rect 22990 28814 23042 28866
rect 7870 28702 7922 28754
rect 19742 28702 19794 28754
rect 21646 28702 21698 28754
rect 21982 28702 22034 28754
rect 26686 28702 26738 28754
rect 2494 28590 2546 28642
rect 3166 28590 3218 28642
rect 4174 28590 4226 28642
rect 4510 28590 4562 28642
rect 5630 28590 5682 28642
rect 5854 28590 5906 28642
rect 6974 28590 7026 28642
rect 9550 28590 9602 28642
rect 9998 28590 10050 28642
rect 14366 28590 14418 28642
rect 18286 28590 18338 28642
rect 18958 28590 19010 28642
rect 19294 28590 19346 28642
rect 23438 28590 23490 28642
rect 25454 28590 25506 28642
rect 28142 28590 28194 28642
rect 2270 28478 2322 28530
rect 2830 28478 2882 28530
rect 3950 28478 4002 28530
rect 4846 28478 4898 28530
rect 4958 28478 5010 28530
rect 14702 28478 14754 28530
rect 23550 28478 23602 28530
rect 4286 28366 4338 28418
rect 6190 28366 6242 28418
rect 12462 28366 12514 28418
rect 15262 28366 15314 28418
rect 15822 28366 15874 28418
rect 14024 28198 14076 28250
rect 14148 28198 14200 28250
rect 14272 28198 14324 28250
rect 14396 28198 14448 28250
rect 14520 28198 14572 28250
rect 14644 28198 14696 28250
rect 14768 28198 14820 28250
rect 14892 28198 14944 28250
rect 15016 28198 15068 28250
rect 15140 28198 15192 28250
rect 34024 28198 34076 28250
rect 34148 28198 34200 28250
rect 34272 28198 34324 28250
rect 34396 28198 34448 28250
rect 34520 28198 34572 28250
rect 34644 28198 34696 28250
rect 34768 28198 34820 28250
rect 34892 28198 34944 28250
rect 35016 28198 35068 28250
rect 35140 28198 35192 28250
rect 1598 28030 1650 28082
rect 2270 28030 2322 28082
rect 10110 28030 10162 28082
rect 12014 28030 12066 28082
rect 15486 28030 15538 28082
rect 16830 28030 16882 28082
rect 17502 28030 17554 28082
rect 17726 28030 17778 28082
rect 17950 28030 18002 28082
rect 18398 28030 18450 28082
rect 18846 28030 18898 28082
rect 23662 28030 23714 28082
rect 25342 28030 25394 28082
rect 29710 28030 29762 28082
rect 6750 27918 6802 27970
rect 9550 27918 9602 27970
rect 12686 27918 12738 27970
rect 13134 27918 13186 27970
rect 14254 27918 14306 27970
rect 14366 27918 14418 27970
rect 14590 27918 14642 27970
rect 15710 27918 15762 27970
rect 20302 27918 20354 27970
rect 30046 27918 30098 27970
rect 30830 27918 30882 27970
rect 31390 27918 31442 27970
rect 31726 27918 31778 27970
rect 4734 27806 4786 27858
rect 5294 27806 5346 27858
rect 5966 27806 6018 27858
rect 6190 27806 6242 27858
rect 6414 27806 6466 27858
rect 7534 27806 7586 27858
rect 13918 27806 13970 27858
rect 15822 27806 15874 27858
rect 17838 27806 17890 27858
rect 19630 27806 19682 27858
rect 20078 27806 20130 27858
rect 20974 27806 21026 27858
rect 21422 27806 21474 27858
rect 30606 27806 30658 27858
rect 5630 27694 5682 27746
rect 7646 27694 7698 27746
rect 8878 27694 8930 27746
rect 11566 27694 11618 27746
rect 12350 27694 12402 27746
rect 15262 27694 15314 27746
rect 16382 27694 16434 27746
rect 24446 27694 24498 27746
rect 25790 27694 25842 27746
rect 5518 27582 5570 27634
rect 9774 27582 9826 27634
rect 19294 27582 19346 27634
rect 30158 27582 30210 27634
rect 4024 27414 4076 27466
rect 4148 27414 4200 27466
rect 4272 27414 4324 27466
rect 4396 27414 4448 27466
rect 4520 27414 4572 27466
rect 4644 27414 4696 27466
rect 4768 27414 4820 27466
rect 4892 27414 4944 27466
rect 5016 27414 5068 27466
rect 5140 27414 5192 27466
rect 24024 27414 24076 27466
rect 24148 27414 24200 27466
rect 24272 27414 24324 27466
rect 24396 27414 24448 27466
rect 24520 27414 24572 27466
rect 24644 27414 24696 27466
rect 24768 27414 24820 27466
rect 24892 27414 24944 27466
rect 25016 27414 25068 27466
rect 25140 27414 25192 27466
rect 3614 27246 3666 27298
rect 4734 27246 4786 27298
rect 6414 27246 6466 27298
rect 7086 27246 7138 27298
rect 7422 27246 7474 27298
rect 8318 27246 8370 27298
rect 8654 27246 8706 27298
rect 19630 27246 19682 27298
rect 25678 27246 25730 27298
rect 25902 27246 25954 27298
rect 26462 27246 26514 27298
rect 3390 27134 3442 27186
rect 5070 27134 5122 27186
rect 6078 27134 6130 27186
rect 9326 27134 9378 27186
rect 9774 27134 9826 27186
rect 13022 27134 13074 27186
rect 13694 27134 13746 27186
rect 14030 27134 14082 27186
rect 15150 27134 15202 27186
rect 16942 27134 16994 27186
rect 17390 27134 17442 27186
rect 26014 27134 26066 27186
rect 26462 27134 26514 27186
rect 2158 27022 2210 27074
rect 4174 27022 4226 27074
rect 4510 27022 4562 27074
rect 4958 27022 5010 27074
rect 5630 27022 5682 27074
rect 6862 27022 6914 27074
rect 2942 26910 2994 26962
rect 3950 26910 4002 26962
rect 2606 26798 2658 26850
rect 8094 27022 8146 27074
rect 18846 27022 18898 27074
rect 22206 27022 22258 27074
rect 22654 27022 22706 27074
rect 29710 27022 29762 27074
rect 29934 27022 29986 27074
rect 30270 27022 30322 27074
rect 30718 27022 30770 27074
rect 33966 27022 34018 27074
rect 5854 26910 5906 26962
rect 14702 26910 14754 26962
rect 19854 26910 19906 26962
rect 20414 26910 20466 26962
rect 24894 26910 24946 26962
rect 29374 26910 29426 26962
rect 33070 26910 33122 26962
rect 3726 26798 3778 26850
rect 5630 26798 5682 26850
rect 19294 26798 19346 26850
rect 29822 26798 29874 26850
rect 14024 26630 14076 26682
rect 14148 26630 14200 26682
rect 14272 26630 14324 26682
rect 14396 26630 14448 26682
rect 14520 26630 14572 26682
rect 14644 26630 14696 26682
rect 14768 26630 14820 26682
rect 14892 26630 14944 26682
rect 15016 26630 15068 26682
rect 15140 26630 15192 26682
rect 34024 26630 34076 26682
rect 34148 26630 34200 26682
rect 34272 26630 34324 26682
rect 34396 26630 34448 26682
rect 34520 26630 34572 26682
rect 34644 26630 34696 26682
rect 34768 26630 34820 26682
rect 34892 26630 34944 26682
rect 35016 26630 35068 26682
rect 35140 26630 35192 26682
rect 3502 26462 3554 26514
rect 3838 26462 3890 26514
rect 4846 26462 4898 26514
rect 7086 26462 7138 26514
rect 7758 26462 7810 26514
rect 8318 26462 8370 26514
rect 21198 26462 21250 26514
rect 21758 26462 21810 26514
rect 23214 26462 23266 26514
rect 6750 26350 6802 26402
rect 22094 26350 22146 26402
rect 22654 26350 22706 26402
rect 26350 26350 26402 26402
rect 26462 26350 26514 26402
rect 30382 26350 30434 26402
rect 30606 26350 30658 26402
rect 4622 26238 4674 26290
rect 5294 26238 5346 26290
rect 6414 26238 6466 26290
rect 6638 26238 6690 26290
rect 7198 26238 7250 26290
rect 18174 26238 18226 26290
rect 18734 26238 18786 26290
rect 26686 26238 26738 26290
rect 30942 26238 30994 26290
rect 4286 26126 4338 26178
rect 23774 26126 23826 26178
rect 26014 26126 26066 26178
rect 29262 26126 29314 26178
rect 29710 26126 29762 26178
rect 3726 26014 3778 26066
rect 4286 26014 4338 26066
rect 4958 26014 5010 26066
rect 5518 26014 5570 26066
rect 5854 26014 5906 26066
rect 6302 26014 6354 26066
rect 22878 26014 22930 26066
rect 29374 26014 29426 26066
rect 29822 26014 29874 26066
rect 31278 26014 31330 26066
rect 4024 25846 4076 25898
rect 4148 25846 4200 25898
rect 4272 25846 4324 25898
rect 4396 25846 4448 25898
rect 4520 25846 4572 25898
rect 4644 25846 4696 25898
rect 4768 25846 4820 25898
rect 4892 25846 4944 25898
rect 5016 25846 5068 25898
rect 5140 25846 5192 25898
rect 24024 25846 24076 25898
rect 24148 25846 24200 25898
rect 24272 25846 24324 25898
rect 24396 25846 24448 25898
rect 24520 25846 24572 25898
rect 24644 25846 24696 25898
rect 24768 25846 24820 25898
rect 24892 25846 24944 25898
rect 25016 25846 25068 25898
rect 25140 25846 25192 25898
rect 5630 25678 5682 25730
rect 5742 25678 5794 25730
rect 5966 25678 6018 25730
rect 9998 25678 10050 25730
rect 23774 25678 23826 25730
rect 34190 25678 34242 25730
rect 4174 25566 4226 25618
rect 5070 25566 5122 25618
rect 7646 25566 7698 25618
rect 8094 25566 8146 25618
rect 14030 25566 14082 25618
rect 21982 25566 22034 25618
rect 29598 25566 29650 25618
rect 30158 25566 30210 25618
rect 6078 25454 6130 25506
rect 14702 25454 14754 25506
rect 26798 25454 26850 25506
rect 27470 25454 27522 25506
rect 29374 25454 29426 25506
rect 30718 25454 30770 25506
rect 31166 25454 31218 25506
rect 4734 25342 4786 25394
rect 10222 25342 10274 25394
rect 10558 25342 10610 25394
rect 14366 25342 14418 25394
rect 14478 25342 14530 25394
rect 27918 25342 27970 25394
rect 6862 25230 6914 25282
rect 9214 25230 9266 25282
rect 9662 25230 9714 25282
rect 13582 25230 13634 25282
rect 15038 25230 15090 25282
rect 22318 25230 22370 25282
rect 24558 25230 24610 25282
rect 28254 25230 28306 25282
rect 33406 25230 33458 25282
rect 14024 25062 14076 25114
rect 14148 25062 14200 25114
rect 14272 25062 14324 25114
rect 14396 25062 14448 25114
rect 14520 25062 14572 25114
rect 14644 25062 14696 25114
rect 14768 25062 14820 25114
rect 14892 25062 14944 25114
rect 15016 25062 15068 25114
rect 15140 25062 15192 25114
rect 34024 25062 34076 25114
rect 34148 25062 34200 25114
rect 34272 25062 34324 25114
rect 34396 25062 34448 25114
rect 34520 25062 34572 25114
rect 34644 25062 34696 25114
rect 34768 25062 34820 25114
rect 34892 25062 34944 25114
rect 35016 25062 35068 25114
rect 35140 25062 35192 25114
rect 1822 24894 1874 24946
rect 3166 24894 3218 24946
rect 8542 24894 8594 24946
rect 12574 24894 12626 24946
rect 13022 24894 13074 24946
rect 18734 24894 18786 24946
rect 26126 24894 26178 24946
rect 26686 24894 26738 24946
rect 28478 24894 28530 24946
rect 29934 24894 29986 24946
rect 10782 24782 10834 24834
rect 14030 24782 14082 24834
rect 14366 24782 14418 24834
rect 15374 24782 15426 24834
rect 19742 24782 19794 24834
rect 20302 24782 20354 24834
rect 24670 24782 24722 24834
rect 25454 24782 25506 24834
rect 27134 24782 27186 24834
rect 27470 24782 27522 24834
rect 2830 24670 2882 24722
rect 3838 24670 3890 24722
rect 8094 24670 8146 24722
rect 8990 24670 9042 24722
rect 9998 24670 10050 24722
rect 10558 24670 10610 24722
rect 13806 24670 13858 24722
rect 15486 24670 15538 24722
rect 19518 24670 19570 24722
rect 26462 24670 26514 24722
rect 26910 24670 26962 24722
rect 27806 24670 27858 24722
rect 28142 24670 28194 24722
rect 28814 24670 28866 24722
rect 29374 24670 29426 24722
rect 29598 24670 29650 24722
rect 30270 24670 30322 24722
rect 2494 24558 2546 24610
rect 5294 24558 5346 24610
rect 11566 24558 11618 24610
rect 16606 24558 16658 24610
rect 18286 24558 18338 24610
rect 25790 24558 25842 24610
rect 27918 24558 27970 24610
rect 30942 24558 30994 24610
rect 31390 24558 31442 24610
rect 31838 24558 31890 24610
rect 9662 24446 9714 24498
rect 13470 24446 13522 24498
rect 19182 24446 19234 24498
rect 25230 24446 25282 24498
rect 26014 24446 26066 24498
rect 27022 24446 27074 24498
rect 4024 24278 4076 24330
rect 4148 24278 4200 24330
rect 4272 24278 4324 24330
rect 4396 24278 4448 24330
rect 4520 24278 4572 24330
rect 4644 24278 4696 24330
rect 4768 24278 4820 24330
rect 4892 24278 4944 24330
rect 5016 24278 5068 24330
rect 5140 24278 5192 24330
rect 24024 24278 24076 24330
rect 24148 24278 24200 24330
rect 24272 24278 24324 24330
rect 24396 24278 24448 24330
rect 24520 24278 24572 24330
rect 24644 24278 24696 24330
rect 24768 24278 24820 24330
rect 24892 24278 24944 24330
rect 25016 24278 25068 24330
rect 25140 24278 25192 24330
rect 11342 24110 11394 24162
rect 19630 24110 19682 24162
rect 30494 24110 30546 24162
rect 30606 24110 30658 24162
rect 6638 23998 6690 24050
rect 24558 23998 24610 24050
rect 27806 23998 27858 24050
rect 31054 23998 31106 24050
rect 2158 23886 2210 23938
rect 7422 23886 7474 23938
rect 7870 23886 7922 23938
rect 8318 23886 8370 23938
rect 11566 23886 11618 23938
rect 13470 23886 13522 23938
rect 13918 23886 13970 23938
rect 23102 23886 23154 23938
rect 24446 23886 24498 23938
rect 24894 23886 24946 23938
rect 25006 23886 25058 23938
rect 25454 23886 25506 23938
rect 29038 23886 29090 23938
rect 29486 23886 29538 23938
rect 30158 23886 30210 23938
rect 30270 23886 30322 23938
rect 2830 23774 2882 23826
rect 4510 23774 4562 23826
rect 6190 23774 6242 23826
rect 11678 23774 11730 23826
rect 18846 23774 18898 23826
rect 19854 23774 19906 23826
rect 20414 23774 20466 23826
rect 22766 23774 22818 23826
rect 1934 23662 1986 23714
rect 2494 23662 2546 23714
rect 3390 23662 3442 23714
rect 4398 23662 4450 23714
rect 5070 23662 5122 23714
rect 10782 23662 10834 23714
rect 11902 23662 11954 23714
rect 12238 23662 12290 23714
rect 16494 23662 16546 23714
rect 17054 23662 17106 23714
rect 17390 23662 17442 23714
rect 17838 23662 17890 23714
rect 19294 23662 19346 23714
rect 21422 23662 21474 23714
rect 21870 23662 21922 23714
rect 22430 23662 22482 23714
rect 22878 23662 22930 23714
rect 24110 23662 24162 23714
rect 24670 23662 24722 23714
rect 28478 23662 28530 23714
rect 29598 23662 29650 23714
rect 29710 23662 29762 23714
rect 31502 23662 31554 23714
rect 31950 23662 32002 23714
rect 14024 23494 14076 23546
rect 14148 23494 14200 23546
rect 14272 23494 14324 23546
rect 14396 23494 14448 23546
rect 14520 23494 14572 23546
rect 14644 23494 14696 23546
rect 14768 23494 14820 23546
rect 14892 23494 14944 23546
rect 15016 23494 15068 23546
rect 15140 23494 15192 23546
rect 34024 23494 34076 23546
rect 34148 23494 34200 23546
rect 34272 23494 34324 23546
rect 34396 23494 34448 23546
rect 34520 23494 34572 23546
rect 34644 23494 34696 23546
rect 34768 23494 34820 23546
rect 34892 23494 34944 23546
rect 35016 23494 35068 23546
rect 35140 23494 35192 23546
rect 3838 23326 3890 23378
rect 4062 23326 4114 23378
rect 5182 23326 5234 23378
rect 15150 23326 15202 23378
rect 21758 23326 21810 23378
rect 28142 23326 28194 23378
rect 31614 23326 31666 23378
rect 1934 23214 1986 23266
rect 2270 23214 2322 23266
rect 5406 23214 5458 23266
rect 13806 23214 13858 23266
rect 16270 23214 16322 23266
rect 16494 23214 16546 23266
rect 20974 23214 21026 23266
rect 25342 23214 25394 23266
rect 27022 23214 27074 23266
rect 2606 23102 2658 23154
rect 4286 23102 4338 23154
rect 5294 23102 5346 23154
rect 5966 23102 6018 23154
rect 11118 23102 11170 23154
rect 11566 23102 11618 23154
rect 14590 23102 14642 23154
rect 15934 23102 15986 23154
rect 18286 23102 18338 23154
rect 18734 23102 18786 23154
rect 21982 23102 22034 23154
rect 26350 23102 26402 23154
rect 30606 23102 30658 23154
rect 31054 23102 31106 23154
rect 3390 22990 3442 23042
rect 3950 22990 4002 23042
rect 8094 22990 8146 23042
rect 17502 22990 17554 23042
rect 23662 22990 23714 23042
rect 26686 22990 26738 23042
rect 4510 22878 4562 22930
rect 15598 22878 15650 22930
rect 27582 22878 27634 22930
rect 4024 22710 4076 22762
rect 4148 22710 4200 22762
rect 4272 22710 4324 22762
rect 4396 22710 4448 22762
rect 4520 22710 4572 22762
rect 4644 22710 4696 22762
rect 4768 22710 4820 22762
rect 4892 22710 4944 22762
rect 5016 22710 5068 22762
rect 5140 22710 5192 22762
rect 24024 22710 24076 22762
rect 24148 22710 24200 22762
rect 24272 22710 24324 22762
rect 24396 22710 24448 22762
rect 24520 22710 24572 22762
rect 24644 22710 24696 22762
rect 24768 22710 24820 22762
rect 24892 22710 24944 22762
rect 25016 22710 25068 22762
rect 25140 22710 25192 22762
rect 4174 22542 4226 22594
rect 13582 22542 13634 22594
rect 13918 22542 13970 22594
rect 28142 22542 28194 22594
rect 29150 22542 29202 22594
rect 3278 22430 3330 22482
rect 11566 22430 11618 22482
rect 20862 22430 20914 22482
rect 21758 22430 21810 22482
rect 23886 22430 23938 22482
rect 27246 22430 27298 22482
rect 29486 22430 29538 22482
rect 30942 22430 30994 22482
rect 31390 22430 31442 22482
rect 2158 22318 2210 22370
rect 4846 22318 4898 22370
rect 5630 22318 5682 22370
rect 6078 22318 6130 22370
rect 11230 22318 11282 22370
rect 12462 22318 12514 22370
rect 12798 22318 12850 22370
rect 15374 22318 15426 22370
rect 15934 22318 15986 22370
rect 23102 22318 23154 22370
rect 23998 22318 24050 22370
rect 24670 22318 24722 22370
rect 25454 22318 25506 22370
rect 27358 22318 27410 22370
rect 29934 22318 29986 22370
rect 30606 22318 30658 22370
rect 2494 22206 2546 22258
rect 4958 22206 5010 22258
rect 11566 22206 11618 22258
rect 12126 22206 12178 22258
rect 14142 22206 14194 22258
rect 14702 22206 14754 22258
rect 21982 22206 22034 22258
rect 22542 22206 22594 22258
rect 24894 22206 24946 22258
rect 25790 22206 25842 22258
rect 30046 22206 30098 22258
rect 1822 22094 1874 22146
rect 2830 22094 2882 22146
rect 3838 22094 3890 22146
rect 8542 22094 8594 22146
rect 9214 22094 9266 22146
rect 9550 22094 9602 22146
rect 9998 22094 10050 22146
rect 11678 22094 11730 22146
rect 11902 22094 11954 22146
rect 12238 22094 12290 22146
rect 18510 22094 18562 22146
rect 19070 22094 19122 22146
rect 19406 22094 19458 22146
rect 20302 22094 20354 22146
rect 21422 22094 21474 22146
rect 23214 22094 23266 22146
rect 23438 22094 23490 22146
rect 29262 22094 29314 22146
rect 30158 22094 30210 22146
rect 14024 21926 14076 21978
rect 14148 21926 14200 21978
rect 14272 21926 14324 21978
rect 14396 21926 14448 21978
rect 14520 21926 14572 21978
rect 14644 21926 14696 21978
rect 14768 21926 14820 21978
rect 14892 21926 14944 21978
rect 15016 21926 15068 21978
rect 15140 21926 15192 21978
rect 34024 21926 34076 21978
rect 34148 21926 34200 21978
rect 34272 21926 34324 21978
rect 34396 21926 34448 21978
rect 34520 21926 34572 21978
rect 34644 21926 34696 21978
rect 34768 21926 34820 21978
rect 34892 21926 34944 21978
rect 35016 21926 35068 21978
rect 35140 21926 35192 21978
rect 4846 21758 4898 21810
rect 5854 21758 5906 21810
rect 8430 21758 8482 21810
rect 8878 21758 8930 21810
rect 13694 21758 13746 21810
rect 6974 21646 7026 21698
rect 8766 21646 8818 21698
rect 12350 21646 12402 21698
rect 15038 21646 15090 21698
rect 15150 21702 15202 21754
rect 15598 21758 15650 21810
rect 23998 21758 24050 21810
rect 25342 21758 25394 21810
rect 31838 21758 31890 21810
rect 16718 21646 16770 21698
rect 26238 21646 26290 21698
rect 28926 21646 28978 21698
rect 29710 21646 29762 21698
rect 1710 21534 1762 21586
rect 2382 21534 2434 21586
rect 6190 21534 6242 21586
rect 6862 21534 6914 21586
rect 7534 21534 7586 21586
rect 9662 21534 9714 21586
rect 10110 21534 10162 21586
rect 15934 21534 15986 21586
rect 16606 21534 16658 21586
rect 17502 21534 17554 21586
rect 21310 21534 21362 21586
rect 21758 21534 21810 21586
rect 25230 21534 25282 21586
rect 27022 21534 27074 21586
rect 28590 21534 28642 21586
rect 29822 21534 29874 21586
rect 14142 21422 14194 21474
rect 14590 21422 14642 21474
rect 5406 21310 5458 21362
rect 8878 21310 8930 21362
rect 13134 21310 13186 21362
rect 15038 21310 15090 21362
rect 24782 21310 24834 21362
rect 28254 21310 28306 21362
rect 4024 21142 4076 21194
rect 4148 21142 4200 21194
rect 4272 21142 4324 21194
rect 4396 21142 4448 21194
rect 4520 21142 4572 21194
rect 4644 21142 4696 21194
rect 4768 21142 4820 21194
rect 4892 21142 4944 21194
rect 5016 21142 5068 21194
rect 5140 21142 5192 21194
rect 24024 21142 24076 21194
rect 24148 21142 24200 21194
rect 24272 21142 24324 21194
rect 24396 21142 24448 21194
rect 24520 21142 24572 21194
rect 24644 21142 24696 21194
rect 24768 21142 24820 21194
rect 24892 21142 24944 21194
rect 25016 21142 25068 21194
rect 25140 21142 25192 21194
rect 4510 20974 4562 21026
rect 20414 20974 20466 21026
rect 21870 20974 21922 21026
rect 22206 20974 22258 21026
rect 33518 20974 33570 21026
rect 1934 20862 1986 20914
rect 6750 20862 6802 20914
rect 10558 20862 10610 20914
rect 12238 20862 12290 20914
rect 12910 20862 12962 20914
rect 15150 20862 15202 20914
rect 15598 20862 15650 20914
rect 25454 20862 25506 20914
rect 27470 20862 27522 20914
rect 4622 20750 4674 20802
rect 6078 20750 6130 20802
rect 8430 20750 8482 20802
rect 9102 20750 9154 20802
rect 10334 20750 10386 20802
rect 11790 20750 11842 20802
rect 12126 20750 12178 20802
rect 20750 20750 20802 20802
rect 21422 20750 21474 20802
rect 23998 20750 24050 20802
rect 24558 20750 24610 20802
rect 24670 20750 24722 20802
rect 25230 20750 25282 20802
rect 27806 20750 27858 20802
rect 28254 20750 28306 20802
rect 29150 20750 29202 20802
rect 29486 20750 29538 20802
rect 30046 20750 30098 20802
rect 30382 20750 30434 20802
rect 2830 20638 2882 20690
rect 3166 20638 3218 20690
rect 6190 20638 6242 20690
rect 9326 20638 9378 20690
rect 10894 20638 10946 20690
rect 22430 20638 22482 20690
rect 22990 20638 23042 20690
rect 29262 20638 29314 20690
rect 32734 20638 32786 20690
rect 2494 20526 2546 20578
rect 5070 20526 5122 20578
rect 5742 20526 5794 20578
rect 6414 20526 6466 20578
rect 8766 20526 8818 20578
rect 9550 20526 9602 20578
rect 9662 20526 9714 20578
rect 13694 20526 13746 20578
rect 14142 20526 14194 20578
rect 20526 20526 20578 20578
rect 23662 20526 23714 20578
rect 23886 20526 23938 20578
rect 14024 20358 14076 20410
rect 14148 20358 14200 20410
rect 14272 20358 14324 20410
rect 14396 20358 14448 20410
rect 14520 20358 14572 20410
rect 14644 20358 14696 20410
rect 14768 20358 14820 20410
rect 14892 20358 14944 20410
rect 15016 20358 15068 20410
rect 15140 20358 15192 20410
rect 34024 20358 34076 20410
rect 34148 20358 34200 20410
rect 34272 20358 34324 20410
rect 34396 20358 34448 20410
rect 34520 20358 34572 20410
rect 34644 20358 34696 20410
rect 34768 20358 34820 20410
rect 34892 20358 34944 20410
rect 35016 20358 35068 20410
rect 35140 20358 35192 20410
rect 6190 20190 6242 20242
rect 10670 20190 10722 20242
rect 11566 20190 11618 20242
rect 11678 20190 11730 20242
rect 1934 20078 1986 20130
rect 10334 20078 10386 20130
rect 10446 20078 10498 20130
rect 12126 20078 12178 20130
rect 12350 20078 12402 20130
rect 12574 20078 12626 20130
rect 13918 20078 13970 20130
rect 14142 20078 14194 20130
rect 18286 20078 18338 20130
rect 18622 20078 18674 20130
rect 18734 20078 18786 20130
rect 25790 20078 25842 20130
rect 26798 20078 26850 20130
rect 31950 20078 32002 20130
rect 9886 19966 9938 20018
rect 11902 19966 11954 20018
rect 12686 19966 12738 20018
rect 14366 19966 14418 20018
rect 14814 19966 14866 20018
rect 18958 19966 19010 20018
rect 23662 19966 23714 20018
rect 24782 19966 24834 20018
rect 25342 19966 25394 20018
rect 28478 19966 28530 20018
rect 29150 19966 29202 20018
rect 29710 19966 29762 20018
rect 30158 19966 30210 20018
rect 30270 19966 30322 20018
rect 30718 19966 30770 20018
rect 2494 19854 2546 19906
rect 5742 19854 5794 19906
rect 10334 19854 10386 19906
rect 14254 19854 14306 19906
rect 23550 19854 23602 19906
rect 27022 19854 27074 19906
rect 29822 19854 29874 19906
rect 30942 19854 30994 19906
rect 31502 19854 31554 19906
rect 24222 19742 24274 19794
rect 30270 19742 30322 19794
rect 4024 19574 4076 19626
rect 4148 19574 4200 19626
rect 4272 19574 4324 19626
rect 4396 19574 4448 19626
rect 4520 19574 4572 19626
rect 4644 19574 4696 19626
rect 4768 19574 4820 19626
rect 4892 19574 4944 19626
rect 5016 19574 5068 19626
rect 5140 19574 5192 19626
rect 24024 19574 24076 19626
rect 24148 19574 24200 19626
rect 24272 19574 24324 19626
rect 24396 19574 24448 19626
rect 24520 19574 24572 19626
rect 24644 19574 24696 19626
rect 24768 19574 24820 19626
rect 24892 19574 24944 19626
rect 25016 19574 25068 19626
rect 25140 19574 25192 19626
rect 2046 19406 2098 19458
rect 2606 19406 2658 19458
rect 23886 19406 23938 19458
rect 24670 19406 24722 19458
rect 26126 19406 26178 19458
rect 26910 19406 26962 19458
rect 2046 19294 2098 19346
rect 14590 19294 14642 19346
rect 24670 19294 24722 19346
rect 28030 19294 28082 19346
rect 2942 19182 2994 19234
rect 3614 19182 3666 19234
rect 14702 19182 14754 19234
rect 15038 19182 15090 19234
rect 18846 19182 18898 19234
rect 18958 19182 19010 19234
rect 20526 19182 20578 19234
rect 25118 19182 25170 19234
rect 25678 19182 25730 19234
rect 26350 19182 26402 19234
rect 27134 19182 27186 19234
rect 27358 19182 27410 19234
rect 27694 19182 27746 19234
rect 27918 19182 27970 19234
rect 28366 19182 28418 19234
rect 29150 19182 29202 19234
rect 32286 19182 32338 19234
rect 32734 19182 32786 19234
rect 19182 19070 19234 19122
rect 19518 19070 19570 19122
rect 19742 19070 19794 19122
rect 20190 19070 20242 19122
rect 20302 19070 20354 19122
rect 26462 19070 26514 19122
rect 26798 19070 26850 19122
rect 2494 18958 2546 19010
rect 3166 18958 3218 19010
rect 3838 18958 3890 19010
rect 14254 18958 14306 19010
rect 14478 18958 14530 19010
rect 17166 18958 17218 19010
rect 19630 18958 19682 19010
rect 24222 18958 24274 19010
rect 28142 18958 28194 19010
rect 29822 18958 29874 19010
rect 14024 18790 14076 18842
rect 14148 18790 14200 18842
rect 14272 18790 14324 18842
rect 14396 18790 14448 18842
rect 14520 18790 14572 18842
rect 14644 18790 14696 18842
rect 14768 18790 14820 18842
rect 14892 18790 14944 18842
rect 15016 18790 15068 18842
rect 15140 18790 15192 18842
rect 34024 18790 34076 18842
rect 34148 18790 34200 18842
rect 34272 18790 34324 18842
rect 34396 18790 34448 18842
rect 34520 18790 34572 18842
rect 34644 18790 34696 18842
rect 34768 18790 34820 18842
rect 34892 18790 34944 18842
rect 35016 18790 35068 18842
rect 35140 18790 35192 18842
rect 15374 18622 15426 18674
rect 16606 18622 16658 18674
rect 20526 18622 20578 18674
rect 27358 18622 27410 18674
rect 27918 18622 27970 18674
rect 29598 18622 29650 18674
rect 3166 18510 3218 18562
rect 12014 18510 12066 18562
rect 12238 18510 12290 18562
rect 13134 18510 13186 18562
rect 13806 18510 13858 18562
rect 15710 18510 15762 18562
rect 21534 18510 21586 18562
rect 26798 18510 26850 18562
rect 29038 18510 29090 18562
rect 2606 18398 2658 18450
rect 2830 18398 2882 18450
rect 13246 18398 13298 18450
rect 13918 18398 13970 18450
rect 14814 18398 14866 18450
rect 15598 18398 15650 18450
rect 16718 18398 16770 18450
rect 17390 18398 17442 18450
rect 18062 18398 18114 18450
rect 21198 18398 21250 18450
rect 21422 18398 21474 18450
rect 21870 18398 21922 18450
rect 22542 18398 22594 18450
rect 23214 18398 23266 18450
rect 28590 18398 28642 18450
rect 29710 18398 29762 18450
rect 30718 18398 30770 18450
rect 28254 18286 28306 18338
rect 30158 18286 30210 18338
rect 11902 18174 11954 18226
rect 21086 18174 21138 18226
rect 23102 18174 23154 18226
rect 4024 18006 4076 18058
rect 4148 18006 4200 18058
rect 4272 18006 4324 18058
rect 4396 18006 4448 18058
rect 4520 18006 4572 18058
rect 4644 18006 4696 18058
rect 4768 18006 4820 18058
rect 4892 18006 4944 18058
rect 5016 18006 5068 18058
rect 5140 18006 5192 18058
rect 24024 18006 24076 18058
rect 24148 18006 24200 18058
rect 24272 18006 24324 18058
rect 24396 18006 24448 18058
rect 24520 18006 24572 18058
rect 24644 18006 24696 18058
rect 24768 18006 24820 18058
rect 24892 18006 24944 18058
rect 25016 18006 25068 18058
rect 25140 18006 25192 18058
rect 4174 17838 4226 17890
rect 10446 17838 10498 17890
rect 13582 17838 13634 17890
rect 9550 17726 9602 17778
rect 17950 17726 18002 17778
rect 19742 17726 19794 17778
rect 29262 17726 29314 17778
rect 4622 17614 4674 17666
rect 5630 17614 5682 17666
rect 6078 17614 6130 17666
rect 9998 17614 10050 17666
rect 11118 17614 11170 17666
rect 11902 17614 11954 17666
rect 16606 17614 16658 17666
rect 17054 17614 17106 17666
rect 19294 17614 19346 17666
rect 19406 17614 19458 17666
rect 20414 17614 20466 17666
rect 20638 17614 20690 17666
rect 21646 17614 21698 17666
rect 22094 17614 22146 17666
rect 22318 17614 22370 17666
rect 22654 17614 22706 17666
rect 23326 17614 23378 17666
rect 23550 17614 23602 17666
rect 23774 17614 23826 17666
rect 4958 17502 5010 17554
rect 9214 17502 9266 17554
rect 12014 17502 12066 17554
rect 12574 17502 12626 17554
rect 18174 17502 18226 17554
rect 18622 17502 18674 17554
rect 22766 17502 22818 17554
rect 2606 17390 2658 17442
rect 2830 17390 2882 17442
rect 3166 17390 3218 17442
rect 3838 17390 3890 17442
rect 8542 17390 8594 17442
rect 10558 17390 10610 17442
rect 10782 17390 10834 17442
rect 11454 17390 11506 17442
rect 12350 17390 12402 17442
rect 14366 17390 14418 17442
rect 17614 17390 17666 17442
rect 21422 17390 21474 17442
rect 22206 17390 22258 17442
rect 22990 17390 23042 17442
rect 23662 17390 23714 17442
rect 24894 17390 24946 17442
rect 28254 17390 28306 17442
rect 14024 17222 14076 17274
rect 14148 17222 14200 17274
rect 14272 17222 14324 17274
rect 14396 17222 14448 17274
rect 14520 17222 14572 17274
rect 14644 17222 14696 17274
rect 14768 17222 14820 17274
rect 14892 17222 14944 17274
rect 15016 17222 15068 17274
rect 15140 17222 15192 17274
rect 34024 17222 34076 17274
rect 34148 17222 34200 17274
rect 34272 17222 34324 17274
rect 34396 17222 34448 17274
rect 34520 17222 34572 17274
rect 34644 17222 34696 17274
rect 34768 17222 34820 17274
rect 34892 17222 34944 17274
rect 35016 17222 35068 17274
rect 35140 17222 35192 17274
rect 2494 17054 2546 17106
rect 7422 17054 7474 17106
rect 8654 17054 8706 17106
rect 10110 17054 10162 17106
rect 18510 17054 18562 17106
rect 20862 17054 20914 17106
rect 22430 17054 22482 17106
rect 23886 17054 23938 17106
rect 24110 17054 24162 17106
rect 25566 17054 25618 17106
rect 26238 17054 26290 17106
rect 26798 17054 26850 17106
rect 1934 16942 1986 16994
rect 3166 16942 3218 16994
rect 4734 16942 4786 16994
rect 8430 16942 8482 16994
rect 9662 16942 9714 16994
rect 10446 16942 10498 16994
rect 10894 16942 10946 16994
rect 11006 16942 11058 16994
rect 11118 16942 11170 16994
rect 13358 16942 13410 16994
rect 15486 16942 15538 16994
rect 16494 16942 16546 16994
rect 16606 16942 16658 16994
rect 19742 16942 19794 16994
rect 20078 16942 20130 16994
rect 22654 16942 22706 16994
rect 23214 16942 23266 16994
rect 23662 16942 23714 16994
rect 25230 16942 25282 16994
rect 26126 16942 26178 16994
rect 2158 16830 2210 16882
rect 2942 16830 2994 16882
rect 4622 16830 4674 16882
rect 5294 16830 5346 16882
rect 5742 16830 5794 16882
rect 6974 16830 7026 16882
rect 7198 16830 7250 16882
rect 8206 16830 8258 16882
rect 8878 16830 8930 16882
rect 9550 16830 9602 16882
rect 12126 16830 12178 16882
rect 14926 16830 14978 16882
rect 15710 16830 15762 16882
rect 17614 16830 17666 16882
rect 20190 16830 20242 16882
rect 20414 16830 20466 16882
rect 21086 16830 21138 16882
rect 21422 16830 21474 16882
rect 22094 16830 22146 16882
rect 23326 16830 23378 16882
rect 24222 16830 24274 16882
rect 25454 16830 25506 16882
rect 25902 16830 25954 16882
rect 3614 16718 3666 16770
rect 3950 16718 4002 16770
rect 6862 16718 6914 16770
rect 18062 16718 18114 16770
rect 19406 16718 19458 16770
rect 22318 16718 22370 16770
rect 1710 16606 1762 16658
rect 1934 16606 1986 16658
rect 7758 16606 7810 16658
rect 7870 16606 7922 16658
rect 8318 16606 8370 16658
rect 14590 16606 14642 16658
rect 16606 16606 16658 16658
rect 19518 16606 19570 16658
rect 20750 16606 20802 16658
rect 23774 16606 23826 16658
rect 26238 16606 26290 16658
rect 4024 16438 4076 16490
rect 4148 16438 4200 16490
rect 4272 16438 4324 16490
rect 4396 16438 4448 16490
rect 4520 16438 4572 16490
rect 4644 16438 4696 16490
rect 4768 16438 4820 16490
rect 4892 16438 4944 16490
rect 5016 16438 5068 16490
rect 5140 16438 5192 16490
rect 24024 16438 24076 16490
rect 24148 16438 24200 16490
rect 24272 16438 24324 16490
rect 24396 16438 24448 16490
rect 24520 16438 24572 16490
rect 24644 16438 24696 16490
rect 24768 16438 24820 16490
rect 24892 16438 24944 16490
rect 25016 16438 25068 16490
rect 25140 16438 25192 16490
rect 3390 16270 3442 16322
rect 6078 16270 6130 16322
rect 13694 16270 13746 16322
rect 21646 16270 21698 16322
rect 26798 16270 26850 16322
rect 30382 16270 30434 16322
rect 4734 16158 4786 16210
rect 7422 16158 7474 16210
rect 7758 16158 7810 16210
rect 9438 16158 9490 16210
rect 11230 16158 11282 16210
rect 13582 16158 13634 16210
rect 14030 16158 14082 16210
rect 14702 16158 14754 16210
rect 15038 16158 15090 16210
rect 23774 16158 23826 16210
rect 29374 16158 29426 16210
rect 3950 16046 4002 16098
rect 5854 16046 5906 16098
rect 6302 16046 6354 16098
rect 7086 16046 7138 16098
rect 8654 16046 8706 16098
rect 12350 16046 12402 16098
rect 12686 16046 12738 16098
rect 17614 16046 17666 16098
rect 24334 16046 24386 16098
rect 24558 16046 24610 16098
rect 24782 16046 24834 16098
rect 25790 16046 25842 16098
rect 29934 16046 29986 16098
rect 30270 16046 30322 16098
rect 4174 15934 4226 15986
rect 12910 15934 12962 15986
rect 21758 15934 21810 15986
rect 25118 15934 25170 15986
rect 1822 15822 1874 15874
rect 3054 15822 3106 15874
rect 5966 15822 6018 15874
rect 14142 15822 14194 15874
rect 17166 15822 17218 15874
rect 22206 15822 22258 15874
rect 22654 15822 22706 15874
rect 24222 15822 24274 15874
rect 24446 15822 24498 15874
rect 25230 15822 25282 15874
rect 25342 15822 25394 15874
rect 14024 15654 14076 15706
rect 14148 15654 14200 15706
rect 14272 15654 14324 15706
rect 14396 15654 14448 15706
rect 14520 15654 14572 15706
rect 14644 15654 14696 15706
rect 14768 15654 14820 15706
rect 14892 15654 14944 15706
rect 15016 15654 15068 15706
rect 15140 15654 15192 15706
rect 34024 15654 34076 15706
rect 34148 15654 34200 15706
rect 34272 15654 34324 15706
rect 34396 15654 34448 15706
rect 34520 15654 34572 15706
rect 34644 15654 34696 15706
rect 34768 15654 34820 15706
rect 34892 15654 34944 15706
rect 35016 15654 35068 15706
rect 35140 15654 35192 15706
rect 4734 15486 4786 15538
rect 5294 15486 5346 15538
rect 5854 15486 5906 15538
rect 6414 15486 6466 15538
rect 8430 15486 8482 15538
rect 8654 15486 8706 15538
rect 9662 15486 9714 15538
rect 9774 15486 9826 15538
rect 10558 15486 10610 15538
rect 12910 15486 12962 15538
rect 13358 15486 13410 15538
rect 21646 15486 21698 15538
rect 28478 15486 28530 15538
rect 29038 15486 29090 15538
rect 29598 15486 29650 15538
rect 5742 15374 5794 15426
rect 6078 15374 6130 15426
rect 7198 15374 7250 15426
rect 7534 15374 7586 15426
rect 9550 15374 9602 15426
rect 13918 15374 13970 15426
rect 23214 15374 23266 15426
rect 23550 15374 23602 15426
rect 30046 15374 30098 15426
rect 1822 15262 1874 15314
rect 2270 15262 2322 15314
rect 6862 15262 6914 15314
rect 7758 15262 7810 15314
rect 8206 15262 8258 15314
rect 8878 15262 8930 15314
rect 10222 15262 10274 15314
rect 11566 15262 11618 15314
rect 12238 15262 12290 15314
rect 12798 15262 12850 15314
rect 13134 15262 13186 15314
rect 13358 15262 13410 15314
rect 18734 15262 18786 15314
rect 19182 15262 19234 15314
rect 22990 15262 23042 15314
rect 25566 15262 25618 15314
rect 25902 15262 25954 15314
rect 7870 15150 7922 15202
rect 11006 15150 11058 15202
rect 12014 15150 12066 15202
rect 14366 15150 14418 15202
rect 22206 15150 22258 15202
rect 6974 15038 7026 15090
rect 8766 15038 8818 15090
rect 11790 15038 11842 15090
rect 12350 15038 12402 15090
rect 22654 15038 22706 15090
rect 4024 14870 4076 14922
rect 4148 14870 4200 14922
rect 4272 14870 4324 14922
rect 4396 14870 4448 14922
rect 4520 14870 4572 14922
rect 4644 14870 4696 14922
rect 4768 14870 4820 14922
rect 4892 14870 4944 14922
rect 5016 14870 5068 14922
rect 5140 14870 5192 14922
rect 24024 14870 24076 14922
rect 24148 14870 24200 14922
rect 24272 14870 24324 14922
rect 24396 14870 24448 14922
rect 24520 14870 24572 14922
rect 24644 14870 24696 14922
rect 24768 14870 24820 14922
rect 24892 14870 24944 14922
rect 25016 14870 25068 14922
rect 25140 14870 25192 14922
rect 4062 14702 4114 14754
rect 21646 14702 21698 14754
rect 22430 14702 22482 14754
rect 23886 14702 23938 14754
rect 5742 14590 5794 14642
rect 6974 14590 7026 14642
rect 7758 14590 7810 14642
rect 11454 14590 11506 14642
rect 12798 14590 12850 14642
rect 13582 14590 13634 14642
rect 17614 14590 17666 14642
rect 18062 14590 18114 14642
rect 18622 14590 18674 14642
rect 19854 14590 19906 14642
rect 21982 14590 22034 14642
rect 4846 14478 4898 14530
rect 7086 14478 7138 14530
rect 8430 14478 8482 14530
rect 9214 14478 9266 14530
rect 9774 14478 9826 14530
rect 11118 14478 11170 14530
rect 11902 14478 11954 14530
rect 12350 14478 12402 14530
rect 19182 14478 19234 14530
rect 20638 14478 20690 14530
rect 26910 14478 26962 14530
rect 27582 14478 27634 14530
rect 4734 14366 4786 14418
rect 8206 14366 8258 14418
rect 8766 14366 8818 14418
rect 9102 14366 9154 14418
rect 9998 14366 10050 14418
rect 10110 14366 10162 14418
rect 10334 14366 10386 14418
rect 15150 14366 15202 14418
rect 18846 14366 18898 14418
rect 18958 14366 19010 14418
rect 20526 14366 20578 14418
rect 3726 14254 3778 14306
rect 6190 14254 6242 14306
rect 9886 14254 9938 14306
rect 19518 14254 19570 14306
rect 22430 14254 22482 14306
rect 24670 14254 24722 14306
rect 27918 14254 27970 14306
rect 28366 14254 28418 14306
rect 14024 14086 14076 14138
rect 14148 14086 14200 14138
rect 14272 14086 14324 14138
rect 14396 14086 14448 14138
rect 14520 14086 14572 14138
rect 14644 14086 14696 14138
rect 14768 14086 14820 14138
rect 14892 14086 14944 14138
rect 15016 14086 15068 14138
rect 15140 14086 15192 14138
rect 34024 14086 34076 14138
rect 34148 14086 34200 14138
rect 34272 14086 34324 14138
rect 34396 14086 34448 14138
rect 34520 14086 34572 14138
rect 34644 14086 34696 14138
rect 34768 14086 34820 14138
rect 34892 14086 34944 14138
rect 35016 14086 35068 14138
rect 35140 14086 35192 14138
rect 5294 13918 5346 13970
rect 8094 13918 8146 13970
rect 10558 13918 10610 13970
rect 11118 13918 11170 13970
rect 12350 13918 12402 13970
rect 15598 13918 15650 13970
rect 16046 13918 16098 13970
rect 16830 13918 16882 13970
rect 25790 13918 25842 13970
rect 25902 13918 25954 13970
rect 26798 13918 26850 13970
rect 27358 13918 27410 13970
rect 9550 13806 9602 13858
rect 9886 13806 9938 13858
rect 11230 13806 11282 13858
rect 18062 13806 18114 13858
rect 18622 13806 18674 13858
rect 20190 13806 20242 13858
rect 21198 13806 21250 13858
rect 21758 13806 21810 13858
rect 7758 13694 7810 13746
rect 9102 13694 9154 13746
rect 10110 13694 10162 13746
rect 10782 13694 10834 13746
rect 11454 13694 11506 13746
rect 14254 13694 14306 13746
rect 14814 13694 14866 13746
rect 17838 13694 17890 13746
rect 20974 13694 21026 13746
rect 26014 13694 26066 13746
rect 26462 13694 26514 13746
rect 26686 13694 26738 13746
rect 8206 13582 8258 13634
rect 9662 13582 9714 13634
rect 12014 13582 12066 13634
rect 14926 13582 14978 13634
rect 17502 13470 17554 13522
rect 20638 13470 20690 13522
rect 26798 13470 26850 13522
rect 4024 13302 4076 13354
rect 4148 13302 4200 13354
rect 4272 13302 4324 13354
rect 4396 13302 4448 13354
rect 4520 13302 4572 13354
rect 4644 13302 4696 13354
rect 4768 13302 4820 13354
rect 4892 13302 4944 13354
rect 5016 13302 5068 13354
rect 5140 13302 5192 13354
rect 24024 13302 24076 13354
rect 24148 13302 24200 13354
rect 24272 13302 24324 13354
rect 24396 13302 24448 13354
rect 24520 13302 24572 13354
rect 24644 13302 24696 13354
rect 24768 13302 24820 13354
rect 24892 13302 24944 13354
rect 25016 13302 25068 13354
rect 25140 13302 25192 13354
rect 3502 13134 3554 13186
rect 7646 13134 7698 13186
rect 9326 13134 9378 13186
rect 9662 13134 9714 13186
rect 14030 13134 14082 13186
rect 19966 13134 20018 13186
rect 23214 13134 23266 13186
rect 24558 13134 24610 13186
rect 4846 13022 4898 13074
rect 5742 13022 5794 13074
rect 8766 13022 8818 13074
rect 9550 13022 9602 13074
rect 22430 13022 22482 13074
rect 26574 13022 26626 13074
rect 4286 12910 4338 12962
rect 6974 12910 7026 12962
rect 7198 12910 7250 12962
rect 8318 12910 8370 12962
rect 10782 12910 10834 12962
rect 11230 12910 11282 12962
rect 11454 12910 11506 12962
rect 15822 12910 15874 12962
rect 16382 12910 16434 12962
rect 16942 12910 16994 12962
rect 24446 12910 24498 12962
rect 27806 12910 27858 12962
rect 4062 12798 4114 12850
rect 7086 12798 7138 12850
rect 8766 12798 8818 12850
rect 8878 12798 8930 12850
rect 10334 12798 10386 12850
rect 12910 12798 12962 12850
rect 14366 12798 14418 12850
rect 14590 12798 14642 12850
rect 23438 12798 23490 12850
rect 23998 12798 24050 12850
rect 3166 12686 3218 12738
rect 9102 12686 9154 12738
rect 11342 12686 11394 12738
rect 13694 12686 13746 12738
rect 15374 12686 15426 12738
rect 15598 12686 15650 12738
rect 15710 12686 15762 12738
rect 19182 12686 19234 12738
rect 20302 12686 20354 12738
rect 22878 12686 22930 12738
rect 14024 12518 14076 12570
rect 14148 12518 14200 12570
rect 14272 12518 14324 12570
rect 14396 12518 14448 12570
rect 14520 12518 14572 12570
rect 14644 12518 14696 12570
rect 14768 12518 14820 12570
rect 14892 12518 14944 12570
rect 15016 12518 15068 12570
rect 15140 12518 15192 12570
rect 34024 12518 34076 12570
rect 34148 12518 34200 12570
rect 34272 12518 34324 12570
rect 34396 12518 34448 12570
rect 34520 12518 34572 12570
rect 34644 12518 34696 12570
rect 34768 12518 34820 12570
rect 34892 12518 34944 12570
rect 35016 12518 35068 12570
rect 35140 12518 35192 12570
rect 4846 12350 4898 12402
rect 6078 12350 6130 12402
rect 8206 12350 8258 12402
rect 8542 12350 8594 12402
rect 8990 12350 9042 12402
rect 10334 12350 10386 12402
rect 10558 12350 10610 12402
rect 10894 12350 10946 12402
rect 13246 12350 13298 12402
rect 13918 12350 13970 12402
rect 17502 12350 17554 12402
rect 20414 12350 20466 12402
rect 28254 12350 28306 12402
rect 6862 12238 6914 12290
rect 1822 12126 1874 12178
rect 2382 12126 2434 12178
rect 6526 12126 6578 12178
rect 6750 12126 6802 12178
rect 7086 12126 7138 12178
rect 7534 12126 7586 12178
rect 7758 12126 7810 12178
rect 10222 12126 10274 12178
rect 16270 12126 16322 12178
rect 16718 12126 16770 12178
rect 19854 12126 19906 12178
rect 27358 12126 27410 12178
rect 7310 12014 7362 12066
rect 17950 12014 18002 12066
rect 22430 12014 22482 12066
rect 5406 11902 5458 11954
rect 25454 11902 25506 11954
rect 4024 11734 4076 11786
rect 4148 11734 4200 11786
rect 4272 11734 4324 11786
rect 4396 11734 4448 11786
rect 4520 11734 4572 11786
rect 4644 11734 4696 11786
rect 4768 11734 4820 11786
rect 4892 11734 4944 11786
rect 5016 11734 5068 11786
rect 5140 11734 5192 11786
rect 24024 11734 24076 11786
rect 24148 11734 24200 11786
rect 24272 11734 24324 11786
rect 24396 11734 24448 11786
rect 24520 11734 24572 11786
rect 24644 11734 24696 11786
rect 24768 11734 24820 11786
rect 24892 11734 24944 11786
rect 25016 11734 25068 11786
rect 25140 11734 25192 11786
rect 3390 11566 3442 11618
rect 3726 11566 3778 11618
rect 6974 11566 7026 11618
rect 11678 11566 11730 11618
rect 25790 11566 25842 11618
rect 5070 11454 5122 11506
rect 7534 11454 7586 11506
rect 17390 11454 17442 11506
rect 26126 11454 26178 11506
rect 4398 11342 4450 11394
rect 6862 11342 6914 11394
rect 7982 11342 8034 11394
rect 8654 11342 8706 11394
rect 13582 11342 13634 11394
rect 13918 11342 13970 11394
rect 22318 11342 22370 11394
rect 22766 11342 22818 11394
rect 4510 11230 4562 11282
rect 6974 11230 7026 11282
rect 17838 11230 17890 11282
rect 5742 11118 5794 11170
rect 10894 11118 10946 11170
rect 12014 11118 12066 11170
rect 12462 11118 12514 11170
rect 16382 11118 16434 11170
rect 17054 11118 17106 11170
rect 25006 11118 25058 11170
rect 26574 11118 26626 11170
rect 14024 10950 14076 11002
rect 14148 10950 14200 11002
rect 14272 10950 14324 11002
rect 14396 10950 14448 11002
rect 14520 10950 14572 11002
rect 14644 10950 14696 11002
rect 14768 10950 14820 11002
rect 14892 10950 14944 11002
rect 15016 10950 15068 11002
rect 15140 10950 15192 11002
rect 34024 10950 34076 11002
rect 34148 10950 34200 11002
rect 34272 10950 34324 11002
rect 34396 10950 34448 11002
rect 34520 10950 34572 11002
rect 34644 10950 34696 11002
rect 34768 10950 34820 11002
rect 34892 10950 34944 11002
rect 35016 10950 35068 11002
rect 35140 10950 35192 11002
rect 4734 10782 4786 10834
rect 5294 10782 5346 10834
rect 5406 10782 5458 10834
rect 5966 10782 6018 10834
rect 9662 10782 9714 10834
rect 10110 10782 10162 10834
rect 13246 10782 13298 10834
rect 14030 10782 14082 10834
rect 14590 10782 14642 10834
rect 15486 10782 15538 10834
rect 15934 10782 15986 10834
rect 22542 10782 22594 10834
rect 23214 10782 23266 10834
rect 23662 10782 23714 10834
rect 15150 10670 15202 10722
rect 15262 10670 15314 10722
rect 23998 10670 24050 10722
rect 1822 10558 1874 10610
rect 2270 10558 2322 10610
rect 8430 10558 8482 10610
rect 8878 10558 8930 10610
rect 10334 10558 10386 10610
rect 11006 10558 11058 10610
rect 19742 10558 19794 10610
rect 20190 10558 20242 10610
rect 4024 10166 4076 10218
rect 4148 10166 4200 10218
rect 4272 10166 4324 10218
rect 4396 10166 4448 10218
rect 4520 10166 4572 10218
rect 4644 10166 4696 10218
rect 4768 10166 4820 10218
rect 4892 10166 4944 10218
rect 5016 10166 5068 10218
rect 5140 10166 5192 10218
rect 24024 10166 24076 10218
rect 24148 10166 24200 10218
rect 24272 10166 24324 10218
rect 24396 10166 24448 10218
rect 24520 10166 24572 10218
rect 24644 10166 24696 10218
rect 24768 10166 24820 10218
rect 24892 10166 24944 10218
rect 25016 10166 25068 10218
rect 25140 10166 25192 10218
rect 6190 9886 6242 9938
rect 27022 9886 27074 9938
rect 28030 9662 28082 9714
rect 5742 9550 5794 9602
rect 9214 9550 9266 9602
rect 14024 9382 14076 9434
rect 14148 9382 14200 9434
rect 14272 9382 14324 9434
rect 14396 9382 14448 9434
rect 14520 9382 14572 9434
rect 14644 9382 14696 9434
rect 14768 9382 14820 9434
rect 14892 9382 14944 9434
rect 15016 9382 15068 9434
rect 15140 9382 15192 9434
rect 34024 9382 34076 9434
rect 34148 9382 34200 9434
rect 34272 9382 34324 9434
rect 34396 9382 34448 9434
rect 34520 9382 34572 9434
rect 34644 9382 34696 9434
rect 34768 9382 34820 9434
rect 34892 9382 34944 9434
rect 35016 9382 35068 9434
rect 35140 9382 35192 9434
rect 18958 9102 19010 9154
rect 28030 9102 28082 9154
rect 29038 9102 29090 9154
rect 18734 8990 18786 9042
rect 19070 8990 19122 9042
rect 25342 8990 25394 9042
rect 25790 8990 25842 9042
rect 29598 8990 29650 9042
rect 22990 8766 23042 8818
rect 28814 8766 28866 8818
rect 4024 8598 4076 8650
rect 4148 8598 4200 8650
rect 4272 8598 4324 8650
rect 4396 8598 4448 8650
rect 4520 8598 4572 8650
rect 4644 8598 4696 8650
rect 4768 8598 4820 8650
rect 4892 8598 4944 8650
rect 5016 8598 5068 8650
rect 5140 8598 5192 8650
rect 24024 8598 24076 8650
rect 24148 8598 24200 8650
rect 24272 8598 24324 8650
rect 24396 8598 24448 8650
rect 24520 8598 24572 8650
rect 24644 8598 24696 8650
rect 24768 8598 24820 8650
rect 24892 8598 24944 8650
rect 25016 8598 25068 8650
rect 25140 8598 25192 8650
rect 19406 8430 19458 8482
rect 27582 8430 27634 8482
rect 7982 8318 8034 8370
rect 25902 8318 25954 8370
rect 26350 8318 26402 8370
rect 27246 8318 27298 8370
rect 17950 8206 18002 8258
rect 18398 8206 18450 8258
rect 19294 8206 19346 8258
rect 22318 8206 22370 8258
rect 22878 8206 22930 8258
rect 28254 8206 28306 8258
rect 17614 8094 17666 8146
rect 18062 8094 18114 8146
rect 18734 8094 18786 8146
rect 18958 8094 19010 8146
rect 19966 8094 20018 8146
rect 20302 8094 20354 8146
rect 28366 8094 28418 8146
rect 5854 7982 5906 8034
rect 17838 7982 17890 8034
rect 18510 7982 18562 8034
rect 19518 7982 19570 8034
rect 19742 7982 19794 8034
rect 20190 7982 20242 8034
rect 25342 7982 25394 8034
rect 14024 7814 14076 7866
rect 14148 7814 14200 7866
rect 14272 7814 14324 7866
rect 14396 7814 14448 7866
rect 14520 7814 14572 7866
rect 14644 7814 14696 7866
rect 14768 7814 14820 7866
rect 14892 7814 14944 7866
rect 15016 7814 15068 7866
rect 15140 7814 15192 7866
rect 34024 7814 34076 7866
rect 34148 7814 34200 7866
rect 34272 7814 34324 7866
rect 34396 7814 34448 7866
rect 34520 7814 34572 7866
rect 34644 7814 34696 7866
rect 34768 7814 34820 7866
rect 34892 7814 34944 7866
rect 35016 7814 35068 7866
rect 35140 7814 35192 7866
rect 4734 7646 4786 7698
rect 6078 7646 6130 7698
rect 15598 7646 15650 7698
rect 16830 7646 16882 7698
rect 20638 7646 20690 7698
rect 21198 7646 21250 7698
rect 21422 7646 21474 7698
rect 7982 7534 8034 7586
rect 8542 7534 8594 7586
rect 11902 7534 11954 7586
rect 24670 7534 24722 7586
rect 26014 7534 26066 7586
rect 27022 7534 27074 7586
rect 27582 7534 27634 7586
rect 1822 7422 1874 7474
rect 2158 7422 2210 7474
rect 6862 7422 6914 7474
rect 7534 7422 7586 7474
rect 8094 7422 8146 7474
rect 8430 7422 8482 7474
rect 8766 7422 8818 7474
rect 14254 7422 14306 7474
rect 14590 7422 14642 7474
rect 15150 7422 15202 7474
rect 17502 7422 17554 7474
rect 18174 7422 18226 7474
rect 26350 7422 26402 7474
rect 27134 7422 27186 7474
rect 5630 7310 5682 7362
rect 6638 7310 6690 7362
rect 9662 7310 9714 7362
rect 10110 7310 10162 7362
rect 21534 7310 21586 7362
rect 5294 7198 5346 7250
rect 6526 7198 6578 7250
rect 7982 7198 8034 7250
rect 11118 7198 11170 7250
rect 4024 7030 4076 7082
rect 4148 7030 4200 7082
rect 4272 7030 4324 7082
rect 4396 7030 4448 7082
rect 4520 7030 4572 7082
rect 4644 7030 4696 7082
rect 4768 7030 4820 7082
rect 4892 7030 4944 7082
rect 5016 7030 5068 7082
rect 5140 7030 5192 7082
rect 24024 7030 24076 7082
rect 24148 7030 24200 7082
rect 24272 7030 24324 7082
rect 24396 7030 24448 7082
rect 24520 7030 24572 7082
rect 24644 7030 24696 7082
rect 24768 7030 24820 7082
rect 24892 7030 24944 7082
rect 25016 7030 25068 7082
rect 25140 7030 25192 7082
rect 5742 6862 5794 6914
rect 6190 6862 6242 6914
rect 6302 6862 6354 6914
rect 6750 6862 6802 6914
rect 6974 6862 7026 6914
rect 8094 6862 8146 6914
rect 21310 6862 21362 6914
rect 4510 6750 4562 6802
rect 15038 6750 15090 6802
rect 21422 6750 21474 6802
rect 26798 6750 26850 6802
rect 2270 6638 2322 6690
rect 2494 6638 2546 6690
rect 4062 6638 4114 6690
rect 5854 6638 5906 6690
rect 7758 6638 7810 6690
rect 8542 6638 8594 6690
rect 9214 6638 9266 6690
rect 9326 6638 9378 6690
rect 9998 6638 10050 6690
rect 17054 6638 17106 6690
rect 17726 6638 17778 6690
rect 22094 6638 22146 6690
rect 22430 6638 22482 6690
rect 2606 6526 2658 6578
rect 2942 6526 2994 6578
rect 3614 6526 3666 6578
rect 6414 6526 6466 6578
rect 7534 6526 7586 6578
rect 7982 6526 8034 6578
rect 12238 6526 12290 6578
rect 13022 6526 13074 6578
rect 13918 6526 13970 6578
rect 16718 6526 16770 6578
rect 16830 6526 16882 6578
rect 25566 6526 25618 6578
rect 27806 6526 27858 6578
rect 3054 6414 3106 6466
rect 3278 6414 3330 6466
rect 5742 6414 5794 6466
rect 8654 6414 8706 6466
rect 8766 6414 8818 6466
rect 16494 6414 16546 6466
rect 20078 6414 20130 6466
rect 20750 6414 20802 6466
rect 25006 6414 25058 6466
rect 26014 6414 26066 6466
rect 14024 6246 14076 6298
rect 14148 6246 14200 6298
rect 14272 6246 14324 6298
rect 14396 6246 14448 6298
rect 14520 6246 14572 6298
rect 14644 6246 14696 6298
rect 14768 6246 14820 6298
rect 14892 6246 14944 6298
rect 15016 6246 15068 6298
rect 15140 6246 15192 6298
rect 34024 6246 34076 6298
rect 34148 6246 34200 6298
rect 34272 6246 34324 6298
rect 34396 6246 34448 6298
rect 34520 6246 34572 6298
rect 34644 6246 34696 6298
rect 34768 6246 34820 6298
rect 34892 6246 34944 6298
rect 35016 6246 35068 6298
rect 35140 6246 35192 6298
rect 7310 6078 7362 6130
rect 7870 6078 7922 6130
rect 8990 6078 9042 6130
rect 12350 6078 12402 6130
rect 13246 6078 13298 6130
rect 13806 6078 13858 6130
rect 17502 6078 17554 6130
rect 18286 6078 18338 6130
rect 18398 6078 18450 6130
rect 18622 6078 18674 6130
rect 28142 6078 28194 6130
rect 28814 6078 28866 6130
rect 2494 5966 2546 6018
rect 3166 5966 3218 6018
rect 3502 5966 3554 6018
rect 8318 5966 8370 6018
rect 17614 5966 17666 6018
rect 2830 5854 2882 5906
rect 4174 5854 4226 5906
rect 4734 5854 4786 5906
rect 8430 5854 8482 5906
rect 8542 5854 8594 5906
rect 9438 5854 9490 5906
rect 9998 5854 10050 5906
rect 16382 5854 16434 5906
rect 16830 5854 16882 5906
rect 17278 5854 17330 5906
rect 18174 5854 18226 5906
rect 24334 5854 24386 5906
rect 25342 5854 25394 5906
rect 25790 5854 25842 5906
rect 2046 5742 2098 5794
rect 3614 5742 3666 5794
rect 22318 5742 22370 5794
rect 2382 5630 2434 5682
rect 13134 5630 13186 5682
rect 4024 5462 4076 5514
rect 4148 5462 4200 5514
rect 4272 5462 4324 5514
rect 4396 5462 4448 5514
rect 4520 5462 4572 5514
rect 4644 5462 4696 5514
rect 4768 5462 4820 5514
rect 4892 5462 4944 5514
rect 5016 5462 5068 5514
rect 5140 5462 5192 5514
rect 24024 5462 24076 5514
rect 24148 5462 24200 5514
rect 24272 5462 24324 5514
rect 24396 5462 24448 5514
rect 24520 5462 24572 5514
rect 24644 5462 24696 5514
rect 24768 5462 24820 5514
rect 24892 5462 24944 5514
rect 25016 5462 25068 5514
rect 25140 5462 25192 5514
rect 6862 5294 6914 5346
rect 22206 5294 22258 5346
rect 5966 5182 6018 5234
rect 11342 5182 11394 5234
rect 13582 5182 13634 5234
rect 14030 5182 14082 5234
rect 21310 5182 21362 5234
rect 25342 5182 25394 5234
rect 5742 5070 5794 5122
rect 5854 5070 5906 5122
rect 6078 5070 6130 5122
rect 6302 5070 6354 5122
rect 9886 5070 9938 5122
rect 10334 5070 10386 5122
rect 10894 5070 10946 5122
rect 20414 5070 20466 5122
rect 22542 5070 22594 5122
rect 15374 4958 15426 5010
rect 7534 4846 7586 4898
rect 14024 4678 14076 4730
rect 14148 4678 14200 4730
rect 14272 4678 14324 4730
rect 14396 4678 14448 4730
rect 14520 4678 14572 4730
rect 14644 4678 14696 4730
rect 14768 4678 14820 4730
rect 14892 4678 14944 4730
rect 15016 4678 15068 4730
rect 15140 4678 15192 4730
rect 34024 4678 34076 4730
rect 34148 4678 34200 4730
rect 34272 4678 34324 4730
rect 34396 4678 34448 4730
rect 34520 4678 34572 4730
rect 34644 4678 34696 4730
rect 34768 4678 34820 4730
rect 34892 4678 34944 4730
rect 35016 4678 35068 4730
rect 35140 4678 35192 4730
rect 4734 4510 4786 4562
rect 6078 4510 6130 4562
rect 6302 4510 6354 4562
rect 6414 4510 6466 4562
rect 6526 4510 6578 4562
rect 8318 4510 8370 4562
rect 8878 4510 8930 4562
rect 9102 4510 9154 4562
rect 12574 4510 12626 4562
rect 16382 4510 16434 4562
rect 26910 4510 26962 4562
rect 5406 4398 5458 4450
rect 7422 4398 7474 4450
rect 8430 4398 8482 4450
rect 8766 4398 8818 4450
rect 18062 4398 18114 4450
rect 23998 4398 24050 4450
rect 24782 4398 24834 4450
rect 25902 4398 25954 4450
rect 1710 4286 1762 4338
rect 2270 4286 2322 4338
rect 6974 4286 7026 4338
rect 8094 4286 8146 4338
rect 9662 4286 9714 4338
rect 10110 4286 10162 4338
rect 13246 4286 13298 4338
rect 13918 4286 13970 4338
rect 20414 4286 20466 4338
rect 20974 4286 21026 4338
rect 21086 4286 21138 4338
rect 21758 4286 21810 4338
rect 25790 4286 25842 4338
rect 7310 4174 7362 4226
rect 25454 4174 25506 4226
rect 13134 4062 13186 4114
rect 16942 4062 16994 4114
rect 17278 4062 17330 4114
rect 26574 4062 26626 4114
rect 4024 3894 4076 3946
rect 4148 3894 4200 3946
rect 4272 3894 4324 3946
rect 4396 3894 4448 3946
rect 4520 3894 4572 3946
rect 4644 3894 4696 3946
rect 4768 3894 4820 3946
rect 4892 3894 4944 3946
rect 5016 3894 5068 3946
rect 5140 3894 5192 3946
rect 24024 3894 24076 3946
rect 24148 3894 24200 3946
rect 24272 3894 24324 3946
rect 24396 3894 24448 3946
rect 24520 3894 24572 3946
rect 24644 3894 24696 3946
rect 24768 3894 24820 3946
rect 24892 3894 24944 3946
rect 25016 3894 25068 3946
rect 25140 3894 25192 3946
rect 19742 3726 19794 3778
rect 5966 3614 6018 3666
rect 6414 3614 6466 3666
rect 8318 3614 8370 3666
rect 16942 3614 16994 3666
rect 19854 3614 19906 3666
rect 21982 3614 22034 3666
rect 13246 3390 13298 3442
rect 13694 3390 13746 3442
rect 16158 3390 16210 3442
rect 17950 3390 18002 3442
rect 18734 3390 18786 3442
rect 19070 3390 19122 3442
rect 20862 3390 20914 3442
rect 14024 3110 14076 3162
rect 14148 3110 14200 3162
rect 14272 3110 14324 3162
rect 14396 3110 14448 3162
rect 14520 3110 14572 3162
rect 14644 3110 14696 3162
rect 14768 3110 14820 3162
rect 14892 3110 14944 3162
rect 15016 3110 15068 3162
rect 15140 3110 15192 3162
rect 34024 3110 34076 3162
rect 34148 3110 34200 3162
rect 34272 3110 34324 3162
rect 34396 3110 34448 3162
rect 34520 3110 34572 3162
rect 34644 3110 34696 3162
rect 34768 3110 34820 3162
rect 34892 3110 34944 3162
rect 35016 3110 35068 3162
rect 35140 3110 35192 3162
<< metal2 >>
rect 9856 99200 9968 100000
rect 29792 99200 29904 100000
rect 4008 96460 5208 96470
rect 4064 96458 4112 96460
rect 4168 96458 4216 96460
rect 4076 96406 4112 96458
rect 4200 96406 4216 96458
rect 4064 96404 4112 96406
rect 4168 96404 4216 96406
rect 4272 96458 4320 96460
rect 4376 96458 4424 96460
rect 4480 96458 4528 96460
rect 4376 96406 4396 96458
rect 4480 96406 4520 96458
rect 4272 96404 4320 96406
rect 4376 96404 4424 96406
rect 4480 96404 4528 96406
rect 4584 96404 4632 96460
rect 4688 96458 4736 96460
rect 4792 96458 4840 96460
rect 4896 96458 4944 96460
rect 4696 96406 4736 96458
rect 4820 96406 4840 96458
rect 4688 96404 4736 96406
rect 4792 96404 4840 96406
rect 4896 96404 4944 96406
rect 5000 96458 5048 96460
rect 5104 96458 5152 96460
rect 5000 96406 5016 96458
rect 5104 96406 5140 96458
rect 5000 96404 5048 96406
rect 5104 96404 5152 96406
rect 4008 96394 5208 96404
rect 1708 95842 1764 95854
rect 1708 95790 1710 95842
rect 1762 95790 1764 95842
rect 1708 95284 1764 95790
rect 1708 95218 1764 95228
rect 4008 94892 5208 94902
rect 4064 94890 4112 94892
rect 4168 94890 4216 94892
rect 4076 94838 4112 94890
rect 4200 94838 4216 94890
rect 4064 94836 4112 94838
rect 4168 94836 4216 94838
rect 4272 94890 4320 94892
rect 4376 94890 4424 94892
rect 4480 94890 4528 94892
rect 4376 94838 4396 94890
rect 4480 94838 4520 94890
rect 4272 94836 4320 94838
rect 4376 94836 4424 94838
rect 4480 94836 4528 94838
rect 4584 94836 4632 94892
rect 4688 94890 4736 94892
rect 4792 94890 4840 94892
rect 4896 94890 4944 94892
rect 4696 94838 4736 94890
rect 4820 94838 4840 94890
rect 4688 94836 4736 94838
rect 4792 94836 4840 94838
rect 4896 94836 4944 94838
rect 5000 94890 5048 94892
rect 5104 94890 5152 94892
rect 5000 94838 5016 94890
rect 5104 94838 5140 94890
rect 5000 94836 5048 94838
rect 5104 94836 5152 94838
rect 4008 94826 5208 94836
rect 1708 94276 1764 94286
rect 1708 94182 1764 94220
rect 9884 94164 9940 99200
rect 29820 97412 29876 99200
rect 29820 97356 30100 97412
rect 24008 96460 25208 96470
rect 24064 96458 24112 96460
rect 24168 96458 24216 96460
rect 24076 96406 24112 96458
rect 24200 96406 24216 96458
rect 24064 96404 24112 96406
rect 24168 96404 24216 96406
rect 24272 96458 24320 96460
rect 24376 96458 24424 96460
rect 24480 96458 24528 96460
rect 24376 96406 24396 96458
rect 24480 96406 24520 96458
rect 24272 96404 24320 96406
rect 24376 96404 24424 96406
rect 24480 96404 24528 96406
rect 24584 96404 24632 96460
rect 24688 96458 24736 96460
rect 24792 96458 24840 96460
rect 24896 96458 24944 96460
rect 24696 96406 24736 96458
rect 24820 96406 24840 96458
rect 24688 96404 24736 96406
rect 24792 96404 24840 96406
rect 24896 96404 24944 96406
rect 25000 96458 25048 96460
rect 25104 96458 25152 96460
rect 25000 96406 25016 96458
rect 25104 96406 25140 96458
rect 25000 96404 25048 96406
rect 25104 96404 25152 96406
rect 24008 96394 25208 96404
rect 30044 95954 30100 97356
rect 30268 96068 30324 96078
rect 30044 95902 30046 95954
rect 30098 95902 30100 95954
rect 30044 95890 30100 95902
rect 30156 96066 30324 96068
rect 30156 96014 30270 96066
rect 30322 96014 30324 96066
rect 30156 96012 30324 96014
rect 29820 95842 29876 95854
rect 29820 95790 29822 95842
rect 29874 95790 29876 95842
rect 29820 95732 29876 95790
rect 30156 95732 30212 96012
rect 30268 96002 30324 96012
rect 14008 95676 15208 95686
rect 14064 95674 14112 95676
rect 14168 95674 14216 95676
rect 14076 95622 14112 95674
rect 14200 95622 14216 95674
rect 14064 95620 14112 95622
rect 14168 95620 14216 95622
rect 14272 95674 14320 95676
rect 14376 95674 14424 95676
rect 14480 95674 14528 95676
rect 14376 95622 14396 95674
rect 14480 95622 14520 95674
rect 14272 95620 14320 95622
rect 14376 95620 14424 95622
rect 14480 95620 14528 95622
rect 14584 95620 14632 95676
rect 14688 95674 14736 95676
rect 14792 95674 14840 95676
rect 14896 95674 14944 95676
rect 14696 95622 14736 95674
rect 14820 95622 14840 95674
rect 14688 95620 14736 95622
rect 14792 95620 14840 95622
rect 14896 95620 14944 95622
rect 15000 95674 15048 95676
rect 15104 95674 15152 95676
rect 15000 95622 15016 95674
rect 15104 95622 15140 95674
rect 15000 95620 15048 95622
rect 15104 95620 15152 95622
rect 14008 95610 15208 95620
rect 29820 95676 30212 95732
rect 34008 95676 35208 95686
rect 24008 94892 25208 94902
rect 24064 94890 24112 94892
rect 24168 94890 24216 94892
rect 24076 94838 24112 94890
rect 24200 94838 24216 94890
rect 24064 94836 24112 94838
rect 24168 94836 24216 94838
rect 24272 94890 24320 94892
rect 24376 94890 24424 94892
rect 24480 94890 24528 94892
rect 24376 94838 24396 94890
rect 24480 94838 24520 94890
rect 24272 94836 24320 94838
rect 24376 94836 24424 94838
rect 24480 94836 24528 94838
rect 24584 94836 24632 94892
rect 24688 94890 24736 94892
rect 24792 94890 24840 94892
rect 24896 94890 24944 94892
rect 24696 94838 24736 94890
rect 24820 94838 24840 94890
rect 24688 94836 24736 94838
rect 24792 94836 24840 94838
rect 24896 94836 24944 94838
rect 25000 94890 25048 94892
rect 25104 94890 25152 94892
rect 25000 94838 25016 94890
rect 25104 94838 25140 94890
rect 25000 94836 25048 94838
rect 25104 94836 25152 94838
rect 24008 94826 25208 94836
rect 9884 94098 9940 94108
rect 12908 94164 12964 94174
rect 1708 93826 1764 93838
rect 1708 93774 1710 93826
rect 1762 93774 1764 93826
rect 1708 93044 1764 93774
rect 4008 93324 5208 93334
rect 4064 93322 4112 93324
rect 4168 93322 4216 93324
rect 4076 93270 4112 93322
rect 4200 93270 4216 93322
rect 4064 93268 4112 93270
rect 4168 93268 4216 93270
rect 4272 93322 4320 93324
rect 4376 93322 4424 93324
rect 4480 93322 4528 93324
rect 4376 93270 4396 93322
rect 4480 93270 4520 93322
rect 4272 93268 4320 93270
rect 4376 93268 4424 93270
rect 4480 93268 4528 93270
rect 4584 93268 4632 93324
rect 4688 93322 4736 93324
rect 4792 93322 4840 93324
rect 4896 93322 4944 93324
rect 4696 93270 4736 93322
rect 4820 93270 4840 93322
rect 4688 93268 4736 93270
rect 4792 93268 4840 93270
rect 4896 93268 4944 93270
rect 5000 93322 5048 93324
rect 5104 93322 5152 93324
rect 5000 93270 5016 93322
rect 5104 93270 5140 93322
rect 5000 93268 5048 93270
rect 5104 93268 5152 93270
rect 4008 93258 5208 93268
rect 1708 92978 1764 92988
rect 1708 92258 1764 92270
rect 1708 92206 1710 92258
rect 1762 92206 1764 92258
rect 1708 91924 1764 92206
rect 1708 91858 1764 91868
rect 4008 91756 5208 91766
rect 4064 91754 4112 91756
rect 4168 91754 4216 91756
rect 4076 91702 4112 91754
rect 4200 91702 4216 91754
rect 4064 91700 4112 91702
rect 4168 91700 4216 91702
rect 4272 91754 4320 91756
rect 4376 91754 4424 91756
rect 4480 91754 4528 91756
rect 4376 91702 4396 91754
rect 4480 91702 4520 91754
rect 4272 91700 4320 91702
rect 4376 91700 4424 91702
rect 4480 91700 4528 91702
rect 4584 91700 4632 91756
rect 4688 91754 4736 91756
rect 4792 91754 4840 91756
rect 4896 91754 4944 91756
rect 4696 91702 4736 91754
rect 4820 91702 4840 91754
rect 4688 91700 4736 91702
rect 4792 91700 4840 91702
rect 4896 91700 4944 91702
rect 5000 91754 5048 91756
rect 5104 91754 5152 91756
rect 5000 91702 5016 91754
rect 5104 91702 5140 91754
rect 5000 91700 5048 91702
rect 5104 91700 5152 91702
rect 4008 91690 5208 91700
rect 1708 91138 1764 91150
rect 1708 91086 1710 91138
rect 1762 91086 1764 91138
rect 1708 90804 1764 91086
rect 1708 90738 1764 90748
rect 4008 90188 5208 90198
rect 4064 90186 4112 90188
rect 4168 90186 4216 90188
rect 4076 90134 4112 90186
rect 4200 90134 4216 90186
rect 4064 90132 4112 90134
rect 4168 90132 4216 90134
rect 4272 90186 4320 90188
rect 4376 90186 4424 90188
rect 4480 90186 4528 90188
rect 4376 90134 4396 90186
rect 4480 90134 4520 90186
rect 4272 90132 4320 90134
rect 4376 90132 4424 90134
rect 4480 90132 4528 90134
rect 4584 90132 4632 90188
rect 4688 90186 4736 90188
rect 4792 90186 4840 90188
rect 4896 90186 4944 90188
rect 4696 90134 4736 90186
rect 4820 90134 4840 90186
rect 4688 90132 4736 90134
rect 4792 90132 4840 90134
rect 4896 90132 4944 90134
rect 5000 90186 5048 90188
rect 5104 90186 5152 90188
rect 5000 90134 5016 90186
rect 5104 90134 5140 90186
rect 5000 90132 5048 90134
rect 5104 90132 5152 90134
rect 4008 90122 5208 90132
rect 1708 89684 1764 89694
rect 1708 89590 1764 89628
rect 1708 89122 1764 89134
rect 1708 89070 1710 89122
rect 1762 89070 1764 89122
rect 1708 88564 1764 89070
rect 12348 89122 12404 89134
rect 12348 89070 12350 89122
rect 12402 89070 12404 89122
rect 9436 89010 9492 89022
rect 9436 88958 9438 89010
rect 9490 88958 9492 89010
rect 8540 88900 8596 88910
rect 8988 88900 9044 88910
rect 9436 88900 9492 88958
rect 8540 88898 9492 88900
rect 8540 88846 8542 88898
rect 8594 88846 8990 88898
rect 9042 88846 9492 88898
rect 8540 88844 9492 88846
rect 9996 89010 10052 89022
rect 9996 88958 9998 89010
rect 10050 88958 10052 89010
rect 8540 88834 8596 88844
rect 4008 88620 5208 88630
rect 4064 88618 4112 88620
rect 4168 88618 4216 88620
rect 4076 88566 4112 88618
rect 4200 88566 4216 88618
rect 4064 88564 4112 88566
rect 4168 88564 4216 88566
rect 4272 88618 4320 88620
rect 4376 88618 4424 88620
rect 4480 88618 4528 88620
rect 4376 88566 4396 88618
rect 4480 88566 4520 88618
rect 4272 88564 4320 88566
rect 4376 88564 4424 88566
rect 4480 88564 4528 88566
rect 4584 88564 4632 88620
rect 4688 88618 4736 88620
rect 4792 88618 4840 88620
rect 4896 88618 4944 88620
rect 4696 88566 4736 88618
rect 4820 88566 4840 88618
rect 4688 88564 4736 88566
rect 4792 88564 4840 88566
rect 4896 88564 4944 88566
rect 5000 88618 5048 88620
rect 5104 88618 5152 88620
rect 5000 88566 5016 88618
rect 5104 88566 5140 88618
rect 5000 88564 5048 88566
rect 5104 88564 5152 88566
rect 4008 88554 5208 88564
rect 1708 88498 1764 88508
rect 1708 88002 1764 88014
rect 1708 87950 1710 88002
rect 1762 87950 1764 88002
rect 1708 87444 1764 87950
rect 8428 88004 8484 88014
rect 8428 87666 8484 87948
rect 8428 87614 8430 87666
rect 8482 87614 8484 87666
rect 8428 87602 8484 87614
rect 8876 88004 8932 88014
rect 8988 88004 9044 88844
rect 9100 88226 9156 88238
rect 9100 88174 9102 88226
rect 9154 88174 9156 88226
rect 9100 88004 9156 88174
rect 9772 88228 9828 88238
rect 9772 88134 9828 88172
rect 8876 88002 9156 88004
rect 8876 87950 8878 88002
rect 8930 87950 9156 88002
rect 8876 87948 9156 87950
rect 1708 87378 1764 87388
rect 5628 87444 5684 87454
rect 5628 87350 5684 87388
rect 6076 87442 6132 87454
rect 6076 87390 6078 87442
rect 6130 87390 6132 87442
rect 4008 87052 5208 87062
rect 4064 87050 4112 87052
rect 4168 87050 4216 87052
rect 4076 86998 4112 87050
rect 4200 86998 4216 87050
rect 4064 86996 4112 86998
rect 4168 86996 4216 86998
rect 4272 87050 4320 87052
rect 4376 87050 4424 87052
rect 4480 87050 4528 87052
rect 4376 86998 4396 87050
rect 4480 86998 4520 87050
rect 4272 86996 4320 86998
rect 4376 86996 4424 86998
rect 4480 86996 4528 86998
rect 4584 86996 4632 87052
rect 4688 87050 4736 87052
rect 4792 87050 4840 87052
rect 4896 87050 4944 87052
rect 4696 86998 4736 87050
rect 4820 86998 4840 87050
rect 4688 86996 4736 86998
rect 4792 86996 4840 86998
rect 4896 86996 4944 86998
rect 5000 87050 5048 87052
rect 5104 87050 5152 87052
rect 5000 86998 5016 87050
rect 5104 86998 5140 87050
rect 5000 86996 5048 86998
rect 5104 86996 5152 86998
rect 4008 86986 5208 86996
rect 6076 86884 6132 87390
rect 6076 86818 6132 86828
rect 6524 87444 6580 87454
rect 1708 86436 1764 86446
rect 1708 86342 1764 86380
rect 1708 85986 1764 85998
rect 1708 85934 1710 85986
rect 1762 85934 1764 85986
rect 1708 85204 1764 85934
rect 4008 85484 5208 85494
rect 4064 85482 4112 85484
rect 4168 85482 4216 85484
rect 4076 85430 4112 85482
rect 4200 85430 4216 85482
rect 4064 85428 4112 85430
rect 4168 85428 4216 85430
rect 4272 85482 4320 85484
rect 4376 85482 4424 85484
rect 4480 85482 4528 85484
rect 4376 85430 4396 85482
rect 4480 85430 4520 85482
rect 4272 85428 4320 85430
rect 4376 85428 4424 85430
rect 4480 85428 4528 85430
rect 4584 85428 4632 85484
rect 4688 85482 4736 85484
rect 4792 85482 4840 85484
rect 4896 85482 4944 85484
rect 4696 85430 4736 85482
rect 4820 85430 4840 85482
rect 4688 85428 4736 85430
rect 4792 85428 4840 85430
rect 4896 85428 4944 85430
rect 5000 85482 5048 85484
rect 5104 85482 5152 85484
rect 5000 85430 5016 85482
rect 5104 85430 5140 85482
rect 5000 85428 5048 85430
rect 5104 85428 5152 85430
rect 4008 85418 5208 85428
rect 1708 85138 1764 85148
rect 4844 85204 4900 85214
rect 4844 85110 4900 85148
rect 5404 85204 5460 85214
rect 3836 85092 3892 85102
rect 1708 84418 1764 84430
rect 1708 84366 1710 84418
rect 1762 84366 1764 84418
rect 1708 84084 1764 84366
rect 3836 84306 3892 85036
rect 3836 84254 3838 84306
rect 3890 84254 3892 84306
rect 3836 84242 3892 84254
rect 4172 84306 4228 84318
rect 4172 84254 4174 84306
rect 4226 84254 4228 84306
rect 4172 84084 4228 84254
rect 1708 84018 1764 84028
rect 3836 84028 4228 84084
rect 3836 83748 3892 84028
rect 4008 83916 5208 83926
rect 4064 83914 4112 83916
rect 4168 83914 4216 83916
rect 4076 83862 4112 83914
rect 4200 83862 4216 83914
rect 4064 83860 4112 83862
rect 4168 83860 4216 83862
rect 4272 83914 4320 83916
rect 4376 83914 4424 83916
rect 4480 83914 4528 83916
rect 4376 83862 4396 83914
rect 4480 83862 4520 83914
rect 4272 83860 4320 83862
rect 4376 83860 4424 83862
rect 4480 83860 4528 83862
rect 4584 83860 4632 83916
rect 4688 83914 4736 83916
rect 4792 83914 4840 83916
rect 4896 83914 4944 83916
rect 4696 83862 4736 83914
rect 4820 83862 4840 83914
rect 4688 83860 4736 83862
rect 4792 83860 4840 83862
rect 4896 83860 4944 83862
rect 5000 83914 5048 83916
rect 5104 83914 5152 83916
rect 5000 83862 5016 83914
rect 5104 83862 5140 83914
rect 5000 83860 5048 83862
rect 5104 83860 5152 83862
rect 4008 83850 5208 83860
rect 3836 83682 3892 83692
rect 3724 83524 3780 83534
rect 4284 83524 4340 83534
rect 3612 83522 3780 83524
rect 3612 83470 3726 83522
rect 3778 83470 3780 83522
rect 3612 83468 3780 83470
rect 1708 83298 1764 83310
rect 1708 83246 1710 83298
rect 1762 83246 1764 83298
rect 1708 82964 1764 83246
rect 1708 82898 1764 82908
rect 2268 83300 2324 83310
rect 1820 82738 1876 82750
rect 1820 82686 1822 82738
rect 1874 82686 1876 82738
rect 1708 81844 1764 81854
rect 1708 81750 1764 81788
rect 1708 81282 1764 81294
rect 1708 81230 1710 81282
rect 1762 81230 1764 81282
rect 1708 80724 1764 81230
rect 1708 80658 1764 80668
rect 1820 80612 1876 82686
rect 2268 82738 2324 83244
rect 3388 83300 3444 83310
rect 3388 83206 3444 83244
rect 2268 82686 2270 82738
rect 2322 82686 2324 82738
rect 2268 82674 2324 82686
rect 3612 82068 3668 83468
rect 3724 83458 3780 83468
rect 3836 83468 4284 83524
rect 3612 82002 3668 82012
rect 1708 80162 1764 80174
rect 1708 80110 1710 80162
rect 1762 80110 1764 80162
rect 1708 79604 1764 80110
rect 1708 79538 1764 79548
rect 1820 79602 1876 80556
rect 1820 79550 1822 79602
rect 1874 79550 1876 79602
rect 1708 78596 1764 78606
rect 1708 78502 1764 78540
rect 1820 78034 1876 79550
rect 2268 79604 2324 79614
rect 2268 79602 3332 79604
rect 2268 79550 2270 79602
rect 2322 79550 3332 79602
rect 2268 79548 3332 79550
rect 2268 79538 2324 79548
rect 3276 79042 3332 79548
rect 3276 78990 3278 79042
rect 3330 78990 3332 79042
rect 3276 78978 3332 78990
rect 3388 78932 3444 78942
rect 3388 78838 3444 78876
rect 1820 77982 1822 78034
rect 1874 77982 1876 78034
rect 1820 77970 1876 77982
rect 2268 78036 2324 78046
rect 2268 78034 3332 78036
rect 2268 77982 2270 78034
rect 2322 77982 3332 78034
rect 2268 77980 3332 77982
rect 2268 77970 2324 77980
rect 3276 77474 3332 77980
rect 3276 77422 3278 77474
rect 3330 77422 3332 77474
rect 3276 77410 3332 77422
rect 3612 77812 3668 77822
rect 3612 77474 3668 77756
rect 3612 77422 3614 77474
rect 3666 77422 3668 77474
rect 3612 77410 3668 77422
rect 1708 77364 1764 77374
rect 1708 77138 1764 77308
rect 1708 77086 1710 77138
rect 1762 77086 1764 77138
rect 1708 77074 1764 77086
rect 3836 77138 3892 83468
rect 4284 83430 4340 83468
rect 5404 83524 5460 85148
rect 6524 85092 6580 87388
rect 8876 87444 8932 87948
rect 9884 87668 9940 87678
rect 9884 87574 9940 87612
rect 8876 87378 8932 87388
rect 9100 87442 9156 87454
rect 9100 87390 9102 87442
rect 9154 87390 9156 87442
rect 7644 86884 7700 86894
rect 7644 86790 7700 86828
rect 7980 86658 8036 86670
rect 7980 86606 7982 86658
rect 8034 86606 8036 86658
rect 7308 86548 7364 86558
rect 7308 86454 7364 86492
rect 7980 86436 8036 86606
rect 8764 86660 8820 86670
rect 7980 86370 8036 86380
rect 8540 86548 8596 86558
rect 8540 86212 8596 86492
rect 8540 86146 8596 86156
rect 7420 85762 7476 85774
rect 7420 85710 7422 85762
rect 7474 85710 7476 85762
rect 7420 85708 7476 85710
rect 8764 85708 8820 86604
rect 9100 86436 9156 87390
rect 9996 86770 10052 88958
rect 12348 88900 12404 89070
rect 10332 88228 10388 88238
rect 10332 87666 10388 88172
rect 10332 87614 10334 87666
rect 10386 87614 10388 87666
rect 10332 87602 10388 87614
rect 10444 88004 10500 88014
rect 9996 86718 9998 86770
rect 10050 86718 10052 86770
rect 9996 86706 10052 86718
rect 9324 86660 9380 86670
rect 9324 86566 9380 86604
rect 9884 86660 9940 86670
rect 9100 86370 9156 86380
rect 9660 86100 9716 86110
rect 9660 86006 9716 86044
rect 9884 85988 9940 86604
rect 10332 86658 10388 86670
rect 10332 86606 10334 86658
rect 10386 86606 10388 86658
rect 10220 86548 10276 86558
rect 10220 86454 10276 86492
rect 10220 86100 10276 86110
rect 10220 86006 10276 86044
rect 9996 85988 10052 85998
rect 9884 85986 10052 85988
rect 9884 85934 9998 85986
rect 10050 85934 10052 85986
rect 9884 85932 10052 85934
rect 9996 85922 10052 85932
rect 6524 84998 6580 85036
rect 6748 85652 7476 85708
rect 8428 85652 8820 85708
rect 10332 85762 10388 86606
rect 10332 85710 10334 85762
rect 10386 85710 10388 85762
rect 10332 85698 10388 85710
rect 6748 84980 6804 85652
rect 5852 84866 5908 84878
rect 5852 84814 5854 84866
rect 5906 84814 5908 84866
rect 5852 84084 5908 84814
rect 6748 84530 6804 84924
rect 6748 84478 6750 84530
rect 6802 84478 6804 84530
rect 6748 84466 6804 84478
rect 6972 85090 7028 85102
rect 6972 85038 6974 85090
rect 7026 85038 7028 85090
rect 6972 84532 7028 85038
rect 6972 84466 7028 84476
rect 7196 85092 7252 85102
rect 5852 84018 5908 84028
rect 6860 84084 6916 84094
rect 5964 83748 6020 83758
rect 5964 83654 6020 83692
rect 6300 83748 6356 83758
rect 6300 83654 6356 83692
rect 5404 83458 5460 83468
rect 5628 83636 5684 83646
rect 4508 83412 4564 83422
rect 4508 83318 4564 83356
rect 5292 83412 5348 83422
rect 5068 83298 5124 83310
rect 5068 83246 5070 83298
rect 5122 83246 5124 83298
rect 4732 82962 4788 82974
rect 4732 82910 4734 82962
rect 4786 82910 4788 82962
rect 4732 82852 4788 82910
rect 4732 82786 4788 82796
rect 5068 82852 5124 83246
rect 5292 82964 5348 83356
rect 5628 82964 5684 83580
rect 6860 83410 6916 84028
rect 6860 83358 6862 83410
rect 6914 83358 6916 83410
rect 6860 83346 6916 83358
rect 7084 83522 7140 83534
rect 7084 83470 7086 83522
rect 7138 83470 7140 83522
rect 7084 83300 7140 83470
rect 7084 83234 7140 83244
rect 6188 82964 6244 82974
rect 5292 82962 5572 82964
rect 5292 82910 5294 82962
rect 5346 82910 5572 82962
rect 5292 82908 5572 82910
rect 5292 82898 5348 82908
rect 5068 82786 5124 82796
rect 5516 82850 5572 82908
rect 5628 82962 5796 82964
rect 5628 82910 5630 82962
rect 5682 82910 5796 82962
rect 5628 82908 5796 82910
rect 5628 82898 5684 82908
rect 5516 82798 5518 82850
rect 5570 82798 5572 82850
rect 5516 82786 5572 82798
rect 5628 82516 5684 82526
rect 5516 82514 5684 82516
rect 5516 82462 5630 82514
rect 5682 82462 5684 82514
rect 5516 82460 5684 82462
rect 5740 82516 5796 82908
rect 6188 82962 6468 82964
rect 6188 82910 6190 82962
rect 6242 82910 6468 82962
rect 6188 82908 6468 82910
rect 6188 82898 6244 82908
rect 6300 82738 6356 82750
rect 6300 82686 6302 82738
rect 6354 82686 6356 82738
rect 6300 82628 6356 82686
rect 6300 82562 6356 82572
rect 5740 82460 6020 82516
rect 4008 82348 5208 82358
rect 4064 82346 4112 82348
rect 4168 82346 4216 82348
rect 4076 82294 4112 82346
rect 4200 82294 4216 82346
rect 4064 82292 4112 82294
rect 4168 82292 4216 82294
rect 4272 82346 4320 82348
rect 4376 82346 4424 82348
rect 4480 82346 4528 82348
rect 4376 82294 4396 82346
rect 4480 82294 4520 82346
rect 4272 82292 4320 82294
rect 4376 82292 4424 82294
rect 4480 82292 4528 82294
rect 4584 82292 4632 82348
rect 4688 82346 4736 82348
rect 4792 82346 4840 82348
rect 4896 82346 4944 82348
rect 4696 82294 4736 82346
rect 4820 82294 4840 82346
rect 4688 82292 4736 82294
rect 4792 82292 4840 82294
rect 4896 82292 4944 82294
rect 5000 82346 5048 82348
rect 5104 82346 5152 82348
rect 5000 82294 5016 82346
rect 5104 82294 5140 82346
rect 5000 82292 5048 82294
rect 5104 82292 5152 82294
rect 4008 82282 5208 82292
rect 4844 82180 4900 82190
rect 4508 82068 4564 82078
rect 4508 81974 4564 82012
rect 4844 81842 4900 82124
rect 4844 81790 4846 81842
rect 4898 81790 4900 81842
rect 4844 81778 4900 81790
rect 4396 81732 4452 81742
rect 4396 81638 4452 81676
rect 4620 81730 4676 81742
rect 4620 81678 4622 81730
rect 4674 81678 4676 81730
rect 4620 81060 4676 81678
rect 4620 80994 4676 81004
rect 5180 81732 5236 81742
rect 5180 81060 5236 81676
rect 5180 81058 5348 81060
rect 5180 81006 5182 81058
rect 5234 81006 5348 81058
rect 5180 81004 5348 81006
rect 5180 80994 5236 81004
rect 4008 80780 5208 80790
rect 4064 80778 4112 80780
rect 4168 80778 4216 80780
rect 4076 80726 4112 80778
rect 4200 80726 4216 80778
rect 4064 80724 4112 80726
rect 4168 80724 4216 80726
rect 4272 80778 4320 80780
rect 4376 80778 4424 80780
rect 4480 80778 4528 80780
rect 4376 80726 4396 80778
rect 4480 80726 4520 80778
rect 4272 80724 4320 80726
rect 4376 80724 4424 80726
rect 4480 80724 4528 80726
rect 4584 80724 4632 80780
rect 4688 80778 4736 80780
rect 4792 80778 4840 80780
rect 4896 80778 4944 80780
rect 4696 80726 4736 80778
rect 4820 80726 4840 80778
rect 4688 80724 4736 80726
rect 4792 80724 4840 80726
rect 4896 80724 4944 80726
rect 5000 80778 5048 80780
rect 5104 80778 5152 80780
rect 5000 80726 5016 80778
rect 5104 80726 5140 80778
rect 5000 80724 5048 80726
rect 5104 80724 5152 80726
rect 4008 80714 5208 80724
rect 4732 79828 4788 79838
rect 4732 79734 4788 79772
rect 4008 79212 5208 79222
rect 4064 79210 4112 79212
rect 4168 79210 4216 79212
rect 4076 79158 4112 79210
rect 4200 79158 4216 79210
rect 4064 79156 4112 79158
rect 4168 79156 4216 79158
rect 4272 79210 4320 79212
rect 4376 79210 4424 79212
rect 4480 79210 4528 79212
rect 4376 79158 4396 79210
rect 4480 79158 4520 79210
rect 4272 79156 4320 79158
rect 4376 79156 4424 79158
rect 4480 79156 4528 79158
rect 4584 79156 4632 79212
rect 4688 79210 4736 79212
rect 4792 79210 4840 79212
rect 4896 79210 4944 79212
rect 4696 79158 4736 79210
rect 4820 79158 4840 79210
rect 4688 79156 4736 79158
rect 4792 79156 4840 79158
rect 4896 79156 4944 79158
rect 5000 79210 5048 79212
rect 5104 79210 5152 79212
rect 5000 79158 5016 79210
rect 5104 79158 5140 79210
rect 5000 79156 5048 79158
rect 5104 79156 5152 79158
rect 4008 79146 5208 79156
rect 4508 78932 4564 78942
rect 5292 78932 5348 81004
rect 5516 80948 5572 82460
rect 5628 82450 5684 82460
rect 5852 82292 5908 82302
rect 5516 80882 5572 80892
rect 5628 82236 5852 82292
rect 5628 81170 5684 82236
rect 5852 82226 5908 82236
rect 5964 82068 6020 82460
rect 6188 82514 6244 82526
rect 6188 82462 6190 82514
rect 6242 82462 6244 82514
rect 6188 82404 6244 82462
rect 6188 82338 6244 82348
rect 6412 82516 6468 82908
rect 5628 81118 5630 81170
rect 5682 81118 5684 81170
rect 5628 80612 5684 81118
rect 5628 80546 5684 80556
rect 5852 82066 6020 82068
rect 5852 82014 5966 82066
rect 6018 82014 6020 82066
rect 5852 82012 6020 82014
rect 5852 80388 5908 82012
rect 5964 82002 6020 82012
rect 6300 82292 6356 82302
rect 6076 81170 6132 81182
rect 6076 81118 6078 81170
rect 6130 81118 6132 81170
rect 5964 80948 6020 80958
rect 5964 80610 6020 80892
rect 5964 80558 5966 80610
rect 6018 80558 6020 80610
rect 5964 80546 6020 80558
rect 6076 80610 6132 81118
rect 6076 80558 6078 80610
rect 6130 80558 6132 80610
rect 6076 80546 6132 80558
rect 6076 80388 6132 80398
rect 5852 80332 6076 80388
rect 5852 79826 5908 80332
rect 6076 80294 6132 80332
rect 5852 79774 5854 79826
rect 5906 79774 5908 79826
rect 5404 79602 5460 79614
rect 5404 79550 5406 79602
rect 5458 79550 5460 79602
rect 5404 79380 5460 79550
rect 5404 79314 5460 79324
rect 5404 78932 5460 78942
rect 5292 78876 5404 78932
rect 4508 78838 4564 78876
rect 5404 78866 5460 78876
rect 4620 78820 4676 78830
rect 5852 78820 5908 79774
rect 6300 79826 6356 82236
rect 6412 82066 6468 82460
rect 6412 82014 6414 82066
rect 6466 82014 6468 82066
rect 6412 82002 6468 82014
rect 6636 82628 6692 82638
rect 6748 82628 6804 82638
rect 6692 82626 6804 82628
rect 6692 82574 6750 82626
rect 6802 82574 6804 82626
rect 6692 82572 6804 82574
rect 6636 81732 6692 82572
rect 6748 82562 6804 82572
rect 7196 82628 7252 85036
rect 8316 84532 8372 84542
rect 8316 84438 8372 84476
rect 8092 84306 8148 84318
rect 8092 84254 8094 84306
rect 8146 84254 8148 84306
rect 7868 84196 7924 84206
rect 8092 84196 8148 84254
rect 7868 84194 8148 84196
rect 7868 84142 7870 84194
rect 7922 84142 8148 84194
rect 7868 84140 8148 84142
rect 7308 84082 7364 84094
rect 7308 84030 7310 84082
rect 7362 84030 7364 84082
rect 7308 83748 7364 84030
rect 7308 83682 7364 83692
rect 7644 83300 7700 83310
rect 7868 83300 7924 84140
rect 8204 83412 8260 83422
rect 8204 83318 8260 83356
rect 8428 83410 8484 85652
rect 10444 85092 10500 87948
rect 12012 88004 12068 88014
rect 12348 88004 12404 88844
rect 12068 87948 12404 88004
rect 12572 88004 12628 88014
rect 12012 87910 12068 87948
rect 11452 87668 11508 87678
rect 10892 87554 10948 87566
rect 10892 87502 10894 87554
rect 10946 87502 10948 87554
rect 10668 87220 10724 87230
rect 10668 87126 10724 87164
rect 10892 86660 10948 87502
rect 11452 87554 11508 87612
rect 11452 87502 11454 87554
rect 11506 87502 11508 87554
rect 11452 87490 11508 87502
rect 12124 87444 12180 87454
rect 12124 87442 12404 87444
rect 12124 87390 12126 87442
rect 12178 87390 12404 87442
rect 12124 87388 12404 87390
rect 12124 87378 12180 87388
rect 12236 86884 12292 86894
rect 12012 86882 12292 86884
rect 12012 86830 12238 86882
rect 12290 86830 12292 86882
rect 12012 86828 12292 86830
rect 12012 86770 12068 86828
rect 12236 86818 12292 86828
rect 12012 86718 12014 86770
rect 12066 86718 12068 86770
rect 12012 86706 12068 86718
rect 10780 86100 10836 86110
rect 10892 86100 10948 86604
rect 10780 86098 10948 86100
rect 10780 86046 10782 86098
rect 10834 86046 10948 86098
rect 10780 86044 10948 86046
rect 11004 86548 11060 86558
rect 10780 86034 10836 86044
rect 10780 85092 10836 85102
rect 10444 85090 10836 85092
rect 10444 85038 10782 85090
rect 10834 85038 10836 85090
rect 10444 85036 10836 85038
rect 9212 84980 9268 84990
rect 9212 84886 9268 84924
rect 10444 84980 10500 85036
rect 10780 85026 10836 85036
rect 10444 84914 10500 84924
rect 9996 84868 10052 84878
rect 9772 84866 10052 84868
rect 9772 84814 9998 84866
rect 10050 84814 10052 84866
rect 9772 84812 10052 84814
rect 9660 84532 9716 84542
rect 8652 84530 9716 84532
rect 8652 84478 9662 84530
rect 9714 84478 9716 84530
rect 8652 84476 9716 84478
rect 8540 84420 8596 84430
rect 8652 84420 8708 84476
rect 8540 84418 8708 84420
rect 8540 84366 8542 84418
rect 8594 84366 8708 84418
rect 8540 84364 8708 84366
rect 8540 84354 8596 84364
rect 8764 84306 8820 84318
rect 8764 84254 8766 84306
rect 8818 84254 8820 84306
rect 8764 83746 8820 84254
rect 8764 83694 8766 83746
rect 8818 83694 8820 83746
rect 8764 83682 8820 83694
rect 8428 83358 8430 83410
rect 8482 83358 8484 83410
rect 7700 83244 7924 83300
rect 8428 83300 8484 83358
rect 7644 83206 7700 83244
rect 8428 83234 8484 83244
rect 8764 83522 8820 83534
rect 8764 83470 8766 83522
rect 8818 83470 8820 83522
rect 8764 83412 8820 83470
rect 8204 82852 8260 82862
rect 7644 82628 7700 82638
rect 7196 82626 7700 82628
rect 7196 82574 7198 82626
rect 7250 82574 7646 82626
rect 7698 82574 7700 82626
rect 7196 82572 7700 82574
rect 7196 82562 7252 82572
rect 7644 82404 7700 82572
rect 7644 82338 7700 82348
rect 6636 81666 6692 81676
rect 8204 81284 8260 82796
rect 8764 82516 8820 83356
rect 9212 83300 9268 83310
rect 9268 83244 9380 83300
rect 9212 83206 9268 83244
rect 8764 82450 8820 82460
rect 8316 81284 8372 81294
rect 8204 81282 8372 81284
rect 8204 81230 8318 81282
rect 8370 81230 8372 81282
rect 8204 81228 8372 81230
rect 6748 80612 6804 80622
rect 6972 80612 7028 80622
rect 6748 80610 7028 80612
rect 6748 80558 6750 80610
rect 6802 80558 6974 80610
rect 7026 80558 7028 80610
rect 6748 80556 7028 80558
rect 6748 80546 6804 80556
rect 6972 80546 7028 80556
rect 7756 80612 7812 80622
rect 7980 80612 8036 80622
rect 7756 80610 8036 80612
rect 7756 80558 7758 80610
rect 7810 80558 7982 80610
rect 8034 80558 8036 80610
rect 7756 80556 8036 80558
rect 7756 80546 7812 80556
rect 7980 80546 8036 80556
rect 6300 79774 6302 79826
rect 6354 79774 6356 79826
rect 4620 78726 4676 78764
rect 5740 78764 5852 78820
rect 5068 78708 5124 78718
rect 5628 78708 5684 78718
rect 5068 78706 5684 78708
rect 5068 78654 5070 78706
rect 5122 78654 5630 78706
rect 5682 78654 5684 78706
rect 5068 78652 5684 78654
rect 5068 78642 5124 78652
rect 5628 78642 5684 78652
rect 4172 78596 4228 78606
rect 4172 78502 4228 78540
rect 4508 78594 4564 78606
rect 4508 78542 4510 78594
rect 4562 78542 4564 78594
rect 4508 78372 4564 78542
rect 4508 78306 4564 78316
rect 4844 78594 4900 78606
rect 4844 78542 4846 78594
rect 4898 78542 4900 78594
rect 4732 78260 4788 78270
rect 4732 78166 4788 78204
rect 4844 77924 4900 78542
rect 4844 77858 4900 77868
rect 5292 78372 5348 78382
rect 5292 78258 5348 78316
rect 5292 78206 5294 78258
rect 5346 78206 5348 78258
rect 4008 77644 5208 77654
rect 4064 77642 4112 77644
rect 4168 77642 4216 77644
rect 4076 77590 4112 77642
rect 4200 77590 4216 77642
rect 4064 77588 4112 77590
rect 4168 77588 4216 77590
rect 4272 77642 4320 77644
rect 4376 77642 4424 77644
rect 4480 77642 4528 77644
rect 4376 77590 4396 77642
rect 4480 77590 4520 77642
rect 4272 77588 4320 77590
rect 4376 77588 4424 77590
rect 4480 77588 4528 77590
rect 4584 77588 4632 77644
rect 4688 77642 4736 77644
rect 4792 77642 4840 77644
rect 4896 77642 4944 77644
rect 4696 77590 4736 77642
rect 4820 77590 4840 77642
rect 4688 77588 4736 77590
rect 4792 77588 4840 77590
rect 4896 77588 4944 77590
rect 5000 77642 5048 77644
rect 5104 77642 5152 77644
rect 5000 77590 5016 77642
rect 5104 77590 5140 77642
rect 5000 77588 5048 77590
rect 5104 77588 5152 77590
rect 4008 77578 5208 77588
rect 3836 77086 3838 77138
rect 3890 77086 3892 77138
rect 3836 76692 3892 77086
rect 4284 77476 4340 77486
rect 4284 77138 4340 77420
rect 5292 77476 5348 78206
rect 5292 77410 5348 77420
rect 5404 78260 5460 78270
rect 5068 77252 5124 77262
rect 5068 77158 5124 77196
rect 4284 77086 4286 77138
rect 4338 77086 4340 77138
rect 4284 77074 4340 77086
rect 3836 76626 3892 76636
rect 4732 76692 4788 76702
rect 4732 76598 4788 76636
rect 5404 76690 5460 78204
rect 5628 77812 5684 77822
rect 5628 77718 5684 77756
rect 5404 76638 5406 76690
rect 5458 76638 5460 76690
rect 5404 76626 5460 76638
rect 5740 77250 5796 78764
rect 5852 78754 5908 78764
rect 6076 79380 6132 79390
rect 6076 78818 6132 79324
rect 6300 79044 6356 79774
rect 6300 78978 6356 78988
rect 6524 80386 6580 80398
rect 6524 80334 6526 80386
rect 6578 80334 6580 80386
rect 6524 79380 6580 80334
rect 7308 80388 7364 80398
rect 7308 80294 7364 80332
rect 6748 80276 6804 80286
rect 6748 79828 6804 80220
rect 8204 80276 8260 81228
rect 8316 81218 8372 81228
rect 9100 80946 9156 80958
rect 9100 80894 9102 80946
rect 9154 80894 9156 80946
rect 8204 80210 8260 80220
rect 8316 80276 8372 80286
rect 8652 80276 8708 80286
rect 8316 80274 8708 80276
rect 8316 80222 8318 80274
rect 8370 80222 8654 80274
rect 8706 80222 8708 80274
rect 8316 80220 8708 80222
rect 8316 80210 8372 80220
rect 8652 80210 8708 80220
rect 8764 80274 8820 80286
rect 8764 80222 8766 80274
rect 8818 80222 8820 80274
rect 6748 79734 6804 79772
rect 7420 80164 7476 80174
rect 7420 79714 7476 80108
rect 8092 80164 8148 80174
rect 8092 80070 8148 80108
rect 7420 79662 7422 79714
rect 7474 79662 7476 79714
rect 7420 79650 7476 79662
rect 7532 79716 7588 79726
rect 7532 79714 8260 79716
rect 7532 79662 7534 79714
rect 7586 79662 8260 79714
rect 7532 79660 8260 79662
rect 7532 79650 7588 79660
rect 8204 79604 8260 79660
rect 8316 79604 8372 79614
rect 8204 79602 8372 79604
rect 8204 79550 8318 79602
rect 8370 79550 8372 79602
rect 8204 79548 8372 79550
rect 6076 78766 6078 78818
rect 6130 78766 6132 78818
rect 5964 78596 6020 78606
rect 5740 77198 5742 77250
rect 5794 77198 5796 77250
rect 1708 76578 1764 76590
rect 1708 76526 1710 76578
rect 1762 76526 1764 76578
rect 1708 76244 1764 76526
rect 1708 76178 1764 76188
rect 5740 76356 5796 77198
rect 5852 78036 5908 78046
rect 5852 77140 5908 77980
rect 5964 78034 6020 78540
rect 5964 77982 5966 78034
rect 6018 77982 6020 78034
rect 5964 77364 6020 77982
rect 6076 77924 6132 78766
rect 6524 78930 6580 79324
rect 7980 79380 8036 79390
rect 7980 79286 8036 79324
rect 6748 79044 6804 79054
rect 7532 79044 7588 79054
rect 6804 78988 6916 79044
rect 6748 78978 6804 78988
rect 6524 78878 6526 78930
rect 6578 78878 6580 78930
rect 6076 77858 6132 77868
rect 6188 78596 6244 78606
rect 6188 78146 6244 78540
rect 6524 78260 6580 78878
rect 6524 78204 6692 78260
rect 6188 78094 6190 78146
rect 6242 78094 6244 78146
rect 5964 77298 6020 77308
rect 6076 77700 6132 77710
rect 5964 77140 6020 77150
rect 5852 77138 6020 77140
rect 5852 77086 5966 77138
rect 6018 77086 6020 77138
rect 5852 77084 6020 77086
rect 4008 76076 5208 76086
rect 4064 76074 4112 76076
rect 4168 76074 4216 76076
rect 4076 76022 4112 76074
rect 4200 76022 4216 76074
rect 4064 76020 4112 76022
rect 4168 76020 4216 76022
rect 4272 76074 4320 76076
rect 4376 76074 4424 76076
rect 4480 76074 4528 76076
rect 4376 76022 4396 76074
rect 4480 76022 4520 76074
rect 4272 76020 4320 76022
rect 4376 76020 4424 76022
rect 4480 76020 4528 76022
rect 4584 76020 4632 76076
rect 4688 76074 4736 76076
rect 4792 76074 4840 76076
rect 4896 76074 4944 76076
rect 4696 76022 4736 76074
rect 4820 76022 4840 76074
rect 4688 76020 4736 76022
rect 4792 76020 4840 76022
rect 4896 76020 4944 76022
rect 5000 76074 5048 76076
rect 5104 76074 5152 76076
rect 5000 76022 5016 76074
rect 5104 76022 5140 76074
rect 5000 76020 5048 76022
rect 5104 76020 5152 76022
rect 4008 76010 5208 76020
rect 4396 75796 4452 75806
rect 4396 75702 4452 75740
rect 5628 75684 5684 75694
rect 5292 75682 5684 75684
rect 5292 75630 5630 75682
rect 5682 75630 5684 75682
rect 5292 75628 5684 75630
rect 1708 75458 1764 75470
rect 4284 75460 4340 75470
rect 1708 75406 1710 75458
rect 1762 75406 1764 75458
rect 1708 75124 1764 75406
rect 1708 75058 1764 75068
rect 3612 75458 4340 75460
rect 3612 75406 4286 75458
rect 4338 75406 4340 75458
rect 3612 75404 4340 75406
rect 3164 74898 3220 74910
rect 3164 74846 3166 74898
rect 3218 74846 3220 74898
rect 1820 74228 1876 74238
rect 1708 73890 1764 73902
rect 1708 73838 1710 73890
rect 1762 73838 1764 73890
rect 1708 72884 1764 73838
rect 1820 73330 1876 74172
rect 3164 74228 3220 74846
rect 3612 74898 3668 75404
rect 4284 75394 4340 75404
rect 3612 74846 3614 74898
rect 3666 74846 3668 74898
rect 3612 74834 3668 74846
rect 4008 74508 5208 74518
rect 4064 74506 4112 74508
rect 4168 74506 4216 74508
rect 4076 74454 4112 74506
rect 4200 74454 4216 74506
rect 4064 74452 4112 74454
rect 4168 74452 4216 74454
rect 4272 74506 4320 74508
rect 4376 74506 4424 74508
rect 4480 74506 4528 74508
rect 4376 74454 4396 74506
rect 4480 74454 4520 74506
rect 4272 74452 4320 74454
rect 4376 74452 4424 74454
rect 4480 74452 4528 74454
rect 4584 74452 4632 74508
rect 4688 74506 4736 74508
rect 4792 74506 4840 74508
rect 4896 74506 4944 74508
rect 4696 74454 4736 74506
rect 4820 74454 4840 74506
rect 4688 74452 4736 74454
rect 4792 74452 4840 74454
rect 4896 74452 4944 74454
rect 5000 74506 5048 74508
rect 5104 74506 5152 74508
rect 5000 74454 5016 74506
rect 5104 74454 5140 74506
rect 5000 74452 5048 74454
rect 5104 74452 5152 74454
rect 4008 74442 5208 74452
rect 3164 74162 3220 74172
rect 4060 74340 4116 74350
rect 3836 74114 3892 74126
rect 3836 74062 3838 74114
rect 3890 74062 3892 74114
rect 2156 74004 2212 74014
rect 2492 74004 2548 74014
rect 2156 73890 2212 73948
rect 2156 73838 2158 73890
rect 2210 73838 2212 73890
rect 2156 73826 2212 73838
rect 2268 73948 2492 74004
rect 1820 73278 1822 73330
rect 1874 73278 1876 73330
rect 1820 73266 1876 73278
rect 2268 73330 2324 73948
rect 2492 73938 2548 73948
rect 3500 74004 3556 74042
rect 3500 73938 3556 73948
rect 2268 73278 2270 73330
rect 2322 73278 2324 73330
rect 2268 73266 2324 73278
rect 1708 72818 1764 72828
rect 3836 72770 3892 74062
rect 4060 74116 4116 74284
rect 4060 74002 4116 74060
rect 4060 73950 4062 74002
rect 4114 73950 4116 74002
rect 4060 73938 4116 73950
rect 4620 74004 4676 74042
rect 4620 73938 4676 73948
rect 5292 74004 5348 75628
rect 5628 75618 5684 75628
rect 5740 75572 5796 76300
rect 5852 75796 5908 75806
rect 5852 75702 5908 75740
rect 5852 75572 5908 75582
rect 5740 75570 5908 75572
rect 5740 75518 5854 75570
rect 5906 75518 5908 75570
rect 5740 75516 5908 75518
rect 5740 74228 5796 74238
rect 5740 73948 5796 74172
rect 4732 73892 4788 73902
rect 4732 73554 4788 73836
rect 4732 73502 4734 73554
rect 4786 73502 4788 73554
rect 4732 73490 4788 73502
rect 5292 73554 5348 73948
rect 5292 73502 5294 73554
rect 5346 73502 5348 73554
rect 5292 73490 5348 73502
rect 5628 73892 5796 73948
rect 5628 73330 5684 73892
rect 5628 73278 5630 73330
rect 5682 73278 5684 73330
rect 5628 73266 5684 73278
rect 4008 72940 5208 72950
rect 4064 72938 4112 72940
rect 4168 72938 4216 72940
rect 4076 72886 4112 72938
rect 4200 72886 4216 72938
rect 4064 72884 4112 72886
rect 4168 72884 4216 72886
rect 4272 72938 4320 72940
rect 4376 72938 4424 72940
rect 4480 72938 4528 72940
rect 4376 72886 4396 72938
rect 4480 72886 4520 72938
rect 4272 72884 4320 72886
rect 4376 72884 4424 72886
rect 4480 72884 4528 72886
rect 4584 72884 4632 72940
rect 4688 72938 4736 72940
rect 4792 72938 4840 72940
rect 4896 72938 4944 72940
rect 4696 72886 4736 72938
rect 4820 72886 4840 72938
rect 4688 72884 4736 72886
rect 4792 72884 4840 72886
rect 4896 72884 4944 72886
rect 5000 72938 5048 72940
rect 5104 72938 5152 72940
rect 5000 72886 5016 72938
rect 5104 72886 5140 72938
rect 5000 72884 5048 72886
rect 5104 72884 5152 72886
rect 4008 72874 5208 72884
rect 3836 72718 3838 72770
rect 3890 72718 3892 72770
rect 3836 72706 3892 72718
rect 4956 72772 5012 72782
rect 3164 72548 3220 72558
rect 1708 72322 1764 72334
rect 1708 72270 1710 72322
rect 1762 72270 1764 72322
rect 1708 71764 1764 72270
rect 1708 71698 1764 71708
rect 2828 70866 2884 70878
rect 2828 70814 2830 70866
rect 2882 70814 2884 70866
rect 1708 70756 1764 70766
rect 1708 70662 1764 70700
rect 2604 70756 2660 70766
rect 2828 70756 2884 70814
rect 3164 70866 3220 72492
rect 4172 72548 4228 72558
rect 4172 72454 4228 72492
rect 4732 72546 4788 72558
rect 4732 72494 4734 72546
rect 4786 72494 4788 72546
rect 4732 72436 4788 72494
rect 4732 72370 4788 72380
rect 4956 72434 5012 72716
rect 4956 72382 4958 72434
rect 5010 72382 5012 72434
rect 4956 72370 5012 72382
rect 5292 72436 5348 72446
rect 5292 71650 5348 72380
rect 5292 71598 5294 71650
rect 5346 71598 5348 71650
rect 4008 71372 5208 71382
rect 4064 71370 4112 71372
rect 4168 71370 4216 71372
rect 4076 71318 4112 71370
rect 4200 71318 4216 71370
rect 4064 71316 4112 71318
rect 4168 71316 4216 71318
rect 4272 71370 4320 71372
rect 4376 71370 4424 71372
rect 4480 71370 4528 71372
rect 4376 71318 4396 71370
rect 4480 71318 4520 71370
rect 4272 71316 4320 71318
rect 4376 71316 4424 71318
rect 4480 71316 4528 71318
rect 4584 71316 4632 71372
rect 4688 71370 4736 71372
rect 4792 71370 4840 71372
rect 4896 71370 4944 71372
rect 4696 71318 4736 71370
rect 4820 71318 4840 71370
rect 4688 71316 4736 71318
rect 4792 71316 4840 71318
rect 4896 71316 4944 71318
rect 5000 71370 5048 71372
rect 5104 71370 5152 71372
rect 5000 71318 5016 71370
rect 5104 71318 5140 71370
rect 5000 71316 5048 71318
rect 5104 71316 5152 71318
rect 4008 71306 5208 71316
rect 3164 70814 3166 70866
rect 3218 70814 3220 70866
rect 3164 70802 3220 70814
rect 2604 70754 2884 70756
rect 2604 70702 2606 70754
rect 2658 70702 2884 70754
rect 2604 70700 2884 70702
rect 1708 70306 1764 70318
rect 1708 70254 1710 70306
rect 1762 70254 1764 70306
rect 1708 69524 1764 70254
rect 1708 69458 1764 69468
rect 1708 68738 1764 68750
rect 1708 68686 1710 68738
rect 1762 68686 1764 68738
rect 1708 68404 1764 68686
rect 1708 68338 1764 68348
rect 1708 67618 1764 67630
rect 1708 67566 1710 67618
rect 1762 67566 1764 67618
rect 1708 67284 1764 67566
rect 2604 67228 2660 70700
rect 4008 69804 5208 69814
rect 4064 69802 4112 69804
rect 4168 69802 4216 69804
rect 4076 69750 4112 69802
rect 4200 69750 4216 69802
rect 4064 69748 4112 69750
rect 4168 69748 4216 69750
rect 4272 69802 4320 69804
rect 4376 69802 4424 69804
rect 4480 69802 4528 69804
rect 4376 69750 4396 69802
rect 4480 69750 4520 69802
rect 4272 69748 4320 69750
rect 4376 69748 4424 69750
rect 4480 69748 4528 69750
rect 4584 69748 4632 69804
rect 4688 69802 4736 69804
rect 4792 69802 4840 69804
rect 4896 69802 4944 69804
rect 4696 69750 4736 69802
rect 4820 69750 4840 69802
rect 4688 69748 4736 69750
rect 4792 69748 4840 69750
rect 4896 69748 4944 69750
rect 5000 69802 5048 69804
rect 5104 69802 5152 69804
rect 5000 69750 5016 69802
rect 5104 69750 5140 69802
rect 5000 69748 5048 69750
rect 5104 69748 5152 69750
rect 4008 69738 5208 69748
rect 5292 69188 5348 71598
rect 5740 69188 5796 69198
rect 5292 69186 5796 69188
rect 5292 69134 5742 69186
rect 5794 69134 5796 69186
rect 5292 69132 5796 69134
rect 3276 68626 3332 68638
rect 3724 68628 3780 68638
rect 3276 68574 3278 68626
rect 3330 68574 3332 68626
rect 1708 67218 1764 67228
rect 2044 67172 2660 67228
rect 3052 67844 3108 67854
rect 1708 66050 1764 66062
rect 1708 65998 1710 66050
rect 1762 65998 1764 66050
rect 1708 65044 1764 65998
rect 1820 65490 1876 65502
rect 1820 65438 1822 65490
rect 1874 65438 1876 65490
rect 1820 65268 1876 65438
rect 1932 65268 1988 65278
rect 1820 65212 1932 65268
rect 1708 64978 1764 64988
rect 1708 64482 1764 64494
rect 1708 64430 1710 64482
rect 1762 64430 1764 64482
rect 1708 63924 1764 64430
rect 1932 63924 1988 65212
rect 1708 63858 1764 63868
rect 1820 63922 1988 63924
rect 1820 63870 1934 63922
rect 1986 63870 1988 63922
rect 1820 63868 1988 63870
rect 1708 62916 1764 62926
rect 1708 62822 1764 62860
rect 1708 62466 1764 62478
rect 1708 62414 1710 62466
rect 1762 62414 1764 62466
rect 1708 61684 1764 62414
rect 1708 61618 1764 61628
rect 1708 61346 1764 61358
rect 1708 61294 1710 61346
rect 1762 61294 1764 61346
rect 1708 60564 1764 61294
rect 1820 60786 1876 63868
rect 1932 63858 1988 63868
rect 1820 60734 1822 60786
rect 1874 60734 1876 60786
rect 1820 60722 1876 60734
rect 1708 60498 1764 60508
rect 1708 59778 1764 59790
rect 1708 59726 1710 59778
rect 1762 59726 1764 59778
rect 1708 59444 1764 59726
rect 1708 59378 1764 59388
rect 2044 55468 2100 67172
rect 2268 66836 2324 66846
rect 2156 66164 2212 66174
rect 2156 66070 2212 66108
rect 2268 65490 2324 66780
rect 2268 65438 2270 65490
rect 2322 65438 2324 65490
rect 2268 65426 2324 65438
rect 2828 64594 2884 64606
rect 2828 64542 2830 64594
rect 2882 64542 2884 64594
rect 2604 64484 2660 64494
rect 2828 64484 2884 64542
rect 2604 64482 2884 64484
rect 2604 64430 2606 64482
rect 2658 64430 2884 64482
rect 2604 64428 2884 64430
rect 2380 63922 2436 63934
rect 2380 63870 2382 63922
rect 2434 63870 2436 63922
rect 2380 63364 2436 63870
rect 2380 63298 2436 63308
rect 2604 61572 2660 64428
rect 1820 55412 1876 55422
rect 1820 54514 1876 55356
rect 1820 54462 1822 54514
rect 1874 54462 1876 54514
rect 1820 51378 1876 54462
rect 1932 55412 2100 55468
rect 2156 61516 2660 61572
rect 1932 51604 1988 55412
rect 2044 52834 2100 52846
rect 2044 52782 2046 52834
rect 2098 52782 2100 52834
rect 2044 52724 2100 52782
rect 2044 52658 2100 52668
rect 1932 51538 1988 51548
rect 1820 51326 1822 51378
rect 1874 51326 1876 51378
rect 1820 51314 1876 51326
rect 2156 50484 2212 61516
rect 2268 61348 2324 61358
rect 2268 60786 2324 61292
rect 2268 60734 2270 60786
rect 2322 60734 2324 60786
rect 2268 60722 2324 60734
rect 2940 58434 2996 58446
rect 2940 58382 2942 58434
rect 2994 58382 2996 58434
rect 2492 58324 2548 58334
rect 2492 58230 2548 58268
rect 2940 58324 2996 58382
rect 2940 58258 2996 58268
rect 2828 57650 2884 57662
rect 2828 57598 2830 57650
rect 2882 57598 2884 57650
rect 2604 57540 2660 57550
rect 2828 57540 2884 57598
rect 2604 57538 2884 57540
rect 2604 57486 2606 57538
rect 2658 57486 2884 57538
rect 2604 57484 2884 57486
rect 2604 57204 2660 57484
rect 2604 57138 2660 57148
rect 2268 56644 2324 56654
rect 2268 54514 2324 56588
rect 2380 56084 2436 56094
rect 2380 55990 2436 56028
rect 2828 56084 2884 56094
rect 2828 55990 2884 56028
rect 3052 55468 3108 67788
rect 3276 65268 3332 68574
rect 3612 68626 3780 68628
rect 3612 68574 3726 68626
rect 3778 68574 3780 68626
rect 3612 68572 3780 68574
rect 3500 67618 3556 67630
rect 3500 67566 3502 67618
rect 3554 67566 3556 67618
rect 3500 66948 3556 67566
rect 3500 66882 3556 66892
rect 3388 66836 3444 66846
rect 3388 66742 3444 66780
rect 3612 66164 3668 68572
rect 3724 68562 3780 68572
rect 4008 68236 5208 68246
rect 4064 68234 4112 68236
rect 4168 68234 4216 68236
rect 4076 68182 4112 68234
rect 4200 68182 4216 68234
rect 4064 68180 4112 68182
rect 4168 68180 4216 68182
rect 4272 68234 4320 68236
rect 4376 68234 4424 68236
rect 4480 68234 4528 68236
rect 4376 68182 4396 68234
rect 4480 68182 4520 68234
rect 4272 68180 4320 68182
rect 4376 68180 4424 68182
rect 4480 68180 4528 68182
rect 4584 68180 4632 68236
rect 4688 68234 4736 68236
rect 4792 68234 4840 68236
rect 4896 68234 4944 68236
rect 4696 68182 4736 68234
rect 4820 68182 4840 68234
rect 4688 68180 4736 68182
rect 4792 68180 4840 68182
rect 4896 68180 4944 68182
rect 5000 68234 5048 68236
rect 5104 68234 5152 68236
rect 5000 68182 5016 68234
rect 5104 68182 5140 68234
rect 5000 68180 5048 68182
rect 5104 68180 5152 68182
rect 4008 68170 5208 68180
rect 4172 67844 4228 67854
rect 4172 67750 4228 67788
rect 4956 67844 5012 67854
rect 5404 67844 5460 69132
rect 5740 69122 5796 69132
rect 5852 68404 5908 75516
rect 5964 75348 6020 77084
rect 6076 77026 6132 77644
rect 6076 76974 6078 77026
rect 6130 76974 6132 77026
rect 6076 75682 6132 76974
rect 6076 75630 6078 75682
rect 6130 75630 6132 75682
rect 6076 75618 6132 75630
rect 6188 75460 6244 78094
rect 6524 77812 6580 77822
rect 6412 77756 6524 77812
rect 6300 77140 6356 77150
rect 6300 77046 6356 77084
rect 6300 75684 6356 75694
rect 6412 75684 6468 77756
rect 6524 77746 6580 77756
rect 6524 77252 6580 77262
rect 6524 76580 6580 77196
rect 6636 77250 6692 78204
rect 6636 77198 6638 77250
rect 6690 77198 6692 77250
rect 6636 77140 6692 77198
rect 6636 77074 6692 77084
rect 6748 78146 6804 78158
rect 6748 78094 6750 78146
rect 6802 78094 6804 78146
rect 6748 77924 6804 78094
rect 6748 77138 6804 77868
rect 6860 77252 6916 78988
rect 7532 78818 7588 78988
rect 7532 78766 7534 78818
rect 7586 78766 7588 78818
rect 7532 78754 7588 78766
rect 8204 78820 8260 78830
rect 8204 78726 8260 78764
rect 7084 78596 7140 78606
rect 8316 78596 8372 79548
rect 8652 79604 8708 79614
rect 8764 79604 8820 80222
rect 9100 80164 9156 80894
rect 9212 80276 9268 80286
rect 9212 80182 9268 80220
rect 9100 80098 9156 80108
rect 8652 79602 8820 79604
rect 8652 79550 8654 79602
rect 8706 79550 8820 79602
rect 8652 79548 8820 79550
rect 8652 79538 8708 79548
rect 8764 79492 8820 79548
rect 8764 79426 8820 79436
rect 7084 78502 7140 78540
rect 8204 78540 8372 78596
rect 7308 78148 7364 78158
rect 7308 78146 7476 78148
rect 7308 78094 7310 78146
rect 7362 78094 7476 78146
rect 7308 78092 7476 78094
rect 7308 78082 7364 78092
rect 7196 78036 7252 78046
rect 6860 77186 6916 77196
rect 6972 78034 7252 78036
rect 6972 77982 7198 78034
rect 7250 77982 7252 78034
rect 6972 77980 7252 77982
rect 6972 77250 7028 77980
rect 7196 77970 7252 77980
rect 7308 77812 7364 77822
rect 7420 77812 7476 78092
rect 7756 78036 7812 78046
rect 7756 77942 7812 77980
rect 7868 77812 7924 77822
rect 7420 77810 8036 77812
rect 7420 77758 7870 77810
rect 7922 77758 8036 77810
rect 7420 77756 8036 77758
rect 7308 77718 7364 77756
rect 7868 77746 7924 77756
rect 6972 77198 6974 77250
rect 7026 77198 7028 77250
rect 6972 77186 7028 77198
rect 7420 77364 7476 77374
rect 6748 77086 6750 77138
rect 6802 77086 6804 77138
rect 6748 77074 6804 77086
rect 7420 77028 7476 77308
rect 7980 77138 8036 77756
rect 8204 77700 8260 78540
rect 8876 78146 8932 78158
rect 8876 78094 8878 78146
rect 8930 78094 8932 78146
rect 8652 78036 8708 78046
rect 8316 77924 8372 77934
rect 8316 77922 8484 77924
rect 8316 77870 8318 77922
rect 8370 77870 8484 77922
rect 8316 77868 8484 77870
rect 8316 77858 8372 77868
rect 8428 77812 8484 77868
rect 8652 77812 8708 77980
rect 8428 77810 8708 77812
rect 8428 77758 8654 77810
rect 8706 77758 8708 77810
rect 8428 77756 8708 77758
rect 8316 77700 8372 77710
rect 8204 77644 8316 77700
rect 8316 77634 8372 77644
rect 7980 77086 7982 77138
rect 8034 77086 8036 77138
rect 7980 77074 8036 77086
rect 7532 77028 7588 77038
rect 7420 77026 7588 77028
rect 7420 76974 7534 77026
rect 7586 76974 7588 77026
rect 7420 76972 7588 76974
rect 7532 76962 7588 76972
rect 8428 77026 8484 77038
rect 8428 76974 8430 77026
rect 8482 76974 8484 77026
rect 6524 76524 6692 76580
rect 6524 76356 6580 76366
rect 6524 76262 6580 76300
rect 6300 75682 6468 75684
rect 6300 75630 6302 75682
rect 6354 75630 6468 75682
rect 6300 75628 6468 75630
rect 6300 75618 6356 75628
rect 6636 75572 6692 76524
rect 6748 76356 6804 76366
rect 6748 75794 6804 76300
rect 6748 75742 6750 75794
rect 6802 75742 6804 75794
rect 6748 75730 6804 75742
rect 6636 75516 7028 75572
rect 6188 75404 6356 75460
rect 6076 75348 6132 75358
rect 5964 75292 6076 75348
rect 6076 75282 6132 75292
rect 6076 75124 6132 75134
rect 6076 75122 6244 75124
rect 6076 75070 6078 75122
rect 6130 75070 6244 75122
rect 6076 75068 6244 75070
rect 6076 75058 6132 75068
rect 6188 74676 6244 75068
rect 6188 74226 6244 74620
rect 6188 74174 6190 74226
rect 6242 74174 6244 74226
rect 6188 74116 6244 74174
rect 6188 74050 6244 74060
rect 6300 73948 6356 75404
rect 6636 75348 6692 75358
rect 6636 74676 6692 75292
rect 6972 75122 7028 75516
rect 6972 75070 6974 75122
rect 7026 75070 7028 75122
rect 6636 74674 6804 74676
rect 6636 74622 6638 74674
rect 6690 74622 6804 74674
rect 6636 74620 6804 74622
rect 6636 74610 6692 74620
rect 6636 74340 6692 74350
rect 6636 74228 6692 74284
rect 6524 74226 6692 74228
rect 6524 74174 6638 74226
rect 6690 74174 6692 74226
rect 6524 74172 6692 74174
rect 6300 73892 6468 73948
rect 6076 73332 6132 73342
rect 6076 73238 6132 73276
rect 5964 72548 6020 72558
rect 5964 72454 6020 72492
rect 6076 72548 6132 72558
rect 6300 72548 6356 72558
rect 6076 72546 6300 72548
rect 6076 72494 6078 72546
rect 6130 72494 6300 72546
rect 6076 72492 6300 72494
rect 6076 72482 6132 72492
rect 6300 72482 6356 72492
rect 6412 72436 6468 73892
rect 6412 72370 6468 72380
rect 6188 70084 6244 70094
rect 6188 69188 6244 70028
rect 4956 67842 5460 67844
rect 4956 67790 4958 67842
rect 5010 67790 5460 67842
rect 4956 67788 5460 67790
rect 5516 68348 5908 68404
rect 6076 69186 6244 69188
rect 6076 69134 6190 69186
rect 6242 69134 6244 69186
rect 6076 69132 6244 69134
rect 4732 67730 4788 67742
rect 4732 67678 4734 67730
rect 4786 67678 4788 67730
rect 3836 67620 3892 67630
rect 3724 67618 3892 67620
rect 3724 67566 3838 67618
rect 3890 67566 3892 67618
rect 3724 67564 3892 67566
rect 3724 67058 3780 67564
rect 3836 67554 3892 67564
rect 3948 67172 4004 67182
rect 3724 67006 3726 67058
rect 3778 67006 3780 67058
rect 3724 66994 3780 67006
rect 3836 67170 4004 67172
rect 3836 67118 3950 67170
rect 4002 67118 4004 67170
rect 3836 67116 4004 67118
rect 3612 66098 3668 66108
rect 3836 66052 3892 67116
rect 3948 67106 4004 67116
rect 4508 67172 4564 67182
rect 4508 67078 4564 67116
rect 4732 66948 4788 67678
rect 4956 67284 5012 67788
rect 4956 67218 5012 67228
rect 5292 67620 5348 67630
rect 4732 66882 4788 66892
rect 4008 66668 5208 66678
rect 4064 66666 4112 66668
rect 4168 66666 4216 66668
rect 4076 66614 4112 66666
rect 4200 66614 4216 66666
rect 4064 66612 4112 66614
rect 4168 66612 4216 66614
rect 4272 66666 4320 66668
rect 4376 66666 4424 66668
rect 4480 66666 4528 66668
rect 4376 66614 4396 66666
rect 4480 66614 4520 66666
rect 4272 66612 4320 66614
rect 4376 66612 4424 66614
rect 4480 66612 4528 66614
rect 4584 66612 4632 66668
rect 4688 66666 4736 66668
rect 4792 66666 4840 66668
rect 4896 66666 4944 66668
rect 4696 66614 4736 66666
rect 4820 66614 4840 66666
rect 4688 66612 4736 66614
rect 4792 66612 4840 66614
rect 4896 66612 4944 66614
rect 5000 66666 5048 66668
rect 5104 66666 5152 66668
rect 5000 66614 5016 66666
rect 5104 66614 5140 66666
rect 5000 66612 5048 66614
rect 5104 66612 5152 66614
rect 4008 66602 5208 66612
rect 5292 66500 5348 67564
rect 5516 67284 5572 68348
rect 5852 68068 5908 68078
rect 5852 67730 5908 68012
rect 5852 67678 5854 67730
rect 5906 67678 5908 67730
rect 5852 67666 5908 67678
rect 5964 67732 6020 67742
rect 6076 67732 6132 69132
rect 6188 69122 6244 69132
rect 5964 67730 6132 67732
rect 5964 67678 5966 67730
rect 6018 67678 6132 67730
rect 5964 67676 6132 67678
rect 6188 68850 6244 68862
rect 6188 68798 6190 68850
rect 6242 68798 6244 68850
rect 5628 67620 5684 67630
rect 5628 67526 5684 67564
rect 5516 67228 5684 67284
rect 5404 67172 5460 67182
rect 5460 67116 5572 67172
rect 5404 67106 5460 67116
rect 5404 66948 5460 66958
rect 5404 66854 5460 66892
rect 4956 66444 5348 66500
rect 4956 66274 5012 66444
rect 5516 66388 5572 67116
rect 4956 66222 4958 66274
rect 5010 66222 5012 66274
rect 4956 66210 5012 66222
rect 5292 66332 5572 66388
rect 4508 66164 4564 66174
rect 4508 66070 4564 66108
rect 4060 66052 4116 66062
rect 3836 66050 4116 66052
rect 3836 65998 4062 66050
rect 4114 65998 4116 66050
rect 3836 65996 4116 65998
rect 4060 65604 4116 65996
rect 4396 66052 4452 66062
rect 4396 65958 4452 65996
rect 4620 66050 4676 66062
rect 4620 65998 4622 66050
rect 4674 65998 4676 66050
rect 4060 65538 4116 65548
rect 4620 65268 4676 65998
rect 4732 65716 4788 65726
rect 4732 65622 4788 65660
rect 5292 65490 5348 66332
rect 5628 65716 5684 67228
rect 5964 67060 6020 67676
rect 5740 67004 6020 67060
rect 6076 67508 6132 67518
rect 6188 67508 6244 68798
rect 6132 67452 6244 67508
rect 6300 67730 6356 67742
rect 6300 67678 6302 67730
rect 6354 67678 6356 67730
rect 6076 67282 6132 67452
rect 6076 67230 6078 67282
rect 6130 67230 6132 67282
rect 5740 66052 5796 67004
rect 6076 66948 6132 67230
rect 6300 67172 6356 67678
rect 6412 67620 6468 67658
rect 6412 67554 6468 67564
rect 6524 67396 6580 74172
rect 6636 74162 6692 74172
rect 6636 72772 6692 72782
rect 6748 72772 6804 74620
rect 6972 74228 7028 75070
rect 7980 74900 8036 74910
rect 7980 74806 8036 74844
rect 7420 74786 7476 74798
rect 7420 74734 7422 74786
rect 7474 74734 7476 74786
rect 7420 74676 7476 74734
rect 7420 74582 7476 74620
rect 8092 74676 8148 74686
rect 7028 74172 7252 74228
rect 6972 74162 7028 74172
rect 7196 74114 7252 74172
rect 7196 74062 7198 74114
rect 7250 74062 7252 74114
rect 7196 74050 7252 74062
rect 7868 74114 7924 74126
rect 7868 74062 7870 74114
rect 7922 74062 7924 74114
rect 7868 73556 7924 74062
rect 7868 73490 7924 73500
rect 6692 72716 6804 72772
rect 7756 73332 7812 73342
rect 6636 72706 6692 72716
rect 7756 72658 7812 73276
rect 7756 72606 7758 72658
rect 7810 72606 7812 72658
rect 7756 72594 7812 72606
rect 7868 72548 7924 72558
rect 7924 72492 8036 72548
rect 7868 72454 7924 72492
rect 7644 72324 7700 72334
rect 7644 72230 7700 72268
rect 6972 70756 7028 70766
rect 6972 69412 7028 70700
rect 7980 70418 8036 72492
rect 8092 72434 8148 74620
rect 8092 72382 8094 72434
rect 8146 72382 8148 72434
rect 8092 72370 8148 72382
rect 8316 74674 8372 74686
rect 8316 74622 8318 74674
rect 8370 74622 8372 74674
rect 8316 73442 8372 74622
rect 8316 73390 8318 73442
rect 8370 73390 8372 73442
rect 8316 72436 8372 73390
rect 8316 72370 8372 72380
rect 7980 70366 7982 70418
rect 8034 70366 8036 70418
rect 7980 70354 8036 70366
rect 8428 70420 8484 76974
rect 8540 76692 8596 76702
rect 8540 75682 8596 76636
rect 8540 75630 8542 75682
rect 8594 75630 8596 75682
rect 8540 75618 8596 75630
rect 8652 74900 8708 77756
rect 8876 77364 8932 78094
rect 9212 78148 9268 78158
rect 9324 78148 9380 83244
rect 9436 82404 9492 82414
rect 9436 82066 9492 82348
rect 9660 82292 9716 84476
rect 9772 84418 9828 84812
rect 9996 84802 10052 84812
rect 10332 84866 10388 84878
rect 10332 84814 10334 84866
rect 10386 84814 10388 84866
rect 9772 84366 9774 84418
rect 9826 84366 9828 84418
rect 9772 84354 9828 84366
rect 10220 83748 10276 83758
rect 9660 82236 10164 82292
rect 9436 82014 9438 82066
rect 9490 82014 9492 82066
rect 9436 82002 9492 82014
rect 9884 81844 9940 81854
rect 9660 81842 9940 81844
rect 9660 81790 9886 81842
rect 9938 81790 9940 81842
rect 9660 81788 9940 81790
rect 9660 81170 9716 81788
rect 9884 81778 9940 81788
rect 9660 81118 9662 81170
rect 9714 81118 9716 81170
rect 9660 80164 9716 81118
rect 9772 81172 9828 81182
rect 9772 80498 9828 81116
rect 9884 81060 9940 81070
rect 9884 80966 9940 81004
rect 9772 80446 9774 80498
rect 9826 80446 9828 80498
rect 9772 80434 9828 80446
rect 9884 80388 9940 80398
rect 9996 80388 10052 82236
rect 10108 81954 10164 82236
rect 10108 81902 10110 81954
rect 10162 81902 10164 81954
rect 10108 81890 10164 81902
rect 10220 81956 10276 83692
rect 10332 82404 10388 84814
rect 10892 83748 10948 83758
rect 10332 82338 10388 82348
rect 10668 82740 10724 82750
rect 10444 82068 10500 82078
rect 10444 81974 10500 82012
rect 10332 81956 10388 81966
rect 10220 81954 10388 81956
rect 10220 81902 10334 81954
rect 10386 81902 10388 81954
rect 10220 81900 10388 81902
rect 10332 81890 10388 81900
rect 10556 81956 10612 81966
rect 10668 81956 10724 82684
rect 10892 82738 10948 83692
rect 10892 82686 10894 82738
rect 10946 82686 10948 82738
rect 10892 82674 10948 82686
rect 11004 82348 11060 86492
rect 11900 86548 11956 86558
rect 11900 86454 11956 86492
rect 10556 81954 10724 81956
rect 10556 81902 10558 81954
rect 10610 81902 10724 81954
rect 10556 81900 10724 81902
rect 10780 82292 11060 82348
rect 11116 86436 11172 86446
rect 11116 82962 11172 86380
rect 12348 85876 12404 87388
rect 12572 87442 12628 87948
rect 12572 87390 12574 87442
rect 12626 87390 12628 87442
rect 12572 87378 12628 87390
rect 12796 88002 12852 88014
rect 12796 87950 12798 88002
rect 12850 87950 12852 88002
rect 12796 87220 12852 87950
rect 12460 86660 12516 86670
rect 12460 86566 12516 86604
rect 12796 86212 12852 87164
rect 12908 86770 12964 94108
rect 14008 94108 15208 94118
rect 14064 94106 14112 94108
rect 14168 94106 14216 94108
rect 14076 94054 14112 94106
rect 14200 94054 14216 94106
rect 14064 94052 14112 94054
rect 14168 94052 14216 94054
rect 14272 94106 14320 94108
rect 14376 94106 14424 94108
rect 14480 94106 14528 94108
rect 14376 94054 14396 94106
rect 14480 94054 14520 94106
rect 14272 94052 14320 94054
rect 14376 94052 14424 94054
rect 14480 94052 14528 94054
rect 14584 94052 14632 94108
rect 14688 94106 14736 94108
rect 14792 94106 14840 94108
rect 14896 94106 14944 94108
rect 14696 94054 14736 94106
rect 14820 94054 14840 94106
rect 14688 94052 14736 94054
rect 14792 94052 14840 94054
rect 14896 94052 14944 94054
rect 15000 94106 15048 94108
rect 15104 94106 15152 94108
rect 15000 94054 15016 94106
rect 15104 94054 15140 94106
rect 15000 94052 15048 94054
rect 15104 94052 15152 94054
rect 14008 94042 15208 94052
rect 24008 93324 25208 93334
rect 24064 93322 24112 93324
rect 24168 93322 24216 93324
rect 24076 93270 24112 93322
rect 24200 93270 24216 93322
rect 24064 93268 24112 93270
rect 24168 93268 24216 93270
rect 24272 93322 24320 93324
rect 24376 93322 24424 93324
rect 24480 93322 24528 93324
rect 24376 93270 24396 93322
rect 24480 93270 24520 93322
rect 24272 93268 24320 93270
rect 24376 93268 24424 93270
rect 24480 93268 24528 93270
rect 24584 93268 24632 93324
rect 24688 93322 24736 93324
rect 24792 93322 24840 93324
rect 24896 93322 24944 93324
rect 24696 93270 24736 93322
rect 24820 93270 24840 93322
rect 24688 93268 24736 93270
rect 24792 93268 24840 93270
rect 24896 93268 24944 93270
rect 25000 93322 25048 93324
rect 25104 93322 25152 93324
rect 25000 93270 25016 93322
rect 25104 93270 25140 93322
rect 25000 93268 25048 93270
rect 25104 93268 25152 93270
rect 24008 93258 25208 93268
rect 14008 92540 15208 92550
rect 14064 92538 14112 92540
rect 14168 92538 14216 92540
rect 14076 92486 14112 92538
rect 14200 92486 14216 92538
rect 14064 92484 14112 92486
rect 14168 92484 14216 92486
rect 14272 92538 14320 92540
rect 14376 92538 14424 92540
rect 14480 92538 14528 92540
rect 14376 92486 14396 92538
rect 14480 92486 14520 92538
rect 14272 92484 14320 92486
rect 14376 92484 14424 92486
rect 14480 92484 14528 92486
rect 14584 92484 14632 92540
rect 14688 92538 14736 92540
rect 14792 92538 14840 92540
rect 14896 92538 14944 92540
rect 14696 92486 14736 92538
rect 14820 92486 14840 92538
rect 14688 92484 14736 92486
rect 14792 92484 14840 92486
rect 14896 92484 14944 92486
rect 15000 92538 15048 92540
rect 15104 92538 15152 92540
rect 15000 92486 15016 92538
rect 15104 92486 15140 92538
rect 15000 92484 15048 92486
rect 15104 92484 15152 92486
rect 14008 92474 15208 92484
rect 24008 91756 25208 91766
rect 24064 91754 24112 91756
rect 24168 91754 24216 91756
rect 24076 91702 24112 91754
rect 24200 91702 24216 91754
rect 24064 91700 24112 91702
rect 24168 91700 24216 91702
rect 24272 91754 24320 91756
rect 24376 91754 24424 91756
rect 24480 91754 24528 91756
rect 24376 91702 24396 91754
rect 24480 91702 24520 91754
rect 24272 91700 24320 91702
rect 24376 91700 24424 91702
rect 24480 91700 24528 91702
rect 24584 91700 24632 91756
rect 24688 91754 24736 91756
rect 24792 91754 24840 91756
rect 24896 91754 24944 91756
rect 24696 91702 24736 91754
rect 24820 91702 24840 91754
rect 24688 91700 24736 91702
rect 24792 91700 24840 91702
rect 24896 91700 24944 91702
rect 25000 91754 25048 91756
rect 25104 91754 25152 91756
rect 25000 91702 25016 91754
rect 25104 91702 25140 91754
rect 25000 91700 25048 91702
rect 25104 91700 25152 91702
rect 24008 91690 25208 91700
rect 14008 90972 15208 90982
rect 14064 90970 14112 90972
rect 14168 90970 14216 90972
rect 14076 90918 14112 90970
rect 14200 90918 14216 90970
rect 14064 90916 14112 90918
rect 14168 90916 14216 90918
rect 14272 90970 14320 90972
rect 14376 90970 14424 90972
rect 14480 90970 14528 90972
rect 14376 90918 14396 90970
rect 14480 90918 14520 90970
rect 14272 90916 14320 90918
rect 14376 90916 14424 90918
rect 14480 90916 14528 90918
rect 14584 90916 14632 90972
rect 14688 90970 14736 90972
rect 14792 90970 14840 90972
rect 14896 90970 14944 90972
rect 14696 90918 14736 90970
rect 14820 90918 14840 90970
rect 14688 90916 14736 90918
rect 14792 90916 14840 90918
rect 14896 90916 14944 90918
rect 15000 90970 15048 90972
rect 15104 90970 15152 90972
rect 15000 90918 15016 90970
rect 15104 90918 15140 90970
rect 15000 90916 15048 90918
rect 15104 90916 15152 90918
rect 14008 90906 15208 90916
rect 24008 90188 25208 90198
rect 24064 90186 24112 90188
rect 24168 90186 24216 90188
rect 24076 90134 24112 90186
rect 24200 90134 24216 90186
rect 24064 90132 24112 90134
rect 24168 90132 24216 90134
rect 24272 90186 24320 90188
rect 24376 90186 24424 90188
rect 24480 90186 24528 90188
rect 24376 90134 24396 90186
rect 24480 90134 24520 90186
rect 24272 90132 24320 90134
rect 24376 90132 24424 90134
rect 24480 90132 24528 90134
rect 24584 90132 24632 90188
rect 24688 90186 24736 90188
rect 24792 90186 24840 90188
rect 24896 90186 24944 90188
rect 24696 90134 24736 90186
rect 24820 90134 24840 90186
rect 24688 90132 24736 90134
rect 24792 90132 24840 90134
rect 24896 90132 24944 90134
rect 25000 90186 25048 90188
rect 25104 90186 25152 90188
rect 25000 90134 25016 90186
rect 25104 90134 25140 90186
rect 25000 90132 25048 90134
rect 25104 90132 25152 90134
rect 24008 90122 25208 90132
rect 13692 89570 13748 89582
rect 13692 89518 13694 89570
rect 13746 89518 13748 89570
rect 13580 88898 13636 88910
rect 13580 88846 13582 88898
rect 13634 88846 13636 88898
rect 13132 88788 13188 88798
rect 13020 88786 13188 88788
rect 13020 88734 13134 88786
rect 13186 88734 13188 88786
rect 13020 88732 13188 88734
rect 13020 86882 13076 88732
rect 13132 88722 13188 88732
rect 13580 88452 13636 88846
rect 13692 88900 13748 89518
rect 14008 89404 15208 89414
rect 14064 89402 14112 89404
rect 14168 89402 14216 89404
rect 14076 89350 14112 89402
rect 14200 89350 14216 89402
rect 14064 89348 14112 89350
rect 14168 89348 14216 89350
rect 14272 89402 14320 89404
rect 14376 89402 14424 89404
rect 14480 89402 14528 89404
rect 14376 89350 14396 89402
rect 14480 89350 14520 89402
rect 14272 89348 14320 89350
rect 14376 89348 14424 89350
rect 14480 89348 14528 89350
rect 14584 89348 14632 89404
rect 14688 89402 14736 89404
rect 14792 89402 14840 89404
rect 14896 89402 14944 89404
rect 14696 89350 14736 89402
rect 14820 89350 14840 89402
rect 14688 89348 14736 89350
rect 14792 89348 14840 89350
rect 14896 89348 14944 89350
rect 15000 89402 15048 89404
rect 15104 89402 15152 89404
rect 15000 89350 15016 89402
rect 15104 89350 15140 89402
rect 15000 89348 15048 89350
rect 15104 89348 15152 89350
rect 14008 89338 15208 89348
rect 13916 88900 13972 88910
rect 13692 88844 13916 88900
rect 13916 88806 13972 88844
rect 14252 88900 14308 88910
rect 13580 88396 14196 88452
rect 13244 88228 13300 88238
rect 13020 86830 13022 86882
rect 13074 86830 13076 86882
rect 13020 86818 13076 86830
rect 13132 88172 13244 88228
rect 12908 86718 12910 86770
rect 12962 86718 12964 86770
rect 12908 86660 12964 86718
rect 12908 86594 12964 86604
rect 12236 84532 12292 84542
rect 12348 84532 12404 85820
rect 12236 84530 12404 84532
rect 12236 84478 12238 84530
rect 12290 84478 12404 84530
rect 12236 84476 12404 84478
rect 12460 86156 12852 86212
rect 12236 84466 12292 84476
rect 11116 82910 11118 82962
rect 11170 82910 11172 82962
rect 10556 81890 10612 81900
rect 10780 81732 10836 82292
rect 11004 82180 11060 82190
rect 11116 82180 11172 82910
rect 11788 84308 11844 84318
rect 11788 84194 11844 84252
rect 11788 84142 11790 84194
rect 11842 84142 11844 84194
rect 11340 82738 11396 82750
rect 11340 82686 11342 82738
rect 11394 82686 11396 82738
rect 11228 82626 11284 82638
rect 11228 82574 11230 82626
rect 11282 82574 11284 82626
rect 11228 82348 11284 82574
rect 11228 82282 11284 82292
rect 11340 82292 11396 82686
rect 11788 82628 11844 84142
rect 11788 82562 11844 82572
rect 12124 83746 12180 83758
rect 12124 83694 12126 83746
rect 12178 83694 12180 83746
rect 11340 82236 11508 82292
rect 11116 82124 11396 82180
rect 11004 81956 11060 82124
rect 11116 81956 11172 81966
rect 11004 81954 11172 81956
rect 11004 81902 11118 81954
rect 11170 81902 11172 81954
rect 11004 81900 11172 81902
rect 11116 81890 11172 81900
rect 11340 81954 11396 82124
rect 11340 81902 11342 81954
rect 11394 81902 11396 81954
rect 11340 81890 11396 81902
rect 11452 81954 11508 82236
rect 11900 82180 11956 82190
rect 11452 81902 11454 81954
rect 11506 81902 11508 81954
rect 10332 81676 10836 81732
rect 10892 81842 10948 81854
rect 10892 81790 10894 81842
rect 10946 81790 10948 81842
rect 10220 81508 10276 81518
rect 10108 80500 10164 80510
rect 10108 80406 10164 80444
rect 9884 80386 10052 80388
rect 9884 80334 9886 80386
rect 9938 80334 10052 80386
rect 9884 80332 10052 80334
rect 9884 80322 9940 80332
rect 9660 80070 9716 80108
rect 9268 78092 9380 78148
rect 9660 79156 9716 79166
rect 9212 78082 9268 78092
rect 9548 78034 9604 78046
rect 9548 77982 9550 78034
rect 9602 77982 9604 78034
rect 8988 77924 9044 77934
rect 9548 77924 9604 77982
rect 8988 77922 9604 77924
rect 8988 77870 8990 77922
rect 9042 77870 9604 77922
rect 8988 77868 9604 77870
rect 9660 77924 9716 79100
rect 8988 77858 9044 77868
rect 8876 77298 8932 77308
rect 9660 77250 9716 77868
rect 9660 77198 9662 77250
rect 9714 77198 9716 77250
rect 9660 77186 9716 77198
rect 9772 78932 9828 78942
rect 10220 78932 10276 81452
rect 10332 81170 10388 81676
rect 10892 81508 10948 81790
rect 11452 81844 11508 81902
rect 11452 81778 11508 81788
rect 11788 81954 11844 81966
rect 11788 81902 11790 81954
rect 11842 81902 11844 81954
rect 11228 81732 11284 81742
rect 10780 81452 10948 81508
rect 11004 81730 11284 81732
rect 11004 81678 11230 81730
rect 11282 81678 11284 81730
rect 11004 81676 11284 81678
rect 10332 81118 10334 81170
rect 10386 81118 10388 81170
rect 10332 80948 10388 81118
rect 10444 81340 10724 81396
rect 10444 81170 10500 81340
rect 10444 81118 10446 81170
rect 10498 81118 10500 81170
rect 10444 81106 10500 81118
rect 10556 81170 10612 81182
rect 10556 81118 10558 81170
rect 10610 81118 10612 81170
rect 10332 80892 10500 80948
rect 10332 80724 10388 80734
rect 10332 80610 10388 80668
rect 10332 80558 10334 80610
rect 10386 80558 10388 80610
rect 10332 80546 10388 80558
rect 10444 80164 10500 80892
rect 10556 80388 10612 81118
rect 10668 81060 10724 81340
rect 10668 80994 10724 81004
rect 10780 80724 10836 81452
rect 10892 81284 10948 81294
rect 11004 81284 11060 81676
rect 11228 81666 11284 81676
rect 10892 81282 11060 81284
rect 10892 81230 10894 81282
rect 10946 81230 11060 81282
rect 10892 81228 11060 81230
rect 10892 81218 10948 81228
rect 11676 81172 11732 81182
rect 11676 81078 11732 81116
rect 11116 80946 11172 80958
rect 11116 80894 11118 80946
rect 11170 80894 11172 80946
rect 11004 80836 11060 80846
rect 10836 80668 10948 80724
rect 10780 80658 10836 80668
rect 10556 80322 10612 80332
rect 10556 80164 10612 80174
rect 10444 80108 10556 80164
rect 10556 80098 10612 80108
rect 10556 79492 10612 79502
rect 10444 79436 10556 79492
rect 10220 78876 10388 78932
rect 9772 76916 9828 78876
rect 9884 78820 9940 78830
rect 9884 78258 9940 78764
rect 9884 78206 9886 78258
rect 9938 78206 9940 78258
rect 9884 78194 9940 78206
rect 9996 78596 10052 78606
rect 9884 78036 9940 78046
rect 9996 78036 10052 78540
rect 9884 78034 10052 78036
rect 9884 77982 9886 78034
rect 9938 77982 10052 78034
rect 9884 77980 10052 77982
rect 10108 78036 10164 78046
rect 9884 77970 9940 77980
rect 10108 77942 10164 77980
rect 10108 77700 10164 77710
rect 10108 77250 10164 77644
rect 10108 77198 10110 77250
rect 10162 77198 10164 77250
rect 10108 77186 10164 77198
rect 9660 76860 9828 76916
rect 9324 76692 9380 76702
rect 8876 75684 8932 75694
rect 8876 75124 8932 75628
rect 8540 74786 8596 74798
rect 8540 74734 8542 74786
rect 8594 74734 8596 74786
rect 8540 73220 8596 74734
rect 8540 73154 8596 73164
rect 8652 72324 8708 74844
rect 8764 75122 8932 75124
rect 8764 75070 8878 75122
rect 8930 75070 8932 75122
rect 8764 75068 8932 75070
rect 8764 73948 8820 75068
rect 8876 75058 8932 75068
rect 8988 74900 9044 74910
rect 8988 74806 9044 74844
rect 8876 74676 8932 74686
rect 8876 74582 8932 74620
rect 8764 73892 9156 73948
rect 9100 73554 9156 73892
rect 9100 73502 9102 73554
rect 9154 73502 9156 73554
rect 9100 73490 9156 73502
rect 8428 70364 8596 70420
rect 7756 70194 7812 70206
rect 7756 70142 7758 70194
rect 7810 70142 7812 70194
rect 7420 70084 7476 70094
rect 7756 70084 7812 70142
rect 8428 70196 8484 70206
rect 8428 70102 8484 70140
rect 7476 70028 7812 70084
rect 7868 70082 7924 70094
rect 7868 70030 7870 70082
rect 7922 70030 7924 70082
rect 7420 69990 7476 70028
rect 7868 69748 7924 70030
rect 7420 69692 7924 69748
rect 6972 69410 7252 69412
rect 6972 69358 6974 69410
rect 7026 69358 7252 69410
rect 6972 69356 7252 69358
rect 6972 69346 7028 69356
rect 7196 68850 7252 69356
rect 7420 69410 7476 69692
rect 7420 69358 7422 69410
rect 7474 69358 7476 69410
rect 7420 69346 7476 69358
rect 7196 68798 7198 68850
rect 7250 68798 7252 68850
rect 6860 68402 6916 68414
rect 6860 68350 6862 68402
rect 6914 68350 6916 68402
rect 6860 68068 6916 68350
rect 6860 68002 6916 68012
rect 6524 67330 6580 67340
rect 6636 67618 6692 67630
rect 6636 67566 6638 67618
rect 6690 67566 6692 67618
rect 6300 67106 6356 67116
rect 6524 67172 6580 67182
rect 5740 65958 5796 65996
rect 5852 66892 6132 66948
rect 5292 65438 5294 65490
rect 5346 65438 5348 65490
rect 5292 65426 5348 65438
rect 5516 65660 5684 65716
rect 3276 65202 3332 65212
rect 3836 65212 4676 65268
rect 3836 64930 3892 65212
rect 4008 65100 5208 65110
rect 4064 65098 4112 65100
rect 4168 65098 4216 65100
rect 4076 65046 4112 65098
rect 4200 65046 4216 65098
rect 4064 65044 4112 65046
rect 4168 65044 4216 65046
rect 4272 65098 4320 65100
rect 4376 65098 4424 65100
rect 4480 65098 4528 65100
rect 4376 65046 4396 65098
rect 4480 65046 4520 65098
rect 4272 65044 4320 65046
rect 4376 65044 4424 65046
rect 4480 65044 4528 65046
rect 4584 65044 4632 65100
rect 4688 65098 4736 65100
rect 4792 65098 4840 65100
rect 4896 65098 4944 65100
rect 4696 65046 4736 65098
rect 4820 65046 4840 65098
rect 4688 65044 4736 65046
rect 4792 65044 4840 65046
rect 4896 65044 4944 65046
rect 5000 65098 5048 65100
rect 5104 65098 5152 65100
rect 5000 65046 5016 65098
rect 5104 65046 5140 65098
rect 5000 65044 5048 65046
rect 5104 65044 5152 65046
rect 4008 65034 5208 65044
rect 3836 64878 3838 64930
rect 3890 64878 3892 64930
rect 3836 64866 3892 64878
rect 3164 64596 3220 64606
rect 3164 64502 3220 64540
rect 3724 64596 3780 64606
rect 3724 64502 3780 64540
rect 4844 64146 4900 64158
rect 4844 64094 4846 64146
rect 4898 64094 4900 64146
rect 4844 64036 4900 64094
rect 4844 63970 4900 63980
rect 5292 64148 5348 64158
rect 4008 63532 5208 63542
rect 4064 63530 4112 63532
rect 4168 63530 4216 63532
rect 4076 63478 4112 63530
rect 4200 63478 4216 63530
rect 4064 63476 4112 63478
rect 4168 63476 4216 63478
rect 4272 63530 4320 63532
rect 4376 63530 4424 63532
rect 4480 63530 4528 63532
rect 4376 63478 4396 63530
rect 4480 63478 4520 63530
rect 4272 63476 4320 63478
rect 4376 63476 4424 63478
rect 4480 63476 4528 63478
rect 4584 63476 4632 63532
rect 4688 63530 4736 63532
rect 4792 63530 4840 63532
rect 4896 63530 4944 63532
rect 4696 63478 4736 63530
rect 4820 63478 4840 63530
rect 4688 63476 4736 63478
rect 4792 63476 4840 63478
rect 4896 63476 4944 63478
rect 5000 63530 5048 63532
rect 5104 63530 5152 63532
rect 5000 63478 5016 63530
rect 5104 63478 5140 63530
rect 5000 63476 5048 63478
rect 5104 63476 5152 63478
rect 4008 63466 5208 63476
rect 3836 63364 3892 63374
rect 3836 63270 3892 63308
rect 4732 63364 4788 63374
rect 4172 63252 4228 63262
rect 4172 63158 4228 63196
rect 3500 63028 3556 63038
rect 3500 57540 3556 62972
rect 4732 63028 4788 63308
rect 4956 63140 5012 63150
rect 4956 63046 5012 63084
rect 4732 62934 4788 62972
rect 4732 62636 5012 62692
rect 4396 62356 4452 62366
rect 4396 62262 4452 62300
rect 4732 62354 4788 62636
rect 4844 62468 4900 62478
rect 4844 62374 4900 62412
rect 4732 62302 4734 62354
rect 4786 62302 4788 62354
rect 4732 62290 4788 62302
rect 4844 62244 4900 62254
rect 4844 62130 4900 62188
rect 4844 62078 4846 62130
rect 4898 62078 4900 62130
rect 4844 62066 4900 62078
rect 4956 62132 5012 62636
rect 5292 62356 5348 64092
rect 5404 63924 5460 63934
rect 5404 63252 5460 63868
rect 5404 63186 5460 63196
rect 5516 63588 5572 65660
rect 5628 65492 5684 65502
rect 5628 65398 5684 65436
rect 5740 65156 5796 65166
rect 5628 65100 5740 65156
rect 5628 64148 5684 65100
rect 5740 65090 5796 65100
rect 5740 64484 5796 64494
rect 5852 64484 5908 66892
rect 6412 66276 6468 66286
rect 5740 64482 5908 64484
rect 5740 64430 5742 64482
rect 5794 64430 5908 64482
rect 5740 64428 5908 64430
rect 5740 64418 5796 64428
rect 5740 64148 5796 64158
rect 5628 64146 5796 64148
rect 5628 64094 5742 64146
rect 5794 64094 5796 64146
rect 5628 64092 5796 64094
rect 5628 63812 5684 64092
rect 5740 64082 5796 64092
rect 5852 64036 5908 64428
rect 5852 63970 5908 63980
rect 6076 66052 6132 66062
rect 5628 63746 5684 63756
rect 5516 63532 5796 63588
rect 5516 62468 5572 63532
rect 5740 63250 5796 63532
rect 5740 63198 5742 63250
rect 5794 63198 5796 63250
rect 5740 63186 5796 63198
rect 6076 63140 6132 65996
rect 6188 65716 6244 65726
rect 6188 65490 6244 65660
rect 6188 65438 6190 65490
rect 6242 65438 6244 65490
rect 6188 65426 6244 65438
rect 6300 65492 6356 65502
rect 6188 64148 6244 64158
rect 6300 64148 6356 65436
rect 6244 64092 6356 64148
rect 6188 64054 6244 64092
rect 6188 63140 6244 63150
rect 6076 63084 6188 63140
rect 6188 63046 6244 63084
rect 5516 62402 5572 62412
rect 5292 62354 5460 62356
rect 5292 62302 5294 62354
rect 5346 62302 5460 62354
rect 5292 62300 5460 62302
rect 5292 62290 5348 62300
rect 5404 62188 5460 62300
rect 5740 62354 5796 62366
rect 5740 62302 5742 62354
rect 5794 62302 5796 62354
rect 4956 62066 5012 62076
rect 5292 62132 5348 62142
rect 5404 62132 5572 62188
rect 4008 61964 5208 61974
rect 4064 61962 4112 61964
rect 4168 61962 4216 61964
rect 4076 61910 4112 61962
rect 4200 61910 4216 61962
rect 4064 61908 4112 61910
rect 4168 61908 4216 61910
rect 4272 61962 4320 61964
rect 4376 61962 4424 61964
rect 4480 61962 4528 61964
rect 4376 61910 4396 61962
rect 4480 61910 4520 61962
rect 4272 61908 4320 61910
rect 4376 61908 4424 61910
rect 4480 61908 4528 61910
rect 4584 61908 4632 61964
rect 4688 61962 4736 61964
rect 4792 61962 4840 61964
rect 4896 61962 4944 61964
rect 4696 61910 4736 61962
rect 4820 61910 4840 61962
rect 4688 61908 4736 61910
rect 4792 61908 4840 61910
rect 4896 61908 4944 61910
rect 5000 61962 5048 61964
rect 5104 61962 5152 61964
rect 5000 61910 5016 61962
rect 5104 61910 5140 61962
rect 5000 61908 5048 61910
rect 5104 61908 5152 61910
rect 4008 61898 5208 61908
rect 4060 61572 4116 61582
rect 4060 61478 4116 61516
rect 4620 61570 4676 61582
rect 4620 61518 4622 61570
rect 4674 61518 4676 61570
rect 3836 61460 3892 61470
rect 3724 61348 3780 61358
rect 3724 61254 3780 61292
rect 3724 58548 3780 58558
rect 3388 57538 3556 57540
rect 3388 57486 3502 57538
rect 3554 57486 3556 57538
rect 3388 57484 3556 57486
rect 3276 56644 3332 56654
rect 3276 56550 3332 56588
rect 3276 55972 3332 55982
rect 3276 55878 3332 55916
rect 3052 55412 3220 55468
rect 2604 55076 2660 55086
rect 2828 55076 2884 55086
rect 2604 55074 2884 55076
rect 2604 55022 2606 55074
rect 2658 55022 2830 55074
rect 2882 55022 2884 55074
rect 2604 55020 2884 55022
rect 2604 54964 2660 55020
rect 2828 55010 2884 55020
rect 2604 54898 2660 54908
rect 2268 54462 2270 54514
rect 2322 54462 2324 54514
rect 2268 54450 2324 54462
rect 2492 53844 2548 53854
rect 2492 53732 2548 53788
rect 2828 53732 2884 53742
rect 2492 53730 2884 53732
rect 2492 53678 2494 53730
rect 2546 53678 2830 53730
rect 2882 53678 2884 53730
rect 2492 53676 2884 53678
rect 2492 53666 2548 53676
rect 2828 53666 2884 53676
rect 2492 52948 2548 52958
rect 2492 52854 2548 52892
rect 2828 52946 2884 52958
rect 2828 52894 2830 52946
rect 2882 52894 2884 52946
rect 2828 52724 2884 52894
rect 2828 52658 2884 52668
rect 3164 52612 3220 55412
rect 3276 55410 3332 55422
rect 3276 55358 3278 55410
rect 3330 55358 3332 55410
rect 3276 55300 3332 55358
rect 3276 55234 3332 55244
rect 3276 53844 3332 53854
rect 3276 53750 3332 53788
rect 3276 53284 3332 53294
rect 3276 52834 3332 53228
rect 3276 52782 3278 52834
rect 3330 52782 3332 52834
rect 3276 52770 3332 52782
rect 2268 51390 2324 51402
rect 2268 51338 2270 51390
rect 2322 51380 2324 51390
rect 2380 51380 2436 51390
rect 2322 51338 2380 51380
rect 2268 51324 2380 51338
rect 2380 51314 2436 51324
rect 2156 50418 2212 50428
rect 2828 49810 2884 49822
rect 2828 49758 2830 49810
rect 2882 49758 2884 49810
rect 2492 49700 2548 49710
rect 2828 49700 2884 49758
rect 2492 49698 2884 49700
rect 2492 49646 2494 49698
rect 2546 49646 2884 49698
rect 2492 49644 2884 49646
rect 3164 49700 3220 52556
rect 3276 51938 3332 51950
rect 3276 51886 3278 51938
rect 3330 51886 3332 51938
rect 3276 51380 3332 51886
rect 3388 51940 3444 57484
rect 3500 57474 3556 57484
rect 3612 58492 3724 58548
rect 3612 57092 3668 58492
rect 3724 58482 3780 58492
rect 3500 57036 3668 57092
rect 3500 53172 3556 57036
rect 3612 56868 3668 56878
rect 3836 56868 3892 61404
rect 4620 61460 4676 61518
rect 4620 61394 4676 61404
rect 4844 61458 4900 61470
rect 4844 61406 4846 61458
rect 4898 61406 4900 61458
rect 4732 61348 4788 61358
rect 4732 61010 4788 61292
rect 4732 60958 4734 61010
rect 4786 60958 4788 61010
rect 4732 60946 4788 60958
rect 4844 61012 4900 61406
rect 5292 61012 5348 62076
rect 4844 61010 5348 61012
rect 4844 60958 5294 61010
rect 5346 60958 5348 61010
rect 4844 60956 5348 60958
rect 5292 60946 5348 60956
rect 4008 60396 5208 60406
rect 4064 60394 4112 60396
rect 4168 60394 4216 60396
rect 4076 60342 4112 60394
rect 4200 60342 4216 60394
rect 4064 60340 4112 60342
rect 4168 60340 4216 60342
rect 4272 60394 4320 60396
rect 4376 60394 4424 60396
rect 4480 60394 4528 60396
rect 4376 60342 4396 60394
rect 4480 60342 4520 60394
rect 4272 60340 4320 60342
rect 4376 60340 4424 60342
rect 4480 60340 4528 60342
rect 4584 60340 4632 60396
rect 4688 60394 4736 60396
rect 4792 60394 4840 60396
rect 4896 60394 4944 60396
rect 4696 60342 4736 60394
rect 4820 60342 4840 60394
rect 4688 60340 4736 60342
rect 4792 60340 4840 60342
rect 4896 60340 4944 60342
rect 5000 60394 5048 60396
rect 5104 60394 5152 60396
rect 5000 60342 5016 60394
rect 5104 60342 5140 60394
rect 5000 60340 5048 60342
rect 5104 60340 5152 60342
rect 4008 60330 5208 60340
rect 5516 60116 5572 62132
rect 5628 61572 5684 61582
rect 5740 61572 5796 62302
rect 5964 61684 6020 61694
rect 5740 61516 5908 61572
rect 5628 61010 5684 61516
rect 5740 61348 5796 61358
rect 5740 61254 5796 61292
rect 5628 60958 5630 61010
rect 5682 60958 5684 61010
rect 5628 60946 5684 60958
rect 5852 60900 5908 61516
rect 5852 60834 5908 60844
rect 5964 60786 6020 61628
rect 5964 60734 5966 60786
rect 6018 60734 6020 60786
rect 5964 60226 6020 60734
rect 5964 60174 5966 60226
rect 6018 60174 6020 60226
rect 5740 60116 5796 60126
rect 5516 60060 5740 60116
rect 5740 60022 5796 60060
rect 4008 58828 5208 58838
rect 4064 58826 4112 58828
rect 4168 58826 4216 58828
rect 4076 58774 4112 58826
rect 4200 58774 4216 58826
rect 4064 58772 4112 58774
rect 4168 58772 4216 58774
rect 4272 58826 4320 58828
rect 4376 58826 4424 58828
rect 4480 58826 4528 58828
rect 4376 58774 4396 58826
rect 4480 58774 4520 58826
rect 4272 58772 4320 58774
rect 4376 58772 4424 58774
rect 4480 58772 4528 58774
rect 4584 58772 4632 58828
rect 4688 58826 4736 58828
rect 4792 58826 4840 58828
rect 4896 58826 4944 58828
rect 4696 58774 4736 58826
rect 4820 58774 4840 58826
rect 4688 58772 4736 58774
rect 4792 58772 4840 58774
rect 4896 58772 4944 58774
rect 5000 58826 5048 58828
rect 5104 58826 5152 58828
rect 5000 58774 5016 58826
rect 5104 58774 5140 58826
rect 5000 58772 5048 58774
rect 5104 58772 5152 58774
rect 4008 58762 5208 58772
rect 3948 58548 4004 58558
rect 3948 58454 4004 58492
rect 4008 57260 5208 57270
rect 4064 57258 4112 57260
rect 4168 57258 4216 57260
rect 4076 57206 4112 57258
rect 4200 57206 4216 57258
rect 4064 57204 4112 57206
rect 4168 57204 4216 57206
rect 4272 57258 4320 57260
rect 4376 57258 4424 57260
rect 4480 57258 4528 57260
rect 4376 57206 4396 57258
rect 4480 57206 4520 57258
rect 4272 57204 4320 57206
rect 4376 57204 4424 57206
rect 4480 57204 4528 57206
rect 4584 57204 4632 57260
rect 4688 57258 4736 57260
rect 4792 57258 4840 57260
rect 4896 57258 4944 57260
rect 4696 57206 4736 57258
rect 4820 57206 4840 57258
rect 4688 57204 4736 57206
rect 4792 57204 4840 57206
rect 4896 57204 4944 57206
rect 5000 57258 5048 57260
rect 5104 57258 5152 57260
rect 5000 57206 5016 57258
rect 5104 57206 5140 57258
rect 5000 57204 5048 57206
rect 5104 57204 5152 57206
rect 4008 57194 5208 57204
rect 4284 56868 4340 56878
rect 3612 56866 3780 56868
rect 3612 56814 3614 56866
rect 3666 56814 3780 56866
rect 3612 56812 3780 56814
rect 3836 56866 4340 56868
rect 3836 56814 4286 56866
rect 4338 56814 4340 56866
rect 3836 56812 4340 56814
rect 3612 56802 3668 56812
rect 3724 56308 3780 56812
rect 4284 56644 4340 56812
rect 4396 56756 4452 56766
rect 4396 56662 4452 56700
rect 5292 56756 5348 56766
rect 4284 56578 4340 56588
rect 4956 56644 5012 56654
rect 4956 56550 5012 56588
rect 4172 56308 4228 56318
rect 3724 56252 3892 56308
rect 3724 56082 3780 56094
rect 3724 56030 3726 56082
rect 3778 56030 3780 56082
rect 3724 55412 3780 56030
rect 3836 55522 3892 56252
rect 4172 56082 4228 56252
rect 4172 56030 4174 56082
rect 4226 56030 4228 56082
rect 4172 56018 4228 56030
rect 4008 55692 5208 55702
rect 4064 55690 4112 55692
rect 4168 55690 4216 55692
rect 4076 55638 4112 55690
rect 4200 55638 4216 55690
rect 4064 55636 4112 55638
rect 4168 55636 4216 55638
rect 4272 55690 4320 55692
rect 4376 55690 4424 55692
rect 4480 55690 4528 55692
rect 4376 55638 4396 55690
rect 4480 55638 4520 55690
rect 4272 55636 4320 55638
rect 4376 55636 4424 55638
rect 4480 55636 4528 55638
rect 4584 55636 4632 55692
rect 4688 55690 4736 55692
rect 4792 55690 4840 55692
rect 4896 55690 4944 55692
rect 4696 55638 4736 55690
rect 4820 55638 4840 55690
rect 4688 55636 4736 55638
rect 4792 55636 4840 55638
rect 4896 55636 4944 55638
rect 5000 55690 5048 55692
rect 5104 55690 5152 55692
rect 5000 55638 5016 55690
rect 5104 55638 5140 55690
rect 5000 55636 5048 55638
rect 5104 55636 5152 55638
rect 4008 55626 5208 55636
rect 3836 55470 3838 55522
rect 3890 55470 3892 55522
rect 3836 55458 3892 55470
rect 3612 55300 3668 55310
rect 3612 53172 3668 55244
rect 3724 54740 3780 55356
rect 4172 55300 4228 55310
rect 3724 54674 3780 54684
rect 3836 55298 4228 55300
rect 3836 55246 4174 55298
rect 4226 55246 4228 55298
rect 3836 55244 4228 55246
rect 3836 53956 3892 55244
rect 4172 55234 4228 55244
rect 4844 55300 4900 55310
rect 4844 55206 4900 55244
rect 4956 55188 5012 55198
rect 4956 55094 5012 55132
rect 4732 54738 4788 54750
rect 4732 54686 4734 54738
rect 4786 54686 4788 54738
rect 4732 54292 4788 54686
rect 5292 54738 5348 56700
rect 5740 56642 5796 56654
rect 5740 56590 5742 56642
rect 5794 56590 5796 56642
rect 5740 56308 5796 56590
rect 5740 56242 5796 56252
rect 5740 55076 5796 55086
rect 5628 54740 5684 54750
rect 5292 54686 5294 54738
rect 5346 54686 5348 54738
rect 5292 54674 5348 54686
rect 5516 54684 5628 54740
rect 4732 54226 4788 54236
rect 4008 54124 5208 54134
rect 4064 54122 4112 54124
rect 4168 54122 4216 54124
rect 4076 54070 4112 54122
rect 4200 54070 4216 54122
rect 4064 54068 4112 54070
rect 4168 54068 4216 54070
rect 4272 54122 4320 54124
rect 4376 54122 4424 54124
rect 4480 54122 4528 54124
rect 4376 54070 4396 54122
rect 4480 54070 4520 54122
rect 4272 54068 4320 54070
rect 4376 54068 4424 54070
rect 4480 54068 4528 54070
rect 4584 54068 4632 54124
rect 4688 54122 4736 54124
rect 4792 54122 4840 54124
rect 4896 54122 4944 54124
rect 4696 54070 4736 54122
rect 4820 54070 4840 54122
rect 4688 54068 4736 54070
rect 4792 54068 4840 54070
rect 4896 54068 4944 54070
rect 5000 54122 5048 54124
rect 5104 54122 5152 54124
rect 5000 54070 5016 54122
rect 5104 54070 5140 54122
rect 5000 54068 5048 54070
rect 5104 54068 5152 54070
rect 4008 54058 5208 54068
rect 3836 53900 4116 53956
rect 4060 53732 4116 53900
rect 3612 53116 3892 53172
rect 3500 53106 3556 53116
rect 3388 51874 3444 51884
rect 3500 52948 3556 52958
rect 3724 52948 3780 52958
rect 3556 52946 3780 52948
rect 3556 52894 3726 52946
rect 3778 52894 3780 52946
rect 3556 52892 3780 52894
rect 3276 51314 3332 51324
rect 3388 51716 3444 51726
rect 3276 49700 3332 49710
rect 3164 49698 3332 49700
rect 3164 49646 3278 49698
rect 3330 49646 3332 49698
rect 3164 49644 3332 49646
rect 2492 49364 2548 49644
rect 3276 49634 3332 49644
rect 2492 49298 2548 49308
rect 3276 48580 3332 48590
rect 2492 48244 2548 48254
rect 2492 48150 2548 48188
rect 2940 48244 2996 48254
rect 2940 48150 2996 48188
rect 3276 48130 3332 48524
rect 3276 48078 3278 48130
rect 3330 48078 3332 48130
rect 3276 48066 3332 48078
rect 3276 47570 3332 47582
rect 3276 47518 3278 47570
rect 3330 47518 3332 47570
rect 3276 47460 3332 47518
rect 3388 47572 3444 51660
rect 3388 47506 3444 47516
rect 3276 47394 3332 47404
rect 2604 47348 2660 47358
rect 2604 47254 2660 47292
rect 3388 47348 3444 47358
rect 2156 47234 2212 47246
rect 2156 47182 2158 47234
rect 2210 47182 2212 47234
rect 2156 47124 2212 47182
rect 2156 47058 2212 47068
rect 2828 47234 2884 47246
rect 2828 47182 2830 47234
rect 2882 47182 2884 47234
rect 2828 47124 2884 47182
rect 2828 47058 2884 47068
rect 1820 46674 1876 46686
rect 1820 46622 1822 46674
rect 1874 46622 1876 46674
rect 1820 43764 1876 46622
rect 2492 46676 2548 46686
rect 2492 46582 2548 46620
rect 2492 46004 2548 46014
rect 3276 46004 3332 46014
rect 2548 45948 2884 46004
rect 2492 45910 2548 45948
rect 2828 45890 2884 45948
rect 3276 45910 3332 45948
rect 2828 45838 2830 45890
rect 2882 45838 2884 45890
rect 2828 45826 2884 45838
rect 3276 45220 3332 45230
rect 2828 45106 2884 45118
rect 2828 45054 2830 45106
rect 2882 45054 2884 45106
rect 2492 44996 2548 45006
rect 2828 44996 2884 45054
rect 2492 44994 2884 44996
rect 2492 44942 2494 44994
rect 2546 44942 2884 44994
rect 2492 44940 2884 44942
rect 3276 44994 3332 45164
rect 3276 44942 3278 44994
rect 3330 44942 3332 44994
rect 2492 44884 2548 44940
rect 3276 44930 3332 44942
rect 2492 44818 2548 44828
rect 1820 43538 1876 43708
rect 1820 43486 1822 43538
rect 1874 43486 1876 43538
rect 1820 40402 1876 43486
rect 2268 44100 2324 44110
rect 2268 43538 2324 44044
rect 3388 43876 3444 47292
rect 3388 43810 3444 43820
rect 2268 43486 2270 43538
rect 2322 43486 2324 43538
rect 2268 43474 2324 43486
rect 3388 43652 3444 43662
rect 3164 42756 3220 42766
rect 2828 42642 2884 42654
rect 2828 42590 2830 42642
rect 2882 42590 2884 42642
rect 2604 42532 2660 42542
rect 2828 42532 2884 42590
rect 3164 42642 3220 42700
rect 3164 42590 3166 42642
rect 3218 42590 3220 42642
rect 3164 42578 3220 42590
rect 2604 42530 2884 42532
rect 2604 42478 2606 42530
rect 2658 42478 2884 42530
rect 2604 42476 2884 42478
rect 2604 41524 2660 42476
rect 2604 41458 2660 41468
rect 3276 41300 3332 41310
rect 3164 41298 3332 41300
rect 3164 41246 3278 41298
rect 3330 41246 3332 41298
rect 3164 41244 3332 41246
rect 2604 40964 2660 40974
rect 2828 40964 2884 40974
rect 2604 40962 2884 40964
rect 2604 40910 2606 40962
rect 2658 40910 2830 40962
rect 2882 40910 2884 40962
rect 2604 40908 2884 40910
rect 1820 40350 1822 40402
rect 1874 40350 1876 40402
rect 1820 35698 1876 40350
rect 2268 40402 2324 40414
rect 2268 40350 2270 40402
rect 2322 40350 2324 40402
rect 2268 39844 2324 40350
rect 2604 40404 2660 40908
rect 2828 40898 2884 40908
rect 2604 40338 2660 40348
rect 2268 39778 2324 39788
rect 3164 39508 3220 41244
rect 3276 41234 3332 41244
rect 3164 39442 3220 39452
rect 3276 39618 3332 39630
rect 3276 39566 3278 39618
rect 3330 39566 3332 39618
rect 2492 39396 2548 39406
rect 2716 39396 2772 39406
rect 2492 39394 2772 39396
rect 2492 39342 2494 39394
rect 2546 39342 2718 39394
rect 2770 39342 2772 39394
rect 2492 39340 2772 39342
rect 2492 39284 2548 39340
rect 2716 39330 2772 39340
rect 2492 39218 2548 39228
rect 3164 39060 3220 39070
rect 3164 38966 3220 39004
rect 3276 38948 3332 39566
rect 3276 38882 3332 38892
rect 2828 38834 2884 38846
rect 2828 38782 2830 38834
rect 2882 38782 2884 38834
rect 2492 38724 2548 38734
rect 2828 38724 2884 38782
rect 2492 38722 2884 38724
rect 2492 38670 2494 38722
rect 2546 38670 2884 38722
rect 2492 38668 2884 38670
rect 3388 38668 3444 43596
rect 3500 42644 3556 52892
rect 3724 52882 3780 52892
rect 3612 52164 3668 52174
rect 3612 52162 3780 52164
rect 3612 52110 3614 52162
rect 3666 52110 3780 52162
rect 3612 52108 3780 52110
rect 3612 52098 3668 52108
rect 3612 51828 3668 51838
rect 3612 49924 3668 51772
rect 3724 50596 3780 52108
rect 3836 50820 3892 53116
rect 4060 53170 4116 53676
rect 4060 53118 4062 53170
rect 4114 53118 4116 53170
rect 4060 53106 4116 53118
rect 5180 53172 5236 53182
rect 5180 53078 5236 53116
rect 5404 52948 5460 52958
rect 5292 52946 5460 52948
rect 5292 52894 5406 52946
rect 5458 52894 5460 52946
rect 5292 52892 5460 52894
rect 4732 52836 4788 52846
rect 4732 52742 4788 52780
rect 4008 52556 5208 52566
rect 4064 52554 4112 52556
rect 4168 52554 4216 52556
rect 4076 52502 4112 52554
rect 4200 52502 4216 52554
rect 4064 52500 4112 52502
rect 4168 52500 4216 52502
rect 4272 52554 4320 52556
rect 4376 52554 4424 52556
rect 4480 52554 4528 52556
rect 4376 52502 4396 52554
rect 4480 52502 4520 52554
rect 4272 52500 4320 52502
rect 4376 52500 4424 52502
rect 4480 52500 4528 52502
rect 4584 52500 4632 52556
rect 4688 52554 4736 52556
rect 4792 52554 4840 52556
rect 4896 52554 4944 52556
rect 4696 52502 4736 52554
rect 4820 52502 4840 52554
rect 4688 52500 4736 52502
rect 4792 52500 4840 52502
rect 4896 52500 4944 52502
rect 5000 52554 5048 52556
rect 5104 52554 5152 52556
rect 5000 52502 5016 52554
rect 5104 52502 5140 52554
rect 5000 52500 5048 52502
rect 5104 52500 5152 52502
rect 4008 52490 5208 52500
rect 4060 52162 4116 52174
rect 4060 52110 4062 52162
rect 4114 52110 4116 52162
rect 4060 51716 4116 52110
rect 5180 52164 5236 52174
rect 5292 52164 5348 52892
rect 5404 52882 5460 52892
rect 5180 52162 5348 52164
rect 5180 52110 5182 52162
rect 5234 52110 5348 52162
rect 5180 52108 5348 52110
rect 5516 52162 5572 54684
rect 5628 54646 5684 54684
rect 5740 54292 5796 55020
rect 5740 54226 5796 54236
rect 5628 53732 5684 53742
rect 5628 53638 5684 53676
rect 5740 53620 5796 53658
rect 5740 53554 5796 53564
rect 5964 53396 6020 60174
rect 6188 60226 6244 60238
rect 6188 60174 6190 60226
rect 6242 60174 6244 60226
rect 6188 60114 6244 60174
rect 6188 60062 6190 60114
rect 6242 60062 6244 60114
rect 6188 60050 6244 60062
rect 6188 59780 6244 59790
rect 6076 57540 6132 57550
rect 6076 57090 6132 57484
rect 6076 57038 6078 57090
rect 6130 57038 6132 57090
rect 6076 57026 6132 57038
rect 6188 55972 6244 59724
rect 6412 56084 6468 66220
rect 6524 62188 6580 67116
rect 6636 66500 6692 67566
rect 6972 67620 7028 67630
rect 6860 66948 6916 66958
rect 6748 66500 6804 66510
rect 6636 66498 6804 66500
rect 6636 66446 6750 66498
rect 6802 66446 6804 66498
rect 6636 66444 6804 66446
rect 6748 66434 6804 66444
rect 6860 63252 6916 66892
rect 6972 66724 7028 67564
rect 6972 66276 7028 66668
rect 6972 66182 7028 66220
rect 7196 65492 7252 68798
rect 7644 68516 7700 68526
rect 7420 68514 7700 68516
rect 7420 68462 7646 68514
rect 7698 68462 7700 68514
rect 7420 68460 7700 68462
rect 7420 67508 7476 68460
rect 7644 68450 7700 68460
rect 8316 68068 8372 68078
rect 8540 68068 8596 70364
rect 8316 68066 8596 68068
rect 8316 68014 8318 68066
rect 8370 68014 8542 68066
rect 8594 68014 8596 68066
rect 8316 68012 8596 68014
rect 8316 68002 8372 68012
rect 7980 67956 8036 67966
rect 7420 67442 7476 67452
rect 7532 67954 8036 67956
rect 7532 67902 7982 67954
rect 8034 67902 8036 67954
rect 7532 67900 8036 67902
rect 7308 66836 7364 66846
rect 7308 66498 7364 66780
rect 7308 66446 7310 66498
rect 7362 66446 7364 66498
rect 7308 66434 7364 66446
rect 7532 66498 7588 67900
rect 7980 67890 8036 67900
rect 7756 67620 7812 67630
rect 8092 67620 8148 67630
rect 7756 67618 8148 67620
rect 7756 67566 7758 67618
rect 7810 67566 8094 67618
rect 8146 67566 8148 67618
rect 7756 67564 8148 67566
rect 7756 67554 7812 67564
rect 8092 66948 8148 67564
rect 7532 66446 7534 66498
rect 7586 66446 7588 66498
rect 7532 66434 7588 66446
rect 7644 66612 7700 66622
rect 7644 66050 7700 66556
rect 8092 66276 8148 66892
rect 8428 67058 8484 67070
rect 8428 67006 8430 67058
rect 8482 67006 8484 67058
rect 8428 66612 8484 67006
rect 8428 66546 8484 66556
rect 8428 66388 8484 66398
rect 8540 66388 8596 68012
rect 8428 66386 8596 66388
rect 8428 66334 8430 66386
rect 8482 66334 8596 66386
rect 8428 66332 8596 66334
rect 8428 66322 8484 66332
rect 8204 66276 8260 66286
rect 7644 65998 7646 66050
rect 7698 65998 7700 66050
rect 7644 65986 7700 65998
rect 7868 66220 8204 66276
rect 7868 65714 7924 66220
rect 8204 66182 8260 66220
rect 7868 65662 7870 65714
rect 7922 65662 7924 65714
rect 7868 65650 7924 65662
rect 7196 65426 7252 65436
rect 8540 65492 8596 65502
rect 7756 65380 7812 65390
rect 7756 64706 7812 65324
rect 8540 64818 8596 65436
rect 8540 64766 8542 64818
rect 8594 64766 8596 64818
rect 8540 64754 8596 64766
rect 7756 64654 7758 64706
rect 7810 64654 7812 64706
rect 7756 64642 7812 64654
rect 8428 64372 8484 64382
rect 8316 63812 8372 63822
rect 7532 63364 7588 63374
rect 7532 63270 7588 63308
rect 6860 63158 6916 63196
rect 7196 63140 7252 63150
rect 7084 63138 7252 63140
rect 7084 63086 7198 63138
rect 7250 63086 7252 63138
rect 7084 63084 7252 63086
rect 7084 62468 7140 63084
rect 7196 63074 7252 63084
rect 8316 63138 8372 63756
rect 8316 63086 8318 63138
rect 8370 63086 8372 63138
rect 8316 63074 8372 63086
rect 7420 62914 7476 62926
rect 7420 62862 7422 62914
rect 7474 62862 7476 62914
rect 7420 62580 7476 62862
rect 7980 62914 8036 62926
rect 7980 62862 7982 62914
rect 8034 62862 8036 62914
rect 7420 62524 7924 62580
rect 6524 62132 6804 62188
rect 6748 61682 6804 62132
rect 6748 61630 6750 61682
rect 6802 61630 6804 61682
rect 6636 61236 6692 61246
rect 6636 60898 6692 61180
rect 6636 60846 6638 60898
rect 6690 60846 6692 60898
rect 6636 60834 6692 60846
rect 6748 60786 6804 61630
rect 7084 61236 7140 62412
rect 7420 62356 7476 62366
rect 7084 61170 7140 61180
rect 7196 62244 7252 62254
rect 7196 60898 7252 62188
rect 7196 60846 7198 60898
rect 7250 60846 7252 60898
rect 7196 60834 7252 60846
rect 6748 60734 6750 60786
rect 6802 60734 6804 60786
rect 6636 60116 6692 60126
rect 6524 58772 6580 58782
rect 6524 57874 6580 58716
rect 6524 57822 6526 57874
rect 6578 57822 6580 57874
rect 6524 56866 6580 57822
rect 6636 56980 6692 60060
rect 6748 60004 6804 60734
rect 7420 60788 7476 62300
rect 7532 60900 7588 60910
rect 7532 60806 7588 60844
rect 7868 60788 7924 62524
rect 7980 61012 8036 62862
rect 8316 62578 8372 62590
rect 8316 62526 8318 62578
rect 8370 62526 8372 62578
rect 8316 62244 8372 62526
rect 8204 61570 8260 61582
rect 8204 61518 8206 61570
rect 8258 61518 8260 61570
rect 7980 60956 8148 61012
rect 7980 60788 8036 60798
rect 7868 60786 8036 60788
rect 7868 60734 7982 60786
rect 8034 60734 8036 60786
rect 7868 60732 8036 60734
rect 7084 60004 7140 60014
rect 6748 59948 7084 60004
rect 7084 59910 7140 59948
rect 7420 58660 7476 60732
rect 7980 60722 8036 60732
rect 7756 60564 7812 60574
rect 8092 60564 8148 60956
rect 7756 60562 8148 60564
rect 7756 60510 7758 60562
rect 7810 60510 8148 60562
rect 7756 60508 8148 60510
rect 8204 60676 8260 61518
rect 8316 61348 8372 62188
rect 8316 61282 8372 61292
rect 7756 60498 7812 60508
rect 7420 58594 7476 58604
rect 7532 58436 7588 58446
rect 7084 58434 7588 58436
rect 7084 58382 7534 58434
rect 7586 58382 7588 58434
rect 7084 58380 7588 58382
rect 7084 57874 7140 58380
rect 7532 58370 7588 58380
rect 7868 58436 7924 60508
rect 8204 58436 8260 60620
rect 7868 58434 8036 58436
rect 7868 58382 7870 58434
rect 7922 58382 8036 58434
rect 7868 58380 8036 58382
rect 7868 58370 7924 58380
rect 7308 58266 7364 58278
rect 7084 57822 7086 57874
rect 7138 57822 7140 57874
rect 6860 57650 6916 57662
rect 6860 57598 6862 57650
rect 6914 57598 6916 57650
rect 6860 57316 6916 57598
rect 6972 57540 7028 57550
rect 6972 57446 7028 57484
rect 6860 57250 6916 57260
rect 7084 57204 7140 57822
rect 7196 58210 7252 58222
rect 7196 58158 7198 58210
rect 7250 58158 7252 58210
rect 7196 57876 7252 58158
rect 7308 58214 7310 58266
rect 7362 58214 7364 58266
rect 7308 58212 7364 58214
rect 7532 58212 7588 58222
rect 7308 58156 7532 58212
rect 7532 58146 7588 58156
rect 7308 57876 7364 57886
rect 7196 57874 7364 57876
rect 7196 57822 7310 57874
rect 7362 57822 7364 57874
rect 7196 57820 7364 57822
rect 7308 57810 7364 57820
rect 7980 57538 8036 58380
rect 7980 57486 7982 57538
rect 8034 57486 8036 57538
rect 7084 57138 7140 57148
rect 7868 57204 7924 57214
rect 7420 56980 7476 56990
rect 6636 56978 7700 56980
rect 6636 56926 7422 56978
rect 7474 56926 7700 56978
rect 6636 56924 7700 56926
rect 6524 56814 6526 56866
rect 6578 56814 6580 56866
rect 6524 56644 6580 56814
rect 6636 56756 6692 56766
rect 6636 56662 6692 56700
rect 6524 56578 6580 56588
rect 6636 56306 6692 56318
rect 6636 56254 6638 56306
rect 6690 56254 6692 56306
rect 6412 56028 6580 56084
rect 6188 55916 6468 55972
rect 6188 55300 6244 55310
rect 6188 55206 6244 55244
rect 6300 54628 6356 54638
rect 6300 54534 6356 54572
rect 6188 54516 6244 54526
rect 6188 54422 6244 54460
rect 6300 54292 6356 54302
rect 5516 52110 5518 52162
rect 5570 52110 5572 52162
rect 5180 52098 5236 52108
rect 4396 52052 4452 52062
rect 4844 52052 4900 52062
rect 4396 52050 4900 52052
rect 4396 51998 4398 52050
rect 4450 51998 4846 52050
rect 4898 51998 4900 52050
rect 4396 51996 4900 51998
rect 4396 51986 4452 51996
rect 4060 51650 4116 51660
rect 4732 51604 4788 51614
rect 4844 51604 4900 51996
rect 4956 52052 5012 52062
rect 4956 51958 5012 51996
rect 5292 51604 5348 51614
rect 4844 51602 5348 51604
rect 4844 51550 5294 51602
rect 5346 51550 5348 51602
rect 4844 51548 5348 51550
rect 4732 51510 4788 51548
rect 5292 51538 5348 51548
rect 4008 50988 5208 50998
rect 4064 50986 4112 50988
rect 4168 50986 4216 50988
rect 4076 50934 4112 50986
rect 4200 50934 4216 50986
rect 4064 50932 4112 50934
rect 4168 50932 4216 50934
rect 4272 50986 4320 50988
rect 4376 50986 4424 50988
rect 4480 50986 4528 50988
rect 4376 50934 4396 50986
rect 4480 50934 4520 50986
rect 4272 50932 4320 50934
rect 4376 50932 4424 50934
rect 4480 50932 4528 50934
rect 4584 50932 4632 50988
rect 4688 50986 4736 50988
rect 4792 50986 4840 50988
rect 4896 50986 4944 50988
rect 4696 50934 4736 50986
rect 4820 50934 4840 50986
rect 4688 50932 4736 50934
rect 4792 50932 4840 50934
rect 4896 50932 4944 50934
rect 5000 50986 5048 50988
rect 5104 50986 5152 50988
rect 5000 50934 5016 50986
rect 5104 50934 5140 50986
rect 5000 50932 5048 50934
rect 5104 50932 5152 50934
rect 4008 50922 5208 50932
rect 3836 50764 4564 50820
rect 3836 50596 3892 50606
rect 3724 50594 3892 50596
rect 3724 50542 3838 50594
rect 3890 50542 3892 50594
rect 3724 50540 3892 50542
rect 3836 50530 3892 50540
rect 4172 50594 4228 50606
rect 4172 50542 4174 50594
rect 4226 50542 4228 50594
rect 4172 50428 4228 50542
rect 3612 46340 3668 49868
rect 3836 50372 4228 50428
rect 4508 50482 4564 50764
rect 5516 50818 5572 52110
rect 5516 50766 5518 50818
rect 5570 50766 5572 50818
rect 5516 50754 5572 50766
rect 5628 53340 6020 53396
rect 6188 53620 6244 53630
rect 4508 50430 4510 50482
rect 4562 50430 4564 50482
rect 3836 48916 3892 50372
rect 4508 50036 4564 50430
rect 4956 50484 5012 50522
rect 4956 50418 5012 50428
rect 5628 50148 5684 53340
rect 5852 53172 5908 53182
rect 5852 52052 5908 53116
rect 6076 53060 6132 53098
rect 6076 52994 6132 53004
rect 5964 52836 6020 52846
rect 5964 52834 6132 52836
rect 5964 52782 5966 52834
rect 6018 52782 6132 52834
rect 5964 52780 6132 52782
rect 5964 52770 6020 52780
rect 6076 52162 6132 52780
rect 6188 52612 6244 53564
rect 6188 52546 6244 52556
rect 6076 52110 6078 52162
rect 6130 52110 6132 52162
rect 6076 52098 6132 52110
rect 5852 51986 5908 51996
rect 6188 51940 6244 51950
rect 6300 51940 6356 54236
rect 6244 51884 6356 51940
rect 6188 51604 6244 51884
rect 6076 51380 6132 51390
rect 5740 50818 5796 50830
rect 5740 50766 5742 50818
rect 5794 50766 5796 50818
rect 5740 50706 5796 50766
rect 5740 50654 5742 50706
rect 5794 50654 5796 50706
rect 5740 50642 5796 50654
rect 6076 50428 6132 51324
rect 6188 50706 6244 51548
rect 6188 50654 6190 50706
rect 6242 50654 6244 50706
rect 6188 50642 6244 50654
rect 6300 51716 6356 51726
rect 5964 50372 6132 50428
rect 5964 50260 6020 50372
rect 5964 50204 6244 50260
rect 5628 50092 6020 50148
rect 4508 49970 4564 49980
rect 5516 50036 5572 50046
rect 5572 49980 5908 50036
rect 5516 49942 5572 49980
rect 4008 49420 5208 49430
rect 4064 49418 4112 49420
rect 4168 49418 4216 49420
rect 4076 49366 4112 49418
rect 4200 49366 4216 49418
rect 4064 49364 4112 49366
rect 4168 49364 4216 49366
rect 4272 49418 4320 49420
rect 4376 49418 4424 49420
rect 4480 49418 4528 49420
rect 4376 49366 4396 49418
rect 4480 49366 4520 49418
rect 4272 49364 4320 49366
rect 4376 49364 4424 49366
rect 4480 49364 4528 49366
rect 4584 49364 4632 49420
rect 4688 49418 4736 49420
rect 4792 49418 4840 49420
rect 4896 49418 4944 49420
rect 4696 49366 4736 49418
rect 4820 49366 4840 49418
rect 4688 49364 4736 49366
rect 4792 49364 4840 49366
rect 4896 49364 4944 49366
rect 5000 49418 5048 49420
rect 5104 49418 5152 49420
rect 5000 49366 5016 49418
rect 5104 49366 5140 49418
rect 5000 49364 5048 49366
rect 5104 49364 5152 49366
rect 4008 49354 5208 49364
rect 3724 47348 3780 47358
rect 3836 47348 3892 48860
rect 5628 48916 5684 48926
rect 5628 48822 5684 48860
rect 5740 48804 5796 48814
rect 5740 48710 5796 48748
rect 5740 48356 5796 48366
rect 5292 48354 5796 48356
rect 5292 48302 5742 48354
rect 5794 48302 5796 48354
rect 5292 48300 5796 48302
rect 4620 48132 4676 48142
rect 4620 48038 4676 48076
rect 4008 47852 5208 47862
rect 4064 47850 4112 47852
rect 4168 47850 4216 47852
rect 4076 47798 4112 47850
rect 4200 47798 4216 47850
rect 4064 47796 4112 47798
rect 4168 47796 4216 47798
rect 4272 47850 4320 47852
rect 4376 47850 4424 47852
rect 4480 47850 4528 47852
rect 4376 47798 4396 47850
rect 4480 47798 4520 47850
rect 4272 47796 4320 47798
rect 4376 47796 4424 47798
rect 4480 47796 4528 47798
rect 4584 47796 4632 47852
rect 4688 47850 4736 47852
rect 4792 47850 4840 47852
rect 4896 47850 4944 47852
rect 4696 47798 4736 47850
rect 4820 47798 4840 47850
rect 4688 47796 4736 47798
rect 4792 47796 4840 47798
rect 4896 47796 4944 47798
rect 5000 47850 5048 47852
rect 5104 47850 5152 47852
rect 5000 47798 5016 47850
rect 5104 47798 5140 47850
rect 5000 47796 5048 47798
rect 5104 47796 5152 47798
rect 4008 47786 5208 47796
rect 4620 47460 4676 47470
rect 4844 47460 4900 47470
rect 5180 47460 5236 47470
rect 5292 47460 5348 48300
rect 5740 48290 5796 48300
rect 4620 47458 5124 47460
rect 4620 47406 4622 47458
rect 4674 47406 4846 47458
rect 4898 47406 5124 47458
rect 4620 47404 5124 47406
rect 4620 47394 4676 47404
rect 4844 47394 4900 47404
rect 4060 47348 4116 47358
rect 3836 47346 4116 47348
rect 3836 47294 4062 47346
rect 4114 47294 4116 47346
rect 3836 47292 4116 47294
rect 3724 47254 3780 47292
rect 4060 47282 4116 47292
rect 4956 47234 5012 47246
rect 4956 47182 4958 47234
rect 5010 47182 5012 47234
rect 4956 47124 5012 47182
rect 5068 47236 5124 47404
rect 5180 47458 5348 47460
rect 5180 47406 5182 47458
rect 5234 47406 5348 47458
rect 5180 47404 5348 47406
rect 5180 47394 5236 47404
rect 5852 47236 5908 49980
rect 5068 47180 5908 47236
rect 4956 47058 5012 47068
rect 4844 47012 4900 47022
rect 4844 46898 4900 46956
rect 5628 47012 5684 47022
rect 4844 46846 4846 46898
rect 4898 46846 4900 46898
rect 4844 46834 4900 46846
rect 5516 46900 5572 46910
rect 3836 46676 3892 46686
rect 3612 46284 3780 46340
rect 3500 42578 3556 42588
rect 3724 42420 3780 46284
rect 3836 46114 3892 46620
rect 4008 46284 5208 46294
rect 4064 46282 4112 46284
rect 4168 46282 4216 46284
rect 4076 46230 4112 46282
rect 4200 46230 4216 46282
rect 4064 46228 4112 46230
rect 4168 46228 4216 46230
rect 4272 46282 4320 46284
rect 4376 46282 4424 46284
rect 4480 46282 4528 46284
rect 4376 46230 4396 46282
rect 4480 46230 4520 46282
rect 4272 46228 4320 46230
rect 4376 46228 4424 46230
rect 4480 46228 4528 46230
rect 4584 46228 4632 46284
rect 4688 46282 4736 46284
rect 4792 46282 4840 46284
rect 4896 46282 4944 46284
rect 4696 46230 4736 46282
rect 4820 46230 4840 46282
rect 4688 46228 4736 46230
rect 4792 46228 4840 46230
rect 4896 46228 4944 46230
rect 5000 46282 5048 46284
rect 5104 46282 5152 46284
rect 5000 46230 5016 46282
rect 5104 46230 5140 46282
rect 5000 46228 5048 46230
rect 5104 46228 5152 46230
rect 4008 46218 5208 46228
rect 3836 46062 3838 46114
rect 3890 46062 3892 46114
rect 3836 46050 3892 46062
rect 4172 45890 4228 45902
rect 4172 45838 4174 45890
rect 4226 45838 4228 45890
rect 4172 45220 4228 45838
rect 4172 45154 4228 45164
rect 4396 45778 4452 45790
rect 4396 45726 4398 45778
rect 4450 45726 4452 45778
rect 4396 44884 4452 45726
rect 4956 45780 5012 45790
rect 4956 45686 5012 45724
rect 5516 45780 5572 46844
rect 5628 46004 5684 46956
rect 5740 46788 5796 47180
rect 5740 46694 5796 46732
rect 5852 46786 5908 46798
rect 5852 46734 5854 46786
rect 5906 46734 5908 46786
rect 5740 46004 5796 46014
rect 5628 46002 5796 46004
rect 5628 45950 5742 46002
rect 5794 45950 5796 46002
rect 5628 45948 5796 45950
rect 5516 45714 5572 45724
rect 5628 45220 5684 45230
rect 5628 45126 5684 45164
rect 4396 44818 4452 44828
rect 5292 44994 5348 45006
rect 5292 44942 5294 44994
rect 5346 44942 5348 44994
rect 5292 44884 5348 44942
rect 5740 44884 5796 45948
rect 5852 45444 5908 46734
rect 5964 46676 6020 50092
rect 6076 47346 6132 47358
rect 6076 47294 6078 47346
rect 6130 47294 6132 47346
rect 6076 46898 6132 47294
rect 6076 46846 6078 46898
rect 6130 46846 6132 46898
rect 6076 46834 6132 46846
rect 5964 46620 6132 46676
rect 5852 45378 5908 45388
rect 6076 44996 6132 46620
rect 6076 44930 6132 44940
rect 5964 44884 6020 44894
rect 5740 44828 5908 44884
rect 5292 44818 5348 44828
rect 4008 44716 5208 44726
rect 4064 44714 4112 44716
rect 4168 44714 4216 44716
rect 4076 44662 4112 44714
rect 4200 44662 4216 44714
rect 4064 44660 4112 44662
rect 4168 44660 4216 44662
rect 4272 44714 4320 44716
rect 4376 44714 4424 44716
rect 4480 44714 4528 44716
rect 4376 44662 4396 44714
rect 4480 44662 4520 44714
rect 4272 44660 4320 44662
rect 4376 44660 4424 44662
rect 4480 44660 4528 44662
rect 4584 44660 4632 44716
rect 4688 44714 4736 44716
rect 4792 44714 4840 44716
rect 4896 44714 4944 44716
rect 4696 44662 4736 44714
rect 4820 44662 4840 44714
rect 4688 44660 4736 44662
rect 4792 44660 4840 44662
rect 4896 44660 4944 44662
rect 5000 44714 5048 44716
rect 5104 44714 5152 44716
rect 5000 44662 5016 44714
rect 5104 44662 5140 44714
rect 5000 44660 5048 44662
rect 5104 44660 5152 44662
rect 4008 44650 5208 44660
rect 5852 44660 5908 44828
rect 5964 44790 6020 44828
rect 5852 44604 6132 44660
rect 4396 44548 4452 44558
rect 4172 44322 4228 44334
rect 4172 44270 4174 44322
rect 4226 44270 4228 44322
rect 3836 44100 3892 44110
rect 3836 44006 3892 44044
rect 4172 43428 4228 44270
rect 4396 44210 4452 44492
rect 4396 44158 4398 44210
rect 4450 44158 4452 44210
rect 4396 44146 4452 44158
rect 4956 44212 5012 44222
rect 4956 44118 5012 44156
rect 5292 44212 5348 44222
rect 4732 43876 4788 43886
rect 4732 43762 4788 43820
rect 4732 43710 4734 43762
rect 4786 43710 4788 43762
rect 4732 43698 4788 43710
rect 5292 43762 5348 44156
rect 6076 43876 6132 44604
rect 5292 43710 5294 43762
rect 5346 43710 5348 43762
rect 5292 43698 5348 43710
rect 5628 43764 5684 43774
rect 4172 43362 4228 43372
rect 5628 43650 5684 43708
rect 6076 43762 6132 43820
rect 6076 43710 6078 43762
rect 6130 43710 6132 43762
rect 6076 43698 6132 43710
rect 5628 43598 5630 43650
rect 5682 43598 5684 43650
rect 4008 43148 5208 43158
rect 4064 43146 4112 43148
rect 4168 43146 4216 43148
rect 4076 43094 4112 43146
rect 4200 43094 4216 43146
rect 4064 43092 4112 43094
rect 4168 43092 4216 43094
rect 4272 43146 4320 43148
rect 4376 43146 4424 43148
rect 4480 43146 4528 43148
rect 4376 43094 4396 43146
rect 4480 43094 4520 43146
rect 4272 43092 4320 43094
rect 4376 43092 4424 43094
rect 4480 43092 4528 43094
rect 4584 43092 4632 43148
rect 4688 43146 4736 43148
rect 4792 43146 4840 43148
rect 4896 43146 4944 43148
rect 4696 43094 4736 43146
rect 4820 43094 4840 43146
rect 4688 43092 4736 43094
rect 4792 43092 4840 43094
rect 4896 43092 4944 43094
rect 5000 43146 5048 43148
rect 5104 43146 5152 43148
rect 5000 43094 5016 43146
rect 5104 43094 5140 43146
rect 5000 43092 5048 43094
rect 5104 43092 5152 43094
rect 4008 43082 5208 43092
rect 3500 42364 3780 42420
rect 5068 42868 5124 42878
rect 5068 42530 5124 42812
rect 5068 42478 5070 42530
rect 5122 42478 5124 42530
rect 3500 39396 3556 42364
rect 5068 41748 5124 42478
rect 5068 41692 5460 41748
rect 4008 41580 5208 41590
rect 4064 41578 4112 41580
rect 4168 41578 4216 41580
rect 4076 41526 4112 41578
rect 4200 41526 4216 41578
rect 4064 41524 4112 41526
rect 4168 41524 4216 41526
rect 4272 41578 4320 41580
rect 4376 41578 4424 41580
rect 4480 41578 4528 41580
rect 4376 41526 4396 41578
rect 4480 41526 4520 41578
rect 4272 41524 4320 41526
rect 4376 41524 4424 41526
rect 4480 41524 4528 41526
rect 4584 41524 4632 41580
rect 4688 41578 4736 41580
rect 4792 41578 4840 41580
rect 4896 41578 4944 41580
rect 4696 41526 4736 41578
rect 4820 41526 4840 41578
rect 4688 41524 4736 41526
rect 4792 41524 4840 41526
rect 4896 41524 4944 41526
rect 5000 41578 5048 41580
rect 5104 41578 5152 41580
rect 5000 41526 5016 41578
rect 5104 41526 5140 41578
rect 5000 41524 5048 41526
rect 5104 41524 5152 41526
rect 4008 41514 5208 41524
rect 5292 40964 5348 40974
rect 4732 40740 4788 40750
rect 4732 40626 4788 40684
rect 4732 40574 4734 40626
rect 4786 40574 4788 40626
rect 4732 40562 4788 40574
rect 5292 40626 5348 40908
rect 5292 40574 5294 40626
rect 5346 40574 5348 40626
rect 3948 40516 4004 40526
rect 3836 40460 3948 40516
rect 3724 39844 3780 39854
rect 3836 39844 3892 40460
rect 3948 40450 4004 40460
rect 4008 40012 5208 40022
rect 4064 40010 4112 40012
rect 4168 40010 4216 40012
rect 4076 39958 4112 40010
rect 4200 39958 4216 40010
rect 4064 39956 4112 39958
rect 4168 39956 4216 39958
rect 4272 40010 4320 40012
rect 4376 40010 4424 40012
rect 4480 40010 4528 40012
rect 4376 39958 4396 40010
rect 4480 39958 4520 40010
rect 4272 39956 4320 39958
rect 4376 39956 4424 39958
rect 4480 39956 4528 39958
rect 4584 39956 4632 40012
rect 4688 40010 4736 40012
rect 4792 40010 4840 40012
rect 4896 40010 4944 40012
rect 4696 39958 4736 40010
rect 4820 39958 4840 40010
rect 4688 39956 4736 39958
rect 4792 39956 4840 39958
rect 4896 39956 4944 39958
rect 5000 40010 5048 40012
rect 5104 40010 5152 40012
rect 5000 39958 5016 40010
rect 5104 39958 5140 40010
rect 5000 39956 5048 39958
rect 5104 39956 5152 39958
rect 4008 39946 5208 39956
rect 4060 39844 4116 39854
rect 5292 39844 5348 40574
rect 3836 39842 4116 39844
rect 3836 39790 4062 39842
rect 4114 39790 4116 39842
rect 3836 39788 4116 39790
rect 3724 39750 3780 39788
rect 4060 39778 4116 39788
rect 4844 39788 5348 39844
rect 4284 39620 4340 39630
rect 4284 39506 4340 39564
rect 4284 39454 4286 39506
rect 4338 39454 4340 39506
rect 4284 39442 4340 39454
rect 4844 39506 4900 39788
rect 4844 39454 4846 39506
rect 4898 39454 4900 39506
rect 4844 39442 4900 39454
rect 3500 39340 3668 39396
rect 2492 38164 2548 38668
rect 3388 38612 3556 38668
rect 2492 38098 2548 38108
rect 3164 37380 3220 37390
rect 3164 37286 3220 37324
rect 2828 37266 2884 37278
rect 2828 37214 2830 37266
rect 2882 37214 2884 37266
rect 2492 37156 2548 37166
rect 2828 37156 2884 37214
rect 2492 37154 2884 37156
rect 2492 37102 2494 37154
rect 2546 37102 2884 37154
rect 2492 37100 2884 37102
rect 2492 37044 2548 37100
rect 2492 36978 2548 36988
rect 2604 36260 2660 36270
rect 2828 36260 2884 36270
rect 2604 36258 2884 36260
rect 2604 36206 2606 36258
rect 2658 36206 2830 36258
rect 2882 36206 2884 36258
rect 2604 36204 2884 36206
rect 2492 35924 2548 35934
rect 2380 35700 2436 35710
rect 1820 35646 1822 35698
rect 1874 35646 1876 35698
rect 1820 34130 1876 35646
rect 2156 35698 2436 35700
rect 2156 35646 2382 35698
rect 2434 35646 2436 35698
rect 2156 35644 2436 35646
rect 2156 35138 2212 35644
rect 2380 35634 2436 35644
rect 2492 35140 2548 35868
rect 2156 35086 2158 35138
rect 2210 35086 2212 35138
rect 2156 35074 2212 35086
rect 2380 35084 2548 35140
rect 1820 34078 1822 34130
rect 1874 34078 1876 34130
rect 1820 32788 1876 34078
rect 2268 34692 2324 34702
rect 2268 34130 2324 34636
rect 2268 34078 2270 34130
rect 2322 34078 2324 34130
rect 2268 34066 2324 34078
rect 2380 33236 2436 35084
rect 2492 34914 2548 34926
rect 2492 34862 2494 34914
rect 2546 34862 2548 34914
rect 2492 33460 2548 34862
rect 2604 34804 2660 36204
rect 2828 36194 2884 36204
rect 3164 36258 3220 36270
rect 3164 36206 3166 36258
rect 3218 36206 3220 36258
rect 3164 35476 3220 36206
rect 3164 35410 3220 35420
rect 3052 35140 3108 35150
rect 3052 34914 3108 35084
rect 3052 34862 3054 34914
rect 3106 34862 3108 34914
rect 3052 34850 3108 34862
rect 2604 34738 2660 34748
rect 3276 34802 3332 34814
rect 3276 34750 3278 34802
rect 3330 34750 3332 34802
rect 3276 34244 3332 34750
rect 3276 34178 3332 34188
rect 2492 33394 2548 33404
rect 2492 33236 2548 33246
rect 2828 33236 2884 33246
rect 2380 33234 2884 33236
rect 2380 33182 2494 33234
rect 2546 33182 2830 33234
rect 2882 33182 2884 33234
rect 2380 33180 2884 33182
rect 2492 33170 2548 33180
rect 2828 33170 2884 33180
rect 3164 33236 3220 33246
rect 3164 33142 3220 33180
rect 1820 29426 1876 32732
rect 3500 31892 3556 38612
rect 3612 32116 3668 39340
rect 5404 38948 5460 41692
rect 5628 39732 5684 43598
rect 5740 43428 5796 43438
rect 5740 42978 5796 43372
rect 5740 42926 5742 42978
rect 5794 42926 5796 42978
rect 5740 42914 5796 42926
rect 6076 42868 6132 42878
rect 6076 42774 6132 42812
rect 6188 41076 6244 50204
rect 6300 47570 6356 51660
rect 6412 48466 6468 55916
rect 6524 54740 6580 56028
rect 6636 55076 6692 56254
rect 6636 55010 6692 55020
rect 6748 54740 6804 56924
rect 7420 56914 7476 56924
rect 7644 56866 7700 56924
rect 7644 56814 7646 56866
rect 7698 56814 7700 56866
rect 7644 56802 7700 56814
rect 7532 56644 7588 56654
rect 7196 55860 7252 55870
rect 7084 55858 7252 55860
rect 7084 55806 7198 55858
rect 7250 55806 7252 55858
rect 7084 55804 7252 55806
rect 7084 55188 7140 55804
rect 7196 55794 7252 55804
rect 7196 55524 7252 55534
rect 7196 55430 7252 55468
rect 7308 55188 7364 55198
rect 7140 55186 7364 55188
rect 7140 55134 7310 55186
rect 7362 55134 7364 55186
rect 7140 55132 7364 55134
rect 7084 55094 7140 55132
rect 6860 55076 6916 55086
rect 6860 54982 6916 55020
rect 6524 54684 6692 54740
rect 6524 54514 6580 54526
rect 6524 54462 6526 54514
rect 6578 54462 6580 54514
rect 6524 54404 6580 54462
rect 6524 54338 6580 54348
rect 6524 53172 6580 53182
rect 6524 53078 6580 53116
rect 6636 51380 6692 54684
rect 6748 54674 6804 54684
rect 7196 54628 7252 54638
rect 6748 54514 6804 54526
rect 7084 54516 7140 54526
rect 6748 54462 6750 54514
rect 6802 54462 6804 54514
rect 6748 54404 6804 54462
rect 6972 54514 7140 54516
rect 6972 54462 7086 54514
rect 7138 54462 7140 54514
rect 6972 54460 7140 54462
rect 6972 54404 7028 54460
rect 7084 54450 7140 54460
rect 7196 54514 7252 54572
rect 7196 54462 7198 54514
rect 7250 54462 7252 54514
rect 6748 54348 7028 54404
rect 7196 54404 7252 54462
rect 7308 54404 7364 55132
rect 7420 54404 7476 54414
rect 7308 54348 7420 54404
rect 7196 54292 7252 54348
rect 7420 54310 7476 54348
rect 6636 51314 6692 51324
rect 6972 54236 7252 54292
rect 6972 53842 7028 54236
rect 6972 53790 6974 53842
rect 7026 53790 7028 53842
rect 6636 50820 6692 50830
rect 6636 50818 6916 50820
rect 6636 50766 6638 50818
rect 6690 50766 6916 50818
rect 6636 50764 6916 50766
rect 6636 50754 6692 50764
rect 6748 50596 6804 50606
rect 6636 50484 6692 50522
rect 6636 50418 6692 50428
rect 6412 48414 6414 48466
rect 6466 48414 6468 48466
rect 6412 48402 6468 48414
rect 6300 47518 6302 47570
rect 6354 47518 6356 47570
rect 6300 47506 6356 47518
rect 6412 46788 6468 46798
rect 6412 45108 6468 46732
rect 6300 45106 6468 45108
rect 6300 45054 6414 45106
rect 6466 45054 6468 45106
rect 6300 45052 6468 45054
rect 6300 42868 6356 45052
rect 6412 45042 6468 45052
rect 6524 45666 6580 45678
rect 6524 45614 6526 45666
rect 6578 45614 6580 45666
rect 6524 45218 6580 45614
rect 6524 45166 6526 45218
rect 6578 45166 6580 45218
rect 6412 44212 6468 44222
rect 6412 44118 6468 44156
rect 6524 44100 6580 45166
rect 6748 44660 6804 50540
rect 6860 49026 6916 50764
rect 6972 50484 7028 53790
rect 6972 50418 7028 50428
rect 7308 53172 7364 53182
rect 7308 51490 7364 53116
rect 7308 51438 7310 51490
rect 7362 51438 7364 51490
rect 7308 50484 7364 51438
rect 7308 50418 7364 50428
rect 7532 50148 7588 56588
rect 7756 56084 7812 56094
rect 7756 55990 7812 56028
rect 7868 55970 7924 57148
rect 7868 55918 7870 55970
rect 7922 55918 7924 55970
rect 7868 55524 7924 55918
rect 7868 55458 7924 55468
rect 7980 57092 8036 57486
rect 7980 55298 8036 57036
rect 7980 55246 7982 55298
rect 8034 55246 8036 55298
rect 7980 55234 8036 55246
rect 8092 58380 8260 58436
rect 8092 55076 8148 58380
rect 8204 58212 8260 58222
rect 8260 58156 8372 58212
rect 8204 58118 8260 58156
rect 8316 57540 8372 58156
rect 8428 57876 8484 64316
rect 8540 64148 8596 64158
rect 8540 63138 8596 64092
rect 8540 63086 8542 63138
rect 8594 63086 8596 63138
rect 8540 63074 8596 63086
rect 8540 60788 8596 60798
rect 8540 60694 8596 60732
rect 8540 57876 8596 57886
rect 8428 57874 8596 57876
rect 8428 57822 8542 57874
rect 8594 57822 8596 57874
rect 8428 57820 8596 57822
rect 8316 57484 8484 57540
rect 8204 57428 8260 57438
rect 8204 57426 8372 57428
rect 8204 57374 8206 57426
rect 8258 57374 8372 57426
rect 8204 57372 8372 57374
rect 8204 57362 8260 57372
rect 8204 57204 8260 57214
rect 8204 56866 8260 57148
rect 8204 56814 8206 56866
rect 8258 56814 8260 56866
rect 8204 56802 8260 56814
rect 8316 56194 8372 57372
rect 8316 56142 8318 56194
rect 8370 56142 8372 56194
rect 7980 55020 8148 55076
rect 8204 55412 8260 55422
rect 7868 54740 7924 54750
rect 7644 54516 7700 54526
rect 7644 54422 7700 54460
rect 7868 53732 7924 54684
rect 7868 53638 7924 53676
rect 7980 50596 8036 55020
rect 8092 54740 8148 54750
rect 8204 54740 8260 55356
rect 8316 55188 8372 56142
rect 8428 56084 8484 57484
rect 8428 56018 8484 56028
rect 8540 55858 8596 57820
rect 8540 55806 8542 55858
rect 8594 55806 8596 55858
rect 8540 55794 8596 55806
rect 8540 55410 8596 55422
rect 8540 55358 8542 55410
rect 8594 55358 8596 55410
rect 8428 55188 8484 55198
rect 8316 55186 8484 55188
rect 8316 55134 8430 55186
rect 8482 55134 8484 55186
rect 8316 55132 8484 55134
rect 8428 55122 8484 55132
rect 8092 54738 8260 54740
rect 8092 54686 8094 54738
rect 8146 54686 8260 54738
rect 8092 54684 8260 54686
rect 8092 54628 8148 54684
rect 8092 54562 8148 54572
rect 8540 54292 8596 55358
rect 8428 54236 8596 54292
rect 8428 51604 8484 54236
rect 8540 54068 8596 54078
rect 8540 53730 8596 54012
rect 8540 53678 8542 53730
rect 8594 53678 8596 53730
rect 8540 53666 8596 53678
rect 8540 51940 8596 51950
rect 8540 51846 8596 51884
rect 8316 51548 8484 51604
rect 8316 50820 8372 51548
rect 8540 51380 8596 51390
rect 8540 51286 8596 51324
rect 8316 50764 8596 50820
rect 8316 50708 8372 50764
rect 7980 50530 8036 50540
rect 8204 50706 8372 50708
rect 8204 50654 8318 50706
rect 8370 50654 8372 50706
rect 8204 50652 8372 50654
rect 8204 50428 8260 50652
rect 8316 50642 8372 50652
rect 7868 50372 8260 50428
rect 8316 50484 8372 50494
rect 8372 50428 8484 50484
rect 8316 50418 8372 50428
rect 7308 50092 7812 50148
rect 7308 50034 7364 50092
rect 7308 49982 7310 50034
rect 7362 49982 7364 50034
rect 7308 49970 7364 49982
rect 7756 49922 7812 50092
rect 7756 49870 7758 49922
rect 7810 49870 7812 49922
rect 7532 49812 7588 49822
rect 7420 49810 7588 49812
rect 7420 49758 7534 49810
rect 7586 49758 7588 49810
rect 7420 49756 7588 49758
rect 7420 49252 7476 49756
rect 7532 49746 7588 49756
rect 6860 48974 6862 49026
rect 6914 48974 6916 49026
rect 6860 48468 6916 48974
rect 6860 48402 6916 48412
rect 7196 49196 7476 49252
rect 7644 49588 7700 49598
rect 7196 48356 7252 49196
rect 7308 49026 7364 49038
rect 7308 48974 7310 49026
rect 7362 48974 7364 49026
rect 7308 48468 7364 48974
rect 7532 48468 7588 48478
rect 7308 48466 7588 48468
rect 7308 48414 7534 48466
rect 7586 48414 7588 48466
rect 7308 48412 7588 48414
rect 7532 48402 7588 48412
rect 7644 48466 7700 49532
rect 7756 48580 7812 49870
rect 7868 49922 7924 50372
rect 7868 49870 7870 49922
rect 7922 49870 7924 49922
rect 7868 49858 7924 49870
rect 7756 48524 8036 48580
rect 7644 48414 7646 48466
rect 7698 48414 7700 48466
rect 7644 48402 7700 48414
rect 7868 48356 7924 48366
rect 7196 48300 7476 48356
rect 6972 48242 7028 48254
rect 6972 48190 6974 48242
rect 7026 48190 7028 48242
rect 6972 47460 7028 48190
rect 7420 48242 7476 48300
rect 7420 48190 7422 48242
rect 7474 48190 7476 48242
rect 7420 48178 7476 48190
rect 7756 48354 7924 48356
rect 7756 48302 7870 48354
rect 7922 48302 7924 48354
rect 7756 48300 7924 48302
rect 7084 47460 7140 47470
rect 6972 47458 7140 47460
rect 6972 47406 7086 47458
rect 7138 47406 7140 47458
rect 6972 47404 7140 47406
rect 7084 47236 7140 47404
rect 7756 47458 7812 48300
rect 7868 48290 7924 48300
rect 7980 48132 8036 48524
rect 8428 48468 8484 50428
rect 8540 49812 8596 50764
rect 8652 50428 8708 72268
rect 8988 70084 9044 70094
rect 8988 69990 9044 70028
rect 8764 68066 8820 68078
rect 8764 68014 8766 68066
rect 8818 68014 8820 68066
rect 8764 67956 8820 68014
rect 8764 67954 9268 67956
rect 8764 67902 8766 67954
rect 8818 67902 9268 67954
rect 8764 67900 9268 67902
rect 8764 67890 8820 67900
rect 9100 67284 9156 67294
rect 9100 67058 9156 67228
rect 9100 67006 9102 67058
rect 9154 67006 9156 67058
rect 9100 66994 9156 67006
rect 8764 66836 8820 66846
rect 8764 66498 8820 66780
rect 8764 66446 8766 66498
rect 8818 66446 8820 66498
rect 8764 66434 8820 66446
rect 9212 66388 9268 67900
rect 8988 66386 9268 66388
rect 8988 66334 9214 66386
rect 9266 66334 9268 66386
rect 8988 66332 9268 66334
rect 8988 65268 9044 66332
rect 9212 66322 9268 66332
rect 9324 65492 9380 76636
rect 9660 75796 9716 76860
rect 9772 76692 9828 76702
rect 9772 76598 9828 76636
rect 10220 76356 10276 76366
rect 9436 75794 9716 75796
rect 9436 75742 9662 75794
rect 9714 75742 9716 75794
rect 9436 75740 9716 75742
rect 9436 74228 9492 75740
rect 9660 75730 9716 75740
rect 10108 76354 10276 76356
rect 10108 76302 10222 76354
rect 10274 76302 10276 76354
rect 10108 76300 10276 76302
rect 10332 76356 10388 78876
rect 10444 77140 10500 79436
rect 10556 79426 10612 79436
rect 10780 79268 10836 79278
rect 10668 78594 10724 78606
rect 10668 78542 10670 78594
rect 10722 78542 10724 78594
rect 10556 78036 10612 78046
rect 10556 77942 10612 77980
rect 10668 77924 10724 78542
rect 10668 77858 10724 77868
rect 10556 77140 10612 77150
rect 10444 77138 10612 77140
rect 10444 77086 10558 77138
rect 10610 77086 10612 77138
rect 10444 77084 10612 77086
rect 10556 77074 10612 77084
rect 10668 76356 10724 76366
rect 10332 76300 10668 76356
rect 10108 75236 10164 76300
rect 10220 76290 10276 76300
rect 10668 76262 10724 76300
rect 9436 72660 9492 74172
rect 9884 75180 10164 75236
rect 10780 75348 10836 79212
rect 10892 79156 10948 80668
rect 11004 79604 11060 80780
rect 11004 79510 11060 79548
rect 10892 79090 10948 79100
rect 11116 79044 11172 80894
rect 11228 80946 11284 80958
rect 11228 80894 11230 80946
rect 11282 80894 11284 80946
rect 11228 80274 11284 80894
rect 11788 80836 11844 81902
rect 11900 81170 11956 82124
rect 12124 81954 12180 83694
rect 12460 83522 12516 86156
rect 13132 85540 13188 88172
rect 13244 88162 13300 88172
rect 13580 88004 13636 88014
rect 13580 87910 13636 87948
rect 13580 86660 13636 86670
rect 13580 86566 13636 86604
rect 13580 86212 13636 86222
rect 13580 86098 13636 86156
rect 13580 86046 13582 86098
rect 13634 86046 13636 86098
rect 12684 85484 13188 85540
rect 13468 85876 13524 85886
rect 12572 84866 12628 84878
rect 12572 84814 12574 84866
rect 12626 84814 12628 84866
rect 12572 84308 12628 84814
rect 12684 84530 12740 85484
rect 12684 84478 12686 84530
rect 12738 84478 12740 84530
rect 12684 84466 12740 84478
rect 13020 84868 13076 84878
rect 12572 84214 12628 84252
rect 12796 84306 12852 84318
rect 12796 84254 12798 84306
rect 12850 84254 12852 84306
rect 12460 83470 12462 83522
rect 12514 83470 12516 83522
rect 12460 83458 12516 83470
rect 12572 83634 12628 83646
rect 12572 83582 12574 83634
rect 12626 83582 12628 83634
rect 12572 82964 12628 83582
rect 12572 82898 12628 82908
rect 12796 82964 12852 84254
rect 13020 84308 13076 84812
rect 13356 84418 13412 84430
rect 13356 84366 13358 84418
rect 13410 84366 13412 84418
rect 13020 84242 13076 84252
rect 13244 84308 13300 84318
rect 13356 84308 13412 84366
rect 13244 84306 13412 84308
rect 13244 84254 13246 84306
rect 13298 84254 13412 84306
rect 13244 84252 13412 84254
rect 13244 84242 13300 84252
rect 13468 83524 13524 85820
rect 13580 85764 13636 86046
rect 13580 85698 13636 85708
rect 13692 85540 13748 88396
rect 13916 88228 13972 88238
rect 13916 88134 13972 88172
rect 14140 88114 14196 88396
rect 14140 88062 14142 88114
rect 14194 88062 14196 88114
rect 14140 88050 14196 88062
rect 14252 88004 14308 88844
rect 24008 88620 25208 88630
rect 24064 88618 24112 88620
rect 24168 88618 24216 88620
rect 24076 88566 24112 88618
rect 24200 88566 24216 88618
rect 24064 88564 24112 88566
rect 24168 88564 24216 88566
rect 24272 88618 24320 88620
rect 24376 88618 24424 88620
rect 24480 88618 24528 88620
rect 24376 88566 24396 88618
rect 24480 88566 24520 88618
rect 24272 88564 24320 88566
rect 24376 88564 24424 88566
rect 24480 88564 24528 88566
rect 24584 88564 24632 88620
rect 24688 88618 24736 88620
rect 24792 88618 24840 88620
rect 24896 88618 24944 88620
rect 24696 88566 24736 88618
rect 24820 88566 24840 88618
rect 24688 88564 24736 88566
rect 24792 88564 24840 88566
rect 24896 88564 24944 88566
rect 25000 88618 25048 88620
rect 25104 88618 25152 88620
rect 25000 88566 25016 88618
rect 25104 88566 25140 88618
rect 25000 88564 25048 88566
rect 25104 88564 25152 88566
rect 24008 88554 25208 88564
rect 14700 88116 14756 88126
rect 14700 88022 14756 88060
rect 15596 88116 15652 88126
rect 14252 87938 14308 87948
rect 14008 87836 15208 87846
rect 14064 87834 14112 87836
rect 14168 87834 14216 87836
rect 14076 87782 14112 87834
rect 14200 87782 14216 87834
rect 14064 87780 14112 87782
rect 14168 87780 14216 87782
rect 14272 87834 14320 87836
rect 14376 87834 14424 87836
rect 14480 87834 14528 87836
rect 14376 87782 14396 87834
rect 14480 87782 14520 87834
rect 14272 87780 14320 87782
rect 14376 87780 14424 87782
rect 14480 87780 14528 87782
rect 14584 87780 14632 87836
rect 14688 87834 14736 87836
rect 14792 87834 14840 87836
rect 14896 87834 14944 87836
rect 14696 87782 14736 87834
rect 14820 87782 14840 87834
rect 14688 87780 14736 87782
rect 14792 87780 14840 87782
rect 14896 87780 14944 87782
rect 15000 87834 15048 87836
rect 15104 87834 15152 87836
rect 15000 87782 15016 87834
rect 15104 87782 15140 87834
rect 15000 87780 15048 87782
rect 15104 87780 15152 87782
rect 14008 87770 15208 87780
rect 15372 87780 15428 87790
rect 15036 87668 15092 87678
rect 15372 87668 15428 87724
rect 15036 87666 15428 87668
rect 15036 87614 15038 87666
rect 15090 87614 15428 87666
rect 15036 87612 15428 87614
rect 15036 87602 15092 87612
rect 15596 87218 15652 88060
rect 17276 88004 17332 88014
rect 16380 87668 16436 87678
rect 16380 87574 16436 87612
rect 16716 87668 16772 87678
rect 15596 87166 15598 87218
rect 15650 87166 15652 87218
rect 14364 86660 14420 86670
rect 14364 86566 14420 86604
rect 15036 86660 15092 86670
rect 15036 86658 15428 86660
rect 15036 86606 15038 86658
rect 15090 86606 15428 86658
rect 15036 86604 15428 86606
rect 15036 86594 15092 86604
rect 14028 86548 14084 86558
rect 13692 85204 13748 85484
rect 13692 85138 13748 85148
rect 13804 86546 14084 86548
rect 13804 86494 14030 86546
rect 14082 86494 14084 86546
rect 13804 86492 14084 86494
rect 13692 84868 13748 84878
rect 13580 84866 13748 84868
rect 13580 84814 13694 84866
rect 13746 84814 13748 84866
rect 13580 84812 13748 84814
rect 13580 84418 13636 84812
rect 13692 84802 13748 84812
rect 13580 84366 13582 84418
rect 13634 84366 13636 84418
rect 13580 84084 13636 84366
rect 13692 84308 13748 84318
rect 13692 84214 13748 84252
rect 13580 84018 13636 84028
rect 13468 83430 13524 83468
rect 13692 83188 13748 83198
rect 12908 82964 12964 82974
rect 12796 82962 12964 82964
rect 12796 82910 12910 82962
rect 12962 82910 12964 82962
rect 12796 82908 12964 82910
rect 12796 82740 12852 82908
rect 12908 82898 12964 82908
rect 13020 82852 13076 82862
rect 13580 82852 13636 82862
rect 13020 82758 13076 82796
rect 13468 82850 13636 82852
rect 13468 82798 13582 82850
rect 13634 82798 13636 82850
rect 13468 82796 13636 82798
rect 12796 82674 12852 82684
rect 12572 82628 12628 82638
rect 12572 82534 12628 82572
rect 13356 82628 13412 82638
rect 13356 82534 13412 82572
rect 12124 81902 12126 81954
rect 12178 81902 12180 81954
rect 12124 81890 12180 81902
rect 12348 82068 12404 82078
rect 12348 81842 12404 82012
rect 12348 81790 12350 81842
rect 12402 81790 12404 81842
rect 12348 81778 12404 81790
rect 13468 81844 13524 82796
rect 13580 82786 13636 82796
rect 13692 82626 13748 83132
rect 13692 82574 13694 82626
rect 13746 82574 13748 82626
rect 13692 82562 13748 82574
rect 13804 82068 13860 86492
rect 14028 86482 14084 86492
rect 14008 86268 15208 86278
rect 14064 86266 14112 86268
rect 14168 86266 14216 86268
rect 14076 86214 14112 86266
rect 14200 86214 14216 86266
rect 14064 86212 14112 86214
rect 14168 86212 14216 86214
rect 14272 86266 14320 86268
rect 14376 86266 14424 86268
rect 14480 86266 14528 86268
rect 14376 86214 14396 86266
rect 14480 86214 14520 86266
rect 14272 86212 14320 86214
rect 14376 86212 14424 86214
rect 14480 86212 14528 86214
rect 14584 86212 14632 86268
rect 14688 86266 14736 86268
rect 14792 86266 14840 86268
rect 14896 86266 14944 86268
rect 14696 86214 14736 86266
rect 14820 86214 14840 86266
rect 14688 86212 14736 86214
rect 14792 86212 14840 86214
rect 14896 86212 14944 86214
rect 15000 86266 15048 86268
rect 15104 86266 15152 86268
rect 15000 86214 15016 86266
rect 15104 86214 15140 86266
rect 15000 86212 15048 86214
rect 15104 86212 15152 86214
rect 14008 86202 15208 86212
rect 15372 86098 15428 86604
rect 15372 86046 15374 86098
rect 15426 86046 15428 86098
rect 15372 86034 15428 86046
rect 14140 85876 14196 85886
rect 14140 85782 14196 85820
rect 14476 85876 14532 85886
rect 14252 85764 14308 85774
rect 14476 85708 14532 85820
rect 15036 85876 15092 85886
rect 14252 85204 14308 85708
rect 14252 85090 14308 85148
rect 14364 85652 14532 85708
rect 14812 85764 14868 85802
rect 15036 85782 15092 85820
rect 15372 85874 15428 85886
rect 15372 85822 15374 85874
rect 15426 85822 15428 85874
rect 14364 85202 14420 85652
rect 14812 85540 14868 85708
rect 15372 85764 15428 85822
rect 15372 85698 15428 85708
rect 14812 85474 14868 85484
rect 14364 85150 14366 85202
rect 14418 85150 14420 85202
rect 14364 85138 14420 85150
rect 14252 85038 14254 85090
rect 14306 85038 14308 85090
rect 14252 85026 14308 85038
rect 13916 84980 13972 84990
rect 13916 84886 13972 84924
rect 14476 84978 14532 84990
rect 14476 84926 14478 84978
rect 14530 84926 14532 84978
rect 14476 84868 14532 84926
rect 14476 84802 14532 84812
rect 14008 84700 15208 84710
rect 14064 84698 14112 84700
rect 14168 84698 14216 84700
rect 14076 84646 14112 84698
rect 14200 84646 14216 84698
rect 14064 84644 14112 84646
rect 14168 84644 14216 84646
rect 14272 84698 14320 84700
rect 14376 84698 14424 84700
rect 14480 84698 14528 84700
rect 14376 84646 14396 84698
rect 14480 84646 14520 84698
rect 14272 84644 14320 84646
rect 14376 84644 14424 84646
rect 14480 84644 14528 84646
rect 14584 84644 14632 84700
rect 14688 84698 14736 84700
rect 14792 84698 14840 84700
rect 14896 84698 14944 84700
rect 14696 84646 14736 84698
rect 14820 84646 14840 84698
rect 14688 84644 14736 84646
rect 14792 84644 14840 84646
rect 14896 84644 14944 84646
rect 15000 84698 15048 84700
rect 15104 84698 15152 84700
rect 15000 84646 15016 84698
rect 15104 84646 15140 84698
rect 15000 84644 15048 84646
rect 15104 84644 15152 84646
rect 14008 84634 15208 84644
rect 14588 84532 14644 84542
rect 14476 84420 14532 84430
rect 14476 84326 14532 84364
rect 14588 84418 14644 84476
rect 15596 84532 15652 87166
rect 16044 87330 16100 87342
rect 16044 87278 16046 87330
rect 16098 87278 16100 87330
rect 16044 87218 16100 87278
rect 16044 87166 16046 87218
rect 16098 87166 16100 87218
rect 16044 86660 16100 87166
rect 16044 86594 16100 86604
rect 15708 85988 15764 85998
rect 16604 85988 16660 85998
rect 15708 85986 16548 85988
rect 15708 85934 15710 85986
rect 15762 85934 16548 85986
rect 15708 85932 16548 85934
rect 15708 85922 15764 85932
rect 16156 85764 16212 85774
rect 16156 85670 16212 85708
rect 16492 85762 16548 85932
rect 16492 85710 16494 85762
rect 16546 85710 16548 85762
rect 16492 85698 16548 85710
rect 15596 84466 15652 84476
rect 14588 84366 14590 84418
rect 14642 84366 14644 84418
rect 14588 84354 14644 84366
rect 15036 84420 15092 84430
rect 15036 84196 15092 84364
rect 16492 84196 16548 84206
rect 15036 84140 15540 84196
rect 14476 84082 14532 84094
rect 14476 84030 14478 84082
rect 14530 84030 14532 84082
rect 14028 83522 14084 83534
rect 14028 83470 14030 83522
rect 14082 83470 14084 83522
rect 14028 83300 14084 83470
rect 14476 83412 14532 84030
rect 14476 83346 14532 83356
rect 15260 83412 15316 83422
rect 15316 83356 15428 83412
rect 15260 83346 15316 83356
rect 14028 83234 14084 83244
rect 14008 83132 15208 83142
rect 14064 83130 14112 83132
rect 14168 83130 14216 83132
rect 14076 83078 14112 83130
rect 14200 83078 14216 83130
rect 14064 83076 14112 83078
rect 14168 83076 14216 83078
rect 14272 83130 14320 83132
rect 14376 83130 14424 83132
rect 14480 83130 14528 83132
rect 14376 83078 14396 83130
rect 14480 83078 14520 83130
rect 14272 83076 14320 83078
rect 14376 83076 14424 83078
rect 14480 83076 14528 83078
rect 14584 83076 14632 83132
rect 14688 83130 14736 83132
rect 14792 83130 14840 83132
rect 14896 83130 14944 83132
rect 14696 83078 14736 83130
rect 14820 83078 14840 83130
rect 14688 83076 14736 83078
rect 14792 83076 14840 83078
rect 14896 83076 14944 83078
rect 15000 83130 15048 83132
rect 15104 83130 15152 83132
rect 15000 83078 15016 83130
rect 15104 83078 15140 83130
rect 15000 83076 15048 83078
rect 15104 83076 15152 83078
rect 14008 83066 15208 83076
rect 15148 82964 15204 82974
rect 14364 82850 14420 82862
rect 14364 82798 14366 82850
rect 14418 82798 14420 82850
rect 14140 82740 14196 82750
rect 14140 82646 14196 82684
rect 13468 81778 13524 81788
rect 13580 82012 13860 82068
rect 12460 81730 12516 81742
rect 12460 81678 12462 81730
rect 12514 81678 12516 81730
rect 11900 81118 11902 81170
rect 11954 81118 11956 81170
rect 11900 81106 11956 81118
rect 12348 81172 12404 81182
rect 12460 81172 12516 81678
rect 12348 81170 12516 81172
rect 12348 81118 12350 81170
rect 12402 81118 12516 81170
rect 12348 81116 12516 81118
rect 12348 81106 12404 81116
rect 12124 81060 12180 81070
rect 12124 80966 12180 81004
rect 13468 81058 13524 81070
rect 13468 81006 13470 81058
rect 13522 81006 13524 81058
rect 12796 80948 12852 80958
rect 12796 80854 12852 80892
rect 11676 80780 11844 80836
rect 11676 80498 11732 80780
rect 11676 80446 11678 80498
rect 11730 80446 11732 80498
rect 11676 80434 11732 80446
rect 11228 80222 11230 80274
rect 11282 80222 11284 80274
rect 11228 79268 11284 80222
rect 11900 80388 11956 80398
rect 11228 79202 11284 79212
rect 11452 80162 11508 80174
rect 11452 80110 11454 80162
rect 11506 80110 11508 80162
rect 11452 79044 11508 80110
rect 11676 80164 11732 80174
rect 11676 80070 11732 80108
rect 11900 79828 11956 80332
rect 12908 80164 12964 80174
rect 12908 79828 12964 80108
rect 13468 80164 13524 81006
rect 13468 80098 13524 80108
rect 12908 79772 13188 79828
rect 11900 79762 11956 79772
rect 11564 79604 11620 79614
rect 12012 79604 12068 79614
rect 11564 79602 11732 79604
rect 11564 79550 11566 79602
rect 11618 79550 11732 79602
rect 11564 79548 11732 79550
rect 11564 79538 11620 79548
rect 11116 78988 11508 79044
rect 11116 77812 11172 78988
rect 11228 78820 11284 78830
rect 11564 78820 11620 78830
rect 11228 78818 11620 78820
rect 11228 78766 11230 78818
rect 11282 78766 11566 78818
rect 11618 78766 11620 78818
rect 11228 78764 11620 78766
rect 11228 78754 11284 78764
rect 11564 78754 11620 78764
rect 11452 78596 11508 78606
rect 11452 78502 11508 78540
rect 11004 77756 11172 77812
rect 11340 77924 11396 77934
rect 11004 75906 11060 77756
rect 11004 75854 11006 75906
rect 11058 75854 11060 75906
rect 11004 75842 11060 75854
rect 11116 76468 11172 76478
rect 10892 75684 10948 75694
rect 10892 75590 10948 75628
rect 9884 75010 9940 75180
rect 9884 74958 9886 75010
rect 9938 74958 9940 75010
rect 9660 73556 9716 73566
rect 9660 73462 9716 73500
rect 9548 73330 9604 73342
rect 9548 73278 9550 73330
rect 9602 73278 9604 73330
rect 9548 73220 9604 73278
rect 9548 73154 9604 73164
rect 9772 73330 9828 73342
rect 9772 73278 9774 73330
rect 9826 73278 9828 73330
rect 9548 72660 9604 72670
rect 9436 72658 9604 72660
rect 9436 72606 9550 72658
rect 9602 72606 9604 72658
rect 9436 72604 9604 72606
rect 9548 72594 9604 72604
rect 9772 72548 9828 73278
rect 9884 73220 9940 74958
rect 9996 75012 10052 75022
rect 9996 74918 10052 74956
rect 10220 74898 10276 74910
rect 10220 74846 10222 74898
rect 10274 74846 10276 74898
rect 9884 73154 9940 73164
rect 10108 73890 10164 73902
rect 10108 73838 10110 73890
rect 10162 73838 10164 73890
rect 10108 73332 10164 73838
rect 9772 72482 9828 72492
rect 9884 72436 9940 72446
rect 10108 72436 10164 73276
rect 10220 73330 10276 74846
rect 10780 74898 10836 75292
rect 10780 74846 10782 74898
rect 10834 74846 10836 74898
rect 10780 74834 10836 74846
rect 10892 75012 10948 75022
rect 10892 74786 10948 74956
rect 10892 74734 10894 74786
rect 10946 74734 10948 74786
rect 10892 74338 10948 74734
rect 10892 74286 10894 74338
rect 10946 74286 10948 74338
rect 10892 74274 10948 74286
rect 10220 73278 10222 73330
rect 10274 73278 10276 73330
rect 10220 73266 10276 73278
rect 11004 73332 11060 73342
rect 11004 73238 11060 73276
rect 10556 73220 10612 73230
rect 10612 73164 10724 73220
rect 10556 73126 10612 73164
rect 9940 72380 10164 72436
rect 9884 72322 9940 72380
rect 9884 72270 9886 72322
rect 9938 72270 9940 72322
rect 9660 70308 9716 70318
rect 9660 70214 9716 70252
rect 9436 70196 9492 70206
rect 9436 70102 9492 70140
rect 9772 70194 9828 70206
rect 9772 70142 9774 70194
rect 9826 70142 9828 70194
rect 9772 70084 9828 70142
rect 9772 70018 9828 70028
rect 9884 69188 9940 72270
rect 10556 70308 10612 70318
rect 10332 70084 10388 70094
rect 10388 70028 10500 70084
rect 10332 69990 10388 70028
rect 10444 69188 10500 70028
rect 10556 69410 10612 70252
rect 10668 69972 10724 73164
rect 10780 73106 10836 73118
rect 10780 73054 10782 73106
rect 10834 73054 10836 73106
rect 10780 70194 10836 73054
rect 11116 73108 11172 76412
rect 11228 74228 11284 74238
rect 11228 74134 11284 74172
rect 11340 73892 11396 77868
rect 11676 77028 11732 79548
rect 11676 76962 11732 76972
rect 11900 79602 12068 79604
rect 11900 79550 12014 79602
rect 12066 79550 12068 79602
rect 11900 79548 12068 79550
rect 11564 76466 11620 76478
rect 11564 76414 11566 76466
rect 11618 76414 11620 76466
rect 11564 75908 11620 76414
rect 11676 75908 11732 75918
rect 11564 75906 11732 75908
rect 11564 75854 11678 75906
rect 11730 75854 11732 75906
rect 11564 75852 11732 75854
rect 11676 75842 11732 75852
rect 11676 75012 11732 75022
rect 11900 75012 11956 79548
rect 12012 79538 12068 79548
rect 13020 79602 13076 79614
rect 13020 79550 13022 79602
rect 13074 79550 13076 79602
rect 12908 79378 12964 79390
rect 12908 79326 12910 79378
rect 12962 79326 12964 79378
rect 12012 78932 12068 78942
rect 12012 78838 12068 78876
rect 12908 78260 12964 79326
rect 12908 78194 12964 78204
rect 12460 78034 12516 78046
rect 12460 77982 12462 78034
rect 12514 77982 12516 78034
rect 12460 77924 12516 77982
rect 12012 77028 12068 77038
rect 12012 76580 12068 76972
rect 12460 76692 12516 77868
rect 13020 77364 13076 79550
rect 13020 77298 13076 77308
rect 12572 77252 12628 77262
rect 12628 77196 12740 77252
rect 12572 77186 12628 77196
rect 12460 76626 12516 76636
rect 12012 75906 12068 76524
rect 12012 75854 12014 75906
rect 12066 75854 12068 75906
rect 12012 75842 12068 75854
rect 12460 76356 12516 76366
rect 12348 75796 12404 75806
rect 11676 75010 11956 75012
rect 11676 74958 11678 75010
rect 11730 74958 11956 75010
rect 11676 74956 11956 74958
rect 12236 75740 12348 75796
rect 11676 74946 11732 74956
rect 12236 74900 12292 75740
rect 12348 75730 12404 75740
rect 12460 75572 12516 76300
rect 12572 75572 12628 75582
rect 11788 74844 12236 74900
rect 11788 74226 11844 74844
rect 12236 74806 12292 74844
rect 12348 75570 12628 75572
rect 12348 75518 12574 75570
rect 12626 75518 12628 75570
rect 12348 75516 12628 75518
rect 12348 74676 12404 75516
rect 12572 75506 12628 75516
rect 12684 75348 12740 77196
rect 13132 76580 13188 79772
rect 13244 79604 13300 79614
rect 13244 79602 13412 79604
rect 13244 79550 13246 79602
rect 13298 79550 13412 79602
rect 13244 79548 13412 79550
rect 13244 79538 13300 79548
rect 13356 79156 13412 79548
rect 13020 76524 13188 76580
rect 13244 78932 13300 78942
rect 12796 75796 12852 75806
rect 12796 75682 12852 75740
rect 12796 75630 12798 75682
rect 12850 75630 12852 75682
rect 12796 75618 12852 75630
rect 12684 75292 12852 75348
rect 12684 75124 12740 75134
rect 12684 75010 12740 75068
rect 12684 74958 12686 75010
rect 12738 74958 12740 75010
rect 12684 74946 12740 74958
rect 12572 74900 12628 74910
rect 11788 74174 11790 74226
rect 11842 74174 11844 74226
rect 11788 73948 11844 74174
rect 11340 73332 11396 73836
rect 11676 73892 11844 73948
rect 12012 74620 12404 74676
rect 12460 74786 12516 74798
rect 12460 74734 12462 74786
rect 12514 74734 12516 74786
rect 11340 73266 11396 73276
rect 11452 73330 11508 73342
rect 11452 73278 11454 73330
rect 11506 73278 11508 73330
rect 11340 73108 11396 73118
rect 11452 73108 11508 73278
rect 11676 73220 11732 73892
rect 11676 73154 11732 73164
rect 11116 73106 11508 73108
rect 11116 73054 11342 73106
rect 11394 73054 11508 73106
rect 11116 73052 11508 73054
rect 11340 73042 11396 73052
rect 11116 70756 11172 70766
rect 11116 70662 11172 70700
rect 10780 70142 10782 70194
rect 10834 70142 10836 70194
rect 10780 70130 10836 70142
rect 11228 70196 11284 70206
rect 11228 70194 11732 70196
rect 11228 70142 11230 70194
rect 11282 70142 11732 70194
rect 11228 70140 11732 70142
rect 11228 70130 11284 70140
rect 10668 69916 11172 69972
rect 10556 69358 10558 69410
rect 10610 69358 10612 69410
rect 10556 69346 10612 69358
rect 9884 69186 10052 69188
rect 9884 69134 9886 69186
rect 9938 69134 10052 69186
rect 9884 69132 10052 69134
rect 9884 69122 9940 69132
rect 9996 68514 10052 69132
rect 10444 68850 10500 69132
rect 10444 68798 10446 68850
rect 10498 68798 10500 68850
rect 10444 68786 10500 68798
rect 9996 68462 9998 68514
rect 10050 68462 10052 68514
rect 9436 67618 9492 67630
rect 9436 67566 9438 67618
rect 9490 67566 9492 67618
rect 9436 67284 9492 67566
rect 9884 67618 9940 67630
rect 9884 67566 9886 67618
rect 9938 67566 9940 67618
rect 9884 67508 9940 67566
rect 9884 67442 9940 67452
rect 9660 67284 9716 67294
rect 9436 67228 9660 67284
rect 9324 65426 9380 65436
rect 9660 67058 9716 67228
rect 9660 67006 9662 67058
rect 9714 67006 9716 67058
rect 8988 64148 9044 65212
rect 8988 64054 9044 64092
rect 9212 65044 9268 65054
rect 9212 63364 9268 64988
rect 9660 63924 9716 67006
rect 9884 66164 9940 66174
rect 9772 66052 9828 66062
rect 9884 66052 9940 66108
rect 9772 66050 9940 66052
rect 9772 65998 9774 66050
rect 9826 65998 9940 66050
rect 9772 65996 9940 65998
rect 9772 65986 9828 65996
rect 9660 63922 9828 63924
rect 9660 63870 9662 63922
rect 9714 63870 9828 63922
rect 9660 63868 9828 63870
rect 9660 63858 9716 63868
rect 8764 63252 8820 63262
rect 8764 63138 8820 63196
rect 8764 63086 8766 63138
rect 8818 63086 8820 63138
rect 8764 63074 8820 63086
rect 8988 63026 9044 63038
rect 8988 62974 8990 63026
rect 9042 62974 9044 63026
rect 8876 62580 8932 62590
rect 8988 62580 9044 62974
rect 8876 62578 9044 62580
rect 8876 62526 8878 62578
rect 8930 62526 9044 62578
rect 8876 62524 9044 62526
rect 8876 62468 8932 62524
rect 8876 62402 8932 62412
rect 8988 62188 9044 62524
rect 8988 62132 9156 62188
rect 8876 61346 8932 61358
rect 8876 61294 8878 61346
rect 8930 61294 8932 61346
rect 8764 58212 8820 58222
rect 8764 58118 8820 58156
rect 8764 56084 8820 56094
rect 8764 55970 8820 56028
rect 8764 55918 8766 55970
rect 8818 55918 8820 55970
rect 8764 55524 8820 55918
rect 8764 55458 8820 55468
rect 8876 54516 8932 61294
rect 9100 61346 9156 62132
rect 9212 61570 9268 63308
rect 9548 63140 9604 63150
rect 9548 63046 9604 63084
rect 9772 62356 9828 63868
rect 9772 62188 9828 62300
rect 9212 61518 9214 61570
rect 9266 61518 9268 61570
rect 9212 61506 9268 61518
rect 9324 62132 9828 62188
rect 9884 63140 9940 65996
rect 9996 65716 10052 68462
rect 10892 68516 10948 68526
rect 10108 67060 10164 67070
rect 10108 67058 10724 67060
rect 10108 67006 10110 67058
rect 10162 67006 10724 67058
rect 10108 67004 10724 67006
rect 10108 66994 10164 67004
rect 10668 66498 10724 67004
rect 10668 66446 10670 66498
rect 10722 66446 10724 66498
rect 10668 66434 10724 66446
rect 10780 66836 10836 66846
rect 10220 66388 10276 66398
rect 10276 66332 10388 66388
rect 10220 66294 10276 66332
rect 9996 65650 10052 65660
rect 9996 65492 10052 65502
rect 9996 64260 10052 65436
rect 10220 65492 10276 65502
rect 10108 65044 10164 65054
rect 10108 64930 10164 64988
rect 10108 64878 10110 64930
rect 10162 64878 10164 64930
rect 10108 64866 10164 64878
rect 9996 64204 10164 64260
rect 9884 62466 9940 63084
rect 9996 63922 10052 63934
rect 9996 63870 9998 63922
rect 10050 63870 10052 63922
rect 9996 62578 10052 63870
rect 10108 63252 10164 64204
rect 10108 63138 10164 63196
rect 10108 63086 10110 63138
rect 10162 63086 10164 63138
rect 10108 63074 10164 63086
rect 10220 62916 10276 65436
rect 9996 62526 9998 62578
rect 10050 62526 10052 62578
rect 9996 62514 10052 62526
rect 10108 62860 10276 62916
rect 9884 62414 9886 62466
rect 9938 62414 9940 62466
rect 9100 61294 9102 61346
rect 9154 61294 9156 61346
rect 8988 60676 9044 60686
rect 8988 60582 9044 60620
rect 9100 60564 9156 61294
rect 9100 60498 9156 60508
rect 9324 59332 9380 62132
rect 9884 61348 9940 62414
rect 9660 60674 9716 60686
rect 9660 60622 9662 60674
rect 9714 60622 9716 60674
rect 9660 60116 9716 60622
rect 9660 60050 9716 60060
rect 9212 58436 9268 58446
rect 9324 58436 9380 59276
rect 9212 58434 9380 58436
rect 9212 58382 9214 58434
rect 9266 58382 9380 58434
rect 9212 58380 9380 58382
rect 9212 58370 9268 58380
rect 9100 57540 9156 57550
rect 9100 57446 9156 57484
rect 9100 55858 9156 55870
rect 9100 55806 9102 55858
rect 9154 55806 9156 55858
rect 8988 54628 9044 54638
rect 8988 54534 9044 54572
rect 8876 54450 8932 54460
rect 9100 50706 9156 55806
rect 9212 54628 9268 54638
rect 9212 52836 9268 54572
rect 9324 52948 9380 58380
rect 9548 58434 9604 58446
rect 9548 58382 9550 58434
rect 9602 58382 9604 58434
rect 9436 58212 9492 58222
rect 9436 57764 9492 58156
rect 9436 56868 9492 57708
rect 9548 56980 9604 58382
rect 9660 57426 9716 57438
rect 9660 57374 9662 57426
rect 9714 57374 9716 57426
rect 9660 57204 9716 57374
rect 9660 57138 9716 57148
rect 9660 56980 9716 56990
rect 9548 56924 9660 56980
rect 9660 56914 9716 56924
rect 9436 56812 9604 56868
rect 9436 52948 9492 52958
rect 9324 52892 9436 52948
rect 9436 52854 9492 52892
rect 9212 52780 9380 52836
rect 9212 51938 9268 51950
rect 9212 51886 9214 51938
rect 9266 51886 9268 51938
rect 9212 51716 9268 51886
rect 9212 51650 9268 51660
rect 9100 50654 9102 50706
rect 9154 50654 9156 50706
rect 9100 50428 9156 50654
rect 8652 50372 8820 50428
rect 8652 50036 8708 50046
rect 8652 49942 8708 49980
rect 8540 49756 8708 49812
rect 8540 49588 8596 49598
rect 8540 49494 8596 49532
rect 8540 48468 8596 48478
rect 8428 48466 8596 48468
rect 8428 48414 8542 48466
rect 8594 48414 8596 48466
rect 8428 48412 8596 48414
rect 8540 48244 8596 48412
rect 8540 48178 8596 48188
rect 7756 47406 7758 47458
rect 7810 47406 7812 47458
rect 7756 47394 7812 47406
rect 7868 48076 8036 48132
rect 6860 46788 6916 46798
rect 6860 46002 6916 46732
rect 6860 45950 6862 46002
rect 6914 45950 6916 46002
rect 6860 45938 6916 45950
rect 6972 46562 7028 46574
rect 6972 46510 6974 46562
rect 7026 46510 7028 46562
rect 6972 45892 7028 46510
rect 7084 46564 7140 47180
rect 7420 47346 7476 47358
rect 7420 47294 7422 47346
rect 7474 47294 7476 47346
rect 7420 46900 7476 47294
rect 7420 46834 7476 46844
rect 7532 47234 7588 47246
rect 7532 47182 7534 47234
rect 7586 47182 7588 47234
rect 7308 46564 7364 46574
rect 7532 46564 7588 47182
rect 7756 46564 7812 46574
rect 7084 46562 7476 46564
rect 7084 46510 7310 46562
rect 7362 46510 7476 46562
rect 7084 46508 7476 46510
rect 7532 46562 7812 46564
rect 7532 46510 7758 46562
rect 7810 46510 7812 46562
rect 7532 46508 7812 46510
rect 7308 46498 7364 46508
rect 7308 45892 7364 45902
rect 6972 45890 7364 45892
rect 6972 45838 7310 45890
rect 7362 45838 7364 45890
rect 6972 45836 7364 45838
rect 6748 44604 6916 44660
rect 6748 44436 6804 44446
rect 6748 44342 6804 44380
rect 6524 44034 6580 44044
rect 6636 44100 6692 44110
rect 6636 44098 6804 44100
rect 6636 44046 6638 44098
rect 6690 44046 6804 44098
rect 6636 44044 6804 44046
rect 6636 44034 6692 44044
rect 6748 43314 6804 44044
rect 6748 43262 6750 43314
rect 6802 43262 6804 43314
rect 6748 43250 6804 43262
rect 6300 42642 6356 42812
rect 6300 42590 6302 42642
rect 6354 42590 6356 42642
rect 6300 42578 6356 42590
rect 6748 42644 6804 42654
rect 6748 42550 6804 42588
rect 5852 41020 6244 41076
rect 5740 40962 5796 40974
rect 5740 40910 5742 40962
rect 5794 40910 5796 40962
rect 5740 40740 5796 40910
rect 5740 40674 5796 40684
rect 5740 40516 5796 40526
rect 5740 40422 5796 40460
rect 5740 39732 5796 39742
rect 5628 39730 5796 39732
rect 5628 39678 5742 39730
rect 5794 39678 5796 39730
rect 5628 39676 5796 39678
rect 5404 38882 5460 38892
rect 4620 38836 4676 38874
rect 4620 38770 4676 38780
rect 5068 38834 5124 38846
rect 5068 38782 5070 38834
rect 5122 38782 5124 38834
rect 5068 38668 5124 38782
rect 5740 38836 5796 39676
rect 5852 38836 5908 41020
rect 6300 40962 6356 40974
rect 6300 40910 6302 40962
rect 6354 40910 6356 40962
rect 6076 40180 6132 40190
rect 6300 40180 6356 40910
rect 6748 40628 6804 40638
rect 6636 40516 6692 40526
rect 6636 40422 6692 40460
rect 6748 40402 6804 40572
rect 6748 40350 6750 40402
rect 6802 40350 6804 40402
rect 6748 40338 6804 40350
rect 6076 40178 6356 40180
rect 6076 40126 6078 40178
rect 6130 40126 6356 40178
rect 6076 40124 6356 40126
rect 6076 39060 6132 40124
rect 6188 39620 6244 39630
rect 6524 39620 6580 39630
rect 6244 39564 6468 39620
rect 6188 39554 6244 39564
rect 6076 38994 6132 39004
rect 6188 39396 6244 39406
rect 5852 38780 6132 38836
rect 5740 38668 5796 38780
rect 5068 38612 5684 38668
rect 5740 38612 6020 38668
rect 4008 38444 5208 38454
rect 4064 38442 4112 38444
rect 4168 38442 4216 38444
rect 4076 38390 4112 38442
rect 4200 38390 4216 38442
rect 4064 38388 4112 38390
rect 4168 38388 4216 38390
rect 4272 38442 4320 38444
rect 4376 38442 4424 38444
rect 4480 38442 4528 38444
rect 4376 38390 4396 38442
rect 4480 38390 4520 38442
rect 4272 38388 4320 38390
rect 4376 38388 4424 38390
rect 4480 38388 4528 38390
rect 4584 38388 4632 38444
rect 4688 38442 4736 38444
rect 4792 38442 4840 38444
rect 4896 38442 4944 38444
rect 4696 38390 4736 38442
rect 4820 38390 4840 38442
rect 4688 38388 4736 38390
rect 4792 38388 4840 38390
rect 4896 38388 4944 38390
rect 5000 38442 5048 38444
rect 5104 38442 5152 38444
rect 5000 38390 5016 38442
rect 5104 38390 5140 38442
rect 5000 38388 5048 38390
rect 5104 38388 5152 38390
rect 4008 38378 5208 38388
rect 5628 38388 5684 38612
rect 5628 38332 5908 38388
rect 5852 38274 5908 38332
rect 5852 38222 5854 38274
rect 5906 38222 5908 38274
rect 5852 38210 5908 38222
rect 4008 36876 5208 36886
rect 4064 36874 4112 36876
rect 4168 36874 4216 36876
rect 4076 36822 4112 36874
rect 4200 36822 4216 36874
rect 4064 36820 4112 36822
rect 4168 36820 4216 36822
rect 4272 36874 4320 36876
rect 4376 36874 4424 36876
rect 4480 36874 4528 36876
rect 4376 36822 4396 36874
rect 4480 36822 4520 36874
rect 4272 36820 4320 36822
rect 4376 36820 4424 36822
rect 4480 36820 4528 36822
rect 4584 36820 4632 36876
rect 4688 36874 4736 36876
rect 4792 36874 4840 36876
rect 4896 36874 4944 36876
rect 4696 36822 4736 36874
rect 4820 36822 4840 36874
rect 4688 36820 4736 36822
rect 4792 36820 4840 36822
rect 4896 36820 4944 36822
rect 5000 36874 5048 36876
rect 5104 36874 5152 36876
rect 5000 36822 5016 36874
rect 5104 36822 5140 36874
rect 5000 36820 5048 36822
rect 5104 36820 5152 36822
rect 4008 36810 5208 36820
rect 4620 36372 4676 36382
rect 4844 36372 4900 36382
rect 4620 36370 4900 36372
rect 4620 36318 4622 36370
rect 4674 36318 4846 36370
rect 4898 36318 4900 36370
rect 4620 36316 4900 36318
rect 4620 36306 4676 36316
rect 4060 36260 4116 36270
rect 4060 35476 4116 36204
rect 4844 36036 4900 36316
rect 5180 36372 5236 36382
rect 5180 36278 5236 36316
rect 5852 36372 5908 36382
rect 5852 36278 5908 36316
rect 4956 36260 5012 36270
rect 4956 36166 5012 36204
rect 4844 35970 4900 35980
rect 4956 35924 5012 35934
rect 4956 35830 5012 35868
rect 5292 35924 5348 35934
rect 3612 32050 3668 32060
rect 3724 35420 4116 35476
rect 3612 31892 3668 31902
rect 3500 31890 3668 31892
rect 3500 31838 3614 31890
rect 3666 31838 3668 31890
rect 3500 31836 3668 31838
rect 2604 31556 2660 31566
rect 2604 31554 2772 31556
rect 2604 31502 2606 31554
rect 2658 31502 2772 31554
rect 2604 31500 2772 31502
rect 2604 31490 2660 31500
rect 2156 31444 2212 31454
rect 2156 31218 2212 31388
rect 2156 31166 2158 31218
rect 2210 31166 2212 31218
rect 2156 31154 2212 31166
rect 2604 30882 2660 30894
rect 2604 30830 2606 30882
rect 2658 30830 2660 30882
rect 2604 30212 2660 30830
rect 2716 30436 2772 31500
rect 2828 31444 2884 31454
rect 2828 31106 2884 31388
rect 2828 31054 2830 31106
rect 2882 31054 2884 31106
rect 2828 31042 2884 31054
rect 3164 31108 3220 31118
rect 3164 31014 3220 31052
rect 3164 30772 3220 30782
rect 2828 30436 2884 30446
rect 2716 30380 2828 30436
rect 2604 30146 2660 30156
rect 2828 30210 2884 30380
rect 2828 30158 2830 30210
rect 2882 30158 2884 30210
rect 2828 30146 2884 30158
rect 3164 30098 3220 30716
rect 3500 30210 3556 31836
rect 3612 31826 3668 31836
rect 3500 30158 3502 30210
rect 3554 30158 3556 30210
rect 3500 30146 3556 30158
rect 3724 30212 3780 35420
rect 4008 35308 5208 35318
rect 4064 35306 4112 35308
rect 4168 35306 4216 35308
rect 4076 35254 4112 35306
rect 4200 35254 4216 35306
rect 4064 35252 4112 35254
rect 4168 35252 4216 35254
rect 4272 35306 4320 35308
rect 4376 35306 4424 35308
rect 4480 35306 4528 35308
rect 4376 35254 4396 35306
rect 4480 35254 4520 35306
rect 4272 35252 4320 35254
rect 4376 35252 4424 35254
rect 4480 35252 4528 35254
rect 4584 35252 4632 35308
rect 4688 35306 4736 35308
rect 4792 35306 4840 35308
rect 4896 35306 4944 35308
rect 4696 35254 4736 35306
rect 4820 35254 4840 35306
rect 4688 35252 4736 35254
rect 4792 35252 4840 35254
rect 4896 35252 4944 35254
rect 5000 35306 5048 35308
rect 5104 35306 5152 35308
rect 5000 35254 5016 35306
rect 5104 35254 5140 35306
rect 5000 35252 5048 35254
rect 5104 35252 5152 35254
rect 4008 35242 5208 35252
rect 4732 35140 4788 35150
rect 4620 35028 4676 35038
rect 4172 34916 4228 34926
rect 4172 34822 4228 34860
rect 3836 34692 3892 34702
rect 3836 34598 3892 34636
rect 4620 34354 4676 34972
rect 4732 34914 4788 35084
rect 5292 35028 5348 35868
rect 5852 35924 5908 35934
rect 5964 35924 6020 38612
rect 5852 35922 6020 35924
rect 5852 35870 5854 35922
rect 5906 35870 6020 35922
rect 5852 35868 6020 35870
rect 5852 35858 5908 35868
rect 4732 34862 4734 34914
rect 4786 34862 4788 34914
rect 4732 34850 4788 34862
rect 5180 34972 5292 35028
rect 4956 34804 5012 34814
rect 4956 34710 5012 34748
rect 4620 34302 4622 34354
rect 4674 34302 4676 34354
rect 4620 34290 4676 34302
rect 5180 33908 5236 34972
rect 5292 34962 5348 34972
rect 5404 35476 5460 35486
rect 5292 34804 5348 34814
rect 5292 34354 5348 34748
rect 5292 34302 5294 34354
rect 5346 34302 5348 34354
rect 5292 34290 5348 34302
rect 5180 33852 5348 33908
rect 4008 33740 5208 33750
rect 4064 33738 4112 33740
rect 4168 33738 4216 33740
rect 4076 33686 4112 33738
rect 4200 33686 4216 33738
rect 4064 33684 4112 33686
rect 4168 33684 4216 33686
rect 4272 33738 4320 33740
rect 4376 33738 4424 33740
rect 4480 33738 4528 33740
rect 4376 33686 4396 33738
rect 4480 33686 4520 33738
rect 4272 33684 4320 33686
rect 4376 33684 4424 33686
rect 4480 33684 4528 33686
rect 4584 33684 4632 33740
rect 4688 33738 4736 33740
rect 4792 33738 4840 33740
rect 4896 33738 4944 33740
rect 4696 33686 4736 33738
rect 4820 33686 4840 33738
rect 4688 33684 4736 33686
rect 4792 33684 4840 33686
rect 4896 33684 4944 33686
rect 5000 33738 5048 33740
rect 5104 33738 5152 33740
rect 5000 33686 5016 33738
rect 5104 33686 5140 33738
rect 5000 33684 5048 33686
rect 5104 33684 5152 33686
rect 4008 33674 5208 33684
rect 4620 33570 4676 33582
rect 4620 33518 4622 33570
rect 4674 33518 4676 33570
rect 4620 33458 4676 33518
rect 5180 33572 5236 33582
rect 5292 33572 5348 33852
rect 5180 33570 5292 33572
rect 5180 33518 5182 33570
rect 5234 33518 5292 33570
rect 5180 33516 5292 33518
rect 5180 33506 5236 33516
rect 5292 33478 5348 33516
rect 5068 33460 5124 33470
rect 4620 33406 4622 33458
rect 4674 33406 4676 33458
rect 4620 33394 4676 33406
rect 4732 33404 5068 33460
rect 4172 33124 4228 33134
rect 4172 33030 4228 33068
rect 4732 32788 4788 33404
rect 5068 33366 5124 33404
rect 5180 33348 5236 33358
rect 5180 33012 5236 33292
rect 5180 32946 5236 32956
rect 4732 32694 4788 32732
rect 3836 32452 3892 32462
rect 3836 30882 3892 32396
rect 5180 32452 5236 32462
rect 5404 32452 5460 35420
rect 5516 35474 5572 35486
rect 5516 35422 5518 35474
rect 5570 35422 5572 35474
rect 5516 34020 5572 35422
rect 6076 35028 6132 38780
rect 6188 38274 6244 39340
rect 6188 38222 6190 38274
rect 6242 38222 6244 38274
rect 6188 38210 6244 38222
rect 6412 37938 6468 39564
rect 6524 39526 6580 39564
rect 6412 37886 6414 37938
rect 6466 37886 6468 37938
rect 6412 36594 6468 37886
rect 6412 36542 6414 36594
rect 6466 36542 6468 36594
rect 6188 36482 6244 36494
rect 6188 36430 6190 36482
rect 6242 36430 6244 36482
rect 6188 36260 6244 36430
rect 6188 35364 6244 36204
rect 6300 35924 6356 35934
rect 6300 35830 6356 35868
rect 6188 35308 6356 35364
rect 5852 34972 6132 35028
rect 5628 34916 5684 34926
rect 5628 34354 5684 34860
rect 5628 34302 5630 34354
rect 5682 34302 5684 34354
rect 5628 34290 5684 34302
rect 5740 34692 5796 34702
rect 5516 33954 5572 33964
rect 5740 33684 5796 34636
rect 5180 32450 5460 32452
rect 5180 32398 5182 32450
rect 5234 32398 5460 32450
rect 5180 32396 5460 32398
rect 5516 33628 5796 33684
rect 5516 32452 5572 33628
rect 5852 33572 5908 34972
rect 6076 34804 6132 34814
rect 6076 34710 6132 34748
rect 6188 34692 6244 34702
rect 6188 34598 6244 34636
rect 6188 34356 6244 34366
rect 5740 33516 5908 33572
rect 5964 33906 6020 33918
rect 5964 33854 5966 33906
rect 6018 33854 6020 33906
rect 5740 33348 5796 33516
rect 5964 33460 6020 33854
rect 5180 32386 5236 32396
rect 4008 32172 5208 32182
rect 4064 32170 4112 32172
rect 4168 32170 4216 32172
rect 4076 32118 4112 32170
rect 4200 32118 4216 32170
rect 4064 32116 4112 32118
rect 4168 32116 4216 32118
rect 4272 32170 4320 32172
rect 4376 32170 4424 32172
rect 4480 32170 4528 32172
rect 4376 32118 4396 32170
rect 4480 32118 4520 32170
rect 4272 32116 4320 32118
rect 4376 32116 4424 32118
rect 4480 32116 4528 32118
rect 4584 32116 4632 32172
rect 4688 32170 4736 32172
rect 4792 32170 4840 32172
rect 4896 32170 4944 32172
rect 4696 32118 4736 32170
rect 4820 32118 4840 32170
rect 4688 32116 4736 32118
rect 4792 32116 4840 32118
rect 4896 32116 4944 32118
rect 5000 32170 5048 32172
rect 5104 32170 5152 32172
rect 5000 32118 5016 32170
rect 5104 32118 5140 32170
rect 5000 32116 5048 32118
rect 5104 32116 5152 32118
rect 4008 32106 5208 32116
rect 5292 31892 5348 32396
rect 5516 32386 5572 32396
rect 5628 33292 5796 33348
rect 5852 33404 6020 33460
rect 5628 32786 5684 33292
rect 5740 33122 5796 33134
rect 5740 33070 5742 33122
rect 5794 33070 5796 33122
rect 5740 33012 5796 33070
rect 5740 32946 5796 32956
rect 5628 32734 5630 32786
rect 5682 32734 5684 32786
rect 5628 32338 5684 32734
rect 5628 32286 5630 32338
rect 5682 32286 5684 32338
rect 5628 32274 5684 32286
rect 5404 31892 5460 31902
rect 5292 31836 5404 31892
rect 5404 31826 5460 31836
rect 5852 31892 5908 33404
rect 6076 33348 6132 33358
rect 5852 31826 5908 31836
rect 5964 33346 6132 33348
rect 5964 33294 6078 33346
rect 6130 33294 6132 33346
rect 5964 33292 6132 33294
rect 5964 33124 6020 33292
rect 6076 33282 6132 33292
rect 5068 31780 5124 31790
rect 5068 31686 5124 31724
rect 5628 31668 5684 31678
rect 5292 31666 5684 31668
rect 5292 31614 5630 31666
rect 5682 31614 5684 31666
rect 5292 31612 5684 31614
rect 4508 31554 4564 31566
rect 4508 31502 4510 31554
rect 4562 31502 4564 31554
rect 4508 30996 4564 31502
rect 4508 30930 4564 30940
rect 3836 30830 3838 30882
rect 3890 30830 3892 30882
rect 3836 30436 3892 30830
rect 4008 30604 5208 30614
rect 4064 30602 4112 30604
rect 4168 30602 4216 30604
rect 4076 30550 4112 30602
rect 4200 30550 4216 30602
rect 4064 30548 4112 30550
rect 4168 30548 4216 30550
rect 4272 30602 4320 30604
rect 4376 30602 4424 30604
rect 4480 30602 4528 30604
rect 4376 30550 4396 30602
rect 4480 30550 4520 30602
rect 4272 30548 4320 30550
rect 4376 30548 4424 30550
rect 4480 30548 4528 30550
rect 4584 30548 4632 30604
rect 4688 30602 4736 30604
rect 4792 30602 4840 30604
rect 4896 30602 4944 30604
rect 4696 30550 4736 30602
rect 4820 30550 4840 30602
rect 4688 30548 4736 30550
rect 4792 30548 4840 30550
rect 4896 30548 4944 30550
rect 5000 30602 5048 30604
rect 5104 30602 5152 30604
rect 5000 30550 5016 30602
rect 5104 30550 5140 30602
rect 5000 30548 5048 30550
rect 5104 30548 5152 30550
rect 4008 30538 5208 30548
rect 3836 30380 4116 30436
rect 3724 30146 3780 30156
rect 4060 30210 4116 30380
rect 4844 30322 4900 30334
rect 4844 30270 4846 30322
rect 4898 30270 4900 30322
rect 4732 30212 4788 30222
rect 4060 30158 4062 30210
rect 4114 30158 4116 30210
rect 3164 30046 3166 30098
rect 3218 30046 3220 30098
rect 3164 30034 3220 30046
rect 3948 30100 4004 30110
rect 2156 29986 2212 29998
rect 2156 29934 2158 29986
rect 2210 29934 2212 29986
rect 2156 29876 2212 29934
rect 2156 29810 2212 29820
rect 2604 29986 2660 29998
rect 2604 29934 2606 29986
rect 2658 29934 2660 29986
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 29362 1876 29374
rect 2044 29540 2100 29550
rect 2044 28644 2100 29484
rect 2268 29426 2324 29438
rect 2268 29374 2270 29426
rect 2322 29374 2324 29426
rect 2156 29204 2212 29214
rect 2156 28756 2212 29148
rect 2268 28980 2324 29374
rect 2492 28980 2548 28990
rect 2268 28924 2492 28980
rect 2492 28914 2548 28924
rect 2156 28700 2548 28756
rect 2044 28588 2324 28644
rect 1596 28532 1652 28542
rect 1596 28082 1652 28476
rect 1596 28030 1598 28082
rect 1650 28030 1652 28082
rect 1596 28018 1652 28030
rect 2268 28530 2324 28588
rect 2268 28478 2270 28530
rect 2322 28478 2324 28530
rect 2268 28082 2324 28478
rect 2268 28030 2270 28082
rect 2322 28030 2324 28082
rect 2268 28018 2324 28030
rect 1820 27972 1876 27982
rect 1708 25844 1764 25854
rect 1708 22932 1764 25788
rect 1820 24948 1876 27916
rect 2156 27076 2212 27086
rect 2380 27076 2436 28700
rect 2492 28642 2548 28700
rect 2492 28590 2494 28642
rect 2546 28590 2548 28642
rect 2492 28578 2548 28590
rect 2156 27074 2436 27076
rect 2156 27022 2158 27074
rect 2210 27022 2436 27074
rect 2156 27020 2436 27022
rect 2156 27010 2212 27020
rect 2604 26850 2660 29934
rect 3276 29988 3332 29998
rect 3164 28868 3220 28906
rect 3164 28802 3220 28812
rect 2828 28644 2884 28654
rect 2828 28530 2884 28588
rect 3164 28644 3220 28654
rect 3276 28644 3332 29932
rect 3724 29988 3780 29998
rect 3724 29894 3780 29932
rect 3948 29652 4004 30044
rect 4060 29876 4116 30158
rect 4620 30156 4732 30212
rect 4060 29810 4116 29820
rect 4508 30098 4564 30110
rect 4508 30046 4510 30098
rect 4562 30046 4564 30098
rect 3836 29428 3892 29438
rect 3164 28642 3332 28644
rect 3164 28590 3166 28642
rect 3218 28590 3332 28642
rect 3164 28588 3332 28590
rect 3500 29316 3556 29326
rect 3500 28866 3556 29260
rect 3500 28814 3502 28866
rect 3554 28814 3556 28866
rect 3164 28578 3220 28588
rect 2828 28478 2830 28530
rect 2882 28478 2884 28530
rect 2828 28466 2884 28478
rect 2940 28420 2996 28430
rect 2940 27076 2996 28364
rect 3388 27300 3444 27310
rect 3500 27300 3556 28814
rect 3836 28868 3892 29372
rect 3948 29204 4004 29596
rect 4508 29428 4564 30046
rect 4620 29650 4676 30156
rect 4732 30146 4788 30156
rect 4620 29598 4622 29650
rect 4674 29598 4676 29650
rect 4620 29540 4676 29598
rect 4620 29474 4676 29484
rect 4732 29986 4788 29998
rect 4732 29934 4734 29986
rect 4786 29934 4788 29986
rect 4508 29362 4564 29372
rect 4732 29316 4788 29934
rect 4732 29250 4788 29260
rect 3948 29138 4004 29148
rect 4844 29204 4900 30270
rect 5180 30324 5236 30334
rect 5180 29204 5236 30268
rect 5292 29650 5348 31612
rect 5628 31602 5684 31612
rect 5516 30996 5572 31006
rect 5516 30902 5572 30940
rect 5852 30212 5908 30222
rect 5852 30118 5908 30156
rect 5292 29598 5294 29650
rect 5346 29598 5348 29650
rect 5292 29586 5348 29598
rect 5404 29708 5796 29764
rect 5180 29148 5348 29204
rect 4844 29138 4900 29148
rect 4008 29036 5208 29046
rect 4064 29034 4112 29036
rect 4168 29034 4216 29036
rect 4076 28982 4112 29034
rect 4200 28982 4216 29034
rect 4064 28980 4112 28982
rect 4168 28980 4216 28982
rect 4272 29034 4320 29036
rect 4376 29034 4424 29036
rect 4480 29034 4528 29036
rect 4376 28982 4396 29034
rect 4480 28982 4520 29034
rect 4272 28980 4320 28982
rect 4376 28980 4424 28982
rect 4480 28980 4528 28982
rect 4584 28980 4632 29036
rect 4688 29034 4736 29036
rect 4792 29034 4840 29036
rect 4896 29034 4944 29036
rect 4696 28982 4736 29034
rect 4820 28982 4840 29034
rect 4688 28980 4736 28982
rect 4792 28980 4840 28982
rect 4896 28980 4944 28982
rect 5000 29034 5048 29036
rect 5104 29034 5152 29036
rect 5000 28982 5016 29034
rect 5104 28982 5140 29034
rect 5000 28980 5048 28982
rect 5104 28980 5152 28982
rect 4008 28970 5208 28980
rect 4172 28868 4228 28878
rect 3836 28812 4116 28868
rect 3836 28644 3892 28654
rect 3724 28588 3836 28644
rect 3612 27300 3668 27310
rect 3500 27298 3668 27300
rect 3500 27246 3614 27298
rect 3666 27246 3668 27298
rect 3500 27244 3668 27246
rect 3388 27186 3444 27244
rect 3612 27234 3668 27244
rect 3388 27134 3390 27186
rect 3442 27134 3444 27186
rect 3388 27122 3444 27134
rect 3724 27076 3780 28588
rect 3836 28578 3892 28588
rect 3948 28532 4004 28542
rect 3948 28438 4004 28476
rect 3836 28420 3892 28430
rect 4060 28420 4116 28812
rect 4172 28642 4228 28812
rect 4732 28868 4788 28878
rect 4172 28590 4174 28642
rect 4226 28590 4228 28642
rect 4172 28578 4228 28590
rect 4508 28644 4564 28654
rect 4508 28550 4564 28588
rect 4284 28420 4340 28430
rect 4060 28418 4340 28420
rect 4060 28366 4286 28418
rect 4338 28366 4340 28418
rect 4060 28364 4340 28366
rect 3836 27300 3892 28364
rect 4284 28354 4340 28364
rect 4732 27858 4788 28812
rect 4956 28868 5012 28878
rect 5292 28868 5348 29148
rect 4956 28866 5348 28868
rect 4956 28814 4958 28866
rect 5010 28814 5348 28866
rect 4956 28812 5348 28814
rect 4956 28802 5012 28812
rect 5404 28756 5460 29708
rect 5628 29538 5684 29550
rect 5628 29486 5630 29538
rect 5682 29486 5684 29538
rect 5068 28700 5460 28756
rect 5516 29202 5572 29214
rect 5516 29150 5518 29202
rect 5570 29150 5572 29202
rect 4844 28532 4900 28542
rect 4844 28438 4900 28476
rect 4956 28532 5012 28542
rect 5068 28532 5124 28700
rect 4956 28530 5124 28532
rect 4956 28478 4958 28530
rect 5010 28478 5124 28530
rect 4956 28476 5124 28478
rect 5180 28532 5236 28542
rect 4732 27806 4734 27858
rect 4786 27806 4788 27858
rect 4732 27794 4788 27806
rect 4956 27636 5012 28476
rect 5180 27636 5236 28476
rect 5516 28420 5572 29150
rect 5628 28644 5684 29486
rect 5740 29540 5796 29708
rect 5852 29540 5908 29550
rect 5740 29538 5908 29540
rect 5740 29486 5854 29538
rect 5906 29486 5908 29538
rect 5740 29484 5908 29486
rect 5852 29474 5908 29484
rect 5628 28642 5796 28644
rect 5628 28590 5630 28642
rect 5682 28590 5796 28642
rect 5628 28588 5796 28590
rect 5628 28578 5684 28588
rect 5516 28354 5572 28364
rect 5516 28196 5572 28206
rect 5292 28140 5516 28196
rect 5292 27858 5348 28140
rect 5292 27806 5294 27858
rect 5346 27806 5348 27858
rect 5292 27794 5348 27806
rect 5180 27580 5348 27636
rect 4956 27570 5012 27580
rect 4008 27468 5208 27478
rect 4064 27466 4112 27468
rect 4168 27466 4216 27468
rect 4076 27414 4112 27466
rect 4200 27414 4216 27466
rect 4064 27412 4112 27414
rect 4168 27412 4216 27414
rect 4272 27466 4320 27468
rect 4376 27466 4424 27468
rect 4480 27466 4528 27468
rect 4376 27414 4396 27466
rect 4480 27414 4520 27466
rect 4272 27412 4320 27414
rect 4376 27412 4424 27414
rect 4480 27412 4528 27414
rect 4584 27412 4632 27468
rect 4688 27466 4736 27468
rect 4792 27466 4840 27468
rect 4896 27466 4944 27468
rect 4696 27414 4736 27466
rect 4820 27414 4840 27466
rect 4688 27412 4736 27414
rect 4792 27412 4840 27414
rect 4896 27412 4944 27414
rect 5000 27466 5048 27468
rect 5104 27466 5152 27468
rect 5000 27414 5016 27466
rect 5104 27414 5140 27466
rect 5000 27412 5048 27414
rect 5104 27412 5152 27414
rect 4008 27402 5208 27412
rect 4284 27300 4340 27310
rect 3836 27244 4228 27300
rect 2940 26962 2996 27020
rect 2940 26910 2942 26962
rect 2994 26910 2996 26962
rect 2940 26898 2996 26910
rect 3500 27020 3780 27076
rect 4172 27074 4228 27244
rect 4172 27022 4174 27074
rect 4226 27022 4228 27074
rect 2604 26798 2606 26850
rect 2658 26798 2660 26850
rect 2604 26516 2660 26798
rect 2604 26450 2660 26460
rect 3164 26852 3220 26862
rect 3052 26068 3108 26078
rect 1820 24946 2212 24948
rect 1820 24894 1822 24946
rect 1874 24894 2212 24946
rect 1820 24892 2212 24894
rect 1820 24882 1876 24892
rect 2044 24612 2100 24622
rect 1932 23716 1988 23726
rect 1708 22866 1764 22876
rect 1820 23714 1988 23716
rect 1820 23662 1934 23714
rect 1986 23662 1988 23714
rect 1820 23660 1988 23662
rect 1820 23492 1876 23660
rect 1932 23650 1988 23660
rect 1708 22484 1764 22494
rect 1820 22484 1876 23436
rect 1764 22428 1876 22484
rect 1932 23268 1988 23278
rect 1708 22418 1764 22428
rect 1820 22146 1876 22158
rect 1820 22094 1822 22146
rect 1874 22094 1876 22146
rect 1708 21588 1764 21598
rect 1708 21494 1764 21532
rect 1820 21364 1876 22094
rect 1820 21298 1876 21308
rect 1932 20914 1988 23212
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20850 1988 20862
rect 2044 20692 2100 24556
rect 2156 23938 2212 24892
rect 2828 24722 2884 24734
rect 2828 24670 2830 24722
rect 2882 24670 2884 24722
rect 2492 24612 2548 24622
rect 2828 24612 2884 24670
rect 2548 24556 2884 24612
rect 2940 24724 2996 24734
rect 2492 24518 2548 24556
rect 2156 23886 2158 23938
rect 2210 23886 2212 23938
rect 2156 23874 2212 23886
rect 2716 23828 2772 23838
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 1820 20636 2100 20692
rect 2156 23604 2212 23614
rect 2156 22370 2212 23548
rect 2268 23266 2324 23278
rect 2268 23214 2270 23266
rect 2322 23214 2324 23266
rect 2268 23156 2324 23214
rect 2268 23090 2324 23100
rect 2156 22318 2158 22370
rect 2210 22318 2212 22370
rect 1708 16658 1764 16670
rect 1708 16606 1710 16658
rect 1762 16606 1764 16658
rect 1708 15876 1764 16606
rect 1820 16212 1876 20636
rect 2156 20188 2212 22318
rect 1932 20132 2212 20188
rect 2268 22932 2324 22942
rect 2268 20188 2324 22876
rect 2380 22820 2436 22830
rect 2380 21586 2436 22764
rect 2492 22596 2548 23662
rect 2492 22530 2548 22540
rect 2604 23154 2660 23166
rect 2604 23102 2606 23154
rect 2658 23102 2660 23154
rect 2604 22484 2660 23102
rect 2716 22596 2772 23772
rect 2828 23826 2884 23838
rect 2828 23774 2830 23826
rect 2882 23774 2884 23826
rect 2828 23492 2884 23774
rect 2828 23426 2884 23436
rect 2716 22540 2884 22596
rect 2604 22428 2772 22484
rect 2492 22372 2548 22382
rect 2492 22258 2548 22316
rect 2716 22260 2772 22428
rect 2828 22372 2884 22540
rect 2828 22306 2884 22316
rect 2492 22206 2494 22258
rect 2546 22206 2548 22258
rect 2492 22194 2548 22206
rect 2604 22204 2772 22260
rect 2380 21534 2382 21586
rect 2434 21534 2436 21586
rect 2380 21522 2436 21534
rect 2604 21364 2660 22204
rect 2828 22148 2884 22158
rect 2604 21298 2660 21308
rect 2716 22146 2884 22148
rect 2716 22094 2830 22146
rect 2882 22094 2884 22146
rect 2716 22092 2884 22094
rect 2492 20580 2548 20590
rect 2716 20580 2772 22092
rect 2828 22082 2884 22092
rect 2492 20578 2772 20580
rect 2492 20526 2494 20578
rect 2546 20526 2772 20578
rect 2492 20524 2772 20526
rect 2828 20690 2884 20702
rect 2828 20638 2830 20690
rect 2882 20638 2884 20690
rect 2492 20244 2548 20524
rect 2268 20132 2436 20188
rect 2492 20178 2548 20188
rect 1932 20130 1988 20132
rect 1932 20078 1934 20130
rect 1986 20078 1988 20130
rect 1932 20066 1988 20078
rect 2044 19458 2100 19470
rect 2044 19406 2046 19458
rect 2098 19406 2100 19458
rect 2044 19346 2100 19406
rect 2044 19294 2046 19346
rect 2098 19294 2100 19346
rect 2044 19282 2100 19294
rect 2380 18788 2436 20132
rect 2492 19908 2548 19918
rect 2828 19908 2884 20638
rect 2492 19906 2884 19908
rect 2492 19854 2494 19906
rect 2546 19854 2884 19906
rect 2492 19852 2884 19854
rect 2492 19236 2548 19852
rect 2604 19460 2660 19470
rect 2940 19460 2996 24668
rect 2604 19458 2996 19460
rect 2604 19406 2606 19458
rect 2658 19406 2996 19458
rect 2604 19404 2996 19406
rect 2604 19394 2660 19404
rect 2492 19170 2548 19180
rect 2828 19236 2884 19246
rect 2492 19012 2548 19022
rect 2828 19012 2884 19180
rect 2940 19234 2996 19404
rect 2940 19182 2942 19234
rect 2994 19182 2996 19234
rect 2940 19170 2996 19182
rect 2492 19010 2884 19012
rect 2492 18958 2494 19010
rect 2546 18958 2884 19010
rect 2492 18956 2884 18958
rect 2492 18946 2548 18956
rect 2380 18732 2660 18788
rect 2604 18452 2660 18732
rect 2828 18452 2884 18462
rect 2604 18450 2884 18452
rect 2604 18398 2606 18450
rect 2658 18398 2830 18450
rect 2882 18398 2884 18450
rect 2604 18396 2884 18398
rect 2604 18386 2660 18396
rect 2828 18386 2884 18396
rect 2604 17444 2660 17454
rect 2828 17444 2884 17454
rect 2604 17442 2884 17444
rect 2604 17390 2606 17442
rect 2658 17390 2830 17442
rect 2882 17390 2884 17442
rect 2604 17388 2884 17390
rect 3052 17444 3108 26012
rect 3164 25508 3220 26796
rect 3500 26514 3556 27020
rect 4172 27010 4228 27022
rect 3948 26964 4004 27002
rect 3948 26898 4004 26908
rect 3724 26850 3780 26862
rect 3724 26798 3726 26850
rect 3778 26798 3780 26850
rect 3500 26462 3502 26514
rect 3554 26462 3556 26514
rect 3500 26450 3556 26462
rect 3612 26628 3668 26638
rect 3164 24946 3220 25452
rect 3164 24894 3166 24946
rect 3218 24894 3220 24946
rect 3164 24882 3220 24894
rect 3276 26292 3332 26302
rect 3164 24724 3220 24734
rect 3164 23268 3220 24668
rect 3276 23548 3332 26236
rect 3500 25732 3556 25742
rect 3388 23716 3444 23726
rect 3388 23622 3444 23660
rect 3276 23482 3332 23492
rect 3164 23212 3332 23268
rect 3276 22482 3332 23212
rect 3388 23044 3444 23054
rect 3388 22950 3444 22988
rect 3276 22430 3278 22482
rect 3330 22430 3332 22482
rect 3276 22418 3332 22430
rect 3500 22372 3556 25676
rect 3612 23268 3668 26572
rect 3724 26516 3780 26798
rect 3836 26516 3892 26526
rect 3724 26460 3836 26516
rect 3836 26422 3892 26460
rect 4284 26178 4340 27244
rect 4732 27300 4788 27310
rect 4732 27206 4788 27244
rect 5068 27188 5124 27198
rect 5068 27094 5124 27132
rect 4508 27074 4564 27086
rect 4508 27022 4510 27074
rect 4562 27022 4564 27074
rect 4508 26964 4564 27022
rect 4508 26898 4564 26908
rect 4844 27076 4900 27086
rect 4844 26514 4900 27020
rect 4844 26462 4846 26514
rect 4898 26462 4900 26514
rect 4844 26450 4900 26462
rect 4956 27074 5012 27086
rect 4956 27022 4958 27074
rect 5010 27022 5012 27074
rect 4620 26292 4676 26302
rect 4956 26292 5012 27022
rect 5292 27076 5348 27580
rect 5292 27010 5348 27020
rect 4676 26236 5012 26292
rect 5292 26516 5348 26526
rect 5292 26290 5348 26460
rect 5292 26238 5294 26290
rect 5346 26238 5348 26290
rect 4620 26198 4676 26236
rect 5292 26226 5348 26238
rect 4284 26126 4286 26178
rect 4338 26126 4340 26178
rect 3612 23202 3668 23212
rect 3724 26066 3780 26078
rect 3724 26014 3726 26066
rect 3778 26014 3780 26066
rect 3500 22316 3668 22372
rect 3164 20692 3220 20702
rect 3164 20598 3220 20636
rect 3612 19236 3668 22316
rect 3612 19142 3668 19180
rect 3164 19012 3220 19022
rect 3164 19010 3332 19012
rect 3164 18958 3166 19010
rect 3218 18958 3332 19010
rect 3164 18956 3332 18958
rect 3164 18946 3220 18956
rect 3164 18562 3220 18574
rect 3164 18510 3166 18562
rect 3218 18510 3220 18562
rect 3164 17668 3220 18510
rect 3276 17892 3332 18956
rect 3276 17826 3332 17836
rect 3164 17612 3332 17668
rect 3164 17444 3220 17454
rect 3052 17442 3220 17444
rect 3052 17390 3166 17442
rect 3218 17390 3220 17442
rect 3052 17388 3220 17390
rect 2492 17108 2548 17118
rect 2492 17014 2548 17052
rect 1932 16996 1988 17006
rect 1932 16902 1988 16940
rect 2156 16882 2212 16894
rect 2156 16830 2158 16882
rect 2210 16830 2212 16882
rect 1932 16660 1988 16670
rect 2156 16660 2212 16830
rect 1932 16658 2212 16660
rect 1932 16606 1934 16658
rect 1986 16606 2212 16658
rect 1932 16604 2212 16606
rect 1932 16594 1988 16604
rect 1820 16156 1988 16212
rect 1820 15876 1876 15886
rect 1708 15874 1876 15876
rect 1708 15822 1822 15874
rect 1874 15822 1876 15874
rect 1708 15820 1876 15822
rect 1708 14644 1764 15820
rect 1820 15810 1876 15820
rect 1708 14578 1764 14588
rect 1820 15314 1876 15326
rect 1820 15262 1822 15314
rect 1874 15262 1876 15314
rect 1820 15204 1876 15262
rect 1820 12178 1876 15148
rect 1932 13524 1988 16156
rect 2604 16100 2660 17388
rect 2828 17378 2884 17388
rect 3164 17378 3220 17388
rect 2940 16996 2996 17006
rect 2940 16882 2996 16940
rect 2940 16830 2942 16882
rect 2994 16830 2996 16882
rect 2940 16818 2996 16830
rect 3164 16994 3220 17006
rect 3164 16942 3166 16994
rect 3218 16942 3220 16994
rect 2604 16034 2660 16044
rect 3052 15876 3108 15886
rect 2268 15874 3108 15876
rect 2268 15822 3054 15874
rect 3106 15822 3108 15874
rect 2268 15820 3108 15822
rect 2268 15314 2324 15820
rect 3052 15810 3108 15820
rect 2268 15262 2270 15314
rect 2322 15262 2324 15314
rect 2268 15250 2324 15262
rect 3164 14756 3220 16942
rect 3276 16772 3332 17612
rect 3612 16772 3668 16782
rect 3276 16706 3332 16716
rect 3388 16770 3668 16772
rect 3388 16718 3614 16770
rect 3666 16718 3668 16770
rect 3388 16716 3668 16718
rect 3388 16322 3444 16716
rect 3612 16706 3668 16716
rect 3724 16548 3780 26014
rect 4284 26066 4340 26126
rect 4284 26014 4286 26066
rect 4338 26014 4340 26066
rect 4284 26002 4340 26014
rect 4956 26068 5012 26106
rect 4956 26002 5012 26012
rect 4008 25900 5208 25910
rect 4064 25898 4112 25900
rect 4168 25898 4216 25900
rect 4076 25846 4112 25898
rect 4200 25846 4216 25898
rect 4064 25844 4112 25846
rect 4168 25844 4216 25846
rect 4272 25898 4320 25900
rect 4376 25898 4424 25900
rect 4480 25898 4528 25900
rect 4376 25846 4396 25898
rect 4480 25846 4520 25898
rect 4272 25844 4320 25846
rect 4376 25844 4424 25846
rect 4480 25844 4528 25846
rect 4584 25844 4632 25900
rect 4688 25898 4736 25900
rect 4792 25898 4840 25900
rect 4896 25898 4944 25900
rect 4696 25846 4736 25898
rect 4820 25846 4840 25898
rect 4688 25844 4736 25846
rect 4792 25844 4840 25846
rect 4896 25844 4944 25846
rect 5000 25898 5048 25900
rect 5104 25898 5152 25900
rect 5000 25846 5016 25898
rect 5104 25846 5140 25898
rect 5000 25844 5048 25846
rect 5104 25844 5152 25846
rect 4008 25834 5208 25844
rect 5404 25732 5460 28140
rect 5516 28130 5572 28140
rect 5740 27860 5796 28588
rect 5852 28642 5908 28654
rect 5852 28590 5854 28642
rect 5906 28590 5908 28642
rect 5852 28532 5908 28590
rect 5964 28532 6020 33068
rect 6188 32676 6244 34300
rect 6300 33572 6356 35308
rect 6412 35140 6468 36542
rect 6412 35074 6468 35084
rect 6524 39060 6580 39070
rect 6412 34692 6468 34702
rect 6412 34598 6468 34636
rect 6524 34468 6580 39004
rect 6524 34402 6580 34412
rect 6636 35252 6692 35262
rect 6524 34244 6580 34254
rect 6412 34188 6524 34244
rect 6412 34130 6468 34188
rect 6524 34178 6580 34188
rect 6636 34242 6692 35196
rect 6636 34190 6638 34242
rect 6690 34190 6692 34242
rect 6636 34178 6692 34190
rect 6748 34914 6804 34926
rect 6748 34862 6750 34914
rect 6802 34862 6804 34914
rect 6412 34078 6414 34130
rect 6466 34078 6468 34130
rect 6412 34066 6468 34078
rect 6524 34020 6580 34030
rect 6300 33516 6468 33572
rect 6188 32620 6356 32676
rect 6188 32452 6244 32462
rect 6188 32358 6244 32396
rect 6076 32338 6132 32350
rect 6076 32286 6078 32338
rect 6130 32286 6132 32338
rect 6076 32004 6132 32286
rect 6188 32004 6244 32014
rect 6076 32002 6244 32004
rect 6076 31950 6190 32002
rect 6242 31950 6244 32002
rect 6076 31948 6244 31950
rect 6076 31780 6132 31948
rect 6188 31938 6244 31948
rect 6076 31714 6132 31724
rect 6076 30324 6132 30334
rect 6076 30230 6132 30268
rect 6076 28532 6132 28542
rect 5964 28476 6076 28532
rect 5852 28466 5908 28476
rect 6076 28466 6132 28476
rect 6188 28420 6244 28430
rect 6188 28326 6244 28364
rect 5628 27748 5684 27758
rect 5516 27636 5572 27646
rect 5516 27300 5572 27580
rect 5516 27234 5572 27244
rect 5628 27074 5684 27692
rect 5628 27022 5630 27074
rect 5682 27022 5684 27074
rect 5628 27010 5684 27022
rect 5740 27076 5796 27804
rect 5964 27858 6020 27870
rect 6188 27860 6244 27870
rect 5964 27806 5966 27858
rect 6018 27806 6020 27858
rect 5964 27412 6020 27806
rect 6076 27858 6244 27860
rect 6076 27806 6190 27858
rect 6242 27806 6244 27858
rect 6076 27804 6244 27806
rect 6076 27748 6132 27804
rect 6188 27794 6244 27804
rect 6076 27682 6132 27692
rect 5964 27346 6020 27356
rect 6188 27636 6244 27646
rect 6076 27188 6132 27198
rect 6076 27094 6132 27132
rect 5740 27010 5796 27020
rect 5852 26962 5908 26974
rect 5852 26910 5854 26962
rect 5906 26910 5908 26962
rect 5628 26850 5684 26862
rect 5628 26798 5630 26850
rect 5682 26798 5684 26850
rect 5068 25676 5460 25732
rect 5516 26066 5572 26078
rect 5516 26014 5518 26066
rect 5570 26014 5572 26066
rect 5516 25732 5572 26014
rect 5628 26068 5684 26798
rect 5628 26002 5684 26012
rect 5740 26852 5796 26862
rect 5628 25732 5684 25742
rect 5516 25730 5684 25732
rect 5516 25678 5630 25730
rect 5682 25678 5684 25730
rect 5516 25676 5684 25678
rect 4172 25620 4228 25630
rect 3836 24724 3892 24734
rect 3836 24630 3892 24668
rect 4172 24500 4228 25564
rect 5068 25618 5124 25676
rect 5068 25566 5070 25618
rect 5122 25566 5124 25618
rect 5068 25554 5124 25566
rect 5404 25620 5460 25676
rect 5628 25666 5684 25676
rect 5740 25730 5796 26796
rect 5852 26516 5908 26910
rect 5852 26450 5908 26460
rect 6076 26628 6132 26638
rect 5740 25678 5742 25730
rect 5794 25678 5796 25730
rect 5740 25666 5796 25678
rect 5852 26066 5908 26078
rect 5852 26014 5854 26066
rect 5906 26014 5908 26066
rect 5404 25554 5460 25564
rect 4732 25396 4788 25406
rect 4732 25302 4788 25340
rect 3836 24444 4228 24500
rect 5292 25284 5348 25294
rect 5292 24610 5348 25228
rect 5292 24558 5294 24610
rect 5346 24558 5348 24610
rect 3836 24164 3892 24444
rect 4008 24332 5208 24342
rect 4064 24330 4112 24332
rect 4168 24330 4216 24332
rect 4076 24278 4112 24330
rect 4200 24278 4216 24330
rect 4064 24276 4112 24278
rect 4168 24276 4216 24278
rect 4272 24330 4320 24332
rect 4376 24330 4424 24332
rect 4480 24330 4528 24332
rect 4376 24278 4396 24330
rect 4480 24278 4520 24330
rect 4272 24276 4320 24278
rect 4376 24276 4424 24278
rect 4480 24276 4528 24278
rect 4584 24276 4632 24332
rect 4688 24330 4736 24332
rect 4792 24330 4840 24332
rect 4896 24330 4944 24332
rect 4696 24278 4736 24330
rect 4820 24278 4840 24330
rect 4688 24276 4736 24278
rect 4792 24276 4840 24278
rect 4896 24276 4944 24278
rect 5000 24330 5048 24332
rect 5104 24330 5152 24332
rect 5000 24278 5016 24330
rect 5104 24278 5140 24330
rect 5000 24276 5048 24278
rect 5104 24276 5152 24278
rect 4008 24266 5208 24276
rect 3836 24108 4004 24164
rect 3836 23492 3892 23502
rect 3836 23378 3892 23436
rect 3836 23326 3838 23378
rect 3890 23326 3892 23378
rect 3836 23314 3892 23326
rect 3948 23268 4004 24108
rect 4508 23828 4564 23838
rect 4508 23734 4564 23772
rect 4396 23716 4452 23726
rect 4060 23714 4452 23716
rect 4060 23662 4398 23714
rect 4450 23662 4452 23714
rect 4060 23660 4452 23662
rect 4060 23378 4116 23660
rect 4396 23650 4452 23660
rect 5068 23714 5124 23726
rect 5068 23662 5070 23714
rect 5122 23662 5124 23714
rect 4508 23604 4564 23614
rect 4060 23326 4062 23378
rect 4114 23326 4116 23378
rect 4060 23314 4116 23326
rect 4284 23492 4564 23548
rect 3948 23202 4004 23212
rect 4284 23154 4340 23492
rect 4284 23102 4286 23154
rect 4338 23102 4340 23154
rect 4284 23090 4340 23102
rect 5068 23156 5124 23662
rect 5180 23492 5236 23502
rect 5180 23378 5236 23436
rect 5180 23326 5182 23378
rect 5234 23326 5236 23378
rect 5180 23314 5236 23326
rect 5292 23156 5348 24558
rect 5068 23154 5348 23156
rect 5068 23102 5294 23154
rect 5346 23102 5348 23154
rect 5068 23100 5348 23102
rect 3948 23042 4004 23054
rect 3948 22990 3950 23042
rect 4002 22990 4004 23042
rect 3948 22932 4004 22990
rect 3948 22866 4004 22876
rect 4508 22932 4564 22970
rect 4508 22866 4564 22876
rect 4008 22764 5208 22774
rect 4064 22762 4112 22764
rect 4168 22762 4216 22764
rect 4076 22710 4112 22762
rect 4200 22710 4216 22762
rect 4064 22708 4112 22710
rect 4168 22708 4216 22710
rect 4272 22762 4320 22764
rect 4376 22762 4424 22764
rect 4480 22762 4528 22764
rect 4376 22710 4396 22762
rect 4480 22710 4520 22762
rect 4272 22708 4320 22710
rect 4376 22708 4424 22710
rect 4480 22708 4528 22710
rect 4584 22708 4632 22764
rect 4688 22762 4736 22764
rect 4792 22762 4840 22764
rect 4896 22762 4944 22764
rect 4696 22710 4736 22762
rect 4820 22710 4840 22762
rect 4688 22708 4736 22710
rect 4792 22708 4840 22710
rect 4896 22708 4944 22710
rect 5000 22762 5048 22764
rect 5104 22762 5152 22764
rect 5000 22710 5016 22762
rect 5104 22710 5140 22762
rect 5000 22708 5048 22710
rect 5104 22708 5152 22710
rect 4008 22698 5208 22708
rect 4172 22596 4228 22606
rect 4172 22502 4228 22540
rect 4844 22370 4900 22382
rect 4844 22318 4846 22370
rect 4898 22318 4900 22370
rect 3836 22146 3892 22158
rect 3836 22094 3838 22146
rect 3890 22094 3892 22146
rect 3836 21700 3892 22094
rect 4844 22148 4900 22318
rect 4844 22082 4900 22092
rect 4956 22258 5012 22270
rect 4956 22206 4958 22258
rect 5010 22206 5012 22258
rect 4844 21812 4900 21822
rect 4844 21718 4900 21756
rect 3836 21634 3892 21644
rect 4956 21364 5012 22206
rect 5292 22148 5348 23100
rect 5404 23268 5460 23278
rect 5404 22820 5460 23212
rect 5852 23156 5908 26014
rect 5964 26068 6020 26078
rect 5964 25730 6020 26012
rect 5964 25678 5966 25730
rect 6018 25678 6020 25730
rect 5964 25666 6020 25678
rect 6076 25732 6132 26572
rect 6188 26292 6244 27580
rect 6300 27076 6356 32620
rect 6412 30434 6468 33516
rect 6524 32674 6580 33964
rect 6748 33460 6804 34862
rect 6860 34132 6916 44604
rect 6972 43764 7028 45836
rect 7196 45444 7252 45454
rect 7196 44100 7252 45388
rect 7308 45332 7364 45836
rect 7308 45266 7364 45276
rect 7308 44994 7364 45006
rect 7308 44942 7310 44994
rect 7362 44942 7364 44994
rect 7308 44772 7364 44942
rect 7308 44706 7364 44716
rect 7308 44436 7364 44446
rect 7308 44322 7364 44380
rect 7308 44270 7310 44322
rect 7362 44270 7364 44322
rect 7308 44258 7364 44270
rect 7420 44212 7476 46508
rect 7756 46450 7812 46508
rect 7756 46398 7758 46450
rect 7810 46398 7812 46450
rect 7756 46386 7812 46398
rect 7644 45892 7700 45902
rect 7532 45890 7700 45892
rect 7532 45838 7646 45890
rect 7698 45838 7700 45890
rect 7532 45836 7700 45838
rect 7532 44434 7588 45836
rect 7644 45826 7700 45836
rect 7644 45332 7700 45342
rect 7644 45330 7812 45332
rect 7644 45278 7646 45330
rect 7698 45278 7812 45330
rect 7644 45276 7812 45278
rect 7644 45266 7700 45276
rect 7644 45108 7700 45118
rect 7644 44772 7700 45052
rect 7644 44706 7700 44716
rect 7644 44548 7700 44558
rect 7756 44548 7812 45276
rect 7644 44546 7812 44548
rect 7644 44494 7646 44546
rect 7698 44494 7812 44546
rect 7644 44492 7812 44494
rect 7644 44482 7700 44492
rect 7868 44436 7924 48076
rect 8092 47236 8148 47246
rect 8092 47142 8148 47180
rect 8204 46562 8260 46574
rect 8204 46510 8206 46562
rect 8258 46510 8260 46562
rect 7980 46450 8036 46462
rect 7980 46398 7982 46450
rect 8034 46398 8036 46450
rect 7980 45108 8036 46398
rect 8204 45444 8260 46510
rect 8204 45378 8260 45388
rect 7980 45042 8036 45052
rect 8204 45108 8260 45118
rect 8428 45108 8484 45118
rect 8652 45108 8708 49756
rect 8764 47684 8820 50372
rect 8876 50372 9156 50428
rect 8876 49588 8932 50372
rect 8876 49586 9044 49588
rect 8876 49534 8878 49586
rect 8930 49534 9044 49586
rect 8876 49532 9044 49534
rect 8876 49522 8932 49532
rect 8988 48132 9044 49532
rect 8988 48038 9044 48076
rect 8764 47618 8820 47628
rect 9100 47348 9156 47358
rect 9100 47254 9156 47292
rect 9100 46564 9156 46574
rect 9100 46470 9156 46508
rect 9324 46004 9380 52780
rect 9548 50428 9604 56812
rect 9660 56532 9716 56542
rect 9660 56306 9716 56476
rect 9660 56254 9662 56306
rect 9714 56254 9716 56306
rect 9660 56242 9716 56254
rect 9660 54290 9716 54302
rect 9660 54238 9662 54290
rect 9714 54238 9716 54290
rect 9660 54068 9716 54238
rect 9660 54002 9716 54012
rect 9772 53732 9828 53742
rect 9772 52274 9828 53676
rect 9772 52222 9774 52274
rect 9826 52222 9828 52274
rect 9772 52210 9828 52222
rect 9660 51940 9716 51950
rect 9660 51268 9716 51884
rect 9660 51266 9828 51268
rect 9660 51214 9662 51266
rect 9714 51214 9828 51266
rect 9660 51212 9828 51214
rect 9660 51202 9716 51212
rect 9436 50372 9604 50428
rect 9436 48580 9492 50372
rect 9660 50036 9716 50046
rect 9660 49942 9716 49980
rect 9772 49700 9828 51212
rect 9772 48802 9828 49644
rect 9772 48750 9774 48802
rect 9826 48750 9828 48802
rect 9772 48738 9828 48750
rect 9436 48514 9492 48524
rect 9884 48468 9940 61292
rect 9996 62244 10052 62254
rect 9996 60676 10052 62188
rect 10108 60900 10164 62860
rect 10220 62354 10276 62366
rect 10220 62302 10222 62354
rect 10274 62302 10276 62354
rect 10220 62132 10276 62302
rect 10332 62188 10388 66332
rect 10668 65492 10724 65502
rect 10668 65398 10724 65436
rect 10780 65156 10836 66780
rect 10668 65100 10836 65156
rect 10444 64820 10500 64830
rect 10444 63812 10500 64764
rect 10668 64818 10724 65100
rect 10668 64766 10670 64818
rect 10722 64766 10724 64818
rect 10668 64754 10724 64766
rect 10892 64596 10948 68460
rect 11004 66500 11060 66510
rect 11004 66406 11060 66444
rect 11116 65940 11172 69916
rect 11676 69634 11732 70140
rect 12012 69860 12068 74620
rect 12460 74340 12516 74734
rect 12124 74284 12516 74340
rect 12572 74338 12628 74844
rect 12572 74286 12574 74338
rect 12626 74286 12628 74338
rect 12124 73330 12180 74284
rect 12572 74274 12628 74286
rect 12236 74116 12292 74126
rect 12796 74116 12852 75292
rect 12908 74898 12964 74910
rect 12908 74846 12910 74898
rect 12962 74846 12964 74898
rect 12908 74338 12964 74846
rect 12908 74286 12910 74338
rect 12962 74286 12964 74338
rect 12908 74274 12964 74286
rect 12236 74114 12852 74116
rect 12236 74062 12238 74114
rect 12290 74062 12852 74114
rect 12236 74060 12852 74062
rect 12236 74050 12292 74060
rect 12124 73278 12126 73330
rect 12178 73278 12180 73330
rect 12124 73266 12180 73278
rect 12796 74002 12852 74060
rect 12796 73950 12798 74002
rect 12850 73950 12852 74002
rect 12012 69804 12180 69860
rect 11676 69582 11678 69634
rect 11730 69582 11732 69634
rect 11676 69570 11732 69582
rect 12012 69636 12068 69646
rect 12012 69542 12068 69580
rect 11900 69300 11956 69310
rect 11788 69244 11900 69300
rect 11228 69188 11284 69198
rect 11284 69132 11732 69188
rect 11228 69094 11284 69132
rect 11676 68738 11732 69132
rect 11788 68850 11844 69244
rect 11900 69234 11956 69244
rect 11788 68798 11790 68850
rect 11842 68798 11844 68850
rect 11788 68786 11844 68798
rect 11676 68686 11678 68738
rect 11730 68686 11732 68738
rect 11676 68674 11732 68686
rect 11900 68740 11956 68750
rect 12124 68740 12180 69804
rect 12236 69298 12292 69310
rect 12236 69246 12238 69298
rect 12290 69246 12292 69298
rect 12236 69188 12292 69246
rect 12236 69122 12292 69132
rect 12572 69300 12628 69310
rect 12796 69300 12852 73950
rect 13020 73780 13076 76524
rect 13020 73714 13076 73724
rect 13132 75012 13188 75022
rect 13132 70420 13188 74956
rect 12572 69298 12852 69300
rect 12572 69246 12574 69298
rect 12626 69246 12852 69298
rect 12572 69244 12852 69246
rect 13020 70364 13188 70420
rect 11900 68738 12180 68740
rect 11900 68686 11902 68738
rect 11954 68686 12180 68738
rect 11900 68684 12180 68686
rect 11452 68514 11508 68526
rect 11452 68462 11454 68514
rect 11506 68462 11508 68514
rect 11228 67620 11284 67630
rect 11228 67060 11284 67564
rect 11452 67284 11508 68462
rect 11900 68516 11956 68684
rect 11900 68450 11956 68460
rect 12236 68626 12292 68638
rect 12236 68574 12238 68626
rect 12290 68574 12292 68626
rect 11452 67218 11508 67228
rect 12236 67284 12292 68574
rect 12572 67620 12628 69244
rect 12908 69188 12964 69198
rect 12908 68626 12964 69132
rect 12908 68574 12910 68626
rect 12962 68574 12964 68626
rect 12908 68562 12964 68574
rect 12572 67554 12628 67564
rect 12236 67218 12292 67228
rect 12572 67282 12628 67294
rect 12572 67230 12574 67282
rect 12626 67230 12628 67282
rect 12572 67172 12628 67230
rect 12460 67116 12572 67172
rect 11676 67060 11732 67070
rect 11228 67004 11508 67060
rect 11228 66164 11284 66174
rect 11284 66108 11396 66164
rect 11228 66070 11284 66108
rect 11116 65884 11284 65940
rect 11116 65492 11172 65502
rect 10444 63746 10500 63756
rect 10668 64540 10948 64596
rect 11004 64818 11060 64830
rect 11004 64766 11006 64818
rect 11058 64766 11060 64818
rect 10444 63364 10500 63374
rect 10444 62466 10500 63308
rect 10444 62414 10446 62466
rect 10498 62414 10500 62466
rect 10444 62402 10500 62414
rect 10332 62132 10500 62188
rect 10220 62066 10276 62076
rect 10332 61572 10388 61582
rect 10332 61478 10388 61516
rect 10108 60844 10276 60900
rect 10108 60676 10164 60686
rect 9996 60620 10108 60676
rect 10108 60582 10164 60620
rect 10220 58548 10276 60844
rect 10220 58482 10276 58492
rect 9996 57426 10052 57438
rect 9996 57374 9998 57426
rect 10050 57374 10052 57426
rect 9996 56868 10052 57374
rect 9996 56802 10052 56812
rect 10444 56644 10500 62132
rect 10556 57764 10612 57774
rect 10556 57670 10612 57708
rect 10108 56308 10164 56318
rect 10108 55970 10164 56252
rect 10108 55918 10110 55970
rect 10162 55918 10164 55970
rect 10108 55524 10164 55918
rect 10444 55972 10500 56588
rect 10556 56642 10612 56654
rect 10556 56590 10558 56642
rect 10610 56590 10612 56642
rect 10556 56532 10612 56590
rect 10556 56466 10612 56476
rect 10668 56196 10724 64540
rect 11004 63364 11060 64766
rect 11116 64594 11172 65436
rect 11116 64542 11118 64594
rect 11170 64542 11172 64594
rect 11116 64530 11172 64542
rect 11228 64372 11284 65884
rect 11340 64932 11396 66108
rect 11340 64838 11396 64876
rect 11004 63298 11060 63308
rect 11116 64316 11284 64372
rect 10892 62916 10948 62926
rect 10892 62356 10948 62860
rect 10892 62290 10948 62300
rect 11116 62188 11172 64316
rect 10892 62132 11172 62188
rect 11228 62354 11284 62366
rect 11228 62302 11230 62354
rect 11282 62302 11284 62354
rect 10780 61348 10836 61358
rect 10780 61254 10836 61292
rect 10444 55906 10500 55916
rect 10556 56140 10724 56196
rect 10780 57650 10836 57662
rect 10780 57598 10782 57650
rect 10834 57598 10836 57650
rect 10780 57540 10836 57598
rect 10780 57204 10836 57484
rect 10556 55636 10612 56140
rect 10108 55458 10164 55468
rect 10332 55580 10612 55636
rect 10668 55972 10724 55982
rect 10108 55298 10164 55310
rect 10108 55246 10110 55298
rect 10162 55246 10164 55298
rect 10108 55188 10164 55246
rect 10220 55188 10276 55198
rect 10108 55132 10220 55188
rect 10108 54964 10164 54974
rect 9996 54740 10052 54750
rect 9996 54514 10052 54684
rect 9996 54462 9998 54514
rect 10050 54462 10052 54514
rect 9996 54450 10052 54462
rect 10108 53172 10164 54908
rect 10108 53106 10164 53116
rect 10220 54404 10276 55132
rect 10108 52946 10164 52958
rect 10108 52894 10110 52946
rect 10162 52894 10164 52946
rect 10108 52276 10164 52894
rect 10108 52210 10164 52220
rect 10220 50036 10276 54348
rect 10332 53844 10388 55580
rect 10668 55188 10724 55916
rect 10668 55122 10724 55132
rect 10780 54852 10836 57148
rect 10332 53284 10388 53788
rect 10668 54796 10836 54852
rect 10892 54852 10948 62132
rect 11228 61908 11284 62302
rect 11452 62188 11508 67004
rect 11676 66388 11732 67004
rect 11676 66162 11732 66332
rect 11676 66110 11678 66162
rect 11730 66110 11732 66162
rect 11676 66098 11732 66110
rect 11788 64932 11844 64942
rect 11788 64818 11844 64876
rect 11788 64766 11790 64818
rect 11842 64766 11844 64818
rect 11788 64754 11844 64766
rect 12236 64932 12292 64942
rect 11228 61842 11284 61852
rect 11340 62132 11508 62188
rect 12012 64484 12068 64494
rect 11004 61572 11060 61582
rect 11340 61572 11396 62132
rect 11004 61236 11060 61516
rect 11228 61516 11396 61572
rect 11452 61682 11508 61694
rect 11452 61630 11454 61682
rect 11506 61630 11508 61682
rect 11452 61572 11508 61630
rect 11788 61572 11844 61582
rect 11452 61570 11844 61572
rect 11452 61518 11790 61570
rect 11842 61518 11844 61570
rect 11452 61516 11844 61518
rect 11116 61458 11172 61470
rect 11116 61406 11118 61458
rect 11170 61406 11172 61458
rect 11116 61348 11172 61406
rect 11116 61282 11172 61292
rect 11004 55076 11060 61180
rect 11116 57204 11172 57214
rect 11116 55410 11172 57148
rect 11116 55358 11118 55410
rect 11170 55358 11172 55410
rect 11116 55346 11172 55358
rect 11004 55010 11060 55020
rect 10892 54796 11172 54852
rect 10668 54514 10724 54796
rect 10668 54462 10670 54514
rect 10722 54462 10724 54514
rect 10668 53620 10724 54462
rect 10780 54628 10836 54638
rect 10780 53732 10836 54572
rect 10780 53676 11060 53732
rect 10668 53554 10724 53564
rect 10892 53508 10948 53518
rect 10892 53414 10948 53452
rect 10332 53228 10500 53284
rect 10220 48804 10276 49980
rect 10332 49700 10388 49710
rect 10332 49606 10388 49644
rect 10332 48804 10388 48814
rect 10220 48802 10388 48804
rect 10220 48750 10334 48802
rect 10386 48750 10388 48802
rect 10220 48748 10388 48750
rect 9884 48412 10164 48468
rect 9996 48244 10052 48254
rect 9996 48150 10052 48188
rect 9884 48132 9940 48142
rect 9884 48038 9940 48076
rect 9772 48018 9828 48030
rect 10108 48020 10164 48412
rect 9772 47966 9774 48018
rect 9826 47966 9828 48018
rect 9436 47234 9492 47246
rect 9436 47182 9438 47234
rect 9490 47182 9492 47234
rect 9436 47124 9492 47182
rect 9436 46676 9492 47068
rect 9436 46610 9492 46620
rect 9324 45938 9380 45948
rect 8204 45106 8372 45108
rect 8204 45054 8206 45106
rect 8258 45054 8372 45106
rect 8204 45052 8372 45054
rect 8204 45042 8260 45052
rect 7980 44882 8036 44894
rect 7980 44830 7982 44882
rect 8034 44830 8036 44882
rect 7980 44548 8036 44830
rect 8204 44548 8260 44558
rect 7980 44546 8260 44548
rect 7980 44494 8206 44546
rect 8258 44494 8260 44546
rect 7980 44492 8260 44494
rect 8204 44482 8260 44492
rect 7532 44382 7534 44434
rect 7586 44382 7588 44434
rect 7532 44370 7588 44382
rect 7756 44380 7924 44436
rect 7420 44156 7700 44212
rect 7196 44044 7364 44100
rect 6972 43698 7028 43708
rect 6972 43428 7028 43438
rect 6972 43426 7140 43428
rect 6972 43374 6974 43426
rect 7026 43374 7140 43426
rect 6972 43372 7140 43374
rect 6972 43362 7028 43372
rect 7084 43314 7140 43372
rect 7084 43262 7086 43314
rect 7138 43262 7140 43314
rect 6972 39396 7028 39406
rect 6972 39302 7028 39340
rect 6972 39060 7028 39070
rect 6972 37938 7028 39004
rect 6972 37886 6974 37938
rect 7026 37886 7028 37938
rect 6972 37874 7028 37886
rect 6860 34066 6916 34076
rect 6972 36596 7028 36606
rect 6972 35924 7028 36540
rect 7084 36484 7140 43262
rect 7196 42644 7252 42654
rect 7196 42194 7252 42588
rect 7196 42142 7198 42194
rect 7250 42142 7252 42194
rect 7196 42130 7252 42142
rect 7196 40740 7252 40750
rect 7196 39060 7252 40684
rect 7308 40178 7364 44044
rect 7308 40126 7310 40178
rect 7362 40126 7364 40178
rect 7308 40114 7364 40126
rect 7420 42868 7476 42878
rect 7420 40628 7476 42812
rect 7420 40068 7476 40572
rect 7532 41188 7588 41198
rect 7532 40962 7588 41132
rect 7532 40910 7534 40962
rect 7586 40910 7588 40962
rect 7532 40292 7588 40910
rect 7532 40226 7588 40236
rect 7420 40012 7588 40068
rect 7308 39620 7364 39630
rect 7364 39564 7476 39620
rect 7308 39526 7364 39564
rect 7308 39060 7364 39070
rect 7196 39058 7364 39060
rect 7196 39006 7310 39058
rect 7362 39006 7364 39058
rect 7196 39004 7364 39006
rect 7308 37828 7364 39004
rect 7308 37762 7364 37772
rect 7084 36418 7140 36428
rect 7420 37380 7476 39564
rect 7084 36036 7140 36046
rect 7084 35924 7140 35980
rect 6972 35922 7140 35924
rect 6972 35870 7086 35922
rect 7138 35870 7140 35922
rect 6972 35868 7140 35870
rect 6972 34244 7028 35868
rect 7084 35858 7140 35868
rect 7420 35812 7476 37324
rect 7532 39506 7588 40012
rect 7532 39454 7534 39506
rect 7586 39454 7588 39506
rect 7532 39172 7588 39454
rect 7532 36596 7588 39116
rect 7532 36530 7588 36540
rect 7532 36260 7588 36270
rect 7644 36260 7700 44156
rect 7756 39284 7812 44380
rect 8092 44324 8148 44334
rect 8092 43764 8148 44268
rect 7980 41188 8036 41198
rect 8092 41188 8148 43708
rect 8316 44324 8372 45052
rect 8428 45106 8708 45108
rect 8428 45054 8430 45106
rect 8482 45054 8708 45106
rect 8428 45052 8708 45054
rect 9660 45108 9716 45118
rect 8428 45042 8484 45052
rect 8540 44548 8596 45052
rect 8876 44994 8932 45006
rect 8876 44942 8878 44994
rect 8930 44942 8932 44994
rect 8876 44548 8932 44942
rect 8540 44546 8932 44548
rect 8540 44494 8542 44546
rect 8594 44494 8932 44546
rect 8540 44492 8932 44494
rect 8540 44482 8596 44492
rect 8204 43428 8260 43438
rect 8204 43334 8260 43372
rect 8204 42868 8260 42878
rect 8316 42868 8372 44268
rect 8764 44322 8820 44334
rect 8764 44270 8766 44322
rect 8818 44270 8820 44322
rect 8764 43762 8820 44270
rect 8876 44100 8932 44492
rect 9660 44434 9716 45052
rect 9660 44382 9662 44434
rect 9714 44382 9716 44434
rect 9660 44324 9716 44382
rect 9212 44100 9268 44110
rect 8876 44098 9380 44100
rect 8876 44046 9214 44098
rect 9266 44046 9380 44098
rect 8876 44044 9380 44046
rect 9212 44034 9268 44044
rect 8764 43710 8766 43762
rect 8818 43710 8820 43762
rect 8764 43698 8820 43710
rect 8540 43538 8596 43550
rect 8540 43486 8542 43538
rect 8594 43486 8596 43538
rect 8540 43428 8596 43486
rect 8204 42866 8372 42868
rect 8204 42814 8206 42866
rect 8258 42814 8372 42866
rect 8204 42812 8372 42814
rect 8428 43372 8540 43428
rect 8204 42644 8260 42812
rect 8428 42644 8484 43372
rect 8540 43362 8596 43372
rect 8876 43316 8932 43326
rect 8652 43314 8932 43316
rect 8652 43262 8878 43314
rect 8930 43262 8932 43314
rect 8652 43260 8932 43262
rect 8540 42868 8596 42878
rect 8540 42774 8596 42812
rect 8652 42756 8708 43260
rect 8876 43250 8932 43260
rect 9212 42980 9268 42990
rect 8876 42868 8932 42878
rect 9100 42868 9156 42878
rect 8932 42866 9156 42868
rect 8932 42814 9102 42866
rect 9154 42814 9156 42866
rect 8932 42812 9156 42814
rect 8876 42802 8932 42812
rect 9100 42802 9156 42812
rect 8652 42700 8820 42756
rect 8428 42588 8596 42644
rect 8204 42578 8260 42588
rect 8428 41972 8484 41982
rect 8428 41878 8484 41916
rect 8036 41132 8148 41188
rect 7980 41122 8036 41132
rect 8092 41074 8148 41132
rect 8316 41860 8372 41870
rect 8316 41186 8372 41804
rect 8316 41134 8318 41186
rect 8370 41134 8372 41186
rect 8316 41122 8372 41134
rect 8540 41188 8596 42588
rect 8652 42532 8708 42542
rect 8652 42438 8708 42476
rect 8652 42196 8708 42206
rect 8764 42196 8820 42700
rect 9212 42754 9268 42924
rect 9212 42702 9214 42754
rect 9266 42702 9268 42754
rect 8988 42532 9044 42542
rect 8652 42194 8820 42196
rect 8652 42142 8654 42194
rect 8706 42142 8820 42194
rect 8652 42140 8820 42142
rect 8876 42530 9044 42532
rect 8876 42478 8990 42530
rect 9042 42478 9044 42530
rect 8876 42476 9044 42478
rect 8652 42130 8708 42140
rect 8876 42082 8932 42476
rect 8988 42466 9044 42476
rect 9212 42196 9268 42702
rect 9212 42130 9268 42140
rect 8876 42030 8878 42082
rect 8930 42030 8932 42082
rect 8540 41186 8820 41188
rect 8540 41134 8542 41186
rect 8594 41134 8820 41186
rect 8540 41132 8820 41134
rect 8540 41122 8596 41132
rect 8092 41022 8094 41074
rect 8146 41022 8148 41074
rect 8092 41010 8148 41022
rect 8204 41076 8260 41086
rect 8204 40982 8260 41020
rect 7980 40964 8036 40974
rect 7980 40870 8036 40908
rect 7980 40628 8036 40638
rect 7980 40534 8036 40572
rect 8764 40628 8820 41132
rect 8876 41076 8932 42030
rect 8988 41972 9044 41982
rect 9212 41972 9268 41982
rect 9324 41972 9380 44044
rect 9660 42868 9716 44268
rect 9660 42754 9716 42812
rect 9660 42702 9662 42754
rect 9714 42702 9716 42754
rect 9660 42690 9716 42702
rect 9660 42532 9716 42542
rect 9660 42082 9716 42476
rect 9660 42030 9662 42082
rect 9714 42030 9716 42082
rect 9660 42018 9716 42030
rect 8988 41970 9156 41972
rect 8988 41918 8990 41970
rect 9042 41918 9156 41970
rect 8988 41916 9156 41918
rect 8988 41906 9044 41916
rect 9100 41188 9156 41916
rect 9268 41916 9380 41972
rect 9548 41970 9604 41982
rect 9548 41918 9550 41970
rect 9602 41918 9604 41970
rect 9212 41906 9268 41916
rect 9548 41298 9604 41918
rect 9772 41860 9828 47966
rect 9996 47964 10164 48020
rect 9884 47684 9940 47694
rect 9884 47590 9940 47628
rect 9996 46900 10052 47964
rect 10220 47908 10276 48748
rect 10332 48738 10388 48748
rect 9548 41246 9550 41298
rect 9602 41246 9604 41298
rect 9548 41234 9604 41246
rect 9660 41804 9772 41860
rect 9436 41188 9492 41198
rect 9100 41186 9492 41188
rect 9100 41134 9438 41186
rect 9490 41134 9492 41186
rect 9100 41132 9492 41134
rect 8988 41076 9044 41086
rect 8876 41074 9268 41076
rect 8876 41022 8990 41074
rect 9042 41022 9268 41074
rect 8876 41020 9268 41022
rect 8988 41010 9044 41020
rect 8876 40628 8932 40638
rect 8820 40626 8932 40628
rect 8820 40574 8878 40626
rect 8930 40574 8932 40626
rect 8820 40572 8932 40574
rect 8764 40534 8820 40572
rect 8876 40562 8932 40572
rect 7868 40516 7924 40526
rect 7868 39506 7924 40460
rect 8316 40516 8372 40526
rect 8316 40422 8372 40460
rect 8204 40178 8260 40190
rect 8204 40126 8206 40178
rect 8258 40126 8260 40178
rect 7868 39454 7870 39506
rect 7922 39454 7924 39506
rect 7868 39442 7924 39454
rect 7980 40068 8036 40078
rect 7756 39228 7924 39284
rect 7868 36596 7924 39228
rect 7980 38668 8036 40012
rect 8092 39060 8148 39070
rect 8092 38966 8148 39004
rect 7980 38612 8148 38668
rect 7868 36540 8036 36596
rect 7588 36204 7700 36260
rect 7868 36372 7924 36382
rect 7532 36166 7588 36204
rect 7868 35922 7924 36316
rect 7868 35870 7870 35922
rect 7922 35870 7924 35922
rect 7868 35858 7924 35870
rect 7196 35756 7476 35812
rect 7196 35028 7252 35756
rect 7196 34962 7252 34972
rect 7420 35588 7476 35598
rect 7756 35588 7812 35598
rect 7308 34916 7364 34954
rect 7308 34850 7364 34860
rect 7084 34804 7140 34814
rect 7084 34354 7140 34748
rect 7084 34302 7086 34354
rect 7138 34302 7140 34354
rect 7084 34290 7140 34302
rect 7308 34468 7364 34478
rect 7308 34354 7364 34412
rect 7308 34302 7310 34354
rect 7362 34302 7364 34354
rect 7308 34290 7364 34302
rect 6972 33908 7028 34188
rect 7420 34242 7476 35532
rect 7420 34190 7422 34242
rect 7474 34190 7476 34242
rect 7420 34178 7476 34190
rect 7532 35586 7812 35588
rect 7532 35534 7758 35586
rect 7810 35534 7812 35586
rect 7532 35532 7812 35534
rect 7196 34132 7252 34142
rect 6636 33236 6692 33246
rect 6636 33142 6692 33180
rect 6524 32622 6526 32674
rect 6578 32622 6580 32674
rect 6524 32610 6580 32622
rect 6636 32674 6692 32686
rect 6636 32622 6638 32674
rect 6690 32622 6692 32674
rect 6636 32452 6692 32622
rect 6636 32386 6692 32396
rect 6412 30382 6414 30434
rect 6466 30382 6468 30434
rect 6412 30370 6468 30382
rect 6524 31892 6580 31902
rect 6412 27860 6468 27870
rect 6412 27766 6468 27804
rect 6412 27300 6468 27310
rect 6412 27206 6468 27244
rect 6300 27010 6356 27020
rect 6412 26292 6468 26302
rect 6188 26290 6468 26292
rect 6188 26238 6414 26290
rect 6466 26238 6468 26290
rect 6188 26236 6468 26238
rect 6412 26226 6468 26236
rect 6300 26066 6356 26078
rect 6524 26068 6580 31836
rect 6748 30882 6804 33404
rect 6860 33852 7028 33908
rect 7084 34020 7140 34030
rect 6860 33346 6916 33852
rect 6860 33294 6862 33346
rect 6914 33294 6916 33346
rect 6860 33012 6916 33294
rect 6860 32946 6916 32956
rect 6860 32788 6916 32798
rect 7084 32788 7140 33964
rect 6860 32786 7140 32788
rect 6860 32734 6862 32786
rect 6914 32734 7140 32786
rect 6860 32732 7140 32734
rect 6860 32722 6916 32732
rect 7196 32116 7252 34076
rect 7532 34132 7588 35532
rect 7756 35522 7812 35532
rect 7644 34692 7700 34702
rect 7644 34468 7700 34636
rect 7644 34402 7700 34412
rect 7532 33346 7588 34076
rect 7532 33294 7534 33346
rect 7586 33294 7588 33346
rect 7420 33236 7476 33246
rect 7532 33236 7588 33294
rect 7476 33180 7588 33236
rect 7644 34244 7700 34254
rect 7420 33170 7476 33180
rect 7532 32452 7588 32462
rect 7532 32358 7588 32396
rect 6748 30830 6750 30882
rect 6802 30830 6804 30882
rect 6748 28196 6804 30830
rect 6972 32060 7252 32116
rect 6748 28130 6804 28140
rect 6860 29540 6916 29550
rect 6748 27972 6804 27982
rect 6860 27972 6916 29484
rect 6748 27970 6916 27972
rect 6748 27918 6750 27970
rect 6802 27918 6916 27970
rect 6748 27916 6916 27918
rect 6972 28642 7028 32060
rect 7532 31892 7588 31902
rect 7420 31836 7532 31892
rect 7308 31554 7364 31566
rect 7308 31502 7310 31554
rect 7362 31502 7364 31554
rect 7308 30996 7364 31502
rect 7308 30930 7364 30940
rect 7308 30212 7364 30222
rect 7420 30212 7476 31836
rect 7532 31826 7588 31836
rect 7644 31556 7700 34188
rect 7868 34020 7924 34058
rect 7868 33954 7924 33964
rect 7980 32788 8036 36540
rect 8092 34130 8148 38556
rect 8204 34244 8260 40126
rect 8764 39620 8820 39630
rect 8652 39172 8708 39182
rect 8652 39058 8708 39116
rect 8652 39006 8654 39058
rect 8706 39006 8708 39058
rect 8652 38994 8708 39006
rect 8316 38836 8372 38846
rect 8372 38780 8484 38836
rect 8316 38770 8372 38780
rect 8428 37826 8484 38780
rect 8652 38276 8708 38286
rect 8428 37774 8430 37826
rect 8482 37774 8484 37826
rect 8428 36596 8484 37774
rect 8428 36530 8484 36540
rect 8540 38220 8652 38276
rect 8316 36484 8372 36494
rect 8316 36258 8372 36428
rect 8316 36206 8318 36258
rect 8370 36206 8372 36258
rect 8316 35812 8372 36206
rect 8428 35812 8484 35822
rect 8316 35810 8484 35812
rect 8316 35758 8430 35810
rect 8482 35758 8484 35810
rect 8316 35756 8484 35758
rect 8428 35700 8484 35756
rect 8428 35634 8484 35644
rect 8204 34178 8260 34188
rect 8428 34356 8484 34366
rect 8092 34078 8094 34130
rect 8146 34078 8148 34130
rect 8092 32900 8148 34078
rect 8428 34130 8484 34300
rect 8428 34078 8430 34130
rect 8482 34078 8484 34130
rect 8428 34066 8484 34078
rect 8204 34020 8260 34030
rect 8204 34018 8372 34020
rect 8204 33966 8206 34018
rect 8258 33966 8372 34018
rect 8204 33964 8372 33966
rect 8204 33954 8260 33964
rect 8316 33348 8372 33964
rect 8540 33908 8596 38220
rect 8652 38210 8708 38220
rect 8764 37378 8820 39564
rect 8988 39396 9044 39406
rect 8988 38724 9044 39340
rect 8988 38658 9044 38668
rect 9212 38668 9268 41020
rect 9324 40628 9380 40638
rect 9324 39732 9380 40572
rect 9436 40516 9492 41132
rect 9660 40964 9716 41804
rect 9772 41794 9828 41804
rect 9884 46844 10052 46900
rect 10108 47852 10276 47908
rect 9660 40908 9828 40964
rect 9548 40516 9604 40526
rect 9436 40514 9604 40516
rect 9436 40462 9550 40514
rect 9602 40462 9604 40514
rect 9436 40460 9604 40462
rect 9548 40450 9604 40460
rect 9660 40402 9716 40414
rect 9660 40350 9662 40402
rect 9714 40350 9716 40402
rect 9436 39732 9492 39742
rect 9324 39730 9492 39732
rect 9324 39678 9438 39730
rect 9490 39678 9492 39730
rect 9324 39676 9492 39678
rect 9436 39666 9492 39676
rect 9660 39620 9716 40350
rect 9660 39554 9716 39564
rect 9772 39618 9828 40908
rect 9772 39566 9774 39618
rect 9826 39566 9828 39618
rect 9772 39554 9828 39566
rect 9436 39394 9492 39406
rect 9436 39342 9438 39394
rect 9490 39342 9492 39394
rect 9436 39060 9492 39342
rect 9548 39396 9604 39406
rect 9548 39302 9604 39340
rect 9436 38994 9492 39004
rect 9212 38612 9828 38668
rect 9660 37940 9716 37950
rect 9100 37938 9716 37940
rect 9100 37886 9662 37938
rect 9714 37886 9716 37938
rect 9100 37884 9716 37886
rect 8876 37828 8932 37838
rect 8932 37772 9044 37828
rect 8876 37734 8932 37772
rect 8764 37326 8766 37378
rect 8818 37326 8820 37378
rect 8764 36594 8820 37326
rect 8764 36542 8766 36594
rect 8818 36542 8820 36594
rect 8764 36530 8820 36542
rect 8876 37378 8932 37390
rect 8876 37326 8878 37378
rect 8930 37326 8932 37378
rect 8764 36372 8820 36382
rect 8764 36278 8820 36316
rect 8876 36148 8932 37326
rect 8988 37268 9044 37772
rect 9100 37490 9156 37884
rect 9660 37874 9716 37884
rect 9100 37438 9102 37490
rect 9154 37438 9156 37490
rect 9100 37426 9156 37438
rect 9772 37826 9828 38612
rect 9884 38276 9940 46844
rect 9996 46676 10052 46686
rect 9996 46582 10052 46620
rect 9996 45666 10052 45678
rect 9996 45614 9998 45666
rect 10050 45614 10052 45666
rect 9996 45220 10052 45614
rect 9996 45154 10052 45164
rect 10108 44324 10164 47852
rect 10444 45892 10500 53228
rect 10780 52948 10836 52958
rect 10556 52724 10612 52734
rect 10556 52274 10612 52668
rect 10556 52222 10558 52274
rect 10610 52222 10612 52274
rect 10556 52210 10612 52222
rect 10780 49810 10836 52892
rect 11004 52836 11060 53676
rect 11004 52770 11060 52780
rect 11004 52276 11060 52286
rect 11004 52182 11060 52220
rect 10892 52052 10948 52062
rect 10892 51958 10948 51996
rect 10780 49758 10782 49810
rect 10834 49758 10836 49810
rect 10780 49746 10836 49758
rect 11004 48468 11060 48478
rect 11004 48374 11060 48412
rect 11116 48244 11172 54796
rect 11228 53284 11284 61516
rect 11788 61506 11844 61516
rect 12012 61570 12068 64428
rect 12236 64482 12292 64876
rect 12236 64430 12238 64482
rect 12290 64430 12292 64482
rect 12236 64372 12292 64430
rect 12236 64306 12292 64316
rect 12460 64146 12516 67116
rect 12572 67106 12628 67116
rect 12796 65378 12852 65390
rect 12796 65326 12798 65378
rect 12850 65326 12852 65378
rect 12796 65268 12852 65326
rect 12796 65202 12852 65212
rect 13020 65156 13076 70364
rect 13244 67620 13300 78876
rect 13356 77252 13412 79100
rect 13580 78932 13636 82012
rect 14364 81956 14420 82798
rect 14476 82740 14532 82750
rect 14476 82646 14532 82684
rect 15148 82292 15204 82908
rect 14476 82068 14532 82078
rect 14476 81974 14532 82012
rect 14364 81890 14420 81900
rect 15036 81956 15092 81966
rect 15148 81956 15204 82236
rect 15036 81954 15204 81956
rect 15036 81902 15038 81954
rect 15090 81902 15204 81954
rect 15036 81900 15204 81902
rect 15260 82852 15316 82862
rect 15260 81954 15316 82796
rect 15372 82740 15428 83356
rect 15372 82674 15428 82684
rect 15484 82626 15540 84140
rect 15932 83524 15988 83534
rect 15932 82962 15988 83468
rect 15932 82910 15934 82962
rect 15986 82910 15988 82962
rect 15484 82574 15486 82626
rect 15538 82574 15540 82626
rect 15484 82514 15540 82574
rect 15708 82852 15764 82862
rect 15484 82462 15486 82514
rect 15538 82462 15540 82514
rect 15484 82450 15540 82462
rect 15596 82516 15652 82526
rect 15260 81902 15262 81954
rect 15314 81902 15316 81954
rect 15036 81890 15092 81900
rect 13692 81844 13748 81854
rect 13692 81750 13748 81788
rect 13804 81844 13860 81854
rect 14028 81844 14084 81854
rect 13804 81842 14028 81844
rect 13804 81790 13806 81842
rect 13858 81790 14028 81842
rect 13804 81788 14028 81790
rect 13804 81778 13860 81788
rect 14028 81778 14084 81788
rect 14812 81844 14868 81882
rect 14812 81778 14868 81788
rect 14700 81732 14756 81770
rect 14700 81666 14756 81676
rect 15260 81732 15316 81902
rect 15260 81666 15316 81676
rect 15372 82180 15428 82190
rect 14008 81564 15208 81574
rect 14064 81562 14112 81564
rect 14168 81562 14216 81564
rect 14076 81510 14112 81562
rect 14200 81510 14216 81562
rect 14064 81508 14112 81510
rect 14168 81508 14216 81510
rect 14272 81562 14320 81564
rect 14376 81562 14424 81564
rect 14480 81562 14528 81564
rect 14376 81510 14396 81562
rect 14480 81510 14520 81562
rect 14272 81508 14320 81510
rect 14376 81508 14424 81510
rect 14480 81508 14528 81510
rect 14584 81508 14632 81564
rect 14688 81562 14736 81564
rect 14792 81562 14840 81564
rect 14896 81562 14944 81564
rect 14696 81510 14736 81562
rect 14820 81510 14840 81562
rect 14688 81508 14736 81510
rect 14792 81508 14840 81510
rect 14896 81508 14944 81510
rect 15000 81562 15048 81564
rect 15104 81562 15152 81564
rect 15000 81510 15016 81562
rect 15104 81510 15140 81562
rect 15000 81508 15048 81510
rect 15104 81508 15152 81510
rect 14008 81498 15208 81508
rect 14700 81396 14756 81406
rect 14140 81172 14196 81182
rect 13916 81060 13972 81070
rect 13916 80500 13972 81004
rect 13356 77186 13412 77196
rect 13468 78876 13636 78932
rect 13692 80444 13916 80500
rect 13692 79602 13748 80444
rect 13916 80406 13972 80444
rect 14140 80386 14196 81116
rect 14140 80334 14142 80386
rect 14194 80334 14196 80386
rect 14140 80322 14196 80334
rect 14364 81058 14420 81070
rect 14364 81006 14366 81058
rect 14418 81006 14420 81058
rect 14364 80388 14420 81006
rect 14588 81060 14644 81070
rect 14364 80322 14420 80332
rect 14476 80612 14532 80622
rect 14476 80386 14532 80556
rect 14476 80334 14478 80386
rect 14530 80334 14532 80386
rect 14476 80322 14532 80334
rect 14588 80386 14644 81004
rect 14588 80334 14590 80386
rect 14642 80334 14644 80386
rect 14588 80322 14644 80334
rect 14700 80500 14756 81340
rect 15372 81394 15428 82124
rect 15372 81342 15374 81394
rect 15426 81342 15428 81394
rect 15372 81330 15428 81342
rect 15484 81842 15540 81854
rect 15484 81790 15486 81842
rect 15538 81790 15540 81842
rect 15484 81396 15540 81790
rect 15484 81330 15540 81340
rect 15036 81284 15092 81294
rect 14700 80386 14756 80444
rect 14700 80334 14702 80386
rect 14754 80334 14756 80386
rect 14700 80322 14756 80334
rect 14812 81170 14868 81182
rect 14812 81118 14814 81170
rect 14866 81118 14868 81170
rect 13692 79550 13694 79602
rect 13746 79550 13748 79602
rect 13692 78932 13748 79550
rect 13804 80274 13860 80286
rect 13804 80222 13806 80274
rect 13858 80222 13860 80274
rect 13804 79492 13860 80222
rect 13916 80164 13972 80202
rect 13916 80098 13972 80108
rect 14812 80164 14868 81118
rect 15036 81170 15092 81228
rect 15260 81284 15316 81294
rect 15260 81190 15316 81228
rect 15484 81172 15540 81182
rect 15036 81118 15038 81170
rect 15090 81118 15092 81170
rect 15036 81106 15092 81118
rect 15372 81170 15540 81172
rect 15372 81118 15486 81170
rect 15538 81118 15540 81170
rect 15372 81116 15540 81118
rect 15372 80724 15428 81116
rect 15484 81106 15540 81116
rect 15148 80668 15428 80724
rect 15148 80610 15204 80668
rect 15148 80558 15150 80610
rect 15202 80558 15204 80610
rect 15148 80546 15204 80558
rect 14812 80098 14868 80108
rect 15372 80388 15428 80398
rect 14008 79996 15208 80006
rect 14064 79994 14112 79996
rect 14168 79994 14216 79996
rect 14076 79942 14112 79994
rect 14200 79942 14216 79994
rect 14064 79940 14112 79942
rect 14168 79940 14216 79942
rect 14272 79994 14320 79996
rect 14376 79994 14424 79996
rect 14480 79994 14528 79996
rect 14376 79942 14396 79994
rect 14480 79942 14520 79994
rect 14272 79940 14320 79942
rect 14376 79940 14424 79942
rect 14480 79940 14528 79942
rect 14584 79940 14632 79996
rect 14688 79994 14736 79996
rect 14792 79994 14840 79996
rect 14896 79994 14944 79996
rect 14696 79942 14736 79994
rect 14820 79942 14840 79994
rect 14688 79940 14736 79942
rect 14792 79940 14840 79942
rect 14896 79940 14944 79942
rect 15000 79994 15048 79996
rect 15104 79994 15152 79996
rect 15000 79942 15016 79994
rect 15104 79942 15140 79994
rect 15000 79940 15048 79942
rect 15104 79940 15152 79942
rect 14008 79930 15208 79940
rect 15260 79828 15316 79838
rect 14140 79716 14196 79726
rect 13804 79398 13860 79436
rect 13916 79714 14196 79716
rect 13916 79662 14142 79714
rect 14194 79662 14196 79714
rect 13916 79660 14196 79662
rect 13916 79042 13972 79660
rect 14140 79650 14196 79660
rect 15148 79714 15204 79726
rect 15148 79662 15150 79714
rect 15202 79662 15204 79714
rect 13916 78990 13918 79042
rect 13970 78990 13972 79042
rect 13916 78978 13972 78990
rect 14252 79604 14308 79614
rect 13356 75796 13412 75806
rect 13356 75122 13412 75740
rect 13356 75070 13358 75122
rect 13410 75070 13412 75122
rect 13356 75058 13412 75070
rect 13468 73948 13524 78876
rect 13692 78866 13748 78876
rect 13916 78818 13972 78830
rect 13916 78766 13918 78818
rect 13970 78766 13972 78818
rect 13580 78706 13636 78718
rect 13580 78654 13582 78706
rect 13634 78654 13636 78706
rect 13580 78596 13636 78654
rect 13916 78708 13972 78766
rect 14252 78818 14308 79548
rect 15148 79492 15204 79662
rect 15260 79602 15316 79772
rect 15260 79550 15262 79602
rect 15314 79550 15316 79602
rect 15260 79538 15316 79550
rect 15148 79426 15204 79436
rect 15372 79044 15428 80332
rect 15596 79828 15652 82460
rect 15596 79762 15652 79772
rect 15708 79380 15764 82796
rect 15932 82404 15988 82910
rect 16268 83300 16324 83310
rect 16268 82852 16324 83244
rect 16492 83298 16548 84140
rect 16492 83246 16494 83298
rect 16546 83246 16548 83298
rect 16492 83234 16548 83246
rect 16268 82758 16324 82796
rect 16492 82738 16548 82750
rect 16492 82686 16494 82738
rect 16546 82686 16548 82738
rect 16044 82516 16100 82526
rect 16044 82514 16436 82516
rect 16044 82462 16046 82514
rect 16098 82462 16436 82514
rect 16044 82460 16436 82462
rect 16044 82450 16100 82460
rect 15820 82292 15988 82348
rect 15820 80388 15876 82292
rect 16380 82068 16436 82460
rect 16492 82292 16548 82686
rect 16492 82226 16548 82236
rect 16380 82012 16548 82068
rect 16156 81954 16212 81966
rect 16156 81902 16158 81954
rect 16210 81902 16212 81954
rect 16156 81844 16212 81902
rect 16268 81956 16324 81966
rect 16268 81862 16324 81900
rect 16156 81778 16212 81788
rect 16380 81730 16436 81742
rect 16380 81678 16382 81730
rect 16434 81678 16436 81730
rect 16380 81620 16436 81678
rect 16492 81732 16548 82012
rect 16604 81954 16660 85932
rect 16716 84196 16772 87612
rect 16940 87332 16996 87342
rect 16940 87218 16996 87276
rect 16940 87166 16942 87218
rect 16994 87166 16996 87218
rect 16940 87154 16996 87166
rect 17276 86434 17332 87948
rect 20412 87668 20468 87678
rect 17388 87442 17444 87454
rect 17388 87390 17390 87442
rect 17442 87390 17444 87442
rect 17388 87332 17444 87390
rect 17948 87444 18004 87454
rect 19404 87444 19460 87454
rect 17948 87442 18452 87444
rect 17948 87390 17950 87442
rect 18002 87390 18452 87442
rect 17948 87388 18452 87390
rect 17948 87378 18004 87388
rect 17388 87266 17444 87276
rect 18396 86882 18452 87388
rect 18396 86830 18398 86882
rect 18450 86830 18452 86882
rect 18396 86818 18452 86830
rect 18732 86658 18788 86670
rect 18732 86606 18734 86658
rect 18786 86606 18788 86658
rect 17276 86382 17278 86434
rect 17330 86382 17332 86434
rect 16828 85764 16884 85774
rect 16828 85670 16884 85708
rect 17276 85764 17332 86382
rect 18060 86434 18116 86446
rect 18060 86382 18062 86434
rect 18114 86382 18116 86434
rect 18060 85988 18116 86382
rect 18060 85922 18116 85932
rect 18284 86100 18340 86110
rect 18172 85764 18228 85774
rect 17276 85762 18228 85764
rect 17276 85710 18174 85762
rect 18226 85710 18228 85762
rect 17276 85708 18228 85710
rect 16716 84130 16772 84140
rect 17052 83300 17108 83310
rect 17052 83206 17108 83244
rect 16716 82964 16772 82974
rect 16716 82962 17108 82964
rect 16716 82910 16718 82962
rect 16770 82910 17108 82962
rect 16716 82908 17108 82910
rect 16716 82898 16772 82908
rect 16828 82740 16884 82750
rect 16828 82646 16884 82684
rect 16716 82404 16772 82414
rect 16716 82292 16772 82348
rect 16716 82236 16996 82292
rect 16604 81902 16606 81954
rect 16658 81902 16660 81954
rect 16604 81890 16660 81902
rect 16716 81956 16772 81966
rect 16492 81638 16548 81676
rect 15932 81564 16436 81620
rect 15932 81282 15988 81564
rect 16492 81508 16548 81518
rect 15932 81230 15934 81282
rect 15986 81230 15988 81282
rect 15932 81218 15988 81230
rect 16044 81396 16100 81406
rect 16044 81170 16100 81340
rect 16044 81118 16046 81170
rect 16098 81118 16100 81170
rect 16044 81106 16100 81118
rect 16492 81172 16548 81452
rect 16716 81396 16772 81900
rect 16940 81954 16996 82236
rect 16940 81902 16942 81954
rect 16994 81902 16996 81954
rect 16940 81890 16996 81902
rect 16716 81330 16772 81340
rect 17052 81844 17108 82908
rect 17052 81284 17108 81788
rect 17052 81218 17108 81228
rect 16492 81078 16548 81116
rect 16716 81172 16772 81182
rect 16716 81078 16772 81116
rect 15820 80294 15876 80332
rect 16268 81058 16324 81070
rect 16268 81006 16270 81058
rect 16322 81006 16324 81058
rect 16268 80386 16324 81006
rect 16268 80334 16270 80386
rect 16322 80334 16324 80386
rect 16268 80322 16324 80334
rect 16380 81060 16436 81070
rect 16380 79492 16436 81004
rect 16380 79426 16436 79436
rect 16716 80948 16772 80958
rect 15708 79324 16100 79380
rect 15372 78978 15428 78988
rect 14252 78766 14254 78818
rect 14306 78766 14308 78818
rect 14252 78754 14308 78766
rect 15596 78820 15652 78830
rect 15596 78818 15764 78820
rect 15596 78766 15598 78818
rect 15650 78766 15764 78818
rect 15596 78764 15764 78766
rect 15596 78754 15652 78764
rect 13916 78642 13972 78652
rect 15484 78706 15540 78718
rect 15484 78654 15486 78706
rect 15538 78654 15540 78706
rect 13580 78530 13636 78540
rect 14008 78428 15208 78438
rect 14064 78426 14112 78428
rect 14168 78426 14216 78428
rect 14076 78374 14112 78426
rect 14200 78374 14216 78426
rect 14064 78372 14112 78374
rect 14168 78372 14216 78374
rect 14272 78426 14320 78428
rect 14376 78426 14424 78428
rect 14480 78426 14528 78428
rect 14376 78374 14396 78426
rect 14480 78374 14520 78426
rect 14272 78372 14320 78374
rect 14376 78372 14424 78374
rect 14480 78372 14528 78374
rect 14584 78372 14632 78428
rect 14688 78426 14736 78428
rect 14792 78426 14840 78428
rect 14896 78426 14944 78428
rect 14696 78374 14736 78426
rect 14820 78374 14840 78426
rect 14688 78372 14736 78374
rect 14792 78372 14840 78374
rect 14896 78372 14944 78374
rect 15000 78426 15048 78428
rect 15104 78426 15152 78428
rect 15000 78374 15016 78426
rect 15104 78374 15140 78426
rect 15000 78372 15048 78374
rect 15104 78372 15152 78374
rect 14008 78362 15208 78372
rect 14700 78260 14756 78270
rect 13580 78148 13636 78158
rect 13580 77922 13636 78092
rect 13580 77870 13582 77922
rect 13634 77870 13636 77922
rect 13580 76468 13636 77870
rect 14588 77364 14644 77374
rect 13804 77252 13860 77262
rect 14028 77252 14084 77262
rect 13804 77158 13860 77196
rect 13916 77196 14028 77252
rect 13916 77028 13972 77196
rect 14028 77186 14084 77196
rect 14588 77250 14644 77308
rect 14588 77198 14590 77250
rect 14642 77198 14644 77250
rect 14588 77186 14644 77198
rect 14700 77138 14756 78204
rect 15260 78260 15316 78270
rect 15484 78260 15540 78654
rect 15260 78258 15540 78260
rect 15260 78206 15262 78258
rect 15314 78206 15540 78258
rect 15260 78204 15540 78206
rect 15260 78194 15316 78204
rect 15148 78036 15204 78046
rect 15372 78036 15428 78046
rect 15148 78034 15316 78036
rect 15148 77982 15150 78034
rect 15202 77982 15316 78034
rect 15148 77980 15316 77982
rect 15148 77970 15204 77980
rect 14700 77086 14702 77138
rect 14754 77086 14756 77138
rect 14700 77074 14756 77086
rect 15260 77140 15316 77980
rect 15428 77980 15540 78036
rect 15372 77942 15428 77980
rect 15484 77250 15540 77980
rect 15484 77198 15486 77250
rect 15538 77198 15540 77250
rect 15484 77186 15540 77198
rect 15596 77922 15652 77934
rect 15596 77870 15598 77922
rect 15650 77870 15652 77922
rect 15372 77140 15428 77150
rect 15260 77084 15372 77140
rect 13804 76972 13972 77028
rect 15148 77028 15204 77066
rect 15372 77046 15428 77084
rect 13804 76692 13860 76972
rect 15148 76962 15204 76972
rect 15372 76916 15428 76926
rect 14008 76860 15208 76870
rect 14064 76858 14112 76860
rect 14168 76858 14216 76860
rect 14076 76806 14112 76858
rect 14200 76806 14216 76858
rect 14064 76804 14112 76806
rect 14168 76804 14216 76806
rect 14272 76858 14320 76860
rect 14376 76858 14424 76860
rect 14480 76858 14528 76860
rect 14376 76806 14396 76858
rect 14480 76806 14520 76858
rect 14272 76804 14320 76806
rect 14376 76804 14424 76806
rect 14480 76804 14528 76806
rect 14584 76804 14632 76860
rect 14688 76858 14736 76860
rect 14792 76858 14840 76860
rect 14896 76858 14944 76860
rect 14696 76806 14736 76858
rect 14820 76806 14840 76858
rect 14688 76804 14736 76806
rect 14792 76804 14840 76806
rect 14896 76804 14944 76806
rect 15000 76858 15048 76860
rect 15104 76858 15152 76860
rect 15000 76806 15016 76858
rect 15104 76806 15140 76858
rect 15000 76804 15048 76806
rect 15104 76804 15152 76806
rect 14008 76794 15208 76804
rect 15372 76692 15428 76860
rect 15596 76804 15652 77870
rect 15596 76738 15652 76748
rect 13804 76690 14532 76692
rect 13804 76638 13806 76690
rect 13858 76638 14532 76690
rect 13804 76636 14532 76638
rect 13804 76626 13860 76636
rect 13580 76402 13636 76412
rect 14476 75794 14532 76636
rect 15260 76636 15428 76692
rect 15708 76692 15764 78764
rect 15820 78596 15876 79324
rect 15820 78034 15876 78540
rect 15820 77982 15822 78034
rect 15874 77982 15876 78034
rect 15820 77970 15876 77982
rect 15932 78930 15988 78942
rect 15932 78878 15934 78930
rect 15986 78878 15988 78930
rect 14588 76580 14644 76590
rect 14588 76486 14644 76524
rect 15260 76578 15316 76636
rect 15708 76626 15764 76636
rect 15260 76526 15262 76578
rect 15314 76526 15316 76578
rect 15260 76514 15316 76526
rect 15820 76580 15876 76590
rect 15820 76486 15876 76524
rect 15372 76468 15428 76478
rect 14476 75742 14478 75794
rect 14530 75742 14532 75794
rect 14476 75572 14532 75742
rect 14476 75506 14532 75516
rect 14700 76354 14756 76366
rect 14700 76302 14702 76354
rect 14754 76302 14756 76354
rect 13804 75460 13860 75470
rect 13468 73892 13748 73948
rect 13580 73780 13636 73790
rect 13580 70980 13636 73724
rect 13580 70914 13636 70924
rect 13580 70420 13636 70430
rect 13580 70326 13636 70364
rect 13356 69410 13412 69422
rect 13356 69358 13358 69410
rect 13410 69358 13412 69410
rect 13356 69076 13412 69358
rect 13580 69188 13636 69198
rect 13580 69094 13636 69132
rect 13356 69010 13412 69020
rect 13580 68852 13636 68862
rect 13244 67554 13300 67564
rect 13468 67732 13524 67742
rect 13468 67508 13524 67676
rect 13356 67452 13524 67508
rect 13244 67172 13300 67182
rect 13020 65090 13076 65100
rect 13132 66834 13188 66846
rect 13132 66782 13134 66834
rect 13186 66782 13188 66834
rect 13132 66500 13188 66782
rect 13132 64708 13188 66444
rect 13244 65714 13300 67116
rect 13244 65662 13246 65714
rect 13298 65662 13300 65714
rect 13244 65650 13300 65662
rect 13356 65380 13412 67452
rect 13468 67284 13524 67294
rect 13468 67170 13524 67228
rect 13468 67118 13470 67170
rect 13522 67118 13524 67170
rect 13468 67106 13524 67118
rect 13580 67060 13636 68796
rect 13580 66994 13636 67004
rect 13692 66836 13748 73892
rect 13804 69748 13860 75404
rect 14700 75460 14756 76302
rect 14924 75796 14980 75806
rect 14924 75702 14980 75740
rect 15372 75796 15428 76412
rect 15932 76466 15988 78878
rect 16044 78818 16100 79324
rect 16044 78766 16046 78818
rect 16098 78766 16100 78818
rect 16044 78754 16100 78766
rect 16268 78706 16324 78718
rect 16268 78654 16270 78706
rect 16322 78654 16324 78706
rect 15932 76414 15934 76466
rect 15986 76414 15988 76466
rect 15932 76402 15988 76414
rect 16044 77140 16100 77150
rect 16044 76356 16100 77084
rect 16268 76804 16324 78654
rect 16380 77924 16436 77934
rect 16380 77830 16436 77868
rect 16380 76804 16436 76814
rect 16268 76748 16380 76804
rect 16380 76738 16436 76748
rect 16380 76468 16436 76478
rect 16436 76412 16548 76468
rect 16380 76374 16436 76412
rect 15372 75794 15540 75796
rect 15372 75742 15374 75794
rect 15426 75742 15540 75794
rect 15372 75740 15540 75742
rect 15372 75730 15428 75740
rect 14700 75394 14756 75404
rect 14008 75292 15208 75302
rect 14064 75290 14112 75292
rect 14168 75290 14216 75292
rect 14076 75238 14112 75290
rect 14200 75238 14216 75290
rect 14064 75236 14112 75238
rect 14168 75236 14216 75238
rect 14272 75290 14320 75292
rect 14376 75290 14424 75292
rect 14480 75290 14528 75292
rect 14376 75238 14396 75290
rect 14480 75238 14520 75290
rect 14272 75236 14320 75238
rect 14376 75236 14424 75238
rect 14480 75236 14528 75238
rect 14584 75236 14632 75292
rect 14688 75290 14736 75292
rect 14792 75290 14840 75292
rect 14896 75290 14944 75292
rect 14696 75238 14736 75290
rect 14820 75238 14840 75290
rect 14688 75236 14736 75238
rect 14792 75236 14840 75238
rect 14896 75236 14944 75238
rect 15000 75290 15048 75292
rect 15104 75290 15152 75292
rect 15000 75238 15016 75290
rect 15104 75238 15140 75290
rect 15000 75236 15048 75238
rect 15104 75236 15152 75238
rect 14008 75226 15208 75236
rect 14252 75124 14308 75134
rect 14252 75030 14308 75068
rect 14364 74898 14420 74910
rect 14364 74846 14366 74898
rect 14418 74846 14420 74898
rect 14364 73892 14420 74846
rect 15260 74786 15316 74798
rect 15260 74734 15262 74786
rect 15314 74734 15316 74786
rect 15260 74674 15316 74734
rect 15260 74622 15262 74674
rect 15314 74622 15316 74674
rect 15260 74610 15316 74622
rect 14364 73826 14420 73836
rect 15372 73892 15428 73902
rect 14008 73724 15208 73734
rect 14064 73722 14112 73724
rect 14168 73722 14216 73724
rect 14076 73670 14112 73722
rect 14200 73670 14216 73722
rect 14064 73668 14112 73670
rect 14168 73668 14216 73670
rect 14272 73722 14320 73724
rect 14376 73722 14424 73724
rect 14480 73722 14528 73724
rect 14376 73670 14396 73722
rect 14480 73670 14520 73722
rect 14272 73668 14320 73670
rect 14376 73668 14424 73670
rect 14480 73668 14528 73670
rect 14584 73668 14632 73724
rect 14688 73722 14736 73724
rect 14792 73722 14840 73724
rect 14896 73722 14944 73724
rect 14696 73670 14736 73722
rect 14820 73670 14840 73722
rect 14688 73668 14736 73670
rect 14792 73668 14840 73670
rect 14896 73668 14944 73670
rect 15000 73722 15048 73724
rect 15104 73722 15152 73724
rect 15000 73670 15016 73722
rect 15104 73670 15140 73722
rect 15000 73668 15048 73670
rect 15104 73668 15152 73670
rect 14008 73658 15208 73668
rect 14364 73556 14420 73566
rect 14364 73462 14420 73500
rect 15148 73556 15204 73566
rect 15372 73556 15428 73836
rect 15148 73554 15428 73556
rect 15148 73502 15150 73554
rect 15202 73502 15428 73554
rect 15148 73500 15428 73502
rect 15484 73892 15540 75740
rect 15708 75684 15764 75694
rect 15708 75590 15764 75628
rect 16044 75682 16100 76300
rect 16044 75630 16046 75682
rect 16098 75630 16100 75682
rect 16044 75618 16100 75630
rect 16156 75684 16212 75694
rect 15932 75458 15988 75470
rect 15932 75406 15934 75458
rect 15986 75406 15988 75458
rect 15708 75124 15764 75134
rect 15708 75030 15764 75068
rect 15932 74228 15988 75406
rect 16156 75122 16212 75628
rect 16492 75682 16548 76412
rect 16492 75630 16494 75682
rect 16546 75630 16548 75682
rect 16492 75618 16548 75630
rect 16268 75572 16324 75582
rect 16268 75570 16436 75572
rect 16268 75518 16270 75570
rect 16322 75518 16436 75570
rect 16268 75516 16436 75518
rect 16268 75506 16324 75516
rect 16156 75070 16158 75122
rect 16210 75070 16212 75122
rect 16156 74674 16212 75070
rect 16380 74788 16436 75516
rect 16492 75124 16548 75134
rect 16548 75068 16660 75124
rect 16492 75058 16548 75068
rect 16604 75010 16660 75068
rect 16604 74958 16606 75010
rect 16658 74958 16660 75010
rect 16604 74946 16660 74958
rect 16492 74788 16548 74798
rect 16380 74786 16548 74788
rect 16380 74734 16494 74786
rect 16546 74734 16548 74786
rect 16380 74732 16548 74734
rect 16492 74722 16548 74732
rect 16156 74622 16158 74674
rect 16210 74622 16212 74674
rect 16156 74610 16212 74622
rect 15932 74172 16436 74228
rect 15820 74114 15876 74126
rect 15820 74062 15822 74114
rect 15874 74062 15876 74114
rect 15820 73948 15876 74062
rect 16380 74114 16436 74172
rect 16380 74062 16382 74114
rect 16434 74062 16436 74114
rect 16380 74050 16436 74062
rect 16716 73948 16772 80892
rect 17276 77252 17332 85708
rect 18172 85698 18228 85708
rect 18172 84868 18228 84878
rect 18172 84774 18228 84812
rect 17500 84196 17556 84206
rect 17500 84102 17556 84140
rect 18284 84194 18340 86044
rect 18620 85764 18676 85774
rect 18620 85670 18676 85708
rect 18732 84530 18788 86606
rect 18956 86546 19012 86558
rect 18956 86494 18958 86546
rect 19010 86494 19012 86546
rect 18956 85764 19012 86494
rect 18956 85698 19012 85708
rect 19404 86546 19460 87388
rect 20412 87332 20468 87612
rect 20412 87266 20468 87276
rect 20524 87556 20580 87566
rect 19404 86494 19406 86546
rect 19458 86494 19460 86546
rect 18732 84478 18734 84530
rect 18786 84478 18788 84530
rect 18732 84466 18788 84478
rect 19292 84868 19348 84878
rect 19292 84418 19348 84812
rect 19292 84366 19294 84418
rect 19346 84366 19348 84418
rect 19292 84354 19348 84366
rect 18284 84142 18286 84194
rect 18338 84142 18340 84194
rect 18284 84084 18340 84142
rect 18284 84018 18340 84028
rect 19068 84084 19124 84094
rect 19068 83990 19124 84028
rect 18732 83748 18788 83758
rect 17612 83524 17668 83534
rect 17836 83524 17892 83534
rect 17388 83522 17668 83524
rect 17388 83470 17614 83522
rect 17666 83470 17668 83522
rect 17388 83468 17668 83470
rect 17388 82850 17444 83468
rect 17612 83458 17668 83468
rect 17724 83522 17892 83524
rect 17724 83470 17838 83522
rect 17890 83470 17892 83522
rect 17724 83468 17892 83470
rect 17388 82798 17390 82850
rect 17442 82798 17444 82850
rect 17388 82786 17444 82798
rect 17500 83298 17556 83310
rect 17500 83246 17502 83298
rect 17554 83246 17556 83298
rect 17500 81954 17556 83246
rect 17612 82740 17668 82750
rect 17612 82646 17668 82684
rect 17500 81902 17502 81954
rect 17554 81902 17556 81954
rect 17500 81890 17556 81902
rect 17724 81508 17780 83468
rect 17836 83458 17892 83468
rect 18284 83524 18340 83534
rect 18284 83430 18340 83468
rect 18396 83412 18452 83422
rect 18396 83318 18452 83356
rect 18732 83410 18788 83692
rect 18732 83358 18734 83410
rect 18786 83358 18788 83410
rect 17836 82738 17892 82750
rect 17836 82686 17838 82738
rect 17890 82686 17892 82738
rect 17836 82516 17892 82686
rect 17836 82450 17892 82460
rect 18732 82516 18788 83358
rect 18732 82450 18788 82460
rect 18844 83692 19236 83748
rect 18844 82626 18900 83692
rect 18844 82574 18846 82626
rect 18898 82574 18900 82626
rect 17724 81442 17780 81452
rect 18060 82292 18116 82302
rect 17388 81172 17444 81182
rect 17388 81078 17444 81116
rect 18060 81060 18116 82236
rect 18844 81732 18900 82574
rect 18060 80966 18116 81004
rect 18284 81284 18340 81294
rect 18284 81170 18340 81228
rect 18284 81118 18286 81170
rect 18338 81118 18340 81170
rect 18284 80612 18340 81118
rect 18844 80948 18900 81676
rect 18844 80882 18900 80892
rect 18956 83524 19012 83534
rect 18956 81956 19012 83468
rect 19180 83522 19236 83692
rect 19180 83470 19182 83522
rect 19234 83470 19236 83522
rect 19180 83458 19236 83470
rect 19404 83522 19460 86494
rect 20076 85876 20132 85886
rect 20076 85782 20132 85820
rect 20300 84868 20356 84878
rect 19628 84418 19684 84430
rect 19628 84366 19630 84418
rect 19682 84366 19684 84418
rect 19628 83748 19684 84366
rect 19628 83682 19684 83692
rect 20300 84308 20356 84812
rect 20300 83634 20356 84252
rect 20524 84308 20580 87500
rect 20972 87444 21028 87454
rect 20972 87350 21028 87388
rect 21308 87442 21364 87454
rect 21308 87390 21310 87442
rect 21362 87390 21364 87442
rect 21308 87332 21364 87390
rect 21308 86100 21364 87276
rect 24008 87052 25208 87062
rect 24064 87050 24112 87052
rect 24168 87050 24216 87052
rect 24076 86998 24112 87050
rect 24200 86998 24216 87050
rect 24064 86996 24112 86998
rect 24168 86996 24216 86998
rect 24272 87050 24320 87052
rect 24376 87050 24424 87052
rect 24480 87050 24528 87052
rect 24376 86998 24396 87050
rect 24480 86998 24520 87050
rect 24272 86996 24320 86998
rect 24376 86996 24424 86998
rect 24480 86996 24528 86998
rect 24584 86996 24632 87052
rect 24688 87050 24736 87052
rect 24792 87050 24840 87052
rect 24896 87050 24944 87052
rect 24696 86998 24736 87050
rect 24820 86998 24840 87050
rect 24688 86996 24736 86998
rect 24792 86996 24840 86998
rect 24896 86996 24944 86998
rect 25000 87050 25048 87052
rect 25104 87050 25152 87052
rect 25000 86998 25016 87050
rect 25104 86998 25140 87050
rect 25000 86996 25048 86998
rect 25104 86996 25152 86998
rect 24008 86986 25208 86996
rect 21308 86034 21364 86044
rect 23100 86098 23156 86110
rect 23100 86046 23102 86098
rect 23154 86046 23156 86098
rect 23100 85988 23156 86046
rect 23100 85922 23156 85932
rect 23996 85988 24052 85998
rect 20636 85876 20692 85886
rect 23884 85876 23940 85886
rect 20636 85874 21476 85876
rect 20636 85822 20638 85874
rect 20690 85822 21476 85874
rect 20636 85820 21476 85822
rect 20636 85810 20692 85820
rect 20748 85540 20804 85550
rect 20748 84980 20804 85484
rect 21420 85314 21476 85820
rect 21420 85262 21422 85314
rect 21474 85262 21476 85314
rect 21420 85250 21476 85262
rect 22540 85764 22596 85774
rect 21756 85092 21812 85102
rect 21756 85090 21924 85092
rect 21756 85038 21758 85090
rect 21810 85038 21924 85090
rect 21756 85036 21924 85038
rect 21756 85026 21812 85036
rect 20748 84886 20804 84924
rect 21868 84532 21924 85036
rect 21980 84980 22036 84990
rect 21980 84886 22036 84924
rect 22540 84978 22596 85708
rect 23660 85764 23716 85774
rect 23660 85670 23716 85708
rect 22540 84926 22542 84978
rect 22594 84926 22596 84978
rect 22092 84532 22148 84542
rect 21868 84530 22148 84532
rect 21868 84478 22094 84530
rect 22146 84478 22148 84530
rect 21868 84476 22148 84478
rect 22092 84466 22148 84476
rect 21084 84418 21140 84430
rect 21084 84366 21086 84418
rect 21138 84366 21140 84418
rect 20972 84308 21028 84318
rect 20524 84306 20692 84308
rect 20524 84254 20526 84306
rect 20578 84254 20692 84306
rect 20524 84252 20692 84254
rect 20524 84242 20580 84252
rect 20636 84196 20692 84252
rect 20972 84214 21028 84252
rect 20636 84130 20692 84140
rect 20300 83582 20302 83634
rect 20354 83582 20356 83634
rect 20300 83570 20356 83582
rect 19404 83470 19406 83522
rect 19458 83470 19460 83522
rect 19404 83458 19460 83470
rect 19068 83412 19124 83422
rect 19068 83318 19124 83356
rect 20636 82516 20692 82526
rect 18956 80946 19012 81900
rect 20076 82180 20132 82190
rect 20636 82180 20692 82460
rect 21084 82516 21140 84366
rect 21084 82422 21140 82460
rect 21756 84196 21812 84206
rect 21756 84082 21812 84140
rect 21756 84030 21758 84082
rect 21810 84030 21812 84082
rect 20076 81732 20132 82124
rect 19964 81730 20132 81732
rect 19964 81678 20078 81730
rect 20130 81678 20132 81730
rect 19964 81676 20132 81678
rect 19292 81170 19348 81182
rect 19292 81118 19294 81170
rect 19346 81118 19348 81170
rect 18956 80894 18958 80946
rect 19010 80894 19012 80946
rect 18956 80882 19012 80894
rect 19180 81060 19236 81070
rect 18284 80546 18340 80556
rect 17500 80500 17556 80510
rect 17500 79826 17556 80444
rect 19180 80500 19236 81004
rect 19292 80948 19348 81118
rect 19292 80882 19348 80892
rect 19404 80612 19460 80622
rect 19404 80518 19460 80556
rect 19180 80434 19236 80444
rect 19964 80498 20020 81676
rect 20076 81666 20132 81676
rect 20300 82178 20692 82180
rect 20300 82126 20638 82178
rect 20690 82126 20692 82178
rect 20300 82124 20692 82126
rect 20076 81060 20132 81070
rect 20076 80966 20132 81004
rect 19964 80446 19966 80498
rect 20018 80446 20020 80498
rect 18844 80276 18900 80286
rect 18844 80162 18900 80220
rect 19964 80276 20020 80446
rect 20020 80220 20244 80276
rect 19964 80210 20020 80220
rect 18844 80110 18846 80162
rect 18898 80110 18900 80162
rect 18844 80098 18900 80110
rect 17500 79774 17502 79826
rect 17554 79774 17556 79826
rect 17500 79762 17556 79774
rect 17276 77186 17332 77196
rect 19964 78930 20020 78942
rect 19964 78878 19966 78930
rect 20018 78878 20020 78930
rect 19964 77252 20020 78878
rect 20188 78484 20244 80220
rect 20300 78818 20356 82124
rect 20636 82114 20692 82124
rect 21420 82180 21476 82190
rect 21420 82066 21476 82124
rect 21420 82014 21422 82066
rect 21474 82014 21476 82066
rect 21420 82002 21476 82014
rect 20524 81058 20580 81070
rect 20524 81006 20526 81058
rect 20578 81006 20580 81058
rect 20524 80948 20580 81006
rect 21756 80948 21812 84030
rect 22316 83636 22372 83646
rect 22372 83580 22484 83636
rect 22316 83570 22372 83580
rect 22428 83300 22484 83580
rect 22540 83524 22596 84926
rect 22988 83524 23044 83534
rect 22540 83522 23044 83524
rect 22540 83470 22990 83522
rect 23042 83470 23044 83522
rect 22540 83468 23044 83470
rect 22988 83458 23044 83468
rect 22540 83300 22596 83310
rect 22428 83244 22540 83300
rect 22540 83206 22596 83244
rect 22652 83300 22708 83310
rect 22876 83300 22932 83310
rect 22652 83298 22820 83300
rect 22652 83246 22654 83298
rect 22706 83246 22820 83298
rect 22652 83244 22820 83246
rect 22652 83234 22708 83244
rect 21868 82850 21924 82862
rect 21868 82798 21870 82850
rect 21922 82798 21924 82850
rect 21868 82180 21924 82798
rect 21868 82114 21924 82124
rect 22092 82516 22148 82526
rect 20580 80892 20916 80948
rect 20524 80854 20580 80892
rect 20636 79490 20692 79502
rect 20636 79438 20638 79490
rect 20690 79438 20692 79490
rect 20636 79378 20692 79438
rect 20636 79326 20638 79378
rect 20690 79326 20692 79378
rect 20636 79314 20692 79326
rect 20300 78766 20302 78818
rect 20354 78766 20356 78818
rect 20300 78754 20356 78766
rect 20748 78708 20804 78718
rect 20748 78614 20804 78652
rect 20188 78418 20244 78428
rect 20300 78260 20356 78270
rect 20300 78166 20356 78204
rect 19964 77186 20020 77196
rect 16828 76916 16884 76926
rect 16828 76690 16884 76860
rect 16828 76638 16830 76690
rect 16882 76638 16884 76690
rect 16828 75684 16884 76638
rect 17388 76916 17444 76926
rect 17388 76580 17444 76860
rect 17724 76692 17780 76702
rect 17388 76578 17668 76580
rect 17388 76526 17390 76578
rect 17442 76526 17668 76578
rect 17388 76524 17668 76526
rect 17388 76514 17444 76524
rect 17500 76354 17556 76366
rect 17500 76302 17502 76354
rect 17554 76302 17556 76354
rect 16828 75010 16884 75628
rect 17164 75684 17220 75694
rect 17500 75684 17556 76302
rect 17164 75682 17556 75684
rect 17164 75630 17166 75682
rect 17218 75630 17556 75682
rect 17164 75628 17556 75630
rect 17164 75618 17220 75628
rect 16828 74958 16830 75010
rect 16882 74958 16884 75010
rect 16828 74946 16884 74958
rect 17612 75012 17668 76524
rect 17724 76578 17780 76636
rect 18732 76692 18788 76702
rect 18732 76598 18788 76636
rect 20300 76692 20356 76702
rect 20300 76598 20356 76636
rect 17724 76526 17726 76578
rect 17778 76526 17780 76578
rect 17724 76514 17780 76526
rect 17836 76466 17892 76478
rect 17836 76414 17838 76466
rect 17890 76414 17892 76466
rect 17836 75122 17892 76414
rect 18396 76466 18452 76478
rect 18396 76414 18398 76466
rect 18450 76414 18452 76466
rect 18284 76356 18340 76366
rect 18284 76262 18340 76300
rect 17836 75070 17838 75122
rect 17890 75070 17892 75122
rect 17836 75058 17892 75070
rect 17724 75012 17780 75022
rect 17612 75010 17780 75012
rect 17612 74958 17726 75010
rect 17778 74958 17780 75010
rect 17612 74956 17780 74958
rect 17724 74946 17780 74956
rect 17948 75010 18004 75022
rect 17948 74958 17950 75010
rect 18002 74958 18004 75010
rect 15596 73892 15876 73948
rect 16604 73892 16772 73948
rect 17948 74788 18004 74958
rect 17948 74004 18004 74732
rect 18396 74340 18452 76414
rect 18844 76468 18900 76478
rect 18844 76374 18900 76412
rect 20188 76468 20244 76478
rect 20188 75906 20244 76412
rect 20748 76356 20804 76366
rect 20748 76262 20804 76300
rect 20188 75854 20190 75906
rect 20242 75854 20244 75906
rect 20188 75842 20244 75854
rect 19404 75460 19460 75470
rect 18508 74788 18564 74798
rect 18508 74694 18564 74732
rect 18396 74274 18452 74284
rect 17948 73938 18004 73948
rect 15484 73890 15652 73892
rect 15484 73838 15598 73890
rect 15650 73838 15652 73890
rect 15484 73836 15652 73838
rect 15148 73490 15204 73500
rect 15484 73220 15540 73836
rect 15596 73826 15652 73836
rect 15372 73218 15540 73220
rect 15372 73166 15486 73218
rect 15538 73166 15540 73218
rect 15372 73164 15540 73166
rect 14008 72156 15208 72166
rect 14064 72154 14112 72156
rect 14168 72154 14216 72156
rect 14076 72102 14112 72154
rect 14200 72102 14216 72154
rect 14064 72100 14112 72102
rect 14168 72100 14216 72102
rect 14272 72154 14320 72156
rect 14376 72154 14424 72156
rect 14480 72154 14528 72156
rect 14376 72102 14396 72154
rect 14480 72102 14520 72154
rect 14272 72100 14320 72102
rect 14376 72100 14424 72102
rect 14480 72100 14528 72102
rect 14584 72100 14632 72156
rect 14688 72154 14736 72156
rect 14792 72154 14840 72156
rect 14896 72154 14944 72156
rect 14696 72102 14736 72154
rect 14820 72102 14840 72154
rect 14688 72100 14736 72102
rect 14792 72100 14840 72102
rect 14896 72100 14944 72102
rect 15000 72154 15048 72156
rect 15104 72154 15152 72156
rect 15000 72102 15016 72154
rect 15104 72102 15140 72154
rect 15000 72100 15048 72102
rect 15104 72100 15152 72102
rect 14008 72090 15208 72100
rect 15372 71988 15428 73164
rect 15484 73154 15540 73164
rect 15932 73556 15988 73566
rect 14812 71932 15428 71988
rect 14812 71090 14868 71932
rect 14812 71038 14814 71090
rect 14866 71038 14868 71090
rect 14812 71026 14868 71038
rect 15260 71092 15316 71102
rect 15260 70868 15316 71036
rect 15932 71092 15988 73500
rect 16044 71092 16100 71102
rect 15988 71090 16100 71092
rect 15988 71038 16046 71090
rect 16098 71038 16100 71090
rect 15988 71036 16100 71038
rect 15932 70998 15988 71036
rect 16044 71026 16100 71036
rect 15260 70802 15316 70812
rect 14008 70588 15208 70598
rect 14064 70586 14112 70588
rect 14168 70586 14216 70588
rect 14076 70534 14112 70586
rect 14200 70534 14216 70586
rect 14064 70532 14112 70534
rect 14168 70532 14216 70534
rect 14272 70586 14320 70588
rect 14376 70586 14424 70588
rect 14480 70586 14528 70588
rect 14376 70534 14396 70586
rect 14480 70534 14520 70586
rect 14272 70532 14320 70534
rect 14376 70532 14424 70534
rect 14480 70532 14528 70534
rect 14584 70532 14632 70588
rect 14688 70586 14736 70588
rect 14792 70586 14840 70588
rect 14896 70586 14944 70588
rect 14696 70534 14736 70586
rect 14820 70534 14840 70586
rect 14688 70532 14736 70534
rect 14792 70532 14840 70534
rect 14896 70532 14944 70534
rect 15000 70586 15048 70588
rect 15104 70586 15152 70588
rect 15000 70534 15016 70586
rect 15104 70534 15140 70586
rect 15000 70532 15048 70534
rect 15104 70532 15152 70534
rect 14008 70522 15208 70532
rect 15036 70420 15092 70430
rect 15036 70196 15092 70364
rect 15148 70420 15204 70430
rect 16604 70420 16660 73892
rect 18732 73890 18788 73902
rect 18732 73838 18734 73890
rect 18786 73838 18788 73890
rect 18284 73556 18340 73566
rect 18284 71986 18340 73500
rect 18732 73556 18788 73838
rect 18732 73490 18788 73500
rect 19404 73892 19460 75404
rect 20524 75460 20580 75470
rect 20524 75366 20580 75404
rect 19516 74340 19572 74350
rect 19516 74246 19572 74284
rect 20860 73948 20916 80892
rect 21308 80892 21812 80948
rect 21980 81732 22036 81742
rect 21980 80948 22036 81676
rect 20972 79490 21028 79502
rect 20972 79438 20974 79490
rect 21026 79438 21028 79490
rect 20972 78708 21028 79438
rect 21308 78708 21364 80892
rect 21980 80882 22036 80892
rect 22092 80836 22148 82460
rect 22428 82516 22484 82526
rect 22428 82066 22484 82460
rect 22428 82014 22430 82066
rect 22482 82014 22484 82066
rect 22428 82002 22484 82014
rect 22764 81842 22820 83244
rect 22876 83206 22932 83244
rect 22764 81790 22766 81842
rect 22818 81790 22820 81842
rect 22764 81778 22820 81790
rect 23884 82740 23940 85820
rect 23996 85764 24052 85932
rect 24556 85876 24612 85886
rect 24556 85782 24612 85820
rect 23996 85670 24052 85708
rect 25340 85764 25396 85774
rect 24008 85484 25208 85494
rect 24064 85482 24112 85484
rect 24168 85482 24216 85484
rect 24076 85430 24112 85482
rect 24200 85430 24216 85482
rect 24064 85428 24112 85430
rect 24168 85428 24216 85430
rect 24272 85482 24320 85484
rect 24376 85482 24424 85484
rect 24480 85482 24528 85484
rect 24376 85430 24396 85482
rect 24480 85430 24520 85482
rect 24272 85428 24320 85430
rect 24376 85428 24424 85430
rect 24480 85428 24528 85430
rect 24584 85428 24632 85484
rect 24688 85482 24736 85484
rect 24792 85482 24840 85484
rect 24896 85482 24944 85484
rect 24696 85430 24736 85482
rect 24820 85430 24840 85482
rect 24688 85428 24736 85430
rect 24792 85428 24840 85430
rect 24896 85428 24944 85430
rect 25000 85482 25048 85484
rect 25104 85482 25152 85484
rect 25000 85430 25016 85482
rect 25104 85430 25140 85482
rect 25000 85428 25048 85430
rect 25104 85428 25152 85430
rect 24008 85418 25208 85428
rect 24008 83916 25208 83926
rect 24064 83914 24112 83916
rect 24168 83914 24216 83916
rect 24076 83862 24112 83914
rect 24200 83862 24216 83914
rect 24064 83860 24112 83862
rect 24168 83860 24216 83862
rect 24272 83914 24320 83916
rect 24376 83914 24424 83916
rect 24480 83914 24528 83916
rect 24376 83862 24396 83914
rect 24480 83862 24520 83914
rect 24272 83860 24320 83862
rect 24376 83860 24424 83862
rect 24480 83860 24528 83862
rect 24584 83860 24632 83916
rect 24688 83914 24736 83916
rect 24792 83914 24840 83916
rect 24896 83914 24944 83916
rect 24696 83862 24736 83914
rect 24820 83862 24840 83914
rect 24688 83860 24736 83862
rect 24792 83860 24840 83862
rect 24896 83860 24944 83862
rect 25000 83914 25048 83916
rect 25104 83914 25152 83916
rect 25000 83862 25016 83914
rect 25104 83862 25140 83914
rect 25000 83860 25048 83862
rect 25104 83860 25152 83862
rect 24008 83850 25208 83860
rect 25340 82962 25396 85708
rect 25340 82910 25342 82962
rect 25394 82910 25396 82962
rect 22316 81732 22372 81742
rect 22204 81730 22372 81732
rect 22204 81678 22318 81730
rect 22370 81678 22372 81730
rect 22204 81676 22372 81678
rect 22204 81058 22260 81676
rect 22316 81666 22372 81676
rect 22540 81732 22596 81742
rect 22540 81638 22596 81676
rect 22540 81170 22596 81182
rect 22540 81118 22542 81170
rect 22594 81118 22596 81170
rect 22204 81006 22206 81058
rect 22258 81006 22260 81058
rect 22204 80994 22260 81006
rect 22316 81060 22372 81070
rect 22316 80966 22372 81004
rect 22540 80836 22596 81118
rect 23660 81060 23716 81070
rect 23660 80966 23716 81004
rect 22092 80780 22596 80836
rect 22092 79602 22148 80780
rect 22092 79550 22094 79602
rect 22146 79550 22148 79602
rect 22092 79538 22148 79550
rect 22204 79490 22260 79502
rect 22204 79438 22206 79490
rect 22258 79438 22260 79490
rect 21420 79380 21476 79390
rect 21420 79378 21588 79380
rect 21420 79326 21422 79378
rect 21474 79326 21588 79378
rect 21420 79324 21588 79326
rect 21420 79314 21476 79324
rect 21532 78820 21588 79324
rect 21532 78764 21924 78820
rect 21420 78708 21476 78718
rect 20972 78706 21476 78708
rect 20972 78654 21422 78706
rect 21474 78654 21476 78706
rect 20972 78652 21476 78654
rect 20972 78484 21028 78494
rect 20972 78258 21028 78428
rect 20972 78206 20974 78258
rect 21026 78206 21028 78258
rect 20972 78194 21028 78206
rect 21196 77252 21252 77262
rect 21196 77158 21252 77196
rect 21308 76578 21364 76590
rect 21308 76526 21310 76578
rect 21362 76526 21364 76578
rect 21308 76356 21364 76526
rect 21308 76290 21364 76300
rect 21420 73948 21476 78652
rect 21868 78706 21924 78764
rect 21868 78654 21870 78706
rect 21922 78654 21924 78706
rect 21868 78596 21924 78654
rect 21756 78540 21924 78596
rect 22204 78818 22260 79438
rect 22652 79492 22708 79502
rect 22652 79490 23268 79492
rect 22652 79438 22654 79490
rect 22706 79438 23268 79490
rect 22652 79436 23268 79438
rect 22652 79426 22708 79436
rect 22204 78766 22206 78818
rect 22258 78766 22260 78818
rect 21756 76692 21812 78540
rect 21980 78484 22036 78494
rect 21756 76578 21812 76636
rect 21756 76526 21758 76578
rect 21810 76526 21812 76578
rect 21756 76514 21812 76526
rect 21868 77252 21924 77262
rect 21868 76468 21924 77196
rect 21980 77138 22036 78428
rect 22204 78260 22260 78766
rect 22988 78708 23044 78718
rect 22988 78614 23044 78652
rect 23212 78706 23268 79436
rect 23324 78932 23380 78942
rect 23324 78930 23492 78932
rect 23324 78878 23326 78930
rect 23378 78878 23492 78930
rect 23324 78876 23492 78878
rect 23324 78866 23380 78876
rect 23212 78654 23214 78706
rect 23266 78654 23268 78706
rect 23212 78642 23268 78654
rect 22540 78596 22596 78606
rect 22540 78594 22932 78596
rect 22540 78542 22542 78594
rect 22594 78542 22932 78594
rect 22540 78540 22932 78542
rect 22540 78530 22596 78540
rect 22876 78260 22932 78540
rect 22876 78204 23380 78260
rect 22204 78194 22260 78204
rect 23324 78034 23380 78204
rect 23324 77982 23326 78034
rect 23378 77982 23380 78034
rect 23324 77970 23380 77982
rect 21980 77086 21982 77138
rect 22034 77086 22036 77138
rect 21980 77074 22036 77086
rect 22316 77252 22372 77262
rect 22316 76690 22372 77196
rect 22316 76638 22318 76690
rect 22370 76638 22372 76690
rect 22316 76626 22372 76638
rect 23436 76580 23492 78876
rect 23884 78260 23940 82684
rect 24108 82738 24164 82750
rect 24108 82686 24110 82738
rect 24162 82686 24164 82738
rect 24108 82516 24164 82686
rect 24556 82740 24612 82750
rect 24556 82646 24612 82684
rect 24108 82450 24164 82460
rect 24008 82348 25208 82358
rect 24064 82346 24112 82348
rect 24168 82346 24216 82348
rect 24076 82294 24112 82346
rect 24200 82294 24216 82346
rect 24064 82292 24112 82294
rect 24168 82292 24216 82294
rect 24272 82346 24320 82348
rect 24376 82346 24424 82348
rect 24480 82346 24528 82348
rect 24376 82294 24396 82346
rect 24480 82294 24520 82346
rect 24272 82292 24320 82294
rect 24376 82292 24424 82294
rect 24480 82292 24528 82294
rect 24584 82292 24632 82348
rect 24688 82346 24736 82348
rect 24792 82346 24840 82348
rect 24896 82346 24944 82348
rect 24696 82294 24736 82346
rect 24820 82294 24840 82346
rect 24688 82292 24736 82294
rect 24792 82292 24840 82294
rect 24896 82292 24944 82294
rect 25000 82346 25048 82348
rect 25104 82346 25152 82348
rect 25000 82294 25016 82346
rect 25104 82294 25140 82346
rect 25000 82292 25048 82294
rect 25104 82292 25152 82294
rect 24008 82282 25208 82292
rect 25340 82180 25396 82910
rect 25788 82740 25844 82750
rect 25788 82646 25844 82684
rect 25340 82114 25396 82124
rect 24008 80780 25208 80790
rect 24064 80778 24112 80780
rect 24168 80778 24216 80780
rect 24076 80726 24112 80778
rect 24200 80726 24216 80778
rect 24064 80724 24112 80726
rect 24168 80724 24216 80726
rect 24272 80778 24320 80780
rect 24376 80778 24424 80780
rect 24480 80778 24528 80780
rect 24376 80726 24396 80778
rect 24480 80726 24520 80778
rect 24272 80724 24320 80726
rect 24376 80724 24424 80726
rect 24480 80724 24528 80726
rect 24584 80724 24632 80780
rect 24688 80778 24736 80780
rect 24792 80778 24840 80780
rect 24896 80778 24944 80780
rect 24696 80726 24736 80778
rect 24820 80726 24840 80778
rect 24688 80724 24736 80726
rect 24792 80724 24840 80726
rect 24896 80724 24944 80726
rect 25000 80778 25048 80780
rect 25104 80778 25152 80780
rect 25000 80726 25016 80778
rect 25104 80726 25140 80778
rect 25000 80724 25048 80726
rect 25104 80724 25152 80726
rect 24008 80714 25208 80724
rect 24008 79212 25208 79222
rect 24064 79210 24112 79212
rect 24168 79210 24216 79212
rect 24076 79158 24112 79210
rect 24200 79158 24216 79210
rect 24064 79156 24112 79158
rect 24168 79156 24216 79158
rect 24272 79210 24320 79212
rect 24376 79210 24424 79212
rect 24480 79210 24528 79212
rect 24376 79158 24396 79210
rect 24480 79158 24520 79210
rect 24272 79156 24320 79158
rect 24376 79156 24424 79158
rect 24480 79156 24528 79158
rect 24584 79156 24632 79212
rect 24688 79210 24736 79212
rect 24792 79210 24840 79212
rect 24896 79210 24944 79212
rect 24696 79158 24736 79210
rect 24820 79158 24840 79210
rect 24688 79156 24736 79158
rect 24792 79156 24840 79158
rect 24896 79156 24944 79158
rect 25000 79210 25048 79212
rect 25104 79210 25152 79212
rect 25000 79158 25016 79210
rect 25104 79158 25140 79210
rect 25000 79156 25048 79158
rect 25104 79156 25152 79158
rect 24008 79146 25208 79156
rect 29820 78988 29876 95676
rect 34064 95674 34112 95676
rect 34168 95674 34216 95676
rect 34076 95622 34112 95674
rect 34200 95622 34216 95674
rect 34064 95620 34112 95622
rect 34168 95620 34216 95622
rect 34272 95674 34320 95676
rect 34376 95674 34424 95676
rect 34480 95674 34528 95676
rect 34376 95622 34396 95674
rect 34480 95622 34520 95674
rect 34272 95620 34320 95622
rect 34376 95620 34424 95622
rect 34480 95620 34528 95622
rect 34584 95620 34632 95676
rect 34688 95674 34736 95676
rect 34792 95674 34840 95676
rect 34896 95674 34944 95676
rect 34696 95622 34736 95674
rect 34820 95622 34840 95674
rect 34688 95620 34736 95622
rect 34792 95620 34840 95622
rect 34896 95620 34944 95622
rect 35000 95674 35048 95676
rect 35104 95674 35152 95676
rect 35000 95622 35016 95674
rect 35104 95622 35140 95674
rect 35000 95620 35048 95622
rect 35104 95620 35152 95622
rect 34008 95610 35208 95620
rect 34008 94108 35208 94118
rect 34064 94106 34112 94108
rect 34168 94106 34216 94108
rect 34076 94054 34112 94106
rect 34200 94054 34216 94106
rect 34064 94052 34112 94054
rect 34168 94052 34216 94054
rect 34272 94106 34320 94108
rect 34376 94106 34424 94108
rect 34480 94106 34528 94108
rect 34376 94054 34396 94106
rect 34480 94054 34520 94106
rect 34272 94052 34320 94054
rect 34376 94052 34424 94054
rect 34480 94052 34528 94054
rect 34584 94052 34632 94108
rect 34688 94106 34736 94108
rect 34792 94106 34840 94108
rect 34896 94106 34944 94108
rect 34696 94054 34736 94106
rect 34820 94054 34840 94106
rect 34688 94052 34736 94054
rect 34792 94052 34840 94054
rect 34896 94052 34944 94054
rect 35000 94106 35048 94108
rect 35104 94106 35152 94108
rect 35000 94054 35016 94106
rect 35104 94054 35140 94106
rect 35000 94052 35048 94054
rect 35104 94052 35152 94054
rect 34008 94042 35208 94052
rect 34008 92540 35208 92550
rect 34064 92538 34112 92540
rect 34168 92538 34216 92540
rect 34076 92486 34112 92538
rect 34200 92486 34216 92538
rect 34064 92484 34112 92486
rect 34168 92484 34216 92486
rect 34272 92538 34320 92540
rect 34376 92538 34424 92540
rect 34480 92538 34528 92540
rect 34376 92486 34396 92538
rect 34480 92486 34520 92538
rect 34272 92484 34320 92486
rect 34376 92484 34424 92486
rect 34480 92484 34528 92486
rect 34584 92484 34632 92540
rect 34688 92538 34736 92540
rect 34792 92538 34840 92540
rect 34896 92538 34944 92540
rect 34696 92486 34736 92538
rect 34820 92486 34840 92538
rect 34688 92484 34736 92486
rect 34792 92484 34840 92486
rect 34896 92484 34944 92486
rect 35000 92538 35048 92540
rect 35104 92538 35152 92540
rect 35000 92486 35016 92538
rect 35104 92486 35140 92538
rect 35000 92484 35048 92486
rect 35104 92484 35152 92486
rect 34008 92474 35208 92484
rect 34008 90972 35208 90982
rect 34064 90970 34112 90972
rect 34168 90970 34216 90972
rect 34076 90918 34112 90970
rect 34200 90918 34216 90970
rect 34064 90916 34112 90918
rect 34168 90916 34216 90918
rect 34272 90970 34320 90972
rect 34376 90970 34424 90972
rect 34480 90970 34528 90972
rect 34376 90918 34396 90970
rect 34480 90918 34520 90970
rect 34272 90916 34320 90918
rect 34376 90916 34424 90918
rect 34480 90916 34528 90918
rect 34584 90916 34632 90972
rect 34688 90970 34736 90972
rect 34792 90970 34840 90972
rect 34896 90970 34944 90972
rect 34696 90918 34736 90970
rect 34820 90918 34840 90970
rect 34688 90916 34736 90918
rect 34792 90916 34840 90918
rect 34896 90916 34944 90918
rect 35000 90970 35048 90972
rect 35104 90970 35152 90972
rect 35000 90918 35016 90970
rect 35104 90918 35140 90970
rect 35000 90916 35048 90918
rect 35104 90916 35152 90918
rect 34008 90906 35208 90916
rect 34008 89404 35208 89414
rect 34064 89402 34112 89404
rect 34168 89402 34216 89404
rect 34076 89350 34112 89402
rect 34200 89350 34216 89402
rect 34064 89348 34112 89350
rect 34168 89348 34216 89350
rect 34272 89402 34320 89404
rect 34376 89402 34424 89404
rect 34480 89402 34528 89404
rect 34376 89350 34396 89402
rect 34480 89350 34520 89402
rect 34272 89348 34320 89350
rect 34376 89348 34424 89350
rect 34480 89348 34528 89350
rect 34584 89348 34632 89404
rect 34688 89402 34736 89404
rect 34792 89402 34840 89404
rect 34896 89402 34944 89404
rect 34696 89350 34736 89402
rect 34820 89350 34840 89402
rect 34688 89348 34736 89350
rect 34792 89348 34840 89350
rect 34896 89348 34944 89350
rect 35000 89402 35048 89404
rect 35104 89402 35152 89404
rect 35000 89350 35016 89402
rect 35104 89350 35140 89402
rect 35000 89348 35048 89350
rect 35104 89348 35152 89350
rect 34008 89338 35208 89348
rect 34008 87836 35208 87846
rect 34064 87834 34112 87836
rect 34168 87834 34216 87836
rect 34076 87782 34112 87834
rect 34200 87782 34216 87834
rect 34064 87780 34112 87782
rect 34168 87780 34216 87782
rect 34272 87834 34320 87836
rect 34376 87834 34424 87836
rect 34480 87834 34528 87836
rect 34376 87782 34396 87834
rect 34480 87782 34520 87834
rect 34272 87780 34320 87782
rect 34376 87780 34424 87782
rect 34480 87780 34528 87782
rect 34584 87780 34632 87836
rect 34688 87834 34736 87836
rect 34792 87834 34840 87836
rect 34896 87834 34944 87836
rect 34696 87782 34736 87834
rect 34820 87782 34840 87834
rect 34688 87780 34736 87782
rect 34792 87780 34840 87782
rect 34896 87780 34944 87782
rect 35000 87834 35048 87836
rect 35104 87834 35152 87836
rect 35000 87782 35016 87834
rect 35104 87782 35140 87834
rect 35000 87780 35048 87782
rect 35104 87780 35152 87782
rect 34008 87770 35208 87780
rect 34008 86268 35208 86278
rect 34064 86266 34112 86268
rect 34168 86266 34216 86268
rect 34076 86214 34112 86266
rect 34200 86214 34216 86266
rect 34064 86212 34112 86214
rect 34168 86212 34216 86214
rect 34272 86266 34320 86268
rect 34376 86266 34424 86268
rect 34480 86266 34528 86268
rect 34376 86214 34396 86266
rect 34480 86214 34520 86266
rect 34272 86212 34320 86214
rect 34376 86212 34424 86214
rect 34480 86212 34528 86214
rect 34584 86212 34632 86268
rect 34688 86266 34736 86268
rect 34792 86266 34840 86268
rect 34896 86266 34944 86268
rect 34696 86214 34736 86266
rect 34820 86214 34840 86266
rect 34688 86212 34736 86214
rect 34792 86212 34840 86214
rect 34896 86212 34944 86214
rect 35000 86266 35048 86268
rect 35104 86266 35152 86268
rect 35000 86214 35016 86266
rect 35104 86214 35140 86266
rect 35000 86212 35048 86214
rect 35104 86212 35152 86214
rect 34008 86202 35208 86212
rect 34008 84700 35208 84710
rect 34064 84698 34112 84700
rect 34168 84698 34216 84700
rect 34076 84646 34112 84698
rect 34200 84646 34216 84698
rect 34064 84644 34112 84646
rect 34168 84644 34216 84646
rect 34272 84698 34320 84700
rect 34376 84698 34424 84700
rect 34480 84698 34528 84700
rect 34376 84646 34396 84698
rect 34480 84646 34520 84698
rect 34272 84644 34320 84646
rect 34376 84644 34424 84646
rect 34480 84644 34528 84646
rect 34584 84644 34632 84700
rect 34688 84698 34736 84700
rect 34792 84698 34840 84700
rect 34896 84698 34944 84700
rect 34696 84646 34736 84698
rect 34820 84646 34840 84698
rect 34688 84644 34736 84646
rect 34792 84644 34840 84646
rect 34896 84644 34944 84646
rect 35000 84698 35048 84700
rect 35104 84698 35152 84700
rect 35000 84646 35016 84698
rect 35104 84646 35140 84698
rect 35000 84644 35048 84646
rect 35104 84644 35152 84646
rect 34008 84634 35208 84644
rect 34008 83132 35208 83142
rect 34064 83130 34112 83132
rect 34168 83130 34216 83132
rect 34076 83078 34112 83130
rect 34200 83078 34216 83130
rect 34064 83076 34112 83078
rect 34168 83076 34216 83078
rect 34272 83130 34320 83132
rect 34376 83130 34424 83132
rect 34480 83130 34528 83132
rect 34376 83078 34396 83130
rect 34480 83078 34520 83130
rect 34272 83076 34320 83078
rect 34376 83076 34424 83078
rect 34480 83076 34528 83078
rect 34584 83076 34632 83132
rect 34688 83130 34736 83132
rect 34792 83130 34840 83132
rect 34896 83130 34944 83132
rect 34696 83078 34736 83130
rect 34820 83078 34840 83130
rect 34688 83076 34736 83078
rect 34792 83076 34840 83078
rect 34896 83076 34944 83078
rect 35000 83130 35048 83132
rect 35104 83130 35152 83132
rect 35000 83078 35016 83130
rect 35104 83078 35140 83130
rect 35000 83076 35048 83078
rect 35104 83076 35152 83078
rect 34008 83066 35208 83076
rect 34008 81564 35208 81574
rect 34064 81562 34112 81564
rect 34168 81562 34216 81564
rect 34076 81510 34112 81562
rect 34200 81510 34216 81562
rect 34064 81508 34112 81510
rect 34168 81508 34216 81510
rect 34272 81562 34320 81564
rect 34376 81562 34424 81564
rect 34480 81562 34528 81564
rect 34376 81510 34396 81562
rect 34480 81510 34520 81562
rect 34272 81508 34320 81510
rect 34376 81508 34424 81510
rect 34480 81508 34528 81510
rect 34584 81508 34632 81564
rect 34688 81562 34736 81564
rect 34792 81562 34840 81564
rect 34896 81562 34944 81564
rect 34696 81510 34736 81562
rect 34820 81510 34840 81562
rect 34688 81508 34736 81510
rect 34792 81508 34840 81510
rect 34896 81508 34944 81510
rect 35000 81562 35048 81564
rect 35104 81562 35152 81564
rect 35000 81510 35016 81562
rect 35104 81510 35140 81562
rect 35000 81508 35048 81510
rect 35104 81508 35152 81510
rect 34008 81498 35208 81508
rect 34008 79996 35208 80006
rect 34064 79994 34112 79996
rect 34168 79994 34216 79996
rect 34076 79942 34112 79994
rect 34200 79942 34216 79994
rect 34064 79940 34112 79942
rect 34168 79940 34216 79942
rect 34272 79994 34320 79996
rect 34376 79994 34424 79996
rect 34480 79994 34528 79996
rect 34376 79942 34396 79994
rect 34480 79942 34520 79994
rect 34272 79940 34320 79942
rect 34376 79940 34424 79942
rect 34480 79940 34528 79942
rect 34584 79940 34632 79996
rect 34688 79994 34736 79996
rect 34792 79994 34840 79996
rect 34896 79994 34944 79996
rect 34696 79942 34736 79994
rect 34820 79942 34840 79994
rect 34688 79940 34736 79942
rect 34792 79940 34840 79942
rect 34896 79940 34944 79942
rect 35000 79994 35048 79996
rect 35104 79994 35152 79996
rect 35000 79942 35016 79994
rect 35104 79942 35140 79994
rect 35000 79940 35048 79942
rect 35104 79940 35152 79942
rect 34008 79930 35208 79940
rect 29596 78932 29876 78988
rect 23884 78036 23940 78204
rect 23436 76514 23492 76524
rect 23548 78034 23940 78036
rect 23548 77982 23886 78034
rect 23938 77982 23940 78034
rect 23548 77980 23940 77982
rect 21980 76468 22036 76478
rect 21868 76466 22036 76468
rect 21868 76414 21982 76466
rect 22034 76414 22036 76466
rect 21868 76412 22036 76414
rect 21980 76402 22036 76412
rect 23548 73948 23604 77980
rect 23884 77970 23940 77980
rect 24332 78484 24388 78494
rect 24332 78258 24388 78428
rect 24332 78206 24334 78258
rect 24386 78206 24388 78258
rect 24332 77812 24388 78206
rect 19852 73892 19908 73902
rect 20860 73892 21028 73948
rect 19404 73890 19908 73892
rect 19404 73838 19854 73890
rect 19906 73838 19908 73890
rect 19404 73836 19908 73838
rect 19404 73556 19460 73836
rect 19852 73826 19908 73836
rect 19404 73490 19460 73500
rect 20636 73444 20692 73454
rect 20636 73350 20692 73388
rect 18284 71934 18286 71986
rect 18338 71934 18340 71986
rect 18284 71922 18340 71934
rect 19852 73106 19908 73118
rect 19852 73054 19854 73106
rect 19906 73054 19908 73106
rect 19852 71876 19908 73054
rect 17724 71538 17780 71550
rect 17724 71486 17726 71538
rect 17778 71486 17780 71538
rect 17724 70588 17780 71486
rect 19292 70980 19348 70990
rect 19292 70886 19348 70924
rect 19404 70868 19460 70878
rect 19852 70868 19908 71820
rect 20748 71764 20804 71774
rect 20300 71762 20804 71764
rect 20300 71710 20750 71762
rect 20802 71710 20804 71762
rect 20300 71708 20804 71710
rect 20300 71202 20356 71708
rect 20748 71698 20804 71708
rect 20300 71150 20302 71202
rect 20354 71150 20356 71202
rect 20300 71138 20356 71150
rect 19964 70980 20020 70990
rect 19964 70978 20132 70980
rect 19964 70926 19966 70978
rect 20018 70926 20132 70978
rect 19964 70924 20132 70926
rect 19964 70914 20020 70924
rect 19404 70866 19908 70868
rect 19404 70814 19406 70866
rect 19458 70814 19908 70866
rect 19404 70812 19908 70814
rect 19404 70802 19460 70812
rect 17724 70532 17892 70588
rect 15148 70418 15876 70420
rect 15148 70366 15150 70418
rect 15202 70366 15876 70418
rect 15148 70364 15876 70366
rect 15148 70354 15204 70364
rect 15036 70140 15428 70196
rect 13804 69682 13860 69692
rect 14252 69970 14308 69982
rect 14252 69918 14254 69970
rect 14306 69918 14308 69970
rect 14252 69636 14308 69918
rect 14252 69570 14308 69580
rect 14812 69636 14868 69646
rect 13804 69412 13860 69422
rect 13804 69410 13972 69412
rect 13804 69358 13806 69410
rect 13858 69358 13972 69410
rect 13804 69356 13972 69358
rect 13804 69346 13860 69356
rect 13916 69188 13972 69356
rect 14028 69300 14084 69310
rect 14028 69206 14084 69244
rect 14812 69298 14868 69580
rect 14924 69524 14980 69534
rect 14924 69430 14980 69468
rect 14812 69246 14814 69298
rect 14866 69246 14868 69298
rect 14812 69234 14868 69246
rect 15036 69298 15092 69310
rect 15036 69246 15038 69298
rect 15090 69246 15092 69298
rect 13916 69122 13972 69132
rect 15036 69188 15092 69246
rect 15036 69122 15092 69132
rect 14008 69020 15208 69030
rect 14064 69018 14112 69020
rect 14168 69018 14216 69020
rect 14076 68966 14112 69018
rect 14200 68966 14216 69018
rect 14064 68964 14112 68966
rect 14168 68964 14216 68966
rect 14272 69018 14320 69020
rect 14376 69018 14424 69020
rect 14480 69018 14528 69020
rect 14376 68966 14396 69018
rect 14480 68966 14520 69018
rect 14272 68964 14320 68966
rect 14376 68964 14424 68966
rect 14480 68964 14528 68966
rect 14584 68964 14632 69020
rect 14688 69018 14736 69020
rect 14792 69018 14840 69020
rect 14896 69018 14944 69020
rect 14696 68966 14736 69018
rect 14820 68966 14840 69018
rect 14688 68964 14736 68966
rect 14792 68964 14840 68966
rect 14896 68964 14944 68966
rect 15000 69018 15048 69020
rect 15104 69018 15152 69020
rect 15000 68966 15016 69018
rect 15104 68966 15140 69018
rect 15000 68964 15048 68966
rect 15104 68964 15152 68966
rect 14008 68954 15208 68964
rect 15372 68850 15428 70140
rect 15596 70194 15652 70206
rect 15596 70142 15598 70194
rect 15650 70142 15652 70194
rect 15484 69970 15540 69982
rect 15484 69918 15486 69970
rect 15538 69918 15540 69970
rect 15484 69412 15540 69918
rect 15596 69524 15652 70142
rect 15596 69458 15652 69468
rect 15708 69636 15764 69646
rect 15484 69346 15540 69356
rect 15596 69300 15652 69310
rect 15708 69300 15764 69580
rect 15820 69524 15876 70364
rect 16380 70418 16660 70420
rect 16380 70366 16606 70418
rect 16658 70366 16660 70418
rect 16380 70364 16660 70366
rect 16044 70308 16100 70318
rect 16044 70214 16100 70252
rect 15932 70194 15988 70206
rect 15932 70142 15934 70194
rect 15986 70142 15988 70194
rect 15932 69636 15988 70142
rect 16268 70194 16324 70206
rect 16268 70142 16270 70194
rect 16322 70142 16324 70194
rect 15932 69580 16212 69636
rect 16156 69524 16212 69580
rect 15820 69468 16100 69524
rect 15596 69298 15764 69300
rect 15596 69246 15598 69298
rect 15650 69246 15764 69298
rect 15596 69244 15764 69246
rect 16044 69298 16100 69468
rect 16044 69246 16046 69298
rect 16098 69246 16100 69298
rect 15372 68798 15374 68850
rect 15426 68798 15428 68850
rect 15372 68786 15428 68798
rect 15484 69186 15540 69198
rect 15484 69134 15486 69186
rect 15538 69134 15540 69186
rect 15260 68740 15316 68750
rect 14812 67956 14868 67966
rect 14812 67954 15092 67956
rect 14812 67902 14814 67954
rect 14866 67902 15092 67954
rect 14812 67900 15092 67902
rect 14812 67890 14868 67900
rect 14476 67844 14532 67854
rect 14476 67750 14532 67788
rect 14028 67732 14084 67742
rect 14028 67638 14084 67676
rect 14252 67730 14308 67742
rect 14252 67678 14254 67730
rect 14306 67678 14308 67730
rect 14252 67620 14308 67678
rect 14588 67732 14644 67742
rect 14644 67676 14756 67732
rect 14588 67666 14644 67676
rect 14252 67554 14308 67564
rect 14700 67618 14756 67676
rect 14700 67566 14702 67618
rect 14754 67566 14756 67618
rect 14700 67554 14756 67566
rect 14812 67620 14868 67658
rect 15036 67620 15092 67900
rect 15260 67842 15316 68684
rect 15260 67790 15262 67842
rect 15314 67790 15316 67842
rect 15260 67778 15316 67790
rect 15036 67564 15428 67620
rect 14812 67554 14868 67564
rect 14008 67452 15208 67462
rect 14064 67450 14112 67452
rect 14168 67450 14216 67452
rect 14076 67398 14112 67450
rect 14200 67398 14216 67450
rect 14064 67396 14112 67398
rect 14168 67396 14216 67398
rect 14272 67450 14320 67452
rect 14376 67450 14424 67452
rect 14480 67450 14528 67452
rect 14376 67398 14396 67450
rect 14480 67398 14520 67450
rect 14272 67396 14320 67398
rect 14376 67396 14424 67398
rect 14480 67396 14528 67398
rect 14584 67396 14632 67452
rect 14688 67450 14736 67452
rect 14792 67450 14840 67452
rect 14896 67450 14944 67452
rect 14696 67398 14736 67450
rect 14820 67398 14840 67450
rect 14688 67396 14736 67398
rect 14792 67396 14840 67398
rect 14896 67396 14944 67398
rect 15000 67450 15048 67452
rect 15104 67450 15152 67452
rect 15000 67398 15016 67450
rect 15104 67398 15140 67450
rect 15000 67396 15048 67398
rect 15104 67396 15152 67398
rect 14008 67386 15208 67396
rect 14924 67284 14980 67294
rect 13916 67172 13972 67182
rect 13916 67078 13972 67116
rect 13244 65324 13412 65380
rect 13468 66780 13748 66836
rect 14924 66946 14980 67228
rect 15260 67060 15316 67070
rect 15372 67060 15428 67564
rect 15484 67170 15540 69134
rect 15596 67732 15652 69244
rect 15820 69188 15876 69198
rect 15820 69094 15876 69132
rect 15596 67666 15652 67676
rect 15708 68964 15764 68974
rect 15708 67282 15764 68908
rect 15932 68850 15988 68862
rect 15932 68798 15934 68850
rect 15986 68798 15988 68850
rect 15820 68740 15876 68750
rect 15932 68740 15988 68798
rect 16044 68852 16100 69246
rect 16044 68786 16100 68796
rect 15876 68684 15988 68740
rect 15820 68674 15876 68684
rect 16156 68628 16212 69468
rect 15708 67230 15710 67282
rect 15762 67230 15764 67282
rect 15708 67218 15764 67230
rect 15932 68572 16212 68628
rect 16268 68628 16324 70142
rect 16380 69298 16436 70364
rect 16604 70354 16660 70364
rect 16492 70196 16548 70206
rect 16716 70196 16772 70206
rect 16548 70140 16660 70196
rect 16492 70130 16548 70140
rect 16380 69246 16382 69298
rect 16434 69246 16436 69298
rect 16380 69234 16436 69246
rect 16492 69412 16548 69422
rect 15484 67118 15486 67170
rect 15538 67118 15540 67170
rect 15484 67106 15540 67118
rect 15932 67172 15988 68572
rect 16268 68562 16324 68572
rect 16492 68740 16548 69356
rect 16492 68626 16548 68684
rect 16492 68574 16494 68626
rect 16546 68574 16548 68626
rect 16492 68562 16548 68574
rect 16604 69076 16660 70140
rect 16716 70102 16772 70140
rect 17500 70194 17556 70206
rect 17500 70142 17502 70194
rect 17554 70142 17556 70194
rect 16156 68402 16212 68414
rect 16156 68350 16158 68402
rect 16210 68350 16212 68402
rect 16156 67620 16212 68350
rect 16156 67554 16212 67564
rect 16268 68068 16324 68078
rect 15260 67058 15428 67060
rect 15260 67006 15262 67058
rect 15314 67006 15428 67058
rect 15260 67004 15428 67006
rect 15260 66994 15316 67004
rect 14924 66894 14926 66946
rect 14978 66894 14980 66946
rect 13244 64932 13300 65324
rect 13468 65156 13524 66780
rect 14924 66612 14980 66894
rect 14924 66556 15428 66612
rect 14008 65884 15208 65894
rect 14064 65882 14112 65884
rect 14168 65882 14216 65884
rect 14076 65830 14112 65882
rect 14200 65830 14216 65882
rect 14064 65828 14112 65830
rect 14168 65828 14216 65830
rect 14272 65882 14320 65884
rect 14376 65882 14424 65884
rect 14480 65882 14528 65884
rect 14376 65830 14396 65882
rect 14480 65830 14520 65882
rect 14272 65828 14320 65830
rect 14376 65828 14424 65830
rect 14480 65828 14528 65830
rect 14584 65828 14632 65884
rect 14688 65882 14736 65884
rect 14792 65882 14840 65884
rect 14896 65882 14944 65884
rect 14696 65830 14736 65882
rect 14820 65830 14840 65882
rect 14688 65828 14736 65830
rect 14792 65828 14840 65830
rect 14896 65828 14944 65830
rect 15000 65882 15048 65884
rect 15104 65882 15152 65884
rect 15000 65830 15016 65882
rect 15104 65830 15140 65882
rect 15000 65828 15048 65830
rect 15104 65828 15152 65830
rect 14008 65818 15208 65828
rect 14028 65604 14084 65614
rect 13916 65602 14084 65604
rect 13916 65550 14030 65602
rect 14082 65550 14084 65602
rect 13916 65548 14084 65550
rect 13580 65490 13636 65502
rect 13580 65438 13582 65490
rect 13634 65438 13636 65490
rect 13580 65380 13636 65438
rect 13580 65314 13636 65324
rect 13804 65490 13860 65502
rect 13804 65438 13806 65490
rect 13858 65438 13860 65490
rect 13804 65156 13860 65438
rect 13916 65268 13972 65548
rect 14028 65538 14084 65548
rect 13916 65202 13972 65212
rect 14028 65380 14084 65390
rect 13468 65100 13636 65156
rect 13244 64866 13300 64876
rect 13188 64652 13300 64708
rect 13132 64642 13188 64652
rect 12572 64594 12628 64606
rect 12572 64542 12574 64594
rect 12626 64542 12628 64594
rect 12572 64484 12628 64542
rect 12572 64418 12628 64428
rect 12908 64594 12964 64606
rect 12908 64542 12910 64594
rect 12962 64542 12964 64594
rect 12460 64094 12462 64146
rect 12514 64094 12516 64146
rect 12348 63250 12404 63262
rect 12348 63198 12350 63250
rect 12402 63198 12404 63250
rect 12348 62916 12404 63198
rect 12460 63028 12516 64094
rect 12516 62972 12740 63028
rect 12460 62962 12516 62972
rect 12348 62850 12404 62860
rect 12012 61518 12014 61570
rect 12066 61518 12068 61570
rect 12012 61506 12068 61518
rect 12124 61908 12180 61918
rect 11340 61346 11396 61358
rect 11340 61294 11342 61346
rect 11394 61294 11396 61346
rect 11340 61236 11396 61294
rect 12124 61346 12180 61852
rect 12124 61294 12126 61346
rect 12178 61294 12180 61346
rect 12124 61282 12180 61294
rect 12348 61458 12404 61470
rect 12348 61406 12350 61458
rect 12402 61406 12404 61458
rect 12348 61348 12404 61406
rect 12348 61282 12404 61292
rect 11340 61170 11396 61180
rect 12684 60676 12740 62972
rect 12908 62580 12964 64542
rect 12908 62514 12964 62524
rect 13132 63924 13188 63934
rect 12796 62468 12852 62478
rect 12796 62132 12852 62412
rect 12796 61794 12852 62076
rect 13132 61908 13188 63868
rect 13244 62356 13300 64652
rect 13468 64596 13524 64606
rect 13468 64502 13524 64540
rect 13580 64372 13636 65100
rect 13804 65090 13860 65100
rect 13916 64932 13972 64942
rect 13916 64706 13972 64876
rect 13916 64654 13918 64706
rect 13970 64654 13972 64706
rect 13916 64642 13972 64654
rect 14028 64706 14084 65324
rect 14476 65380 14532 65390
rect 14476 65378 14756 65380
rect 14476 65326 14478 65378
rect 14530 65326 14756 65378
rect 14476 65324 14756 65326
rect 14476 65314 14532 65324
rect 14140 65266 14196 65278
rect 14140 65214 14142 65266
rect 14194 65214 14196 65266
rect 14140 65156 14196 65214
rect 14140 65090 14196 65100
rect 14028 64654 14030 64706
rect 14082 64654 14084 64706
rect 14028 64642 14084 64654
rect 14588 64708 14644 64718
rect 14476 64594 14532 64606
rect 14476 64542 14478 64594
rect 14530 64542 14532 64594
rect 13468 64316 13636 64372
rect 13692 64482 13748 64494
rect 13692 64430 13694 64482
rect 13746 64430 13748 64482
rect 13244 62290 13300 62300
rect 13356 62468 13412 62478
rect 12796 61742 12798 61794
rect 12850 61742 12852 61794
rect 12796 61730 12852 61742
rect 12908 61852 13132 61908
rect 12908 61570 12964 61852
rect 13132 61842 13188 61852
rect 12908 61518 12910 61570
rect 12962 61518 12964 61570
rect 12908 61506 12964 61518
rect 11676 60116 11732 60126
rect 12684 60116 12740 60620
rect 13356 60564 13412 62412
rect 13468 60788 13524 64316
rect 13692 64036 13748 64430
rect 13580 63980 13748 64036
rect 13804 64482 13860 64494
rect 13804 64430 13806 64482
rect 13858 64430 13860 64482
rect 13580 63476 13636 63980
rect 13692 63810 13748 63822
rect 13692 63758 13694 63810
rect 13746 63758 13748 63810
rect 13692 63700 13748 63758
rect 13804 63812 13860 64430
rect 14476 64484 14532 64542
rect 14588 64594 14644 64652
rect 14588 64542 14590 64594
rect 14642 64542 14644 64594
rect 14588 64530 14644 64542
rect 14700 64596 14756 65324
rect 14812 64932 14868 64942
rect 14812 64706 14868 64876
rect 14812 64654 14814 64706
rect 14866 64654 14868 64706
rect 14812 64642 14868 64654
rect 14700 64530 14756 64540
rect 15372 64596 15428 66556
rect 15932 66386 15988 67116
rect 15932 66334 15934 66386
rect 15986 66334 15988 66386
rect 15932 66322 15988 66334
rect 16268 67058 16324 68012
rect 16492 67732 16548 67742
rect 16492 67638 16548 67676
rect 16268 67006 16270 67058
rect 16322 67006 16324 67058
rect 16268 66386 16324 67006
rect 16604 67060 16660 69020
rect 16828 69970 16884 69982
rect 16828 69918 16830 69970
rect 16882 69918 16884 69970
rect 16716 68516 16772 68526
rect 16716 67732 16772 68460
rect 16716 67666 16772 67676
rect 16716 67060 16772 67070
rect 16604 67004 16716 67060
rect 16716 66966 16772 67004
rect 16268 66334 16270 66386
rect 16322 66334 16324 66386
rect 16268 66322 16324 66334
rect 15820 65380 15876 65390
rect 15372 64530 15428 64540
rect 15484 64818 15540 64830
rect 15484 64766 15486 64818
rect 15538 64766 15540 64818
rect 14476 64418 14532 64428
rect 14008 64316 15208 64326
rect 14064 64314 14112 64316
rect 14168 64314 14216 64316
rect 14076 64262 14112 64314
rect 14200 64262 14216 64314
rect 14064 64260 14112 64262
rect 14168 64260 14216 64262
rect 14272 64314 14320 64316
rect 14376 64314 14424 64316
rect 14480 64314 14528 64316
rect 14376 64262 14396 64314
rect 14480 64262 14520 64314
rect 14272 64260 14320 64262
rect 14376 64260 14424 64262
rect 14480 64260 14528 64262
rect 14584 64260 14632 64316
rect 14688 64314 14736 64316
rect 14792 64314 14840 64316
rect 14896 64314 14944 64316
rect 14696 64262 14736 64314
rect 14820 64262 14840 64314
rect 14688 64260 14736 64262
rect 14792 64260 14840 64262
rect 14896 64260 14944 64262
rect 15000 64314 15048 64316
rect 15104 64314 15152 64316
rect 15000 64262 15016 64314
rect 15104 64262 15140 64314
rect 15000 64260 15048 64262
rect 15104 64260 15152 64262
rect 14008 64250 15208 64260
rect 15372 64260 15428 64270
rect 14700 64148 14756 64158
rect 14700 64034 14756 64092
rect 14700 63982 14702 64034
rect 14754 63982 14756 64034
rect 14700 63970 14756 63982
rect 15260 64148 15316 64158
rect 13804 63746 13860 63756
rect 13916 63924 13972 63934
rect 13916 63810 13972 63868
rect 15260 63922 15316 64092
rect 15260 63870 15262 63922
rect 15314 63870 15316 63922
rect 15260 63858 15316 63870
rect 13916 63758 13918 63810
rect 13970 63758 13972 63810
rect 13916 63746 13972 63758
rect 14924 63812 14980 63822
rect 13692 63634 13748 63644
rect 14252 63700 14308 63710
rect 14252 63606 14308 63644
rect 13804 63588 13860 63598
rect 13804 63476 13860 63532
rect 13580 63410 13636 63420
rect 13692 63420 13860 63476
rect 13580 63252 13636 63262
rect 13580 63158 13636 63196
rect 13580 63028 13636 63038
rect 13580 62578 13636 62972
rect 13580 62526 13582 62578
rect 13634 62526 13636 62578
rect 13580 62132 13636 62526
rect 13580 62066 13636 62076
rect 13580 61572 13636 61582
rect 13692 61572 13748 63420
rect 14924 63138 14980 63756
rect 14924 63086 14926 63138
rect 14978 63086 14980 63138
rect 14924 63074 14980 63086
rect 14476 63028 14532 63038
rect 14028 62916 14084 62954
rect 14476 62934 14532 62972
rect 15260 63028 15316 63038
rect 15260 62934 15316 62972
rect 14028 62850 14084 62860
rect 14008 62748 15208 62758
rect 14064 62746 14112 62748
rect 14168 62746 14216 62748
rect 13804 62692 13860 62702
rect 14076 62694 14112 62746
rect 14200 62694 14216 62746
rect 14064 62692 14112 62694
rect 14168 62692 14216 62694
rect 14272 62746 14320 62748
rect 14376 62746 14424 62748
rect 14480 62746 14528 62748
rect 14376 62694 14396 62746
rect 14480 62694 14520 62746
rect 14272 62692 14320 62694
rect 14376 62692 14424 62694
rect 14480 62692 14528 62694
rect 14584 62692 14632 62748
rect 14688 62746 14736 62748
rect 14792 62746 14840 62748
rect 14896 62746 14944 62748
rect 14696 62694 14736 62746
rect 14820 62694 14840 62746
rect 14688 62692 14736 62694
rect 14792 62692 14840 62694
rect 14896 62692 14944 62694
rect 15000 62746 15048 62748
rect 15104 62746 15152 62748
rect 15000 62694 15016 62746
rect 15104 62694 15140 62746
rect 15000 62692 15048 62694
rect 15104 62692 15152 62694
rect 14008 62682 15208 62692
rect 13804 62188 13860 62636
rect 14364 62580 14420 62590
rect 14364 62486 14420 62524
rect 14588 62468 14644 62478
rect 14644 62412 14868 62468
rect 14588 62402 14644 62412
rect 14812 62354 14868 62412
rect 14812 62302 14814 62354
rect 14866 62302 14868 62354
rect 14812 62290 14868 62302
rect 14924 62356 14980 62366
rect 13916 62244 13972 62254
rect 13804 62132 13972 62188
rect 13580 61570 13748 61572
rect 13580 61518 13582 61570
rect 13634 61518 13748 61570
rect 13580 61516 13748 61518
rect 13804 61684 13860 61694
rect 13804 61570 13860 61628
rect 13804 61518 13806 61570
rect 13858 61518 13860 61570
rect 13580 61506 13636 61516
rect 13804 61506 13860 61518
rect 13692 61348 13748 61358
rect 13916 61348 13972 62132
rect 14588 62244 14644 62282
rect 14924 62262 14980 62300
rect 15372 62356 15428 64204
rect 15484 63250 15540 64766
rect 15596 64708 15652 64718
rect 15596 64706 15764 64708
rect 15596 64654 15598 64706
rect 15650 64654 15764 64706
rect 15596 64652 15764 64654
rect 15596 64642 15652 64652
rect 15596 63924 15652 63934
rect 15596 63830 15652 63868
rect 15484 63198 15486 63250
rect 15538 63198 15540 63250
rect 15484 63186 15540 63198
rect 15708 62692 15764 64652
rect 15372 62262 15428 62300
rect 15484 62636 15764 62692
rect 15820 63700 15876 65324
rect 16156 64932 16212 64942
rect 16156 64838 16212 64876
rect 16044 64706 16100 64718
rect 16044 64654 16046 64706
rect 16098 64654 16100 64706
rect 16044 64146 16100 64654
rect 16716 64484 16772 64494
rect 16044 64094 16046 64146
rect 16098 64094 16100 64146
rect 16044 64082 16100 64094
rect 16492 64428 16716 64484
rect 16156 64036 16212 64046
rect 16156 63942 16212 63980
rect 14588 62020 14644 62188
rect 14588 61954 14644 61964
rect 15036 62244 15092 62254
rect 14924 61684 14980 61722
rect 14924 61618 14980 61628
rect 15036 61570 15092 62188
rect 15372 62020 15428 62030
rect 15372 61682 15428 61964
rect 15372 61630 15374 61682
rect 15426 61630 15428 61682
rect 15372 61618 15428 61630
rect 15484 61684 15540 62636
rect 15708 62468 15764 62478
rect 15708 62244 15764 62412
rect 15820 62466 15876 63644
rect 15932 63138 15988 63150
rect 15932 63086 15934 63138
rect 15986 63086 15988 63138
rect 15932 62580 15988 63086
rect 16380 63138 16436 63150
rect 16380 63086 16382 63138
rect 16434 63086 16436 63138
rect 16380 63028 16436 63086
rect 15932 62514 15988 62524
rect 16268 62580 16324 62590
rect 16380 62580 16436 62972
rect 16268 62578 16436 62580
rect 16268 62526 16270 62578
rect 16322 62526 16436 62578
rect 16268 62524 16436 62526
rect 16268 62514 16324 62524
rect 15820 62414 15822 62466
rect 15874 62414 15876 62466
rect 15820 62402 15876 62414
rect 16380 62468 16436 62524
rect 16380 62402 16436 62412
rect 16044 62356 16100 62366
rect 15708 62188 15876 62244
rect 15596 62132 15652 62142
rect 15596 62130 15764 62132
rect 15596 62078 15598 62130
rect 15650 62078 15764 62130
rect 15596 62076 15764 62078
rect 15596 62066 15652 62076
rect 15596 61908 15652 61918
rect 15596 61794 15652 61852
rect 15596 61742 15598 61794
rect 15650 61742 15652 61794
rect 15596 61730 15652 61742
rect 15484 61618 15540 61628
rect 15708 61572 15764 62076
rect 15820 61794 15876 62188
rect 16044 62188 16100 62300
rect 15820 61742 15822 61794
rect 15874 61742 15876 61794
rect 15820 61730 15876 61742
rect 15932 62130 15988 62142
rect 16044 62132 16436 62188
rect 15932 62078 15934 62130
rect 15986 62078 15988 62130
rect 15036 61518 15038 61570
rect 15090 61518 15092 61570
rect 15036 61506 15092 61518
rect 15596 61516 15764 61572
rect 13580 61292 13692 61348
rect 13580 61010 13636 61292
rect 13692 61282 13748 61292
rect 13804 61292 13972 61348
rect 14924 61458 14980 61470
rect 14924 61406 14926 61458
rect 14978 61406 14980 61458
rect 14924 61348 14980 61406
rect 14924 61292 15428 61348
rect 13580 60958 13582 61010
rect 13634 60958 13636 61010
rect 13580 60946 13636 60958
rect 13692 61012 13748 61022
rect 13804 61012 13860 61292
rect 14008 61180 15208 61190
rect 14064 61178 14112 61180
rect 14168 61178 14216 61180
rect 14076 61126 14112 61178
rect 14200 61126 14216 61178
rect 14064 61124 14112 61126
rect 14168 61124 14216 61126
rect 14272 61178 14320 61180
rect 14376 61178 14424 61180
rect 14480 61178 14528 61180
rect 14376 61126 14396 61178
rect 14480 61126 14520 61178
rect 14272 61124 14320 61126
rect 14376 61124 14424 61126
rect 14480 61124 14528 61126
rect 14584 61124 14632 61180
rect 14688 61178 14736 61180
rect 14792 61178 14840 61180
rect 14896 61178 14944 61180
rect 14696 61126 14736 61178
rect 14820 61126 14840 61178
rect 14688 61124 14736 61126
rect 14792 61124 14840 61126
rect 14896 61124 14944 61126
rect 15000 61178 15048 61180
rect 15104 61178 15152 61180
rect 15000 61126 15016 61178
rect 15104 61126 15140 61178
rect 15000 61124 15048 61126
rect 15104 61124 15152 61126
rect 14008 61114 15208 61124
rect 13692 61010 13860 61012
rect 13692 60958 13694 61010
rect 13746 60958 13860 61010
rect 13692 60956 13860 60958
rect 13692 60946 13748 60956
rect 13468 60732 13748 60788
rect 13468 60564 13524 60574
rect 13356 60562 13524 60564
rect 13356 60510 13470 60562
rect 13522 60510 13524 60562
rect 13356 60508 13524 60510
rect 13468 60498 13524 60508
rect 13580 60564 13636 60574
rect 12796 60116 12852 60126
rect 11676 59444 11732 60060
rect 12348 60114 12852 60116
rect 12348 60062 12798 60114
rect 12850 60062 12852 60114
rect 12348 60060 12852 60062
rect 11676 59442 12068 59444
rect 11676 59390 11678 59442
rect 11730 59390 12068 59442
rect 11676 59388 12068 59390
rect 11676 59378 11732 59388
rect 11340 59106 11396 59118
rect 11340 59054 11342 59106
rect 11394 59054 11396 59106
rect 11340 57652 11396 59054
rect 11900 57762 11956 57774
rect 11900 57710 11902 57762
rect 11954 57710 11956 57762
rect 11340 57586 11396 57596
rect 11788 57652 11844 57662
rect 11788 57558 11844 57596
rect 11900 57316 11956 57710
rect 11788 57260 11956 57316
rect 11564 57204 11620 57214
rect 11340 56868 11396 56878
rect 11340 56774 11396 56812
rect 11564 56866 11620 57148
rect 11676 56980 11732 56990
rect 11676 56886 11732 56924
rect 11564 56814 11566 56866
rect 11618 56814 11620 56866
rect 11564 56802 11620 56814
rect 11340 56644 11396 56654
rect 11340 54628 11396 56588
rect 11788 56196 11844 57260
rect 11900 57092 11956 57102
rect 11900 56866 11956 57036
rect 11900 56814 11902 56866
rect 11954 56814 11956 56866
rect 11900 56802 11956 56814
rect 11788 56130 11844 56140
rect 11452 56082 11508 56094
rect 11452 56030 11454 56082
rect 11506 56030 11508 56082
rect 11452 55076 11508 56030
rect 11676 56084 11732 56094
rect 11676 55990 11732 56028
rect 11900 55972 11956 55982
rect 11788 55970 11956 55972
rect 11788 55918 11902 55970
rect 11954 55918 11956 55970
rect 11788 55916 11956 55918
rect 11676 55524 11732 55534
rect 11452 55010 11508 55020
rect 11564 55076 11620 55086
rect 11676 55076 11732 55468
rect 11788 55522 11844 55916
rect 11900 55906 11956 55916
rect 12012 55636 12068 59388
rect 12124 58212 12180 58222
rect 12348 58212 12404 60060
rect 12796 60050 12852 60060
rect 13580 59444 13636 60508
rect 13580 59378 13636 59388
rect 13020 59332 13076 59342
rect 13020 59238 13076 59276
rect 12572 59220 12628 59230
rect 12124 58210 12404 58212
rect 12124 58158 12126 58210
rect 12178 58158 12404 58210
rect 12124 58156 12404 58158
rect 12460 59106 12516 59118
rect 12460 59054 12462 59106
rect 12514 59054 12516 59106
rect 12460 58548 12516 59054
rect 12124 58146 12180 58156
rect 12124 56980 12180 56990
rect 12124 56866 12180 56924
rect 12124 56814 12126 56866
rect 12178 56814 12180 56866
rect 12124 56802 12180 56814
rect 11788 55470 11790 55522
rect 11842 55470 11844 55522
rect 11788 55458 11844 55470
rect 11900 55580 12068 55636
rect 12236 56532 12292 58156
rect 11564 55074 11732 55076
rect 11564 55022 11566 55074
rect 11618 55022 11732 55074
rect 11564 55020 11732 55022
rect 11564 55010 11620 55020
rect 11340 54562 11396 54572
rect 11564 54740 11620 54750
rect 11452 54404 11508 54414
rect 11452 53732 11508 54348
rect 11452 53666 11508 53676
rect 11564 53730 11620 54684
rect 11564 53678 11566 53730
rect 11618 53678 11620 53730
rect 11564 53666 11620 53678
rect 11676 53508 11732 55020
rect 11900 54738 11956 55580
rect 11900 54686 11902 54738
rect 11954 54686 11956 54738
rect 11900 54674 11956 54686
rect 12012 55076 12068 55086
rect 11228 53218 11284 53228
rect 11340 53452 11732 53508
rect 11228 52500 11284 52510
rect 11228 52162 11284 52444
rect 11228 52110 11230 52162
rect 11282 52110 11284 52162
rect 11228 52098 11284 52110
rect 11228 49812 11284 49822
rect 11228 49718 11284 49756
rect 11228 49364 11284 49374
rect 11228 49138 11284 49308
rect 11228 49086 11230 49138
rect 11282 49086 11284 49138
rect 11228 49074 11284 49086
rect 10780 48188 11172 48244
rect 10108 44258 10164 44268
rect 10220 45836 10500 45892
rect 10668 47460 10724 47470
rect 10108 44098 10164 44110
rect 10108 44046 10110 44098
rect 10162 44046 10164 44098
rect 10108 43764 10164 44046
rect 9996 43426 10052 43438
rect 9996 43374 9998 43426
rect 10050 43374 10052 43426
rect 9996 43092 10052 43374
rect 9996 43026 10052 43036
rect 9996 42868 10052 42878
rect 9996 42084 10052 42812
rect 10108 42866 10164 43708
rect 10108 42814 10110 42866
rect 10162 42814 10164 42866
rect 10108 42802 10164 42814
rect 9996 41186 10052 42028
rect 9996 41134 9998 41186
rect 10050 41134 10052 41186
rect 9996 41122 10052 41134
rect 10108 42196 10164 42206
rect 10108 40964 10164 42140
rect 10220 41300 10276 45836
rect 10556 45108 10612 45118
rect 10444 44994 10500 45006
rect 10444 44942 10446 44994
rect 10498 44942 10500 44994
rect 10444 44882 10500 44942
rect 10444 44830 10446 44882
rect 10498 44830 10500 44882
rect 10444 44818 10500 44830
rect 10556 44434 10612 45052
rect 10668 44884 10724 47404
rect 10780 46898 10836 48188
rect 11340 47796 11396 53452
rect 11564 53284 11620 53294
rect 11452 52276 11508 52286
rect 11452 52162 11508 52220
rect 11452 52110 11454 52162
rect 11506 52110 11508 52162
rect 11452 52098 11508 52110
rect 11564 50428 11620 53228
rect 11788 52724 11844 52734
rect 11844 52668 11956 52724
rect 11788 52658 11844 52668
rect 11788 52276 11844 52286
rect 11788 52182 11844 52220
rect 11900 52050 11956 52668
rect 11900 51998 11902 52050
rect 11954 51998 11956 52050
rect 11900 51986 11956 51998
rect 10780 46846 10782 46898
rect 10834 46846 10836 46898
rect 10780 46834 10836 46846
rect 10892 47740 11396 47796
rect 11452 50372 11620 50428
rect 11676 51940 11732 51950
rect 11676 51602 11732 51884
rect 11676 51550 11678 51602
rect 11730 51550 11732 51602
rect 11676 50428 11732 51550
rect 11676 50372 11844 50428
rect 10892 45892 10948 47740
rect 11004 47458 11060 47470
rect 11004 47406 11006 47458
rect 11058 47406 11060 47458
rect 11004 46676 11060 47406
rect 11228 47348 11284 47358
rect 11228 47254 11284 47292
rect 11452 47012 11508 50372
rect 11676 49812 11732 49822
rect 11564 49364 11620 49374
rect 11564 49026 11620 49308
rect 11676 49138 11732 49756
rect 11788 49364 11844 50372
rect 11788 49298 11844 49308
rect 11676 49086 11678 49138
rect 11730 49086 11732 49138
rect 11676 49074 11732 49086
rect 11564 48974 11566 49026
rect 11618 48974 11620 49026
rect 11564 48962 11620 48974
rect 11788 48804 11844 48814
rect 11788 48710 11844 48748
rect 11004 46610 11060 46620
rect 11340 46956 11508 47012
rect 11676 48244 11732 48254
rect 10780 45890 10948 45892
rect 10780 45838 10894 45890
rect 10946 45838 10948 45890
rect 10780 45836 10948 45838
rect 10780 45108 10836 45836
rect 10892 45826 10948 45836
rect 11340 45556 11396 46956
rect 11116 45500 11396 45556
rect 11452 46786 11508 46798
rect 11452 46734 11454 46786
rect 11506 46734 11508 46786
rect 11452 46564 11508 46734
rect 11452 45778 11508 46508
rect 11452 45726 11454 45778
rect 11506 45726 11508 45778
rect 10892 45444 10948 45454
rect 10892 45330 10948 45388
rect 10892 45278 10894 45330
rect 10946 45278 10948 45330
rect 10892 45266 10948 45278
rect 10780 45042 10836 45052
rect 10668 44828 10836 44884
rect 10556 44382 10558 44434
rect 10610 44382 10612 44434
rect 10556 44212 10612 44382
rect 10612 44156 10724 44212
rect 10556 44146 10612 44156
rect 10668 43762 10724 44156
rect 10668 43710 10670 43762
rect 10722 43710 10724 43762
rect 10668 43540 10724 43710
rect 10668 43474 10724 43484
rect 10780 43316 10836 44828
rect 11004 44436 11060 44446
rect 10556 43260 10836 43316
rect 10892 44380 11004 44436
rect 10220 41234 10276 41244
rect 10332 42754 10388 42766
rect 10332 42702 10334 42754
rect 10386 42702 10388 42754
rect 10332 42196 10388 42702
rect 10556 42532 10612 43260
rect 10668 42868 10724 42878
rect 10668 42866 10836 42868
rect 10668 42814 10670 42866
rect 10722 42814 10836 42866
rect 10668 42812 10836 42814
rect 10668 42802 10724 42812
rect 10780 42644 10836 42812
rect 10892 42756 10948 44380
rect 11004 44370 11060 44380
rect 11004 44100 11060 44110
rect 11004 44006 11060 44044
rect 11116 43652 11172 45500
rect 11340 45332 11396 45342
rect 11340 45238 11396 45276
rect 11452 44882 11508 45726
rect 11452 44830 11454 44882
rect 11506 44830 11508 44882
rect 11452 44548 11508 44830
rect 11452 44492 11620 44548
rect 11340 44210 11396 44222
rect 11340 44158 11342 44210
rect 11394 44158 11396 44210
rect 11340 44100 11396 44158
rect 11452 44212 11508 44222
rect 11452 44118 11508 44156
rect 11340 44034 11396 44044
rect 11116 43586 11172 43596
rect 11452 43538 11508 43550
rect 11452 43486 11454 43538
rect 11506 43486 11508 43538
rect 11004 43428 11060 43438
rect 11452 43428 11508 43486
rect 11004 43426 11396 43428
rect 11004 43374 11006 43426
rect 11058 43374 11396 43426
rect 11004 43372 11396 43374
rect 11004 43362 11060 43372
rect 10892 42700 11284 42756
rect 10780 42588 11172 42644
rect 10556 42476 10836 42532
rect 10556 42196 10612 42206
rect 10332 42194 10612 42196
rect 10332 42142 10558 42194
rect 10610 42142 10612 42194
rect 10332 42140 10612 42142
rect 9996 40908 10164 40964
rect 9996 40516 10052 40908
rect 9996 40402 10052 40460
rect 9996 40350 9998 40402
rect 10050 40350 10052 40402
rect 9996 39732 10052 40350
rect 9996 39618 10052 39676
rect 9996 39566 9998 39618
rect 10050 39566 10052 39618
rect 9996 39554 10052 39566
rect 10332 38668 10388 42140
rect 10556 42130 10612 42140
rect 10668 41860 10724 41870
rect 10668 41188 10724 41804
rect 10668 41094 10724 41132
rect 10556 41076 10612 41086
rect 10556 40982 10612 41020
rect 10780 40964 10836 42476
rect 10892 42084 10948 42094
rect 10948 42028 11060 42084
rect 10892 42018 10948 42028
rect 9884 38210 9940 38220
rect 9996 38612 10388 38668
rect 10668 40908 10836 40964
rect 10668 38668 10724 40908
rect 11004 40628 11060 42028
rect 11116 41412 11172 42588
rect 11116 41318 11172 41356
rect 11116 40628 11172 40638
rect 11004 40626 11172 40628
rect 11004 40574 11118 40626
rect 11170 40574 11172 40626
rect 11004 40572 11172 40574
rect 11116 40562 11172 40572
rect 11228 40404 11284 42700
rect 11340 41410 11396 43372
rect 11452 43362 11508 43372
rect 11564 42532 11620 44492
rect 11676 44436 11732 48188
rect 12012 47068 12068 55020
rect 12236 54404 12292 56476
rect 12348 57652 12404 57662
rect 12348 55412 12404 57596
rect 12460 57428 12516 58492
rect 12572 57874 12628 59164
rect 13580 59108 13636 59118
rect 13468 59106 13636 59108
rect 13468 59054 13582 59106
rect 13634 59054 13636 59106
rect 13468 59052 13636 59054
rect 12684 58210 12740 58222
rect 12684 58158 12686 58210
rect 12738 58158 12740 58210
rect 12684 57988 12740 58158
rect 12684 57932 12964 57988
rect 12572 57822 12574 57874
rect 12626 57822 12628 57874
rect 12572 57810 12628 57822
rect 12460 57362 12516 57372
rect 12684 57762 12740 57774
rect 12684 57710 12686 57762
rect 12738 57710 12740 57762
rect 12460 56980 12516 56990
rect 12460 56886 12516 56924
rect 12572 56644 12628 56654
rect 12460 56642 12628 56644
rect 12460 56590 12574 56642
rect 12626 56590 12628 56642
rect 12460 56588 12628 56590
rect 12460 56308 12516 56588
rect 12572 56578 12628 56588
rect 12460 55860 12516 56252
rect 12460 55794 12516 55804
rect 12572 56420 12628 56430
rect 12572 56082 12628 56364
rect 12684 56308 12740 57710
rect 12796 57652 12852 57662
rect 12796 57558 12852 57596
rect 12796 57428 12852 57438
rect 12796 57090 12852 57372
rect 12796 57038 12798 57090
rect 12850 57038 12852 57090
rect 12796 57026 12852 57038
rect 12684 56242 12740 56252
rect 12572 56030 12574 56082
rect 12626 56030 12628 56082
rect 12572 55524 12628 56030
rect 12908 56084 12964 57932
rect 13468 57092 13524 59052
rect 13580 59042 13636 59052
rect 13580 58548 13636 58558
rect 13580 58454 13636 58492
rect 12908 56018 12964 56028
rect 13132 57036 13524 57092
rect 13580 57092 13636 57102
rect 13132 56868 13188 57036
rect 13580 56998 13636 57036
rect 13692 56868 13748 60732
rect 14008 59612 15208 59622
rect 14064 59610 14112 59612
rect 14168 59610 14216 59612
rect 14076 59558 14112 59610
rect 14200 59558 14216 59610
rect 14064 59556 14112 59558
rect 14168 59556 14216 59558
rect 14272 59610 14320 59612
rect 14376 59610 14424 59612
rect 14480 59610 14528 59612
rect 14376 59558 14396 59610
rect 14480 59558 14520 59610
rect 14272 59556 14320 59558
rect 14376 59556 14424 59558
rect 14480 59556 14528 59558
rect 14584 59556 14632 59612
rect 14688 59610 14736 59612
rect 14792 59610 14840 59612
rect 14896 59610 14944 59612
rect 14696 59558 14736 59610
rect 14820 59558 14840 59610
rect 14688 59556 14736 59558
rect 14792 59556 14840 59558
rect 14896 59556 14944 59558
rect 15000 59610 15048 59612
rect 15104 59610 15152 59612
rect 15000 59558 15016 59610
rect 15104 59558 15140 59610
rect 15000 59556 15048 59558
rect 15104 59556 15152 59558
rect 14008 59546 15208 59556
rect 13916 59444 13972 59454
rect 13916 58436 13972 59388
rect 14924 59444 14980 59454
rect 14028 59218 14084 59230
rect 14028 59166 14030 59218
rect 14082 59166 14084 59218
rect 14028 58884 14084 59166
rect 14476 59220 14532 59230
rect 14812 59220 14868 59230
rect 14476 59218 14868 59220
rect 14476 59166 14478 59218
rect 14530 59166 14814 59218
rect 14866 59166 14868 59218
rect 14476 59164 14868 59166
rect 14476 59154 14532 59164
rect 14812 59154 14868 59164
rect 14700 58996 14756 59006
rect 14700 58902 14756 58940
rect 14028 58818 14084 58828
rect 13916 58370 13972 58380
rect 14812 58436 14868 58446
rect 14812 58342 14868 58380
rect 14924 58212 14980 59388
rect 15372 59444 15428 61292
rect 15372 59378 15428 59388
rect 15036 59332 15092 59342
rect 15036 59330 15316 59332
rect 15036 59278 15038 59330
rect 15090 59278 15316 59330
rect 15036 59276 15316 59278
rect 15036 59266 15092 59276
rect 15260 58546 15316 59276
rect 15372 59220 15428 59230
rect 15372 59126 15428 59164
rect 15260 58494 15262 58546
rect 15314 58494 15316 58546
rect 15260 58482 15316 58494
rect 15036 58434 15092 58446
rect 15036 58382 15038 58434
rect 15090 58382 15092 58434
rect 15036 58324 15092 58382
rect 15036 58258 15092 58268
rect 14924 58146 14980 58156
rect 14008 58044 15208 58054
rect 14064 58042 14112 58044
rect 14168 58042 14216 58044
rect 14076 57990 14112 58042
rect 14200 57990 14216 58042
rect 14064 57988 14112 57990
rect 14168 57988 14216 57990
rect 14272 58042 14320 58044
rect 14376 58042 14424 58044
rect 14480 58042 14528 58044
rect 14376 57990 14396 58042
rect 14480 57990 14520 58042
rect 14272 57988 14320 57990
rect 14376 57988 14424 57990
rect 14480 57988 14528 57990
rect 14584 57988 14632 58044
rect 14688 58042 14736 58044
rect 14792 58042 14840 58044
rect 14896 58042 14944 58044
rect 14696 57990 14736 58042
rect 14820 57990 14840 58042
rect 14688 57988 14736 57990
rect 14792 57988 14840 57990
rect 14896 57988 14944 57990
rect 15000 58042 15048 58044
rect 15104 58042 15152 58044
rect 15000 57990 15016 58042
rect 15104 57990 15140 58042
rect 15000 57988 15048 57990
rect 15104 57988 15152 57990
rect 14008 57978 15208 57988
rect 15596 57988 15652 61516
rect 15932 61236 15988 62078
rect 16268 61346 16324 61358
rect 16268 61294 16270 61346
rect 16322 61294 16324 61346
rect 15932 61180 16100 61236
rect 15932 61012 15988 61022
rect 15932 60786 15988 60956
rect 15932 60734 15934 60786
rect 15986 60734 15988 60786
rect 15932 60722 15988 60734
rect 16044 60340 16100 61180
rect 16268 61012 16324 61294
rect 16268 60946 16324 60956
rect 16380 60786 16436 62132
rect 16380 60734 16382 60786
rect 16434 60734 16436 60786
rect 16380 60722 16436 60734
rect 16492 60788 16548 64428
rect 16716 64390 16772 64428
rect 16828 63476 16884 69918
rect 17500 69522 17556 70142
rect 17500 69470 17502 69522
rect 17554 69470 17556 69522
rect 17500 69458 17556 69470
rect 17724 70194 17780 70206
rect 17724 70142 17726 70194
rect 17778 70142 17780 70194
rect 16940 69410 16996 69422
rect 16940 69358 16942 69410
rect 16994 69358 16996 69410
rect 16940 68628 16996 69358
rect 17388 69412 17444 69422
rect 17388 69318 17444 69356
rect 17724 68964 17780 70142
rect 17836 70084 17892 70532
rect 17836 70018 17892 70028
rect 18172 70306 18228 70318
rect 18172 70254 18174 70306
rect 18226 70254 18228 70306
rect 17948 69412 18004 69422
rect 17724 68898 17780 68908
rect 17836 69300 17892 69310
rect 16940 68562 16996 68572
rect 17052 68852 17108 68862
rect 17052 66052 17108 68796
rect 17500 68628 17556 68638
rect 17500 68534 17556 68572
rect 17724 68628 17780 68638
rect 17836 68628 17892 69244
rect 17724 68626 17892 68628
rect 17724 68574 17726 68626
rect 17778 68574 17892 68626
rect 17724 68572 17892 68574
rect 17948 69298 18004 69356
rect 17948 69246 17950 69298
rect 18002 69246 18004 69298
rect 17724 68562 17780 68572
rect 17948 68516 18004 69246
rect 18172 68964 18228 70254
rect 18620 70306 18676 70318
rect 18620 70254 18622 70306
rect 18674 70254 18676 70306
rect 18508 70196 18564 70206
rect 18508 70102 18564 70140
rect 18620 69636 18676 70254
rect 19404 70084 19460 70094
rect 19460 70028 19572 70084
rect 19404 69990 19460 70028
rect 18172 68898 18228 68908
rect 18284 69580 18676 69636
rect 18284 68850 18340 69580
rect 18956 69524 19012 69534
rect 18396 69412 18452 69422
rect 18396 69318 18452 69356
rect 18956 69410 19012 69468
rect 18956 69358 18958 69410
rect 19010 69358 19012 69410
rect 18956 69346 19012 69358
rect 18508 69300 18564 69310
rect 18508 69206 18564 69244
rect 18732 69298 18788 69310
rect 18732 69246 18734 69298
rect 18786 69246 18788 69298
rect 18732 69076 18788 69246
rect 19404 69188 19460 69198
rect 19404 69094 19460 69132
rect 18732 69010 18788 69020
rect 19516 68964 19572 70028
rect 19740 69188 19796 69198
rect 19404 68908 19572 68964
rect 19628 69186 19796 69188
rect 19628 69134 19742 69186
rect 19794 69134 19796 69186
rect 19628 69132 19796 69134
rect 18284 68798 18286 68850
rect 18338 68798 18340 68850
rect 18284 68786 18340 68798
rect 19068 68852 19124 68862
rect 19068 68758 19124 68796
rect 17948 68422 18004 68460
rect 18172 68628 18228 68638
rect 17388 67844 17444 67854
rect 17276 67842 17444 67844
rect 17276 67790 17390 67842
rect 17442 67790 17444 67842
rect 17276 67788 17444 67790
rect 17164 67060 17220 67070
rect 17276 67060 17332 67788
rect 17388 67778 17444 67788
rect 17948 67732 18004 67742
rect 17724 67730 18004 67732
rect 17724 67678 17950 67730
rect 18002 67678 18004 67730
rect 17724 67676 18004 67678
rect 17220 67004 17332 67060
rect 17388 67620 17444 67630
rect 17612 67620 17668 67630
rect 17388 67058 17444 67564
rect 17388 67006 17390 67058
rect 17442 67006 17444 67058
rect 17164 66994 17220 67004
rect 17388 66994 17444 67006
rect 17500 67618 17668 67620
rect 17500 67566 17614 67618
rect 17666 67566 17668 67618
rect 17500 67564 17668 67566
rect 17164 66276 17220 66286
rect 17164 66182 17220 66220
rect 17164 66052 17220 66062
rect 17052 65996 17164 66052
rect 17164 65268 17220 65996
rect 17164 64818 17220 65212
rect 17164 64766 17166 64818
rect 17218 64766 17220 64818
rect 17164 64754 17220 64766
rect 17276 64708 17332 64718
rect 17276 64146 17332 64652
rect 17276 64094 17278 64146
rect 17330 64094 17332 64146
rect 17276 64082 17332 64094
rect 16828 63420 17220 63476
rect 16828 63252 16884 63262
rect 16828 63250 16996 63252
rect 16828 63198 16830 63250
rect 16882 63198 16996 63250
rect 16828 63196 16996 63198
rect 16828 63186 16884 63196
rect 16828 63028 16884 63038
rect 16828 62934 16884 62972
rect 16604 62916 16660 62926
rect 16604 62580 16660 62860
rect 16716 62580 16772 62590
rect 16604 62578 16772 62580
rect 16604 62526 16718 62578
rect 16770 62526 16772 62578
rect 16604 62524 16772 62526
rect 16716 62514 16772 62524
rect 16940 62244 16996 63196
rect 17052 62914 17108 62926
rect 17052 62862 17054 62914
rect 17106 62862 17108 62914
rect 17052 62356 17108 62862
rect 17164 62916 17220 63420
rect 17276 63252 17332 63262
rect 17276 63138 17332 63196
rect 17276 63086 17278 63138
rect 17330 63086 17332 63138
rect 17276 63074 17332 63086
rect 17164 62860 17332 62916
rect 17052 62290 17108 62300
rect 17164 62692 17220 62702
rect 16940 62178 16996 62188
rect 16828 62132 16884 62142
rect 16828 61684 16884 62076
rect 17164 61794 17220 62636
rect 17164 61742 17166 61794
rect 17218 61742 17220 61794
rect 17164 61730 17220 61742
rect 16940 61684 16996 61694
rect 16828 61628 16940 61684
rect 16940 61590 16996 61628
rect 16492 60722 16548 60732
rect 16156 60564 16212 60574
rect 16156 60470 16212 60508
rect 16492 60562 16548 60574
rect 16492 60510 16494 60562
rect 16546 60510 16548 60562
rect 16044 60284 16324 60340
rect 16044 59218 16100 59230
rect 16044 59166 16046 59218
rect 16098 59166 16100 59218
rect 15708 58324 15764 58334
rect 15708 58230 15764 58268
rect 15596 57932 15764 57988
rect 15036 57876 15092 57886
rect 14252 57762 14308 57774
rect 14252 57710 14254 57762
rect 14306 57710 14308 57762
rect 13804 57652 13860 57662
rect 14252 57652 14308 57710
rect 13804 57650 14308 57652
rect 13804 57598 13806 57650
rect 13858 57598 14308 57650
rect 13804 57596 14308 57598
rect 13804 57586 13860 57596
rect 13132 56082 13188 56812
rect 13580 56812 13748 56868
rect 13804 57428 13860 57438
rect 13132 56030 13134 56082
rect 13186 56030 13188 56082
rect 13132 56018 13188 56030
rect 13468 56754 13524 56766
rect 13468 56702 13470 56754
rect 13522 56702 13524 56754
rect 13468 56084 13524 56702
rect 13468 56018 13524 56028
rect 13244 55972 13300 55982
rect 13244 55970 13412 55972
rect 13244 55918 13246 55970
rect 13298 55918 13412 55970
rect 13244 55916 13412 55918
rect 13244 55906 13300 55916
rect 13020 55748 13076 55758
rect 12572 55458 12628 55468
rect 12908 55522 12964 55534
rect 12908 55470 12910 55522
rect 12962 55470 12964 55522
rect 12348 55188 12404 55356
rect 12460 55188 12516 55198
rect 12348 55132 12460 55188
rect 12460 55094 12516 55132
rect 12908 54516 12964 55470
rect 13020 55410 13076 55692
rect 13020 55358 13022 55410
rect 13074 55358 13076 55410
rect 13020 55346 13076 55358
rect 13020 54516 13076 54526
rect 12908 54514 13076 54516
rect 12908 54462 13022 54514
rect 13074 54462 13076 54514
rect 12908 54460 13076 54462
rect 13356 54516 13412 55916
rect 13468 54516 13524 54526
rect 13356 54514 13524 54516
rect 13356 54462 13470 54514
rect 13522 54462 13524 54514
rect 13356 54460 13524 54462
rect 13020 54450 13076 54460
rect 13468 54450 13524 54460
rect 12348 54404 12404 54414
rect 12236 54402 12404 54404
rect 12236 54350 12350 54402
rect 12402 54350 12404 54402
rect 12236 54348 12404 54350
rect 12236 53732 12292 53742
rect 12236 53638 12292 53676
rect 12348 53508 12404 54348
rect 13244 54290 13300 54302
rect 13244 54238 13246 54290
rect 13298 54238 13300 54290
rect 12908 53844 12964 53854
rect 13244 53844 13300 54238
rect 12908 53842 13300 53844
rect 12908 53790 12910 53842
rect 12962 53790 13300 53842
rect 12908 53788 13300 53790
rect 13468 54180 13524 54190
rect 13468 53842 13524 54124
rect 13580 54068 13636 56812
rect 13692 55970 13748 55982
rect 13692 55918 13694 55970
rect 13746 55918 13748 55970
rect 13692 55748 13748 55918
rect 13692 55682 13748 55692
rect 13804 55412 13860 57372
rect 14252 57428 14308 57596
rect 14364 57652 14420 57662
rect 14364 57558 14420 57596
rect 14252 57362 14308 57372
rect 14252 56868 14308 56878
rect 14252 56774 14308 56812
rect 14364 56756 14420 56766
rect 14364 56662 14420 56700
rect 15036 56642 15092 57820
rect 15372 57652 15428 57662
rect 15372 57650 15652 57652
rect 15372 57598 15374 57650
rect 15426 57598 15652 57650
rect 15372 57596 15652 57598
rect 15372 57586 15428 57596
rect 15260 57538 15316 57550
rect 15260 57486 15262 57538
rect 15314 57486 15316 57538
rect 15260 56754 15316 57486
rect 15372 57092 15428 57102
rect 15372 56866 15428 57036
rect 15372 56814 15374 56866
rect 15426 56814 15428 56866
rect 15372 56802 15428 56814
rect 15260 56702 15262 56754
rect 15314 56702 15316 56754
rect 15260 56690 15316 56702
rect 15036 56590 15038 56642
rect 15090 56590 15092 56642
rect 15036 56578 15092 56590
rect 14008 56476 15208 56486
rect 14064 56474 14112 56476
rect 14168 56474 14216 56476
rect 14076 56422 14112 56474
rect 14200 56422 14216 56474
rect 14064 56420 14112 56422
rect 14168 56420 14216 56422
rect 14272 56474 14320 56476
rect 14376 56474 14424 56476
rect 14480 56474 14528 56476
rect 14376 56422 14396 56474
rect 14480 56422 14520 56474
rect 14272 56420 14320 56422
rect 14376 56420 14424 56422
rect 14480 56420 14528 56422
rect 14584 56420 14632 56476
rect 14688 56474 14736 56476
rect 14792 56474 14840 56476
rect 14896 56474 14944 56476
rect 14696 56422 14736 56474
rect 14820 56422 14840 56474
rect 14688 56420 14736 56422
rect 14792 56420 14840 56422
rect 14896 56420 14944 56422
rect 15000 56474 15048 56476
rect 15104 56474 15152 56476
rect 15000 56422 15016 56474
rect 15104 56422 15140 56474
rect 15000 56420 15048 56422
rect 15104 56420 15152 56422
rect 14008 56410 15208 56420
rect 14028 56308 14084 56318
rect 13692 55356 13860 55412
rect 13916 56196 13972 56206
rect 13692 54740 13748 55356
rect 13916 55298 13972 56140
rect 14028 55410 14084 56252
rect 15036 56196 15092 56206
rect 15036 56082 15092 56140
rect 15036 56030 15038 56082
rect 15090 56030 15092 56082
rect 15036 56018 15092 56030
rect 14252 55972 14308 55982
rect 14252 55878 14308 55916
rect 14588 55972 14644 55982
rect 14588 55878 14644 55916
rect 15484 55970 15540 55982
rect 15484 55918 15486 55970
rect 15538 55918 15540 55970
rect 14588 55748 14644 55758
rect 14588 55522 14644 55692
rect 15484 55748 15540 55918
rect 15484 55682 15540 55692
rect 14588 55470 14590 55522
rect 14642 55470 14644 55522
rect 14588 55458 14644 55470
rect 14028 55358 14030 55410
rect 14082 55358 14084 55410
rect 14028 55346 14084 55358
rect 14252 55412 14308 55422
rect 13916 55246 13918 55298
rect 13970 55246 13972 55298
rect 13916 55234 13972 55246
rect 14252 55298 14308 55356
rect 14252 55246 14254 55298
rect 14306 55246 14308 55298
rect 14252 55234 14308 55246
rect 14028 55188 14084 55198
rect 14084 55132 14196 55188
rect 14028 55122 14084 55132
rect 14140 55074 14196 55132
rect 14140 55022 14142 55074
rect 14194 55022 14196 55074
rect 14140 55010 14196 55022
rect 15036 55076 15092 55114
rect 15484 55076 15540 55086
rect 15036 55010 15092 55020
rect 15372 55020 15484 55076
rect 14008 54908 15208 54918
rect 14064 54906 14112 54908
rect 14168 54906 14216 54908
rect 14076 54854 14112 54906
rect 14200 54854 14216 54906
rect 14064 54852 14112 54854
rect 14168 54852 14216 54854
rect 14272 54906 14320 54908
rect 14376 54906 14424 54908
rect 14480 54906 14528 54908
rect 14376 54854 14396 54906
rect 14480 54854 14520 54906
rect 14272 54852 14320 54854
rect 14376 54852 14424 54854
rect 14480 54852 14528 54854
rect 14584 54852 14632 54908
rect 14688 54906 14736 54908
rect 14792 54906 14840 54908
rect 14896 54906 14944 54908
rect 14696 54854 14736 54906
rect 14820 54854 14840 54906
rect 14688 54852 14736 54854
rect 14792 54852 14840 54854
rect 14896 54852 14944 54854
rect 15000 54906 15048 54908
rect 15104 54906 15152 54908
rect 15000 54854 15016 54906
rect 15104 54854 15140 54906
rect 15000 54852 15048 54854
rect 15104 54852 15152 54854
rect 14008 54842 15208 54852
rect 13692 54674 13748 54684
rect 14364 54740 14420 54750
rect 13692 54292 13748 54330
rect 13692 54226 13748 54236
rect 13804 54290 13860 54302
rect 13804 54238 13806 54290
rect 13858 54238 13860 54290
rect 13580 54012 13748 54068
rect 13468 53790 13470 53842
rect 13522 53790 13524 53842
rect 12908 53778 12964 53788
rect 13468 53778 13524 53790
rect 12348 53172 12404 53452
rect 12796 53730 12852 53742
rect 12796 53678 12798 53730
rect 12850 53678 12852 53730
rect 12796 53284 12852 53678
rect 12796 53228 13188 53284
rect 12572 53172 12628 53182
rect 12348 53170 12628 53172
rect 12348 53118 12574 53170
rect 12626 53118 12628 53170
rect 12348 53116 12628 53118
rect 12572 53060 12628 53116
rect 13132 53172 13188 53228
rect 13132 53170 13412 53172
rect 13132 53118 13134 53170
rect 13186 53118 13412 53170
rect 13132 53116 13412 53118
rect 13132 53106 13188 53116
rect 12572 52994 12628 53004
rect 13356 53058 13412 53116
rect 13356 53006 13358 53058
rect 13410 53006 13412 53058
rect 13356 52994 13412 53006
rect 13580 53060 13636 53070
rect 13468 52722 13524 52734
rect 13468 52670 13470 52722
rect 13522 52670 13524 52722
rect 13468 52500 13524 52670
rect 13468 52434 13524 52444
rect 12124 52164 12180 52174
rect 12124 52070 12180 52108
rect 12572 52164 12628 52174
rect 12572 52070 12628 52108
rect 13468 52052 13524 52062
rect 13468 50148 13524 51996
rect 13244 50092 13524 50148
rect 13580 51938 13636 53004
rect 13580 51886 13582 51938
rect 13634 51886 13636 51938
rect 13580 50372 13636 51886
rect 12908 49252 12964 49262
rect 12236 49028 12292 49038
rect 12572 49028 12628 49038
rect 12236 49026 12628 49028
rect 12236 48974 12238 49026
rect 12290 48974 12574 49026
rect 12626 48974 12628 49026
rect 12236 48972 12628 48974
rect 12236 48962 12292 48972
rect 12572 48962 12628 48972
rect 12908 49026 12964 49196
rect 12908 48974 12910 49026
rect 12962 48974 12964 49026
rect 12796 48916 12852 48926
rect 12796 48822 12852 48860
rect 12124 48242 12180 48254
rect 12124 48190 12126 48242
rect 12178 48190 12180 48242
rect 12124 47572 12180 48190
rect 12124 47506 12180 47516
rect 12348 47234 12404 47246
rect 12348 47182 12350 47234
rect 12402 47182 12404 47234
rect 12348 47068 12404 47182
rect 12908 47068 12964 48974
rect 13244 47908 13300 50092
rect 13468 49924 13524 49934
rect 13580 49924 13636 50316
rect 13468 49922 13636 49924
rect 13468 49870 13470 49922
rect 13522 49870 13636 49922
rect 13468 49868 13636 49870
rect 13468 49700 13524 49868
rect 13468 49028 13524 49644
rect 13356 48972 13524 49028
rect 13692 49028 13748 54012
rect 13804 53956 13860 54238
rect 13804 53890 13860 53900
rect 13916 54068 13972 54078
rect 13916 53732 13972 54012
rect 14364 53842 14420 54684
rect 15036 54516 15092 54526
rect 15036 54180 15092 54460
rect 15036 54114 15092 54124
rect 15260 54402 15316 54414
rect 15260 54350 15262 54402
rect 15314 54350 15316 54402
rect 14476 53956 14532 53966
rect 14812 53956 14868 53966
rect 14532 53954 14868 53956
rect 14532 53902 14814 53954
rect 14866 53902 14868 53954
rect 14532 53900 14868 53902
rect 14476 53890 14532 53900
rect 14812 53890 14868 53900
rect 15036 53956 15092 53966
rect 14364 53790 14366 53842
rect 14418 53790 14420 53842
rect 14364 53778 14420 53790
rect 15036 53842 15092 53900
rect 15036 53790 15038 53842
rect 15090 53790 15092 53842
rect 15036 53778 15092 53790
rect 13804 53730 13972 53732
rect 13804 53678 13918 53730
rect 13970 53678 13972 53730
rect 13804 53676 13972 53678
rect 13804 53172 13860 53676
rect 13916 53666 13972 53676
rect 15036 53620 15092 53630
rect 15036 53526 15092 53564
rect 15260 53508 15316 54350
rect 15372 54404 15428 55020
rect 15484 54982 15540 55020
rect 15372 54338 15428 54348
rect 15596 54402 15652 57596
rect 15596 54350 15598 54402
rect 15650 54350 15652 54402
rect 15596 54338 15652 54350
rect 15708 54180 15764 57932
rect 16044 57876 16100 59166
rect 16156 58324 16212 58334
rect 16156 58230 16212 58268
rect 16044 57810 16100 57820
rect 15820 57650 15876 57662
rect 15820 57598 15822 57650
rect 15874 57598 15876 57650
rect 15820 57092 15876 57598
rect 15820 57026 15876 57036
rect 15932 55970 15988 55982
rect 15932 55918 15934 55970
rect 15986 55918 15988 55970
rect 15932 55188 15988 55918
rect 15932 55122 15988 55132
rect 16044 55410 16100 55422
rect 16044 55358 16046 55410
rect 16098 55358 16100 55410
rect 16044 55076 16100 55358
rect 16044 55010 16100 55020
rect 15484 54124 15764 54180
rect 15372 53956 15428 53966
rect 15484 53956 15540 54124
rect 15372 53954 15540 53956
rect 15372 53902 15374 53954
rect 15426 53902 15540 53954
rect 15372 53900 15540 53902
rect 15372 53890 15428 53900
rect 15596 53842 15652 53854
rect 15596 53790 15598 53842
rect 15650 53790 15652 53842
rect 15260 53452 15540 53508
rect 14008 53340 15208 53350
rect 14064 53338 14112 53340
rect 14168 53338 14216 53340
rect 14076 53286 14112 53338
rect 14200 53286 14216 53338
rect 14064 53284 14112 53286
rect 14168 53284 14216 53286
rect 14272 53338 14320 53340
rect 14376 53338 14424 53340
rect 14480 53338 14528 53340
rect 14376 53286 14396 53338
rect 14480 53286 14520 53338
rect 14272 53284 14320 53286
rect 14376 53284 14424 53286
rect 14480 53284 14528 53286
rect 14584 53284 14632 53340
rect 14688 53338 14736 53340
rect 14792 53338 14840 53340
rect 14896 53338 14944 53340
rect 14696 53286 14736 53338
rect 14820 53286 14840 53338
rect 14688 53284 14736 53286
rect 14792 53284 14840 53286
rect 14896 53284 14944 53286
rect 15000 53338 15048 53340
rect 15104 53338 15152 53340
rect 15000 53286 15016 53338
rect 15104 53286 15140 53338
rect 15000 53284 15048 53286
rect 15104 53284 15152 53286
rect 14008 53274 15208 53284
rect 13804 53116 14084 53172
rect 13916 52948 13972 52958
rect 13804 52892 13916 52948
rect 13804 50036 13860 52892
rect 13916 52854 13972 52892
rect 14028 52052 14084 53116
rect 14140 52948 14196 52958
rect 14140 52724 14196 52892
rect 14140 52658 14196 52668
rect 14700 52834 14756 52846
rect 14700 52782 14702 52834
rect 14754 52782 14756 52834
rect 14028 51986 14084 51996
rect 14364 52052 14420 52062
rect 14700 52052 14756 52782
rect 14420 51996 14756 52052
rect 15372 52052 15428 52062
rect 14364 51986 14420 51996
rect 14008 51772 15208 51782
rect 14064 51770 14112 51772
rect 14168 51770 14216 51772
rect 14076 51718 14112 51770
rect 14200 51718 14216 51770
rect 14064 51716 14112 51718
rect 14168 51716 14216 51718
rect 14272 51770 14320 51772
rect 14376 51770 14424 51772
rect 14480 51770 14528 51772
rect 14376 51718 14396 51770
rect 14480 51718 14520 51770
rect 14272 51716 14320 51718
rect 14376 51716 14424 51718
rect 14480 51716 14528 51718
rect 14584 51716 14632 51772
rect 14688 51770 14736 51772
rect 14792 51770 14840 51772
rect 14896 51770 14944 51772
rect 14696 51718 14736 51770
rect 14820 51718 14840 51770
rect 14688 51716 14736 51718
rect 14792 51716 14840 51718
rect 14896 51716 14944 51718
rect 15000 51770 15048 51772
rect 15104 51770 15152 51772
rect 15000 51718 15016 51770
rect 15104 51718 15140 51770
rect 15000 51716 15048 51718
rect 15104 51716 15152 51718
rect 14008 51706 15208 51716
rect 14252 51604 14308 51614
rect 14252 51510 14308 51548
rect 14812 51492 14868 51502
rect 14812 51490 15204 51492
rect 14812 51438 14814 51490
rect 14866 51438 15204 51490
rect 14812 51436 15204 51438
rect 14812 51426 14868 51436
rect 14364 51266 14420 51278
rect 14364 51214 14366 51266
rect 14418 51214 14420 51266
rect 13916 50372 13972 50382
rect 13916 50278 13972 50316
rect 14364 50372 14420 51214
rect 15148 51044 15204 51436
rect 15372 51378 15428 51996
rect 15372 51326 15374 51378
rect 15426 51326 15428 51378
rect 15372 51314 15428 51326
rect 15484 51940 15540 53452
rect 15484 51156 15540 51884
rect 15596 51490 15652 53790
rect 16268 52052 16324 60284
rect 16380 58324 16436 58334
rect 16380 57650 16436 58268
rect 16380 57598 16382 57650
rect 16434 57598 16436 57650
rect 16380 56866 16436 57598
rect 16380 56814 16382 56866
rect 16434 56814 16436 56866
rect 16380 56802 16436 56814
rect 16380 56420 16436 56430
rect 16380 56082 16436 56364
rect 16380 56030 16382 56082
rect 16434 56030 16436 56082
rect 16380 56018 16436 56030
rect 16380 55300 16436 55310
rect 16380 55206 16436 55244
rect 16268 51986 16324 51996
rect 16268 51492 16324 51502
rect 15596 51438 15598 51490
rect 15650 51438 15652 51490
rect 15596 51426 15652 51438
rect 16044 51490 16324 51492
rect 16044 51438 16270 51490
rect 16322 51438 16324 51490
rect 16044 51436 16324 51438
rect 15484 51090 15540 51100
rect 15708 51378 15764 51390
rect 15708 51326 15710 51378
rect 15762 51326 15764 51378
rect 15148 50988 15316 51044
rect 15148 50820 15204 50830
rect 14812 50594 14868 50606
rect 14812 50542 14814 50594
rect 14866 50542 14868 50594
rect 14812 50484 14868 50542
rect 15148 50594 15204 50764
rect 15260 50706 15316 50988
rect 15708 50932 15764 51326
rect 15260 50654 15262 50706
rect 15314 50654 15316 50706
rect 15260 50642 15316 50654
rect 15372 50876 15764 50932
rect 15148 50542 15150 50594
rect 15202 50542 15204 50594
rect 15148 50530 15204 50542
rect 14812 50418 14868 50428
rect 14364 50306 14420 50316
rect 14008 50204 15208 50214
rect 14064 50202 14112 50204
rect 14168 50202 14216 50204
rect 14076 50150 14112 50202
rect 14200 50150 14216 50202
rect 14064 50148 14112 50150
rect 14168 50148 14216 50150
rect 14272 50202 14320 50204
rect 14376 50202 14424 50204
rect 14480 50202 14528 50204
rect 14376 50150 14396 50202
rect 14480 50150 14520 50202
rect 14272 50148 14320 50150
rect 14376 50148 14424 50150
rect 14480 50148 14528 50150
rect 14584 50148 14632 50204
rect 14688 50202 14736 50204
rect 14792 50202 14840 50204
rect 14896 50202 14944 50204
rect 14696 50150 14736 50202
rect 14820 50150 14840 50202
rect 14688 50148 14736 50150
rect 14792 50148 14840 50150
rect 14896 50148 14944 50150
rect 15000 50202 15048 50204
rect 15104 50202 15152 50204
rect 15000 50150 15016 50202
rect 15104 50150 15140 50202
rect 15000 50148 15048 50150
rect 15104 50148 15152 50150
rect 14008 50138 15208 50148
rect 14588 50036 14644 50046
rect 15372 50036 15428 50876
rect 13804 50034 14644 50036
rect 13804 49982 14590 50034
rect 14642 49982 14644 50034
rect 13804 49980 14644 49982
rect 14588 49970 14644 49980
rect 15036 49980 15428 50036
rect 15484 50596 15540 50606
rect 15932 50596 15988 50606
rect 15540 50594 15988 50596
rect 15540 50542 15934 50594
rect 15986 50542 15988 50594
rect 15540 50540 15988 50542
rect 14252 49700 14308 49710
rect 14252 49586 14308 49644
rect 14252 49534 14254 49586
rect 14306 49534 14308 49586
rect 13916 49028 13972 49038
rect 13692 48972 13860 49028
rect 13356 48132 13412 48972
rect 13580 48916 13636 48926
rect 13356 48066 13412 48076
rect 13468 48914 13636 48916
rect 13468 48862 13582 48914
rect 13634 48862 13636 48914
rect 13468 48860 13636 48862
rect 13244 47852 13412 47908
rect 12012 47012 12292 47068
rect 11788 46676 11844 46686
rect 11844 46620 11956 46676
rect 11788 46582 11844 46620
rect 11788 45892 11844 45902
rect 11788 45444 11844 45836
rect 11788 45378 11844 45388
rect 11788 45220 11844 45230
rect 11788 45126 11844 45164
rect 11676 44370 11732 44380
rect 11676 44098 11732 44110
rect 11676 44046 11678 44098
rect 11730 44046 11732 44098
rect 11676 43428 11732 44046
rect 11788 43428 11844 43438
rect 11676 43426 11844 43428
rect 11676 43374 11790 43426
rect 11842 43374 11844 43426
rect 11676 43372 11844 43374
rect 11788 43362 11844 43372
rect 11676 42980 11732 42990
rect 11676 42754 11732 42924
rect 11676 42702 11678 42754
rect 11730 42702 11732 42754
rect 11676 42690 11732 42702
rect 11340 41358 11342 41410
rect 11394 41358 11396 41410
rect 11340 41346 11396 41358
rect 11452 42476 11620 42532
rect 11452 41188 11508 42476
rect 11900 42420 11956 46620
rect 12236 44436 12292 47012
rect 12348 47012 12964 47068
rect 13244 47012 13300 47022
rect 12348 46004 12404 47012
rect 13132 46562 13188 46574
rect 13132 46510 13134 46562
rect 13186 46510 13188 46562
rect 12348 46002 12740 46004
rect 12348 45950 12350 46002
rect 12402 45950 12740 46002
rect 12348 45948 12740 45950
rect 12348 45938 12404 45948
rect 12684 45332 12740 45948
rect 13132 45892 13188 46510
rect 13132 45826 13188 45836
rect 13132 45332 13188 45342
rect 12684 45330 13188 45332
rect 12684 45278 12686 45330
rect 12738 45278 13134 45330
rect 13186 45278 13188 45330
rect 12684 45276 13188 45278
rect 12684 45266 12740 45276
rect 13132 45108 13188 45276
rect 13132 45042 13188 45052
rect 12908 44436 12964 44446
rect 12236 44434 12852 44436
rect 12236 44382 12238 44434
rect 12290 44382 12852 44434
rect 12236 44380 12852 44382
rect 12236 44370 12292 44380
rect 12572 44100 12628 44110
rect 12348 43650 12404 43662
rect 12348 43598 12350 43650
rect 12402 43598 12404 43650
rect 12348 43540 12404 43598
rect 12348 43474 12404 43484
rect 12572 43538 12628 44044
rect 12572 43486 12574 43538
rect 12626 43486 12628 43538
rect 12236 43316 12292 43326
rect 12012 43314 12292 43316
rect 12012 43262 12238 43314
rect 12290 43262 12292 43314
rect 12012 43260 12292 43262
rect 12012 42754 12068 43260
rect 12236 43250 12292 43260
rect 12572 42868 12628 43486
rect 12796 43650 12852 44380
rect 13244 44436 13300 46956
rect 13356 46228 13412 47852
rect 13468 47234 13524 48860
rect 13580 48850 13636 48860
rect 13692 48804 13748 48814
rect 13692 48710 13748 48748
rect 13580 48692 13636 48702
rect 13580 48244 13636 48636
rect 13580 48188 13748 48244
rect 13580 47572 13636 47582
rect 13580 47478 13636 47516
rect 13692 47458 13748 48188
rect 13692 47406 13694 47458
rect 13746 47406 13748 47458
rect 13692 47394 13748 47406
rect 13468 47182 13470 47234
rect 13522 47182 13524 47234
rect 13468 46450 13524 47182
rect 13580 47348 13636 47358
rect 13580 46564 13636 47292
rect 13804 46900 13860 48972
rect 13916 48934 13972 48972
rect 14252 49026 14308 49534
rect 15036 49140 15092 49980
rect 15372 49812 15428 49822
rect 15484 49812 15540 50540
rect 15932 50530 15988 50540
rect 15932 50428 15988 50438
rect 15372 49810 15540 49812
rect 15372 49758 15374 49810
rect 15426 49758 15540 49810
rect 15372 49756 15540 49758
rect 15708 50372 15764 50382
rect 15372 49746 15428 49756
rect 15708 49700 15764 50316
rect 15932 50036 15988 50372
rect 15708 49606 15764 49644
rect 15820 49980 15988 50036
rect 15820 49252 15876 49980
rect 15932 49810 15988 49822
rect 15932 49758 15934 49810
rect 15986 49758 15988 49810
rect 15932 49700 15988 49758
rect 15932 49634 15988 49644
rect 15708 49196 15876 49252
rect 15148 49140 15204 49150
rect 15036 49138 15204 49140
rect 15036 49086 15150 49138
rect 15202 49086 15204 49138
rect 15036 49084 15204 49086
rect 15148 49074 15204 49084
rect 14252 48974 14254 49026
rect 14306 48974 14308 49026
rect 14252 48916 14308 48974
rect 14252 48850 14308 48860
rect 14700 49026 14756 49038
rect 14700 48974 14702 49026
rect 14754 48974 14756 49026
rect 14700 48916 14756 48974
rect 14700 48850 14756 48860
rect 15372 49028 15428 49038
rect 15372 48804 15428 48972
rect 15596 49026 15652 49038
rect 15596 48974 15598 49026
rect 15650 48974 15652 49026
rect 15596 48804 15652 48974
rect 14008 48636 15208 48646
rect 14064 48634 14112 48636
rect 14168 48634 14216 48636
rect 14076 48582 14112 48634
rect 14200 48582 14216 48634
rect 14064 48580 14112 48582
rect 14168 48580 14216 48582
rect 14272 48634 14320 48636
rect 14376 48634 14424 48636
rect 14480 48634 14528 48636
rect 14376 48582 14396 48634
rect 14480 48582 14520 48634
rect 14272 48580 14320 48582
rect 14376 48580 14424 48582
rect 14480 48580 14528 48582
rect 14584 48580 14632 48636
rect 14688 48634 14736 48636
rect 14792 48634 14840 48636
rect 14896 48634 14944 48636
rect 14696 48582 14736 48634
rect 14820 48582 14840 48634
rect 14688 48580 14736 48582
rect 14792 48580 14840 48582
rect 14896 48580 14944 48582
rect 15000 48634 15048 48636
rect 15104 48634 15152 48636
rect 15000 48582 15016 48634
rect 15104 48582 15140 48634
rect 15000 48580 15048 48582
rect 15104 48580 15152 48582
rect 14008 48570 15208 48580
rect 14588 48466 14644 48478
rect 14588 48414 14590 48466
rect 14642 48414 14644 48466
rect 14588 48132 14644 48414
rect 15148 48468 15204 48478
rect 15372 48468 15428 48748
rect 15148 48466 15428 48468
rect 15148 48414 15150 48466
rect 15202 48414 15428 48466
rect 15148 48412 15428 48414
rect 15484 48748 15596 48804
rect 15484 48466 15540 48748
rect 15596 48738 15652 48748
rect 15484 48414 15486 48466
rect 15538 48414 15540 48466
rect 15148 48402 15204 48412
rect 15484 48402 15540 48414
rect 14588 48066 14644 48076
rect 15372 48132 15428 48142
rect 13916 47460 13972 47470
rect 13916 47346 13972 47404
rect 13916 47294 13918 47346
rect 13970 47294 13972 47346
rect 13916 47282 13972 47294
rect 14700 47458 14756 47470
rect 14700 47406 14702 47458
rect 14754 47406 14756 47458
rect 14700 47236 14756 47406
rect 14700 47170 14756 47180
rect 15372 47236 15428 48076
rect 15596 47236 15652 47246
rect 15372 47234 15652 47236
rect 15372 47182 15598 47234
rect 15650 47182 15652 47234
rect 15372 47180 15652 47182
rect 14008 47068 15208 47078
rect 14064 47066 14112 47068
rect 14168 47066 14216 47068
rect 14076 47014 14112 47066
rect 14200 47014 14216 47066
rect 14064 47012 14112 47014
rect 14168 47012 14216 47014
rect 14272 47066 14320 47068
rect 14376 47066 14424 47068
rect 14480 47066 14528 47068
rect 14376 47014 14396 47066
rect 14480 47014 14520 47066
rect 14272 47012 14320 47014
rect 14376 47012 14424 47014
rect 14480 47012 14528 47014
rect 14584 47012 14632 47068
rect 14688 47066 14736 47068
rect 14792 47066 14840 47068
rect 14896 47066 14944 47068
rect 14696 47014 14736 47066
rect 14820 47014 14840 47066
rect 14688 47012 14736 47014
rect 14792 47012 14840 47014
rect 14896 47012 14944 47014
rect 15000 47066 15048 47068
rect 15104 47066 15152 47068
rect 15000 47014 15016 47066
rect 15104 47014 15140 47066
rect 15000 47012 15048 47014
rect 15104 47012 15152 47014
rect 14008 47002 15208 47012
rect 13916 46900 13972 46910
rect 13804 46844 13916 46900
rect 13916 46834 13972 46844
rect 15372 46898 15428 47180
rect 15596 47170 15652 47180
rect 15372 46846 15374 46898
rect 15426 46846 15428 46898
rect 15372 46834 15428 46846
rect 13580 46562 13748 46564
rect 13580 46510 13582 46562
rect 13634 46510 13748 46562
rect 13580 46508 13748 46510
rect 13580 46498 13636 46508
rect 13468 46398 13470 46450
rect 13522 46398 13524 46450
rect 13468 46340 13524 46398
rect 13468 46284 13636 46340
rect 13356 46172 13524 46228
rect 13468 44660 13524 46172
rect 13580 45666 13636 46284
rect 13580 45614 13582 45666
rect 13634 45614 13636 45666
rect 13580 44884 13636 45614
rect 13692 45778 13748 46508
rect 14028 46562 14084 46574
rect 14028 46510 14030 46562
rect 14082 46510 14084 46562
rect 14028 46450 14084 46510
rect 14028 46398 14030 46450
rect 14082 46398 14084 46450
rect 14028 46386 14084 46398
rect 14476 46562 14532 46574
rect 14476 46510 14478 46562
rect 14530 46510 14532 46562
rect 14476 46450 14532 46510
rect 14476 46398 14478 46450
rect 14530 46398 14532 46450
rect 14476 46386 14532 46398
rect 13804 45892 13860 45902
rect 13804 45798 13860 45836
rect 13692 45726 13694 45778
rect 13746 45726 13748 45778
rect 13692 45556 13748 45726
rect 15372 45666 15428 45678
rect 15372 45614 15374 45666
rect 15426 45614 15428 45666
rect 13692 45500 13860 45556
rect 13692 45332 13748 45342
rect 13804 45332 13860 45500
rect 14008 45500 15208 45510
rect 14064 45498 14112 45500
rect 14168 45498 14216 45500
rect 14076 45446 14112 45498
rect 14200 45446 14216 45498
rect 14064 45444 14112 45446
rect 14168 45444 14216 45446
rect 14272 45498 14320 45500
rect 14376 45498 14424 45500
rect 14480 45498 14528 45500
rect 14376 45446 14396 45498
rect 14480 45446 14520 45498
rect 14272 45444 14320 45446
rect 14376 45444 14424 45446
rect 14480 45444 14528 45446
rect 14584 45444 14632 45500
rect 14688 45498 14736 45500
rect 14792 45498 14840 45500
rect 14896 45498 14944 45500
rect 14696 45446 14736 45498
rect 14820 45446 14840 45498
rect 14688 45444 14736 45446
rect 14792 45444 14840 45446
rect 14896 45444 14944 45446
rect 15000 45498 15048 45500
rect 15104 45498 15152 45500
rect 15000 45446 15016 45498
rect 15104 45446 15140 45498
rect 15000 45444 15048 45446
rect 15104 45444 15152 45446
rect 14008 45434 15208 45444
rect 14140 45332 14196 45342
rect 13804 45276 13972 45332
rect 13692 45238 13748 45276
rect 13804 45108 13860 45118
rect 13692 44884 13748 44894
rect 13580 44828 13692 44884
rect 13692 44818 13748 44828
rect 13804 44772 13860 45052
rect 13804 44706 13860 44716
rect 13468 44604 13636 44660
rect 13468 44436 13524 44446
rect 13244 44380 13412 44436
rect 12908 44342 12964 44380
rect 13356 44100 13412 44380
rect 13468 44322 13524 44380
rect 13468 44270 13470 44322
rect 13522 44270 13524 44322
rect 13468 44258 13524 44270
rect 13356 44044 13524 44100
rect 12796 43598 12798 43650
rect 12850 43598 12852 43650
rect 12796 43428 12852 43598
rect 13356 43428 13412 43438
rect 12684 42868 12740 42878
rect 12572 42866 12740 42868
rect 12572 42814 12686 42866
rect 12738 42814 12740 42866
rect 12572 42812 12740 42814
rect 12684 42802 12740 42812
rect 12012 42702 12014 42754
rect 12066 42702 12068 42754
rect 12012 42690 12068 42702
rect 12124 42644 12180 42654
rect 12796 42644 12852 43372
rect 12124 42642 12628 42644
rect 12124 42590 12126 42642
rect 12178 42590 12628 42642
rect 12124 42588 12628 42590
rect 12124 42578 12180 42588
rect 11900 42364 12292 42420
rect 11564 41972 11620 41982
rect 11564 41878 11620 41916
rect 11340 41132 11508 41188
rect 11900 41410 11956 41422
rect 11900 41358 11902 41410
rect 11954 41358 11956 41410
rect 11340 40740 11396 41132
rect 11788 41074 11844 41086
rect 11788 41022 11790 41074
rect 11842 41022 11844 41074
rect 11452 40964 11508 40974
rect 11452 40962 11732 40964
rect 11452 40910 11454 40962
rect 11506 40910 11732 40962
rect 11452 40908 11732 40910
rect 11452 40898 11508 40908
rect 11340 40684 11508 40740
rect 11228 40402 11396 40404
rect 11228 40350 11230 40402
rect 11282 40350 11396 40402
rect 11228 40348 11396 40350
rect 11228 40338 11284 40348
rect 10780 39732 10836 39742
rect 10780 39638 10836 39676
rect 11228 39732 11284 39742
rect 11228 39060 11284 39676
rect 11228 38994 11284 39004
rect 11340 38836 11396 40348
rect 11340 38742 11396 38780
rect 10668 38612 11284 38668
rect 9996 38052 10052 38612
rect 9772 37774 9774 37826
rect 9826 37774 9828 37826
rect 8988 37212 9156 37268
rect 8988 36484 9044 36494
rect 8988 36390 9044 36428
rect 8764 36092 8932 36148
rect 8652 35812 8708 35822
rect 8652 35718 8708 35756
rect 8764 35810 8820 36092
rect 8764 35758 8766 35810
rect 8818 35758 8820 35810
rect 8652 35588 8708 35598
rect 8652 35494 8708 35532
rect 8764 35364 8820 35758
rect 9100 35924 9156 37212
rect 9548 36372 9604 36382
rect 9548 36278 9604 36316
rect 9772 36258 9828 37774
rect 9772 36206 9774 36258
rect 9826 36206 9828 36258
rect 9772 36194 9828 36206
rect 9884 37996 10052 38052
rect 9884 37380 9940 37996
rect 9996 37828 10052 37838
rect 9996 37826 10276 37828
rect 9996 37774 9998 37826
rect 10050 37774 10276 37826
rect 9996 37772 10276 37774
rect 9996 37762 10052 37772
rect 9996 37380 10052 37390
rect 9884 37378 10052 37380
rect 9884 37326 9998 37378
rect 10050 37326 10052 37378
rect 9884 37324 10052 37326
rect 8764 35298 8820 35308
rect 8988 35698 9044 35710
rect 8988 35646 8990 35698
rect 9042 35646 9044 35698
rect 8988 34804 9044 35646
rect 9100 35308 9156 35868
rect 9660 35812 9716 35822
rect 9660 35718 9716 35756
rect 9772 35810 9828 35822
rect 9772 35758 9774 35810
rect 9826 35758 9828 35810
rect 9548 35698 9604 35710
rect 9548 35646 9550 35698
rect 9602 35646 9604 35698
rect 9548 35476 9604 35646
rect 9548 35410 9604 35420
rect 9100 35252 9492 35308
rect 8652 34132 8708 34142
rect 8988 34132 9044 34748
rect 8652 34130 9044 34132
rect 8652 34078 8654 34130
rect 8706 34078 9044 34130
rect 8652 34076 9044 34078
rect 9436 34692 9492 35196
rect 9772 34916 9828 35758
rect 9884 35810 9940 37324
rect 9996 37314 10052 37324
rect 10220 37266 10276 37772
rect 10220 37214 10222 37266
rect 10274 37214 10276 37266
rect 10220 37202 10276 37214
rect 10444 37156 10500 37166
rect 10332 36484 10388 36494
rect 10108 36372 10164 36382
rect 9884 35758 9886 35810
rect 9938 35758 9940 35810
rect 9884 35140 9940 35758
rect 9996 36370 10164 36372
rect 9996 36318 10110 36370
rect 10162 36318 10164 36370
rect 9996 36316 10164 36318
rect 9996 35810 10052 36316
rect 10108 36306 10164 36316
rect 9996 35758 9998 35810
rect 10050 35758 10052 35810
rect 9996 35364 10052 35758
rect 10332 35476 10388 36428
rect 10332 35410 10388 35420
rect 10052 35308 10276 35364
rect 9996 35298 10052 35308
rect 10220 35140 10276 35308
rect 10332 35140 10388 35150
rect 9940 35084 10052 35140
rect 10220 35138 10388 35140
rect 10220 35086 10334 35138
rect 10386 35086 10388 35138
rect 10220 35084 10388 35086
rect 9884 35074 9940 35084
rect 9548 34692 9604 34702
rect 9436 34690 9604 34692
rect 9436 34638 9550 34690
rect 9602 34638 9604 34690
rect 9436 34636 9604 34638
rect 8652 34066 8708 34076
rect 8316 33282 8372 33292
rect 8428 33852 8596 33908
rect 8652 33908 8708 33918
rect 8316 33124 8372 33134
rect 8316 33030 8372 33068
rect 8092 32844 8372 32900
rect 7980 32732 8260 32788
rect 7980 32564 8036 32574
rect 7980 31892 8036 32508
rect 7980 31826 8036 31836
rect 7980 31556 8036 31566
rect 7644 31554 8036 31556
rect 7644 31502 7982 31554
rect 8034 31502 8036 31554
rect 7644 31500 8036 31502
rect 7364 30156 7476 30212
rect 7532 30324 7588 30334
rect 7644 30324 7700 30334
rect 7588 30322 7700 30324
rect 7588 30270 7646 30322
rect 7698 30270 7700 30322
rect 7588 30268 7700 30270
rect 7308 30118 7364 30156
rect 7084 29652 7140 29662
rect 7084 29426 7140 29596
rect 7084 29374 7086 29426
rect 7138 29374 7140 29426
rect 7084 29362 7140 29374
rect 7420 29316 7476 29326
rect 7308 29260 7420 29316
rect 6972 28590 6974 28642
rect 7026 28590 7028 28642
rect 6748 27906 6804 27916
rect 6748 27636 6804 27646
rect 6636 26852 6692 26862
rect 6636 26290 6692 26796
rect 6748 26402 6804 27580
rect 6972 27300 7028 28590
rect 6972 27234 7028 27244
rect 7084 28644 7140 28654
rect 7084 27298 7140 28588
rect 7084 27246 7086 27298
rect 7138 27246 7140 27298
rect 6748 26350 6750 26402
rect 6802 26350 6804 26402
rect 6748 26338 6804 26350
rect 6860 27074 6916 27086
rect 6860 27022 6862 27074
rect 6914 27022 6916 27074
rect 6636 26238 6638 26290
rect 6690 26238 6692 26290
rect 6636 26226 6692 26238
rect 6300 26014 6302 26066
rect 6354 26014 6356 26066
rect 6076 25676 6244 25732
rect 6076 25508 6132 25518
rect 6076 25414 6132 25452
rect 6188 25284 6244 25676
rect 6300 25508 6356 26014
rect 6300 25442 6356 25452
rect 6412 26012 6580 26068
rect 6188 25228 6356 25284
rect 6188 23826 6244 23838
rect 6188 23774 6190 23826
rect 6242 23774 6244 23826
rect 6188 23492 6244 23774
rect 6188 23426 6244 23436
rect 5964 23156 6020 23166
rect 5852 23154 6020 23156
rect 5852 23102 5966 23154
rect 6018 23102 6020 23154
rect 5852 23100 6020 23102
rect 5964 23090 6020 23100
rect 5404 22764 5572 22820
rect 5404 22148 5460 22158
rect 5292 22092 5404 22148
rect 5404 22082 5460 22092
rect 4956 21308 5348 21364
rect 4008 21196 5208 21206
rect 4064 21194 4112 21196
rect 4168 21194 4216 21196
rect 4076 21142 4112 21194
rect 4200 21142 4216 21194
rect 4064 21140 4112 21142
rect 4168 21140 4216 21142
rect 4272 21194 4320 21196
rect 4376 21194 4424 21196
rect 4480 21194 4528 21196
rect 4376 21142 4396 21194
rect 4480 21142 4520 21194
rect 4272 21140 4320 21142
rect 4376 21140 4424 21142
rect 4480 21140 4528 21142
rect 4584 21140 4632 21196
rect 4688 21194 4736 21196
rect 4792 21194 4840 21196
rect 4896 21194 4944 21196
rect 4696 21142 4736 21194
rect 4820 21142 4840 21194
rect 4688 21140 4736 21142
rect 4792 21140 4840 21142
rect 4896 21140 4944 21142
rect 5000 21194 5048 21196
rect 5104 21194 5152 21196
rect 5000 21142 5016 21194
rect 5104 21142 5140 21194
rect 5000 21140 5048 21142
rect 5104 21140 5152 21142
rect 4008 21130 5208 21140
rect 4508 21028 4564 21038
rect 4508 20934 4564 20972
rect 4620 20804 4676 20814
rect 4620 20710 4676 20748
rect 5068 20580 5124 20590
rect 5292 20580 5348 21308
rect 5404 21362 5460 21374
rect 5404 21310 5406 21362
rect 5458 21310 5460 21362
rect 5404 20804 5460 21310
rect 5404 20738 5460 20748
rect 5516 20692 5572 22764
rect 5516 20626 5572 20636
rect 5628 22370 5684 22382
rect 6076 22372 6132 22382
rect 5628 22318 5630 22370
rect 5682 22318 5684 22370
rect 5628 21588 5684 22318
rect 5852 22370 6132 22372
rect 5852 22318 6078 22370
rect 6130 22318 6132 22370
rect 5852 22316 6132 22318
rect 5852 21810 5908 22316
rect 6076 22306 6132 22316
rect 5852 21758 5854 21810
rect 5906 21758 5908 21810
rect 5852 21746 5908 21758
rect 6076 22148 6132 22158
rect 5124 20524 5348 20580
rect 5068 20486 5124 20524
rect 5628 19908 5684 21532
rect 6076 21476 6132 22092
rect 6188 21700 6244 21710
rect 6188 21586 6244 21644
rect 6188 21534 6190 21586
rect 6242 21534 6244 21586
rect 6188 21522 6244 21534
rect 5852 21420 6132 21476
rect 5740 20580 5796 20590
rect 5852 20580 5908 21420
rect 6300 21364 6356 25228
rect 6412 23940 6468 26012
rect 6860 25508 6916 27022
rect 7084 27076 7140 27246
rect 7308 27300 7364 29260
rect 7420 29250 7476 29260
rect 7532 27858 7588 30268
rect 7644 30258 7700 30268
rect 7980 30324 8036 31500
rect 7868 30212 7924 30222
rect 7868 30098 7924 30156
rect 7868 30046 7870 30098
rect 7922 30046 7924 30098
rect 7756 29988 7812 29998
rect 7756 29894 7812 29932
rect 7868 28754 7924 30046
rect 7868 28702 7870 28754
rect 7922 28702 7924 28754
rect 7868 28644 7924 28702
rect 7868 28578 7924 28588
rect 7532 27806 7534 27858
rect 7586 27806 7588 27858
rect 7532 27794 7588 27806
rect 7644 27746 7700 27758
rect 7644 27694 7646 27746
rect 7698 27694 7700 27746
rect 7420 27300 7476 27310
rect 7308 27298 7476 27300
rect 7308 27246 7422 27298
rect 7474 27246 7476 27298
rect 7308 27244 7476 27246
rect 7420 27234 7476 27244
rect 7084 27010 7140 27020
rect 7308 26964 7364 26974
rect 7084 26852 7140 26862
rect 7084 26514 7140 26796
rect 7084 26462 7086 26514
rect 7138 26462 7140 26514
rect 7084 26450 7140 26462
rect 7196 26292 7252 26302
rect 7196 26198 7252 26236
rect 6748 25452 6916 25508
rect 7196 25956 7252 25966
rect 6636 24724 6692 24734
rect 6636 24050 6692 24668
rect 6636 23998 6638 24050
rect 6690 23998 6692 24050
rect 6412 23884 6580 23940
rect 6412 23604 6468 23614
rect 6412 23492 6468 23548
rect 6412 21588 6468 23436
rect 6412 21522 6468 21532
rect 5740 20578 5908 20580
rect 5740 20526 5742 20578
rect 5794 20526 5908 20578
rect 5740 20524 5908 20526
rect 5740 20514 5796 20524
rect 5740 19908 5796 19918
rect 5628 19906 5796 19908
rect 5628 19854 5742 19906
rect 5794 19854 5796 19906
rect 5628 19852 5796 19854
rect 4008 19628 5208 19638
rect 4064 19626 4112 19628
rect 4168 19626 4216 19628
rect 4076 19574 4112 19626
rect 4200 19574 4216 19626
rect 4064 19572 4112 19574
rect 4168 19572 4216 19574
rect 4272 19626 4320 19628
rect 4376 19626 4424 19628
rect 4480 19626 4528 19628
rect 4376 19574 4396 19626
rect 4480 19574 4520 19626
rect 4272 19572 4320 19574
rect 4376 19572 4424 19574
rect 4480 19572 4528 19574
rect 4584 19572 4632 19628
rect 4688 19626 4736 19628
rect 4792 19626 4840 19628
rect 4896 19626 4944 19628
rect 4696 19574 4736 19626
rect 4820 19574 4840 19626
rect 4688 19572 4736 19574
rect 4792 19572 4840 19574
rect 4896 19572 4944 19574
rect 5000 19626 5048 19628
rect 5104 19626 5152 19628
rect 5000 19574 5016 19626
rect 5104 19574 5140 19626
rect 5000 19572 5048 19574
rect 5104 19572 5152 19574
rect 4008 19562 5208 19572
rect 3836 19010 3892 19022
rect 3836 18958 3838 19010
rect 3890 18958 3892 19010
rect 3836 17780 3892 18958
rect 4008 18060 5208 18070
rect 4064 18058 4112 18060
rect 4168 18058 4216 18060
rect 4076 18006 4112 18058
rect 4200 18006 4216 18058
rect 4064 18004 4112 18006
rect 4168 18004 4216 18006
rect 4272 18058 4320 18060
rect 4376 18058 4424 18060
rect 4480 18058 4528 18060
rect 4376 18006 4396 18058
rect 4480 18006 4520 18058
rect 4272 18004 4320 18006
rect 4376 18004 4424 18006
rect 4480 18004 4528 18006
rect 4584 18004 4632 18060
rect 4688 18058 4736 18060
rect 4792 18058 4840 18060
rect 4896 18058 4944 18060
rect 4696 18006 4736 18058
rect 4820 18006 4840 18058
rect 4688 18004 4736 18006
rect 4792 18004 4840 18006
rect 4896 18004 4944 18006
rect 5000 18058 5048 18060
rect 5104 18058 5152 18060
rect 5000 18006 5016 18058
rect 5104 18006 5140 18058
rect 5000 18004 5048 18006
rect 5104 18004 5152 18006
rect 4008 17994 5208 18004
rect 4172 17892 4228 17902
rect 4172 17798 4228 17836
rect 3836 17714 3892 17724
rect 4620 17666 4676 17678
rect 4620 17614 4622 17666
rect 4674 17614 4676 17666
rect 3388 16270 3390 16322
rect 3442 16270 3444 16322
rect 3388 16258 3444 16270
rect 3500 16492 3780 16548
rect 3836 17442 3892 17454
rect 3836 17390 3838 17442
rect 3890 17390 3892 17442
rect 3500 15148 3556 16492
rect 3164 14690 3220 14700
rect 3388 15092 3556 15148
rect 1932 13458 1988 13468
rect 3164 12740 3220 12750
rect 1820 12126 1822 12178
rect 1874 12126 1876 12178
rect 1820 10610 1876 12126
rect 1820 10558 1822 10610
rect 1874 10558 1876 10610
rect 1820 7474 1876 10558
rect 2268 12738 3220 12740
rect 2268 12686 3166 12738
rect 3218 12686 3220 12738
rect 2268 12684 3220 12686
rect 2268 10610 2324 12684
rect 3164 12674 3220 12684
rect 2380 12178 2436 12190
rect 2380 12126 2382 12178
rect 2434 12126 2436 12178
rect 2380 11620 2436 12126
rect 3388 11844 3444 15092
rect 3724 14306 3780 14318
rect 3724 14254 3726 14306
rect 3778 14254 3780 14306
rect 3724 14196 3780 14254
rect 3500 14140 3780 14196
rect 3500 13186 3556 14140
rect 3500 13134 3502 13186
rect 3554 13134 3556 13186
rect 3500 13122 3556 13134
rect 3612 13972 3668 13982
rect 3388 11788 3556 11844
rect 2380 11554 2436 11564
rect 3388 11620 3444 11630
rect 3388 11526 3444 11564
rect 2268 10558 2270 10610
rect 2322 10558 2324 10610
rect 2268 10546 2324 10558
rect 3500 8036 3556 11788
rect 1820 7422 1822 7474
rect 1874 7422 1876 7474
rect 1708 4340 1764 4350
rect 1820 4340 1876 7422
rect 2156 7474 2212 7486
rect 2156 7422 2158 7474
rect 2210 7422 2212 7474
rect 2156 6020 2212 7422
rect 3500 6916 3556 7980
rect 3500 6850 3556 6860
rect 3612 6804 3668 13916
rect 3724 11620 3780 11630
rect 3836 11620 3892 17390
rect 4620 16884 4676 17614
rect 5628 17666 5684 19852
rect 5740 19842 5796 19852
rect 5628 17614 5630 17666
rect 5682 17614 5684 17666
rect 4956 17556 5012 17566
rect 4956 17462 5012 17500
rect 4620 16790 4676 16828
rect 4732 16994 4788 17006
rect 4732 16942 4734 16994
rect 4786 16942 4788 16994
rect 3948 16772 4004 16782
rect 3948 16678 4004 16716
rect 4732 16660 4788 16942
rect 5292 16884 5348 16894
rect 5404 16884 5460 16894
rect 5292 16882 5404 16884
rect 5292 16830 5294 16882
rect 5346 16830 5404 16882
rect 5292 16828 5404 16830
rect 5292 16818 5348 16828
rect 4732 16594 4788 16604
rect 4008 16492 5208 16502
rect 4064 16490 4112 16492
rect 4168 16490 4216 16492
rect 4076 16438 4112 16490
rect 4200 16438 4216 16490
rect 4064 16436 4112 16438
rect 4168 16436 4216 16438
rect 4272 16490 4320 16492
rect 4376 16490 4424 16492
rect 4480 16490 4528 16492
rect 4376 16438 4396 16490
rect 4480 16438 4520 16490
rect 4272 16436 4320 16438
rect 4376 16436 4424 16438
rect 4480 16436 4528 16438
rect 4584 16436 4632 16492
rect 4688 16490 4736 16492
rect 4792 16490 4840 16492
rect 4896 16490 4944 16492
rect 4696 16438 4736 16490
rect 4820 16438 4840 16490
rect 4688 16436 4736 16438
rect 4792 16436 4840 16438
rect 4896 16436 4944 16438
rect 5000 16490 5048 16492
rect 5104 16490 5152 16492
rect 5000 16438 5016 16490
rect 5104 16438 5140 16490
rect 5000 16436 5048 16438
rect 5104 16436 5152 16438
rect 4008 16426 5208 16436
rect 3948 16212 4004 16222
rect 3948 16098 4004 16156
rect 4732 16212 4788 16222
rect 4732 16118 4788 16156
rect 3948 16046 3950 16098
rect 4002 16046 4004 16098
rect 3948 16034 4004 16046
rect 4172 15988 4228 15998
rect 4172 15894 4228 15932
rect 5292 15988 5348 15998
rect 4732 15652 4788 15662
rect 4732 15538 4788 15596
rect 4732 15486 4734 15538
rect 4786 15486 4788 15538
rect 4732 15474 4788 15486
rect 5292 15538 5348 15932
rect 5292 15486 5294 15538
rect 5346 15486 5348 15538
rect 5292 15474 5348 15486
rect 5404 15148 5460 16828
rect 5292 15092 5460 15148
rect 5628 15204 5684 17614
rect 5740 16884 5796 16894
rect 5852 16884 5908 20524
rect 5796 16828 5908 16884
rect 5964 21308 6356 21364
rect 5740 16790 5796 16828
rect 5852 16660 5908 16670
rect 5852 16100 5908 16604
rect 5964 16324 6020 21308
rect 6076 20804 6132 20814
rect 6076 20710 6132 20748
rect 6188 20692 6244 20702
rect 6244 20636 6356 20692
rect 6188 20598 6244 20636
rect 6188 20244 6244 20254
rect 6188 20150 6244 20188
rect 6300 18564 6356 20636
rect 6412 20578 6468 20590
rect 6412 20526 6414 20578
rect 6466 20526 6468 20578
rect 6412 18788 6468 20526
rect 6412 18722 6468 18732
rect 6300 18508 6468 18564
rect 6076 17666 6132 17678
rect 6076 17614 6078 17666
rect 6130 17614 6132 17666
rect 6076 16772 6132 17614
rect 6076 16706 6132 16716
rect 6188 16884 6244 16894
rect 5964 16258 6020 16268
rect 6076 16324 6132 16334
rect 6188 16324 6244 16828
rect 6076 16322 6244 16324
rect 6076 16270 6078 16322
rect 6130 16270 6244 16322
rect 6076 16268 6244 16270
rect 6076 16258 6132 16268
rect 5852 16098 6244 16100
rect 5852 16046 5854 16098
rect 5906 16046 6244 16098
rect 5852 16044 6244 16046
rect 5852 16034 5908 16044
rect 5740 15988 5796 15998
rect 5740 15426 5796 15932
rect 5964 15874 6020 15886
rect 5964 15822 5966 15874
rect 6018 15822 6020 15874
rect 5852 15540 5908 15550
rect 5852 15446 5908 15484
rect 5740 15374 5742 15426
rect 5794 15374 5796 15426
rect 5740 15362 5796 15374
rect 5628 15092 5796 15148
rect 4008 14924 5208 14934
rect 4064 14922 4112 14924
rect 4168 14922 4216 14924
rect 4076 14870 4112 14922
rect 4200 14870 4216 14922
rect 4064 14868 4112 14870
rect 4168 14868 4216 14870
rect 4272 14922 4320 14924
rect 4376 14922 4424 14924
rect 4480 14922 4528 14924
rect 4376 14870 4396 14922
rect 4480 14870 4520 14922
rect 4272 14868 4320 14870
rect 4376 14868 4424 14870
rect 4480 14868 4528 14870
rect 4584 14868 4632 14924
rect 4688 14922 4736 14924
rect 4792 14922 4840 14924
rect 4896 14922 4944 14924
rect 4696 14870 4736 14922
rect 4820 14870 4840 14922
rect 4688 14868 4736 14870
rect 4792 14868 4840 14870
rect 4896 14868 4944 14870
rect 5000 14922 5048 14924
rect 5104 14922 5152 14924
rect 5000 14870 5016 14922
rect 5104 14870 5140 14922
rect 5000 14868 5048 14870
rect 5104 14868 5152 14870
rect 4008 14858 5208 14868
rect 4060 14756 4116 14766
rect 4060 14662 4116 14700
rect 5292 14644 5348 15092
rect 4844 14588 5348 14644
rect 4844 14530 4900 14588
rect 4844 14478 4846 14530
rect 4898 14478 4900 14530
rect 4844 14466 4900 14478
rect 4732 14420 4788 14430
rect 4732 14326 4788 14364
rect 5292 13970 5348 14588
rect 5740 14642 5796 15092
rect 5740 14590 5742 14642
rect 5794 14590 5796 14642
rect 5740 14578 5796 14590
rect 5964 14532 6020 15822
rect 6076 15428 6132 15438
rect 6076 15334 6132 15372
rect 6188 14644 6244 16044
rect 6300 16098 6356 16110
rect 6300 16046 6302 16098
rect 6354 16046 6356 16098
rect 6300 15148 6356 16046
rect 6412 15540 6468 18508
rect 6412 15446 6468 15484
rect 6300 15092 6468 15148
rect 6188 14588 6356 14644
rect 5964 14466 6020 14476
rect 5292 13918 5294 13970
rect 5346 13918 5348 13970
rect 5292 13906 5348 13918
rect 5740 14308 5796 14318
rect 4008 13356 5208 13366
rect 4064 13354 4112 13356
rect 4168 13354 4216 13356
rect 4076 13302 4112 13354
rect 4200 13302 4216 13354
rect 4064 13300 4112 13302
rect 4168 13300 4216 13302
rect 4272 13354 4320 13356
rect 4376 13354 4424 13356
rect 4480 13354 4528 13356
rect 4376 13302 4396 13354
rect 4480 13302 4520 13354
rect 4272 13300 4320 13302
rect 4376 13300 4424 13302
rect 4480 13300 4528 13302
rect 4584 13300 4632 13356
rect 4688 13354 4736 13356
rect 4792 13354 4840 13356
rect 4896 13354 4944 13356
rect 4696 13302 4736 13354
rect 4820 13302 4840 13354
rect 4688 13300 4736 13302
rect 4792 13300 4840 13302
rect 4896 13300 4944 13302
rect 5000 13354 5048 13356
rect 5104 13354 5152 13356
rect 5000 13302 5016 13354
rect 5104 13302 5140 13354
rect 5000 13300 5048 13302
rect 5104 13300 5152 13302
rect 4008 13290 5208 13300
rect 4284 13076 4340 13086
rect 4284 12962 4340 13020
rect 4844 13076 4900 13086
rect 4844 12982 4900 13020
rect 5740 13074 5796 14252
rect 6188 14308 6244 14318
rect 6188 14214 6244 14252
rect 5740 13022 5742 13074
rect 5794 13022 5796 13074
rect 4284 12910 4286 12962
rect 4338 12910 4340 12962
rect 4284 12898 4340 12910
rect 4060 12850 4116 12862
rect 4060 12798 4062 12850
rect 4114 12798 4116 12850
rect 4060 12180 4116 12798
rect 4844 12404 4900 12414
rect 4844 12310 4900 12348
rect 5740 12404 5796 13022
rect 6300 13076 6356 14588
rect 6412 14532 6468 15092
rect 6524 14756 6580 23884
rect 6636 23492 6692 23998
rect 6636 23426 6692 23436
rect 6636 23268 6692 23278
rect 6748 23268 6804 25452
rect 6860 25284 6916 25294
rect 6860 25190 6916 25228
rect 7196 25284 7252 25900
rect 7196 25218 7252 25228
rect 6692 23212 6804 23268
rect 6636 23202 6692 23212
rect 7308 22484 7364 26908
rect 7644 25956 7700 27694
rect 7980 26908 8036 30268
rect 8092 29540 8148 29550
rect 8092 29446 8148 29484
rect 7868 26852 8036 26908
rect 8092 27972 8148 27982
rect 8092 27074 8148 27916
rect 8092 27022 8094 27074
rect 8146 27022 8148 27074
rect 7756 26516 7812 26526
rect 7756 26422 7812 26460
rect 7644 25890 7700 25900
rect 7644 25732 7700 25742
rect 7868 25732 7924 26852
rect 8092 26516 8148 27022
rect 8092 26450 8148 26460
rect 7644 25620 7700 25676
rect 7420 25618 7700 25620
rect 7420 25566 7646 25618
rect 7698 25566 7700 25618
rect 7420 25564 7700 25566
rect 7420 23938 7476 25564
rect 7644 25554 7700 25564
rect 7756 25676 7924 25732
rect 7420 23886 7422 23938
rect 7474 23886 7476 23938
rect 7420 23874 7476 23886
rect 7756 23044 7812 25676
rect 8092 25620 8148 25630
rect 7868 25564 8092 25620
rect 7868 23938 7924 25564
rect 8092 25526 8148 25564
rect 8204 24948 8260 32732
rect 8316 32452 8372 32844
rect 8316 32386 8372 32396
rect 8316 29316 8372 29326
rect 8428 29316 8484 33852
rect 8316 29314 8484 29316
rect 8316 29262 8318 29314
rect 8370 29262 8484 29314
rect 8316 29260 8484 29262
rect 8540 31554 8596 31566
rect 8540 31502 8542 31554
rect 8594 31502 8596 31554
rect 8540 30210 8596 31502
rect 8540 30158 8542 30210
rect 8594 30158 8596 30210
rect 8540 29426 8596 30158
rect 8540 29374 8542 29426
rect 8594 29374 8596 29426
rect 8316 29250 8372 29260
rect 8316 28420 8372 28430
rect 8316 27298 8372 28364
rect 8540 27972 8596 29374
rect 8540 27906 8596 27916
rect 8652 27748 8708 33852
rect 9324 33124 9380 33134
rect 9436 33124 9492 34636
rect 9548 34626 9604 34636
rect 9548 34132 9604 34142
rect 9772 34132 9828 34860
rect 9884 34356 9940 34394
rect 9884 34290 9940 34300
rect 9604 34076 9828 34132
rect 9884 34132 9940 34142
rect 9996 34132 10052 35084
rect 10332 35074 10388 35084
rect 10444 34916 10500 37100
rect 10556 37044 10612 37054
rect 10556 37042 10724 37044
rect 10556 36990 10558 37042
rect 10610 36990 10724 37042
rect 10556 36988 10724 36990
rect 10556 36978 10612 36988
rect 9884 34130 10052 34132
rect 9884 34078 9886 34130
rect 9938 34078 10052 34130
rect 9884 34076 10052 34078
rect 10108 34860 10500 34916
rect 9548 34038 9604 34076
rect 9884 34066 9940 34076
rect 9380 33068 9492 33124
rect 9324 33058 9380 33068
rect 8876 31892 8932 31902
rect 8876 31798 8932 31836
rect 9996 31892 10052 31902
rect 9996 31780 10052 31836
rect 9660 31778 10052 31780
rect 9660 31726 9998 31778
rect 10050 31726 10052 31778
rect 9660 31724 10052 31726
rect 9660 31218 9716 31724
rect 9996 31714 10052 31724
rect 9660 31166 9662 31218
rect 9714 31166 9716 31218
rect 8988 30996 9044 31006
rect 8988 30902 9044 30940
rect 9660 30996 9716 31166
rect 9660 30930 9716 30940
rect 8876 30098 8932 30110
rect 8876 30046 8878 30098
rect 8930 30046 8932 30098
rect 8876 29540 8932 30046
rect 8876 29474 8932 29484
rect 9772 29988 9828 29998
rect 9772 29426 9828 29932
rect 9772 29374 9774 29426
rect 9826 29374 9828 29426
rect 9772 29362 9828 29374
rect 9996 29988 10052 29998
rect 9660 29316 9716 29326
rect 9660 29222 9716 29260
rect 9884 28756 9940 28766
rect 9548 28644 9604 28654
rect 9548 28550 9604 28588
rect 9548 27972 9604 27982
rect 9604 27916 9716 27972
rect 9548 27878 9604 27916
rect 8316 27246 8318 27298
rect 8370 27246 8372 27298
rect 8316 27234 8372 27246
rect 8540 27692 8708 27748
rect 8876 27746 8932 27758
rect 8876 27694 8878 27746
rect 8930 27694 8932 27746
rect 8316 27076 8372 27086
rect 8316 26514 8372 27020
rect 8316 26462 8318 26514
rect 8370 26462 8372 26514
rect 8316 26450 8372 26462
rect 7868 23886 7870 23938
rect 7922 23886 7924 23938
rect 7868 23874 7924 23886
rect 7980 24892 8260 24948
rect 8540 24946 8596 27692
rect 8652 27524 8708 27534
rect 8652 27298 8708 27468
rect 8652 27246 8654 27298
rect 8706 27246 8708 27298
rect 8652 27234 8708 27246
rect 8876 27076 8932 27694
rect 9324 27300 9380 27310
rect 9324 27186 9380 27244
rect 9324 27134 9326 27186
rect 9378 27134 9380 27186
rect 9324 27122 9380 27134
rect 9660 27188 9716 27916
rect 9884 27748 9940 28700
rect 9996 28642 10052 29932
rect 9996 28590 9998 28642
rect 10050 28590 10052 28642
rect 9996 28578 10052 28590
rect 10108 28082 10164 34860
rect 10556 34804 10612 34814
rect 10556 34710 10612 34748
rect 10668 34356 10724 36988
rect 10892 36596 10948 36606
rect 10892 36502 10948 36540
rect 10892 35476 10948 35486
rect 10892 35382 10948 35420
rect 10892 35140 10948 35150
rect 10892 35046 10948 35084
rect 11116 34916 11172 34926
rect 11116 34822 11172 34860
rect 10556 34244 10612 34254
rect 10668 34244 10724 34300
rect 11228 34804 11284 38612
rect 11452 37156 11508 40684
rect 11676 40404 11732 40908
rect 11788 40628 11844 41022
rect 11788 40562 11844 40572
rect 11788 40404 11844 40414
rect 11676 40402 11844 40404
rect 11676 40350 11790 40402
rect 11842 40350 11844 40402
rect 11676 40348 11844 40350
rect 11788 40338 11844 40348
rect 11452 37062 11508 37100
rect 11564 38836 11620 38846
rect 11340 36372 11396 36382
rect 11340 36278 11396 36316
rect 11228 34354 11284 34748
rect 11228 34302 11230 34354
rect 11282 34302 11284 34354
rect 11228 34290 11284 34302
rect 10556 34242 10724 34244
rect 10556 34190 10558 34242
rect 10610 34190 10724 34242
rect 10556 34188 10724 34190
rect 10556 34178 10612 34188
rect 10220 34132 10276 34142
rect 10444 34132 10500 34142
rect 10220 34130 10500 34132
rect 10220 34078 10222 34130
rect 10274 34078 10446 34130
rect 10498 34078 10500 34130
rect 10220 34076 10500 34078
rect 10220 34066 10276 34076
rect 10444 34066 10500 34076
rect 10780 34020 10836 34030
rect 10556 33348 10612 33358
rect 10556 33254 10612 33292
rect 10220 31780 10276 31790
rect 10220 30324 10276 31724
rect 10780 30434 10836 33964
rect 11564 33460 11620 38780
rect 11900 38834 11956 41358
rect 12012 41188 12068 41198
rect 12012 41094 12068 41132
rect 11900 38782 11902 38834
rect 11954 38782 11956 38834
rect 11900 38770 11956 38782
rect 11676 37826 11732 37838
rect 11676 37774 11678 37826
rect 11730 37774 11732 37826
rect 11676 37380 11732 37774
rect 12236 37492 12292 42364
rect 12348 41412 12404 41422
rect 12348 41318 12404 41356
rect 12572 41410 12628 42588
rect 12684 42084 12740 42094
rect 12796 42084 12852 42588
rect 12684 42082 12852 42084
rect 12684 42030 12686 42082
rect 12738 42030 12852 42082
rect 12684 42028 12852 42030
rect 13244 43372 13356 43428
rect 12684 42018 12740 42028
rect 12572 41358 12574 41410
rect 12626 41358 12628 41410
rect 12572 41346 12628 41358
rect 12348 37492 12404 37502
rect 12236 37490 12404 37492
rect 12236 37438 12350 37490
rect 12402 37438 12404 37490
rect 12236 37436 12404 37438
rect 11676 37324 12068 37380
rect 12012 37268 12068 37324
rect 12236 37268 12292 37278
rect 12012 37212 12236 37268
rect 11900 37154 11956 37166
rect 11900 37102 11902 37154
rect 11954 37102 11956 37154
rect 11900 36706 11956 37102
rect 11900 36654 11902 36706
rect 11954 36654 11956 36706
rect 11900 36642 11956 36654
rect 12124 36596 12180 36606
rect 12012 36594 12180 36596
rect 12012 36542 12126 36594
rect 12178 36542 12180 36594
rect 12012 36540 12180 36542
rect 11900 36484 11956 36494
rect 12012 36484 12068 36540
rect 12124 36530 12180 36540
rect 11900 36482 12068 36484
rect 11900 36430 11902 36482
rect 11954 36430 12068 36482
rect 11900 36428 12068 36430
rect 11900 36418 11956 36428
rect 12124 36372 12180 36382
rect 11900 35700 11956 35710
rect 12124 35700 12180 36316
rect 11900 35698 12180 35700
rect 11900 35646 11902 35698
rect 11954 35646 12180 35698
rect 11900 35644 12180 35646
rect 11900 35634 11956 35644
rect 12012 35364 12068 35644
rect 11788 34916 11844 34926
rect 11676 34804 11732 34814
rect 11676 34710 11732 34748
rect 11676 34020 11732 34030
rect 11788 34020 11844 34860
rect 11732 33964 11844 34020
rect 11676 33926 11732 33964
rect 12012 33460 12068 35308
rect 12124 34356 12180 34366
rect 12124 34262 12180 34300
rect 12236 33908 12292 37212
rect 12236 33842 12292 33852
rect 12348 36594 12404 37436
rect 12572 37380 12628 37390
rect 12572 37286 12628 37324
rect 12908 37378 12964 37390
rect 12908 37326 12910 37378
rect 12962 37326 12964 37378
rect 12796 37266 12852 37278
rect 12796 37214 12798 37266
rect 12850 37214 12852 37266
rect 12796 37156 12852 37214
rect 12796 37090 12852 37100
rect 12348 36542 12350 36594
rect 12402 36542 12404 36594
rect 11228 33458 11956 33460
rect 11228 33406 11566 33458
rect 11618 33406 11956 33458
rect 11228 33404 11956 33406
rect 11228 33346 11284 33404
rect 11564 33394 11620 33404
rect 11228 33294 11230 33346
rect 11282 33294 11284 33346
rect 11228 33282 11284 33294
rect 11900 32788 11956 33404
rect 12012 33366 12068 33404
rect 12012 32788 12068 32798
rect 11900 32786 12292 32788
rect 11900 32734 12014 32786
rect 12066 32734 12292 32786
rect 11900 32732 12292 32734
rect 11900 31892 11956 32732
rect 12012 32722 12068 32732
rect 12236 32562 12292 32732
rect 12236 32510 12238 32562
rect 12290 32510 12292 32562
rect 12236 32498 12292 32510
rect 10780 30382 10782 30434
rect 10834 30382 10836 30434
rect 10780 30370 10836 30382
rect 11564 31890 11956 31892
rect 11564 31838 11902 31890
rect 11954 31838 11956 31890
rect 11564 31836 11956 31838
rect 10220 30210 10276 30268
rect 10220 30158 10222 30210
rect 10274 30158 10276 30210
rect 10220 30146 10276 30158
rect 10332 30100 10388 30110
rect 10332 29538 10388 30044
rect 11340 29988 11396 29998
rect 11340 29894 11396 29932
rect 10780 29652 10836 29662
rect 10780 29558 10836 29596
rect 10332 29486 10334 29538
rect 10386 29486 10388 29538
rect 10332 29474 10388 29486
rect 11564 29426 11620 31836
rect 11900 31826 11956 31836
rect 11676 30212 11732 30222
rect 11676 30118 11732 30156
rect 12236 30100 12292 30110
rect 12012 30098 12292 30100
rect 12012 30046 12238 30098
rect 12290 30046 12292 30098
rect 12012 30044 12292 30046
rect 11564 29374 11566 29426
rect 11618 29374 11620 29426
rect 11564 28644 11620 29374
rect 11900 29428 11956 29438
rect 11900 29334 11956 29372
rect 11564 28578 11620 28588
rect 10108 28030 10110 28082
rect 10162 28030 10164 28082
rect 10108 28018 10164 28030
rect 12012 28082 12068 30044
rect 12236 30034 12292 30044
rect 12348 29652 12404 36542
rect 12908 36706 12964 37326
rect 13244 37268 13300 43372
rect 13356 43334 13412 43372
rect 13468 40628 13524 44044
rect 13580 42980 13636 44604
rect 13916 44548 13972 45276
rect 14140 45108 14196 45276
rect 14924 45332 14980 45342
rect 15372 45332 15428 45614
rect 14924 45330 15428 45332
rect 14924 45278 14926 45330
rect 14978 45278 15428 45330
rect 14924 45276 15428 45278
rect 14924 45266 14980 45276
rect 14140 45014 14196 45052
rect 14364 45108 14420 45118
rect 13580 42886 13636 42924
rect 13692 44492 13972 44548
rect 14028 44994 14084 45006
rect 14028 44942 14030 44994
rect 14082 44942 14084 44994
rect 13468 40562 13524 40572
rect 13580 42644 13636 42654
rect 13580 40292 13636 42588
rect 13580 40226 13636 40236
rect 13356 38724 13412 38734
rect 13692 38668 13748 44492
rect 14028 44322 14084 44942
rect 14364 44772 14420 45052
rect 14476 45106 14532 45118
rect 14476 45054 14478 45106
rect 14530 45054 14532 45106
rect 14476 44996 14532 45054
rect 15148 45108 15204 45118
rect 15148 45014 15204 45052
rect 15372 45108 15428 45276
rect 14812 44996 14868 45006
rect 14476 44994 14868 44996
rect 14476 44942 14814 44994
rect 14866 44942 14868 44994
rect 14476 44940 14868 44942
rect 14812 44930 14868 44940
rect 14364 44706 14420 44716
rect 15372 44772 15428 45052
rect 15372 44706 15428 44716
rect 15484 44996 15540 45006
rect 14028 44270 14030 44322
rect 14082 44270 14084 44322
rect 14028 44258 14084 44270
rect 14008 43932 15208 43942
rect 14064 43930 14112 43932
rect 14168 43930 14216 43932
rect 14076 43878 14112 43930
rect 14200 43878 14216 43930
rect 14064 43876 14112 43878
rect 14168 43876 14216 43878
rect 14272 43930 14320 43932
rect 14376 43930 14424 43932
rect 14480 43930 14528 43932
rect 14376 43878 14396 43930
rect 14480 43878 14520 43930
rect 14272 43876 14320 43878
rect 14376 43876 14424 43878
rect 14480 43876 14528 43878
rect 14584 43876 14632 43932
rect 14688 43930 14736 43932
rect 14792 43930 14840 43932
rect 14896 43930 14944 43932
rect 14696 43878 14736 43930
rect 14820 43878 14840 43930
rect 14688 43876 14736 43878
rect 14792 43876 14840 43878
rect 14896 43876 14944 43878
rect 15000 43930 15048 43932
rect 15104 43930 15152 43932
rect 15000 43878 15016 43930
rect 15104 43878 15140 43930
rect 15000 43876 15048 43878
rect 15104 43876 15152 43878
rect 14008 43866 15208 43876
rect 13916 43652 13972 43662
rect 13916 43558 13972 43596
rect 14252 43652 14308 43662
rect 14252 43558 14308 43596
rect 15484 43652 15540 44940
rect 15484 43558 15540 43596
rect 14140 43538 14196 43550
rect 14140 43486 14142 43538
rect 14194 43486 14196 43538
rect 14140 43428 14196 43486
rect 14476 43540 14532 43550
rect 14476 43446 14532 43484
rect 14028 42978 14084 42990
rect 14028 42926 14030 42978
rect 14082 42926 14084 42978
rect 14028 42866 14084 42926
rect 14028 42814 14030 42866
rect 14082 42814 14084 42866
rect 14028 42802 14084 42814
rect 13804 42644 13860 42654
rect 13804 42194 13860 42588
rect 14140 42644 14196 43372
rect 14140 42578 14196 42588
rect 14008 42364 15208 42374
rect 14064 42362 14112 42364
rect 14168 42362 14216 42364
rect 14076 42310 14112 42362
rect 14200 42310 14216 42362
rect 14064 42308 14112 42310
rect 14168 42308 14216 42310
rect 14272 42362 14320 42364
rect 14376 42362 14424 42364
rect 14480 42362 14528 42364
rect 14376 42310 14396 42362
rect 14480 42310 14520 42362
rect 14272 42308 14320 42310
rect 14376 42308 14424 42310
rect 14480 42308 14528 42310
rect 14584 42308 14632 42364
rect 14688 42362 14736 42364
rect 14792 42362 14840 42364
rect 14896 42362 14944 42364
rect 14696 42310 14736 42362
rect 14820 42310 14840 42362
rect 14688 42308 14736 42310
rect 14792 42308 14840 42310
rect 14896 42308 14944 42310
rect 15000 42362 15048 42364
rect 15104 42362 15152 42364
rect 15000 42310 15016 42362
rect 15104 42310 15140 42362
rect 15000 42308 15048 42310
rect 15104 42308 15152 42310
rect 14008 42298 15208 42308
rect 13804 42142 13806 42194
rect 13858 42142 13860 42194
rect 13804 42130 13860 42142
rect 14008 40796 15208 40806
rect 14064 40794 14112 40796
rect 14168 40794 14216 40796
rect 14076 40742 14112 40794
rect 14200 40742 14216 40794
rect 14064 40740 14112 40742
rect 14168 40740 14216 40742
rect 14272 40794 14320 40796
rect 14376 40794 14424 40796
rect 14480 40794 14528 40796
rect 14376 40742 14396 40794
rect 14480 40742 14520 40794
rect 14272 40740 14320 40742
rect 14376 40740 14424 40742
rect 14480 40740 14528 40742
rect 14584 40740 14632 40796
rect 14688 40794 14736 40796
rect 14792 40794 14840 40796
rect 14896 40794 14944 40796
rect 14696 40742 14736 40794
rect 14820 40742 14840 40794
rect 14688 40740 14736 40742
rect 14792 40740 14840 40742
rect 14896 40740 14944 40742
rect 15000 40794 15048 40796
rect 15104 40794 15152 40796
rect 15000 40742 15016 40794
rect 15104 40742 15140 40794
rect 15000 40740 15048 40742
rect 15104 40740 15152 40742
rect 14008 40730 15208 40740
rect 13804 40628 13860 40638
rect 13804 39060 13860 40572
rect 14140 40628 14196 40638
rect 14140 40534 14196 40572
rect 15148 40628 15204 40638
rect 14924 40404 14980 40414
rect 14924 39730 14980 40348
rect 15036 40402 15092 40414
rect 15036 40350 15038 40402
rect 15090 40350 15092 40402
rect 15036 40292 15092 40350
rect 15036 40226 15092 40236
rect 15148 39842 15204 40572
rect 15148 39790 15150 39842
rect 15202 39790 15204 39842
rect 15148 39778 15204 39790
rect 15484 40290 15540 40302
rect 15484 40238 15486 40290
rect 15538 40238 15540 40290
rect 14924 39678 14926 39730
rect 14978 39678 14980 39730
rect 14924 39666 14980 39678
rect 14008 39228 15208 39238
rect 14064 39226 14112 39228
rect 14168 39226 14216 39228
rect 14076 39174 14112 39226
rect 14200 39174 14216 39226
rect 14064 39172 14112 39174
rect 14168 39172 14216 39174
rect 14272 39226 14320 39228
rect 14376 39226 14424 39228
rect 14480 39226 14528 39228
rect 14376 39174 14396 39226
rect 14480 39174 14520 39226
rect 14272 39172 14320 39174
rect 14376 39172 14424 39174
rect 14480 39172 14528 39174
rect 14584 39172 14632 39228
rect 14688 39226 14736 39228
rect 14792 39226 14840 39228
rect 14896 39226 14944 39228
rect 14696 39174 14736 39226
rect 14820 39174 14840 39226
rect 14688 39172 14736 39174
rect 14792 39172 14840 39174
rect 14896 39172 14944 39174
rect 15000 39226 15048 39228
rect 15104 39226 15152 39228
rect 15000 39174 15016 39226
rect 15104 39174 15140 39226
rect 15000 39172 15048 39174
rect 15104 39172 15152 39174
rect 14008 39162 15208 39172
rect 14140 39060 14196 39070
rect 13804 39058 14196 39060
rect 13804 39006 14142 39058
rect 14194 39006 14196 39058
rect 13804 39004 14196 39006
rect 14140 38994 14196 39004
rect 14924 39060 14980 39070
rect 14924 38966 14980 39004
rect 15484 39058 15540 40238
rect 15484 39006 15486 39058
rect 15538 39006 15540 39058
rect 15484 38836 15540 39006
rect 15484 38770 15540 38780
rect 13356 37490 13412 38668
rect 13356 37438 13358 37490
rect 13410 37438 13412 37490
rect 13356 37426 13412 37438
rect 13580 38612 13748 38668
rect 15708 38668 15764 49196
rect 15820 49028 15876 49038
rect 15820 48934 15876 48972
rect 15932 48244 15988 48254
rect 15932 48150 15988 48188
rect 16044 46002 16100 51436
rect 16268 51426 16324 51436
rect 16156 50594 16212 50606
rect 16156 50542 16158 50594
rect 16210 50542 16212 50594
rect 16156 49028 16212 50542
rect 16492 50428 16548 60510
rect 16604 60564 16660 60574
rect 16660 60508 16772 60564
rect 16604 60498 16660 60508
rect 16604 58324 16660 58334
rect 16604 58230 16660 58268
rect 16716 55524 16772 60508
rect 17276 59444 17332 62860
rect 17276 59378 17332 59388
rect 17500 59220 17556 67564
rect 17612 67554 17668 67564
rect 17612 67172 17668 67182
rect 17724 67172 17780 67676
rect 17948 67666 18004 67676
rect 18060 67282 18116 67294
rect 18060 67230 18062 67282
rect 18114 67230 18116 67282
rect 17668 67116 17780 67172
rect 17948 67170 18004 67182
rect 17948 67118 17950 67170
rect 18002 67118 18004 67170
rect 17612 67078 17668 67116
rect 17948 67060 18004 67118
rect 17948 66994 18004 67004
rect 17836 66836 17892 66846
rect 17612 66052 17668 66062
rect 17612 65958 17668 65996
rect 17836 65378 17892 66780
rect 18060 66276 18116 67230
rect 18172 66500 18228 68572
rect 18396 68628 18452 68638
rect 18396 68626 18676 68628
rect 18396 68574 18398 68626
rect 18450 68574 18676 68626
rect 18396 68572 18676 68574
rect 18396 68562 18452 68572
rect 18172 66434 18228 66444
rect 17836 65326 17838 65378
rect 17890 65326 17892 65378
rect 17612 64484 17668 64494
rect 17836 64484 17892 65326
rect 17612 64482 17892 64484
rect 17612 64430 17614 64482
rect 17666 64430 17892 64482
rect 17612 64428 17892 64430
rect 17948 66220 18116 66276
rect 18172 66276 18228 66286
rect 17612 63924 17668 64428
rect 17948 64148 18004 66220
rect 18060 66052 18116 66062
rect 18172 66052 18228 66220
rect 18508 66164 18564 66174
rect 18508 66070 18564 66108
rect 18060 66050 18228 66052
rect 18060 65998 18062 66050
rect 18114 65998 18228 66050
rect 18060 65996 18228 65998
rect 18060 65986 18116 65996
rect 18284 65378 18340 65390
rect 18284 65326 18286 65378
rect 18338 65326 18340 65378
rect 18172 65268 18228 65278
rect 17612 63858 17668 63868
rect 17836 64092 18004 64148
rect 18060 65156 18116 65166
rect 17724 61684 17780 61694
rect 17724 61346 17780 61628
rect 17724 61294 17726 61346
rect 17778 61294 17780 61346
rect 17724 61282 17780 61294
rect 17276 59164 17556 59220
rect 17164 58436 17220 58446
rect 17164 58342 17220 58380
rect 16828 57540 16884 57550
rect 16828 56868 16884 57484
rect 16828 56802 16884 56812
rect 16828 56644 16884 56654
rect 16828 56550 16884 56588
rect 17052 56084 17108 56094
rect 16940 56028 17052 56084
rect 16828 55970 16884 55982
rect 16828 55918 16830 55970
rect 16882 55918 16884 55970
rect 16828 55860 16884 55918
rect 16828 55794 16884 55804
rect 16940 55636 16996 56028
rect 17052 56018 17108 56028
rect 17276 55748 17332 59164
rect 17836 58828 17892 64092
rect 18060 64036 18116 65100
rect 18172 64818 18228 65212
rect 18172 64766 18174 64818
rect 18226 64766 18228 64818
rect 18172 64754 18228 64766
rect 18284 64708 18340 65326
rect 18284 64484 18340 64652
rect 18284 64418 18340 64428
rect 18508 64484 18564 64494
rect 17948 63980 18116 64036
rect 17948 63922 18004 63980
rect 17948 63870 17950 63922
rect 18002 63870 18004 63922
rect 17948 63858 18004 63870
rect 18284 63924 18340 63934
rect 18060 63810 18116 63822
rect 18060 63758 18062 63810
rect 18114 63758 18116 63810
rect 18060 63362 18116 63758
rect 18060 63310 18062 63362
rect 18114 63310 18116 63362
rect 18060 63298 18116 63310
rect 18172 63026 18228 63038
rect 18172 62974 18174 63026
rect 18226 62974 18228 63026
rect 18172 62692 18228 62974
rect 18172 62626 18228 62636
rect 18284 62468 18340 63868
rect 18172 62412 18340 62468
rect 17388 58772 17892 58828
rect 18060 59106 18116 59118
rect 18060 59054 18062 59106
rect 18114 59054 18116 59106
rect 18060 58828 18116 59054
rect 18172 58828 18228 62412
rect 18508 59668 18564 64428
rect 18620 61908 18676 68572
rect 18732 68626 18788 68638
rect 18732 68574 18734 68626
rect 18786 68574 18788 68626
rect 18732 66948 18788 68574
rect 19180 68626 19236 68638
rect 19180 68574 19182 68626
rect 19234 68574 19236 68626
rect 19180 68180 19236 68574
rect 19180 67396 19236 68124
rect 18732 66882 18788 66892
rect 18956 67340 19236 67396
rect 19404 68626 19460 68908
rect 19404 68574 19406 68626
rect 19458 68574 19460 68626
rect 18956 67058 19012 67340
rect 19404 67172 19460 68574
rect 19516 68628 19572 68638
rect 19628 68628 19684 69132
rect 19740 69122 19796 69132
rect 19740 68852 19796 68862
rect 19740 68738 19796 68796
rect 19964 68740 20020 68750
rect 19740 68686 19742 68738
rect 19794 68686 19796 68738
rect 19740 68674 19796 68686
rect 19852 68738 20020 68740
rect 19852 68686 19966 68738
rect 20018 68686 20020 68738
rect 19852 68684 20020 68686
rect 19572 68572 19684 68628
rect 19516 68562 19572 68572
rect 19628 67620 19684 67630
rect 19628 67618 19796 67620
rect 19628 67566 19630 67618
rect 19682 67566 19796 67618
rect 19628 67564 19796 67566
rect 19628 67554 19684 67564
rect 19404 67106 19460 67116
rect 18956 67006 18958 67058
rect 19010 67006 19012 67058
rect 18732 66276 18788 66286
rect 18956 66276 19012 67006
rect 19068 67058 19124 67070
rect 19068 67006 19070 67058
rect 19122 67006 19124 67058
rect 19068 66500 19124 67006
rect 19180 67060 19236 67070
rect 19180 66836 19236 67004
rect 19180 66770 19236 66780
rect 19628 67058 19684 67070
rect 19628 67006 19630 67058
rect 19682 67006 19684 67058
rect 19628 66724 19684 67006
rect 19740 66948 19796 67564
rect 19852 67282 19908 68684
rect 19964 68674 20020 68684
rect 20076 68514 20132 70924
rect 20636 68628 20692 68638
rect 20636 68626 20916 68628
rect 20636 68574 20638 68626
rect 20690 68574 20916 68626
rect 20636 68572 20916 68574
rect 20636 68562 20692 68572
rect 20076 68462 20078 68514
rect 20130 68462 20132 68514
rect 20076 68450 20132 68462
rect 20748 68402 20804 68414
rect 20748 68350 20750 68402
rect 20802 68350 20804 68402
rect 20748 68068 20804 68350
rect 20748 68002 20804 68012
rect 20636 67842 20692 67854
rect 20636 67790 20638 67842
rect 20690 67790 20692 67842
rect 19852 67230 19854 67282
rect 19906 67230 19908 67282
rect 19852 67218 19908 67230
rect 19964 67618 20020 67630
rect 19964 67566 19966 67618
rect 20018 67566 20020 67618
rect 19964 66948 20020 67566
rect 20076 67620 20132 67630
rect 20076 67526 20132 67564
rect 20188 67620 20244 67630
rect 20188 67618 20356 67620
rect 20188 67566 20190 67618
rect 20242 67566 20356 67618
rect 20188 67564 20356 67566
rect 20188 67554 20244 67564
rect 19740 66892 20020 66948
rect 19516 66668 19684 66724
rect 19292 66500 19348 66510
rect 19068 66444 19236 66500
rect 19180 66386 19236 66444
rect 19180 66334 19182 66386
rect 19234 66334 19236 66386
rect 19068 66276 19124 66286
rect 18956 66274 19124 66276
rect 18956 66222 19070 66274
rect 19122 66222 19124 66274
rect 18956 66220 19124 66222
rect 18732 65714 18788 66220
rect 18732 65662 18734 65714
rect 18786 65662 18788 65714
rect 18732 65650 18788 65662
rect 19068 65602 19124 66220
rect 19180 66276 19236 66334
rect 19180 66210 19236 66220
rect 19068 65550 19070 65602
rect 19122 65550 19124 65602
rect 18956 65380 19012 65390
rect 18956 65156 19012 65324
rect 19068 65268 19124 65550
rect 19068 65202 19124 65212
rect 19180 65492 19236 65502
rect 18732 65100 19012 65156
rect 18732 64818 18788 65100
rect 19180 65044 19236 65436
rect 18732 64766 18734 64818
rect 18786 64766 18788 64818
rect 18732 64754 18788 64766
rect 18844 64988 19236 65044
rect 18844 62188 18900 64988
rect 19292 64932 19348 66444
rect 19516 66052 19572 66668
rect 19516 65986 19572 65996
rect 19628 66498 19684 66510
rect 19628 66446 19630 66498
rect 19682 66446 19684 66498
rect 19628 65490 19684 66446
rect 19964 66164 20020 66892
rect 20188 66946 20244 66958
rect 20188 66894 20190 66946
rect 20242 66894 20244 66946
rect 20188 66276 20244 66894
rect 20188 66210 20244 66220
rect 19964 66098 20020 66108
rect 19628 65438 19630 65490
rect 19682 65438 19684 65490
rect 19628 65426 19684 65438
rect 20300 65492 20356 67564
rect 20636 66498 20692 67790
rect 20636 66446 20638 66498
rect 20690 66446 20692 66498
rect 20636 66434 20692 66446
rect 20636 66276 20692 66286
rect 20636 66162 20692 66220
rect 20636 66110 20638 66162
rect 20690 66110 20692 66162
rect 20636 66098 20692 66110
rect 20748 66164 20804 66174
rect 20300 65426 20356 65436
rect 20412 65716 20468 65726
rect 19740 65380 19796 65390
rect 19740 65286 19796 65324
rect 20076 65380 20132 65390
rect 19964 65266 20020 65278
rect 19964 65214 19966 65266
rect 20018 65214 20020 65266
rect 19180 64876 19348 64932
rect 19516 65156 19572 65166
rect 18956 64706 19012 64718
rect 18956 64654 18958 64706
rect 19010 64654 19012 64706
rect 18956 63924 19012 64654
rect 18956 63858 19012 63868
rect 19068 62914 19124 62926
rect 19068 62862 19070 62914
rect 19122 62862 19124 62914
rect 19068 62468 19124 62862
rect 19068 62402 19124 62412
rect 18844 62132 19012 62188
rect 18620 61852 18900 61908
rect 18060 58772 18228 58828
rect 17388 58212 17444 58772
rect 17500 58436 17556 58446
rect 17500 58434 17892 58436
rect 17500 58382 17502 58434
rect 17554 58382 17892 58434
rect 17500 58380 17892 58382
rect 17500 58370 17556 58380
rect 17724 58212 17780 58222
rect 17388 58156 17556 58212
rect 17388 56978 17444 56990
rect 17388 56926 17390 56978
rect 17442 56926 17444 56978
rect 17388 56644 17444 56926
rect 17388 56578 17444 56588
rect 17388 56084 17444 56094
rect 17388 55990 17444 56028
rect 17276 55692 17444 55748
rect 16156 48962 16212 48972
rect 16380 50372 16548 50428
rect 16604 55468 16772 55524
rect 16828 55580 16996 55636
rect 16044 45950 16046 46002
rect 16098 45950 16100 46002
rect 16044 45938 16100 45950
rect 16380 45892 16436 50372
rect 16604 49922 16660 55468
rect 16828 55410 16884 55580
rect 16828 55358 16830 55410
rect 16882 55358 16884 55410
rect 16828 55346 16884 55358
rect 16828 53844 16884 53854
rect 16828 50706 16884 53788
rect 16828 50654 16830 50706
rect 16882 50654 16884 50706
rect 16828 50642 16884 50654
rect 17276 51154 17332 51166
rect 17276 51102 17278 51154
rect 17330 51102 17332 51154
rect 17276 50484 17332 51102
rect 17388 50596 17444 55692
rect 17388 50530 17444 50540
rect 17276 50418 17332 50428
rect 17500 50428 17556 58156
rect 17612 57652 17668 57662
rect 17612 56866 17668 57596
rect 17724 57538 17780 58156
rect 17724 57486 17726 57538
rect 17778 57486 17780 57538
rect 17724 57204 17780 57486
rect 17836 57426 17892 58380
rect 17836 57374 17838 57426
rect 17890 57374 17892 57426
rect 17836 57362 17892 57374
rect 18060 58322 18116 58334
rect 18060 58270 18062 58322
rect 18114 58270 18116 58322
rect 17724 57138 17780 57148
rect 17612 56814 17614 56866
rect 17666 56814 17668 56866
rect 17612 56802 17668 56814
rect 18060 56756 18116 58270
rect 18172 58324 18228 58772
rect 18172 58258 18228 58268
rect 18284 59612 18564 59668
rect 18284 57652 18340 59612
rect 18396 59444 18452 59454
rect 18396 59350 18452 59388
rect 18508 59332 18564 59342
rect 18508 59330 18676 59332
rect 18508 59278 18510 59330
rect 18562 59278 18676 59330
rect 18508 59276 18676 59278
rect 18508 59266 18564 59276
rect 18508 58436 18564 58446
rect 18508 58342 18564 58380
rect 18396 58324 18452 58334
rect 18396 58230 18452 58268
rect 18620 58212 18676 59276
rect 18732 59220 18788 59230
rect 18732 59126 18788 59164
rect 18844 58660 18900 61852
rect 18844 58594 18900 58604
rect 18956 58884 19012 62132
rect 19068 59778 19124 59790
rect 19068 59726 19070 59778
rect 19122 59726 19124 59778
rect 19068 59556 19124 59726
rect 19068 59490 19124 59500
rect 18956 58548 19012 58828
rect 19068 59218 19124 59230
rect 19068 59166 19070 59218
rect 19122 59166 19124 59218
rect 19068 58772 19124 59166
rect 19068 58706 19124 58716
rect 18956 58492 19124 58548
rect 19068 58434 19124 58492
rect 19068 58382 19070 58434
rect 19122 58382 19124 58434
rect 18844 58322 18900 58334
rect 18844 58270 18846 58322
rect 18898 58270 18900 58322
rect 18732 58212 18788 58222
rect 18620 58210 18788 58212
rect 18620 58158 18734 58210
rect 18786 58158 18788 58210
rect 18620 58156 18788 58158
rect 18732 58146 18788 58156
rect 18844 58212 18900 58270
rect 18172 57596 18340 57652
rect 18396 58100 18452 58110
rect 18172 57540 18228 57596
rect 18172 57446 18228 57484
rect 18284 57426 18340 57438
rect 18284 57374 18286 57426
rect 18338 57374 18340 57426
rect 18060 56690 18116 56700
rect 18172 56754 18228 56766
rect 18172 56702 18174 56754
rect 18226 56702 18228 56754
rect 18172 56196 18228 56702
rect 17612 56140 18228 56196
rect 17612 56082 17668 56140
rect 17612 56030 17614 56082
rect 17666 56030 17668 56082
rect 17612 56018 17668 56030
rect 17836 55858 17892 55870
rect 17836 55806 17838 55858
rect 17890 55806 17892 55858
rect 17836 55748 17892 55806
rect 18060 55860 18116 55870
rect 18060 55766 18116 55804
rect 17836 55682 17892 55692
rect 18284 54852 18340 57374
rect 18396 57428 18452 58044
rect 18844 57988 18900 58156
rect 19068 58100 19124 58382
rect 19068 58034 19124 58044
rect 18620 57932 18900 57988
rect 18620 57652 18676 57932
rect 19180 57876 19236 64876
rect 19516 64594 19572 65100
rect 19516 64542 19518 64594
rect 19570 64542 19572 64594
rect 19516 64530 19572 64542
rect 19964 65044 20020 65214
rect 19292 64484 19348 64494
rect 19292 64390 19348 64428
rect 19628 64482 19684 64494
rect 19628 64430 19630 64482
rect 19682 64430 19684 64482
rect 19516 63922 19572 63934
rect 19516 63870 19518 63922
rect 19570 63870 19572 63922
rect 19516 63140 19572 63870
rect 19628 63810 19684 64430
rect 19964 64036 20020 64988
rect 19964 63970 20020 63980
rect 19964 63812 20020 63822
rect 19628 63758 19630 63810
rect 19682 63758 19684 63810
rect 19628 63746 19684 63758
rect 19740 63810 20020 63812
rect 19740 63758 19966 63810
rect 20018 63758 20020 63810
rect 19740 63756 20020 63758
rect 19516 63084 19684 63140
rect 19404 63028 19460 63038
rect 19404 62934 19460 62972
rect 19516 62914 19572 62926
rect 19516 62862 19518 62914
rect 19570 62862 19572 62914
rect 19404 62580 19460 62590
rect 19292 62468 19348 62478
rect 19292 62374 19348 62412
rect 19292 59890 19348 59902
rect 19292 59838 19294 59890
rect 19346 59838 19348 59890
rect 19292 58884 19348 59838
rect 19292 58818 19348 58828
rect 19404 58828 19460 62524
rect 19516 62356 19572 62862
rect 19516 62290 19572 62300
rect 19628 62692 19684 63084
rect 19628 60114 19684 62636
rect 19740 62354 19796 63756
rect 19964 63746 20020 63756
rect 20076 63140 20132 65324
rect 20188 65266 20244 65278
rect 20188 65214 20190 65266
rect 20242 65214 20244 65266
rect 20188 64708 20244 65214
rect 20300 65268 20356 65278
rect 20300 65174 20356 65212
rect 20412 65044 20468 65660
rect 20524 65490 20580 65502
rect 20524 65438 20526 65490
rect 20578 65438 20580 65490
rect 20524 65156 20580 65438
rect 20748 65156 20804 66108
rect 20860 65716 20916 68572
rect 20972 67284 21028 73892
rect 21308 73892 21476 73948
rect 23436 73892 23604 73948
rect 23884 77756 24388 77812
rect 25228 78484 25284 78494
rect 25228 77812 25284 78428
rect 25340 78260 25396 78270
rect 25396 78204 25732 78260
rect 25340 78166 25396 78204
rect 25228 77756 25396 77812
rect 20972 67218 21028 67228
rect 21196 71762 21252 71774
rect 21196 71710 21198 71762
rect 21250 71710 21252 71762
rect 21196 71652 21252 71710
rect 20972 67060 21028 67070
rect 21196 67060 21252 71596
rect 20972 67058 21252 67060
rect 20972 67006 20974 67058
rect 21026 67006 21252 67058
rect 20972 67004 21252 67006
rect 20972 66994 21028 67004
rect 21308 66388 21364 73892
rect 21532 73556 21588 73566
rect 21532 72770 21588 73500
rect 21532 72718 21534 72770
rect 21586 72718 21588 72770
rect 21532 71202 21588 72718
rect 21756 73332 21812 73342
rect 21756 71986 21812 73276
rect 22876 73332 22932 73342
rect 22876 73238 22932 73276
rect 23436 73330 23492 73892
rect 23436 73278 23438 73330
rect 23490 73278 23492 73330
rect 21756 71934 21758 71986
rect 21810 71934 21812 71986
rect 21756 71922 21812 71934
rect 23436 73220 23492 73278
rect 22316 71874 22372 71886
rect 22316 71822 22318 71874
rect 22370 71822 22372 71874
rect 22316 71764 22372 71822
rect 22652 71876 22708 71886
rect 22652 71782 22708 71820
rect 21532 71150 21534 71202
rect 21586 71150 21588 71202
rect 21532 71138 21588 71150
rect 21980 71708 22372 71764
rect 21420 70980 21476 70990
rect 21420 70886 21476 70924
rect 21868 70756 21924 70766
rect 21980 70756 22036 71708
rect 23436 71652 23492 73164
rect 23884 73444 23940 77756
rect 24008 77644 25208 77654
rect 24064 77642 24112 77644
rect 24168 77642 24216 77644
rect 24076 77590 24112 77642
rect 24200 77590 24216 77642
rect 24064 77588 24112 77590
rect 24168 77588 24216 77590
rect 24272 77642 24320 77644
rect 24376 77642 24424 77644
rect 24480 77642 24528 77644
rect 24376 77590 24396 77642
rect 24480 77590 24520 77642
rect 24272 77588 24320 77590
rect 24376 77588 24424 77590
rect 24480 77588 24528 77590
rect 24584 77588 24632 77644
rect 24688 77642 24736 77644
rect 24792 77642 24840 77644
rect 24896 77642 24944 77644
rect 24696 77590 24736 77642
rect 24820 77590 24840 77642
rect 24688 77588 24736 77590
rect 24792 77588 24840 77590
rect 24896 77588 24944 77590
rect 25000 77642 25048 77644
rect 25104 77642 25152 77644
rect 25000 77590 25016 77642
rect 25104 77590 25140 77642
rect 25000 77588 25048 77590
rect 25104 77588 25152 77590
rect 24008 77578 25208 77588
rect 24780 77364 24836 77374
rect 24220 77252 24276 77262
rect 24220 77158 24276 77196
rect 24780 77250 24836 77308
rect 24780 77198 24782 77250
rect 24834 77198 24836 77250
rect 24780 77186 24836 77198
rect 25228 77252 25284 77262
rect 25340 77252 25396 77756
rect 25676 77364 25732 78204
rect 25676 77270 25732 77308
rect 25228 77250 25396 77252
rect 25228 77198 25230 77250
rect 25282 77198 25396 77250
rect 25228 77196 25396 77198
rect 25228 77186 25284 77196
rect 24008 76076 25208 76086
rect 24064 76074 24112 76076
rect 24168 76074 24216 76076
rect 24076 76022 24112 76074
rect 24200 76022 24216 76074
rect 24064 76020 24112 76022
rect 24168 76020 24216 76022
rect 24272 76074 24320 76076
rect 24376 76074 24424 76076
rect 24480 76074 24528 76076
rect 24376 76022 24396 76074
rect 24480 76022 24520 76074
rect 24272 76020 24320 76022
rect 24376 76020 24424 76022
rect 24480 76020 24528 76022
rect 24584 76020 24632 76076
rect 24688 76074 24736 76076
rect 24792 76074 24840 76076
rect 24896 76074 24944 76076
rect 24696 76022 24736 76074
rect 24820 76022 24840 76074
rect 24688 76020 24736 76022
rect 24792 76020 24840 76022
rect 24896 76020 24944 76022
rect 25000 76074 25048 76076
rect 25104 76074 25152 76076
rect 25000 76022 25016 76074
rect 25104 76022 25140 76074
rect 25000 76020 25048 76022
rect 25104 76020 25152 76022
rect 24008 76010 25208 76020
rect 24008 74508 25208 74518
rect 24064 74506 24112 74508
rect 24168 74506 24216 74508
rect 24076 74454 24112 74506
rect 24200 74454 24216 74506
rect 24064 74452 24112 74454
rect 24168 74452 24216 74454
rect 24272 74506 24320 74508
rect 24376 74506 24424 74508
rect 24480 74506 24528 74508
rect 24376 74454 24396 74506
rect 24480 74454 24520 74506
rect 24272 74452 24320 74454
rect 24376 74452 24424 74454
rect 24480 74452 24528 74454
rect 24584 74452 24632 74508
rect 24688 74506 24736 74508
rect 24792 74506 24840 74508
rect 24896 74506 24944 74508
rect 24696 74454 24736 74506
rect 24820 74454 24840 74506
rect 24688 74452 24736 74454
rect 24792 74452 24840 74454
rect 24896 74452 24944 74454
rect 25000 74506 25048 74508
rect 25104 74506 25152 74508
rect 25000 74454 25016 74506
rect 25104 74454 25140 74506
rect 25000 74452 25048 74454
rect 25104 74452 25152 74454
rect 24008 74442 25208 74452
rect 23884 73218 23940 73388
rect 23884 73166 23886 73218
rect 23938 73166 23940 73218
rect 21868 70754 22036 70756
rect 21868 70702 21870 70754
rect 21922 70702 22036 70754
rect 21868 70700 22036 70702
rect 22092 71538 22148 71550
rect 22092 71486 22094 71538
rect 22146 71486 22148 71538
rect 21420 68180 21476 68190
rect 21420 68066 21476 68124
rect 21420 68014 21422 68066
rect 21474 68014 21476 68066
rect 21420 68002 21476 68014
rect 21532 67620 21588 67630
rect 21588 67564 21812 67620
rect 21532 67554 21588 67564
rect 21532 67172 21588 67182
rect 21420 67058 21476 67070
rect 21420 67006 21422 67058
rect 21474 67006 21476 67058
rect 21420 66498 21476 67006
rect 21420 66446 21422 66498
rect 21474 66446 21476 66498
rect 21420 66434 21476 66446
rect 21196 66332 21364 66388
rect 20972 65716 21028 65726
rect 20860 65714 21028 65716
rect 20860 65662 20974 65714
rect 21026 65662 21028 65714
rect 20860 65660 21028 65662
rect 20972 65650 21028 65660
rect 20860 65490 20916 65502
rect 20860 65438 20862 65490
rect 20914 65438 20916 65490
rect 20860 65380 20916 65438
rect 21196 65492 21252 66332
rect 21196 65426 21252 65436
rect 21308 66164 21364 66174
rect 21308 65490 21364 66108
rect 21308 65438 21310 65490
rect 21362 65438 21364 65490
rect 21308 65426 21364 65438
rect 21532 65716 21588 67116
rect 21756 66498 21812 67564
rect 21756 66446 21758 66498
rect 21810 66446 21812 66498
rect 21756 66434 21812 66446
rect 21868 66164 21924 70700
rect 21980 66164 22036 66174
rect 21868 66162 22036 66164
rect 21868 66110 21982 66162
rect 22034 66110 22036 66162
rect 21868 66108 22036 66110
rect 21532 65490 21588 65660
rect 21532 65438 21534 65490
rect 21586 65438 21588 65490
rect 21532 65426 21588 65438
rect 20860 65314 20916 65324
rect 21980 65378 22036 66108
rect 21980 65326 21982 65378
rect 22034 65326 22036 65378
rect 21084 65268 21140 65278
rect 21084 65174 21140 65212
rect 20748 65100 20916 65156
rect 20524 65090 20580 65100
rect 20300 64988 20468 65044
rect 20300 64818 20356 64988
rect 20300 64766 20302 64818
rect 20354 64766 20356 64818
rect 20300 64754 20356 64766
rect 20188 63476 20244 64652
rect 20412 63924 20468 63934
rect 20412 63830 20468 63868
rect 20188 63420 20468 63476
rect 20300 63140 20356 63150
rect 19964 63138 20132 63140
rect 19964 63086 20078 63138
rect 20130 63086 20132 63138
rect 19964 63084 20132 63086
rect 19852 63026 19908 63038
rect 19852 62974 19854 63026
rect 19906 62974 19908 63026
rect 19852 62692 19908 62974
rect 19852 62626 19908 62636
rect 19740 62302 19742 62354
rect 19794 62302 19796 62354
rect 19740 62290 19796 62302
rect 19852 62356 19908 62366
rect 19964 62356 20020 63084
rect 20076 63074 20132 63084
rect 20188 63138 20356 63140
rect 20188 63086 20302 63138
rect 20354 63086 20356 63138
rect 20188 63084 20356 63086
rect 19852 62354 20020 62356
rect 19852 62302 19854 62354
rect 19906 62302 20020 62354
rect 19852 62300 20020 62302
rect 20076 62916 20132 62926
rect 20076 62354 20132 62860
rect 20188 62578 20244 63084
rect 20300 63074 20356 63084
rect 20188 62526 20190 62578
rect 20242 62526 20244 62578
rect 20188 62514 20244 62526
rect 20300 62804 20356 62814
rect 20412 62804 20468 63420
rect 20356 62748 20468 62804
rect 20524 63138 20580 63150
rect 20524 63086 20526 63138
rect 20578 63086 20580 63138
rect 20300 62468 20356 62748
rect 20076 62302 20078 62354
rect 20130 62302 20132 62354
rect 19852 62290 19908 62300
rect 20076 62290 20132 62302
rect 20188 62356 20244 62366
rect 20188 61570 20244 62300
rect 20300 62354 20356 62412
rect 20524 62468 20580 63086
rect 20636 63028 20692 63038
rect 20636 62934 20692 62972
rect 20748 63026 20804 63038
rect 20748 62974 20750 63026
rect 20802 62974 20804 63026
rect 20748 62804 20804 62974
rect 20748 62738 20804 62748
rect 20524 62402 20580 62412
rect 20300 62302 20302 62354
rect 20354 62302 20356 62354
rect 20300 62290 20356 62302
rect 20860 62188 20916 65100
rect 20188 61518 20190 61570
rect 20242 61518 20244 61570
rect 20188 61506 20244 61518
rect 20636 62132 20916 62188
rect 20972 62354 21028 62366
rect 20972 62302 20974 62354
rect 21026 62302 21028 62354
rect 19628 60062 19630 60114
rect 19682 60062 19684 60114
rect 19628 59220 19684 60062
rect 20524 60116 20580 60126
rect 20636 60116 20692 62132
rect 20860 61572 20916 61582
rect 20972 61572 21028 62302
rect 21532 62354 21588 62366
rect 21532 62302 21534 62354
rect 21586 62302 21588 62354
rect 21420 61796 21476 61806
rect 21532 61796 21588 62302
rect 21420 61794 21588 61796
rect 21420 61742 21422 61794
rect 21474 61742 21588 61794
rect 21420 61740 21588 61742
rect 21420 61730 21476 61740
rect 21756 61572 21812 61582
rect 20860 61570 21028 61572
rect 20860 61518 20862 61570
rect 20914 61518 21028 61570
rect 20860 61516 21028 61518
rect 20860 61506 20916 61516
rect 20972 60676 21028 61516
rect 21532 61570 21812 61572
rect 21532 61518 21758 61570
rect 21810 61518 21812 61570
rect 21532 61516 21812 61518
rect 21420 61348 21476 61358
rect 21420 61010 21476 61292
rect 21420 60958 21422 61010
rect 21474 60958 21476 61010
rect 21420 60946 21476 60958
rect 20972 60674 21140 60676
rect 20972 60622 20974 60674
rect 21026 60622 21140 60674
rect 20972 60620 21140 60622
rect 20972 60610 21028 60620
rect 20860 60564 20916 60574
rect 20580 60060 20692 60116
rect 20524 60022 20580 60060
rect 20188 59778 20244 59790
rect 20188 59726 20190 59778
rect 20242 59726 20244 59778
rect 19740 59556 19796 59566
rect 19740 59442 19796 59500
rect 20188 59556 20244 59726
rect 19740 59390 19742 59442
rect 19794 59390 19796 59442
rect 19740 59378 19796 59390
rect 19852 59444 19908 59454
rect 19852 59350 19908 59388
rect 19628 59164 19908 59220
rect 19516 59108 19572 59118
rect 19516 59014 19572 59052
rect 19852 58828 19908 59164
rect 19404 58772 19684 58828
rect 19628 58660 19684 58772
rect 19740 58772 19908 58828
rect 19964 59218 20020 59230
rect 19964 59166 19966 59218
rect 20018 59166 20020 59218
rect 19740 58706 19796 58716
rect 19628 58594 19684 58604
rect 19404 58548 19460 58558
rect 19068 57820 19236 57876
rect 19292 58434 19348 58446
rect 19292 58382 19294 58434
rect 19346 58382 19348 58434
rect 19292 57874 19348 58382
rect 19404 58100 19460 58492
rect 19516 58434 19572 58446
rect 19516 58382 19518 58434
rect 19570 58382 19572 58434
rect 19516 58324 19572 58382
rect 19852 58436 19908 58446
rect 19964 58436 20020 59166
rect 20188 58996 20244 59500
rect 20636 59442 20692 60060
rect 20636 59390 20638 59442
rect 20690 59390 20692 59442
rect 20636 59378 20692 59390
rect 20748 60562 20916 60564
rect 20748 60510 20862 60562
rect 20914 60510 20916 60562
rect 20748 60508 20916 60510
rect 20748 59442 20804 60508
rect 20860 60498 20916 60508
rect 20748 59390 20750 59442
rect 20802 59390 20804 59442
rect 20748 59378 20804 59390
rect 20188 58930 20244 58940
rect 20412 59218 20468 59230
rect 20412 59166 20414 59218
rect 20466 59166 20468 59218
rect 20300 58436 20356 58446
rect 19908 58380 20020 58436
rect 20188 58380 20300 58436
rect 19852 58342 19908 58380
rect 20076 58324 20132 58334
rect 19516 58268 19796 58324
rect 19740 58212 19796 58268
rect 19964 58322 20132 58324
rect 19964 58270 20078 58322
rect 20130 58270 20132 58322
rect 19964 58268 20132 58270
rect 19964 58212 20020 58268
rect 20076 58258 20132 58268
rect 20188 58322 20244 58380
rect 20188 58270 20190 58322
rect 20242 58270 20244 58322
rect 20188 58258 20244 58270
rect 19740 58156 20020 58212
rect 19404 58044 19572 58100
rect 19292 57822 19294 57874
rect 19346 57822 19348 57874
rect 18620 57586 18676 57596
rect 18844 57762 18900 57774
rect 18844 57710 18846 57762
rect 18898 57710 18900 57762
rect 18508 57428 18564 57438
rect 18396 57426 18564 57428
rect 18396 57374 18510 57426
rect 18562 57374 18564 57426
rect 18396 57372 18564 57374
rect 18508 57362 18564 57372
rect 18620 57428 18676 57438
rect 18620 56866 18676 57372
rect 18620 56814 18622 56866
rect 18674 56814 18676 56866
rect 18620 56802 18676 56814
rect 18508 56308 18564 56318
rect 18508 56214 18564 56252
rect 18844 56196 18900 57710
rect 18620 56140 18900 56196
rect 18956 56308 19012 56318
rect 18396 55188 18452 55198
rect 18396 55094 18452 55132
rect 18284 54796 18452 54852
rect 18284 54514 18340 54526
rect 18284 54462 18286 54514
rect 18338 54462 18340 54514
rect 18172 54180 18228 54190
rect 18172 53842 18228 54124
rect 18284 54068 18340 54462
rect 18284 54002 18340 54012
rect 18172 53790 18174 53842
rect 18226 53790 18228 53842
rect 18172 53778 18228 53790
rect 18284 53730 18340 53742
rect 18284 53678 18286 53730
rect 18338 53678 18340 53730
rect 18284 53060 18340 53678
rect 18284 51378 18340 53004
rect 18284 51326 18286 51378
rect 18338 51326 18340 51378
rect 18284 51314 18340 51326
rect 17612 51268 17668 51278
rect 17612 51154 17668 51212
rect 17836 51268 17892 51278
rect 18172 51268 18228 51278
rect 17836 51266 18116 51268
rect 17836 51214 17838 51266
rect 17890 51214 18116 51266
rect 17836 51212 18116 51214
rect 17836 51202 17892 51212
rect 17612 51102 17614 51154
rect 17666 51102 17668 51154
rect 17612 51090 17668 51102
rect 17500 50372 18004 50428
rect 16604 49870 16606 49922
rect 16658 49870 16660 49922
rect 16604 49858 16660 49870
rect 16492 49812 16548 49822
rect 16492 49138 16548 49756
rect 17948 49810 18004 50372
rect 18060 49922 18116 51212
rect 18172 51174 18228 51212
rect 18172 50594 18228 50606
rect 18172 50542 18174 50594
rect 18226 50542 18228 50594
rect 18172 50034 18228 50542
rect 18396 50428 18452 54796
rect 18620 53954 18676 56140
rect 18844 55970 18900 55982
rect 18844 55918 18846 55970
rect 18898 55918 18900 55970
rect 18844 55300 18900 55918
rect 18844 55234 18900 55244
rect 18956 55298 19012 56252
rect 18956 55246 18958 55298
rect 19010 55246 19012 55298
rect 18956 55234 19012 55246
rect 18732 55188 18788 55198
rect 18732 55094 18788 55132
rect 18844 55074 18900 55086
rect 18844 55022 18846 55074
rect 18898 55022 18900 55074
rect 18732 54516 18788 54526
rect 18844 54516 18900 55022
rect 18732 54514 18900 54516
rect 18732 54462 18734 54514
rect 18786 54462 18900 54514
rect 18732 54460 18900 54462
rect 18732 54450 18788 54460
rect 18620 53902 18622 53954
rect 18674 53902 18676 53954
rect 18620 53890 18676 53902
rect 18956 53620 19012 53630
rect 18956 53170 19012 53564
rect 18956 53118 18958 53170
rect 19010 53118 19012 53170
rect 18956 52836 19012 53118
rect 18956 52770 19012 52780
rect 18620 50708 18676 50718
rect 19068 50708 19124 57820
rect 19292 57810 19348 57822
rect 19180 57650 19236 57662
rect 19180 57598 19182 57650
rect 19234 57598 19236 57650
rect 19180 57540 19236 57598
rect 19404 57652 19460 57662
rect 19404 57558 19460 57596
rect 19516 57540 19572 58044
rect 19964 57764 20020 58156
rect 20300 57764 20356 58380
rect 20412 58434 20468 59166
rect 20412 58382 20414 58434
rect 20466 58382 20468 58434
rect 20412 58370 20468 58382
rect 20524 59220 20580 59230
rect 20524 57876 20580 59164
rect 20860 59218 20916 59230
rect 20860 59166 20862 59218
rect 20914 59166 20916 59218
rect 20636 59108 20692 59118
rect 20636 58210 20692 59052
rect 20748 58996 20804 59006
rect 20748 58434 20804 58940
rect 20860 58884 20916 59166
rect 20860 58818 20916 58828
rect 20748 58382 20750 58434
rect 20802 58382 20804 58434
rect 20748 58370 20804 58382
rect 20636 58158 20638 58210
rect 20690 58158 20692 58210
rect 20636 58100 20692 58158
rect 20636 58044 20916 58100
rect 20636 57876 20692 57886
rect 20524 57874 20692 57876
rect 20524 57822 20638 57874
rect 20690 57822 20692 57874
rect 20524 57820 20692 57822
rect 20636 57810 20692 57820
rect 20300 57708 20468 57764
rect 19740 57650 19796 57662
rect 19740 57598 19742 57650
rect 19794 57598 19796 57650
rect 19516 57484 19684 57540
rect 19180 57474 19236 57484
rect 19516 56866 19572 56878
rect 19516 56814 19518 56866
rect 19570 56814 19572 56866
rect 19516 55300 19572 56814
rect 19628 56642 19684 57484
rect 19740 57428 19796 57598
rect 19740 57362 19796 57372
rect 19740 56756 19796 56766
rect 19740 56662 19796 56700
rect 19628 56590 19630 56642
rect 19682 56590 19684 56642
rect 19628 56578 19684 56590
rect 19852 56420 19908 56430
rect 19964 56420 20020 57708
rect 19908 56364 20020 56420
rect 20076 57650 20132 57662
rect 20076 57598 20078 57650
rect 20130 57598 20132 57650
rect 19852 56354 19908 56364
rect 20076 56308 20132 57598
rect 20300 57428 20356 57438
rect 20076 56242 20132 56252
rect 20188 57426 20356 57428
rect 20188 57374 20302 57426
rect 20354 57374 20356 57426
rect 20188 57372 20356 57374
rect 19516 55234 19572 55244
rect 19292 55186 19348 55198
rect 19292 55134 19294 55186
rect 19346 55134 19348 55186
rect 19292 53954 19348 55134
rect 19292 53902 19294 53954
rect 19346 53902 19348 53954
rect 19292 53890 19348 53902
rect 19628 55188 19684 55198
rect 19628 53956 19684 55132
rect 19628 53862 19684 53900
rect 19964 54068 20020 54078
rect 19404 53620 19460 53630
rect 19404 53526 19460 53564
rect 19852 52612 19908 52622
rect 19852 52274 19908 52556
rect 19852 52222 19854 52274
rect 19906 52222 19908 52274
rect 19852 52210 19908 52222
rect 19964 52164 20020 54012
rect 20076 53956 20132 53966
rect 20076 53842 20132 53900
rect 20076 53790 20078 53842
rect 20130 53790 20132 53842
rect 20076 53778 20132 53790
rect 20188 53844 20244 57372
rect 20300 57362 20356 57372
rect 20300 57204 20356 57214
rect 20300 56754 20356 57148
rect 20412 56866 20468 57708
rect 20748 57652 20804 57662
rect 20524 57540 20580 57550
rect 20524 57446 20580 57484
rect 20748 56980 20804 57596
rect 20412 56814 20414 56866
rect 20466 56814 20468 56866
rect 20412 56802 20468 56814
rect 20636 56924 20804 56980
rect 20300 56702 20302 56754
rect 20354 56702 20356 56754
rect 20300 56690 20356 56702
rect 20636 56306 20692 56924
rect 20636 56254 20638 56306
rect 20690 56254 20692 56306
rect 20636 56242 20692 56254
rect 20748 56196 20804 56206
rect 20748 56102 20804 56140
rect 20300 56084 20356 56094
rect 20300 55188 20356 56028
rect 20860 55972 20916 58044
rect 20860 55906 20916 55916
rect 21084 57650 21140 60620
rect 21532 60562 21588 61516
rect 21756 61506 21812 61516
rect 21980 61458 22036 65326
rect 21980 61406 21982 61458
rect 22034 61406 22036 61458
rect 21980 61348 22036 61406
rect 21980 61282 22036 61292
rect 21532 60510 21534 60562
rect 21586 60510 21588 60562
rect 21532 60498 21588 60510
rect 21532 59778 21588 59790
rect 21532 59726 21534 59778
rect 21586 59726 21588 59778
rect 21308 59218 21364 59230
rect 21308 59166 21310 59218
rect 21362 59166 21364 59218
rect 21308 58996 21364 59166
rect 21532 59220 21588 59726
rect 22092 59444 22148 71486
rect 22316 71202 22372 71214
rect 22316 71150 22318 71202
rect 22370 71150 22372 71202
rect 22316 71090 22372 71150
rect 22316 71038 22318 71090
rect 22370 71038 22372 71090
rect 22316 71026 22372 71038
rect 22204 70532 22260 70542
rect 23436 70532 23492 71596
rect 23548 72548 23604 72558
rect 23884 72548 23940 73166
rect 24332 73220 24388 73230
rect 24332 73126 24388 73164
rect 24008 72940 25208 72950
rect 24064 72938 24112 72940
rect 24168 72938 24216 72940
rect 24076 72886 24112 72938
rect 24200 72886 24216 72938
rect 24064 72884 24112 72886
rect 24168 72884 24216 72886
rect 24272 72938 24320 72940
rect 24376 72938 24424 72940
rect 24480 72938 24528 72940
rect 24376 72886 24396 72938
rect 24480 72886 24520 72938
rect 24272 72884 24320 72886
rect 24376 72884 24424 72886
rect 24480 72884 24528 72886
rect 24584 72884 24632 72940
rect 24688 72938 24736 72940
rect 24792 72938 24840 72940
rect 24896 72938 24944 72940
rect 24696 72886 24736 72938
rect 24820 72886 24840 72938
rect 24688 72884 24736 72886
rect 24792 72884 24840 72886
rect 24896 72884 24944 72886
rect 25000 72938 25048 72940
rect 25104 72938 25152 72940
rect 25000 72886 25016 72938
rect 25104 72886 25140 72938
rect 25000 72884 25048 72886
rect 25104 72884 25152 72886
rect 24008 72874 25208 72884
rect 23548 72546 23940 72548
rect 23548 72494 23550 72546
rect 23602 72494 23940 72546
rect 23548 72492 23940 72494
rect 23548 72324 23604 72492
rect 23548 70756 23604 72268
rect 24332 72324 24388 72334
rect 24332 72230 24388 72268
rect 27804 71764 27860 71774
rect 27468 71762 27860 71764
rect 27468 71710 27806 71762
rect 27858 71710 27860 71762
rect 27468 71708 27860 71710
rect 27468 71652 27524 71708
rect 27804 71698 27860 71708
rect 27356 71650 27524 71652
rect 27356 71598 27470 71650
rect 27522 71598 27524 71650
rect 27356 71596 27524 71598
rect 24008 71372 25208 71382
rect 24064 71370 24112 71372
rect 24168 71370 24216 71372
rect 24076 71318 24112 71370
rect 24200 71318 24216 71370
rect 24064 71316 24112 71318
rect 24168 71316 24216 71318
rect 24272 71370 24320 71372
rect 24376 71370 24424 71372
rect 24480 71370 24528 71372
rect 24376 71318 24396 71370
rect 24480 71318 24520 71370
rect 24272 71316 24320 71318
rect 24376 71316 24424 71318
rect 24480 71316 24528 71318
rect 24584 71316 24632 71372
rect 24688 71370 24736 71372
rect 24792 71370 24840 71372
rect 24896 71370 24944 71372
rect 24696 71318 24736 71370
rect 24820 71318 24840 71370
rect 24688 71316 24736 71318
rect 24792 71316 24840 71318
rect 24896 71316 24944 71318
rect 25000 71370 25048 71372
rect 25104 71370 25152 71372
rect 25000 71318 25016 71370
rect 25104 71318 25140 71370
rect 25000 71316 25048 71318
rect 25104 71316 25152 71318
rect 24008 71306 25208 71316
rect 25676 71090 25732 71102
rect 25676 71038 25678 71090
rect 25730 71038 25732 71090
rect 24220 70980 24276 70990
rect 24220 70886 24276 70924
rect 25116 70980 25172 70990
rect 25116 70886 25172 70924
rect 23548 70690 23604 70700
rect 23884 70532 23940 70542
rect 23436 70476 23884 70532
rect 22204 67730 22260 70476
rect 22204 67678 22206 67730
rect 22258 67678 22260 67730
rect 22204 67666 22260 67678
rect 23772 70084 23828 70094
rect 23772 68628 23828 70028
rect 23884 69410 23940 70476
rect 25676 70532 25732 71038
rect 27356 70980 27412 71596
rect 27468 71586 27524 71596
rect 25732 70476 25956 70532
rect 25676 70466 25732 70476
rect 25116 70194 25172 70206
rect 25116 70142 25118 70194
rect 25170 70142 25172 70194
rect 24668 70084 24724 70094
rect 24668 69990 24724 70028
rect 25116 70084 25172 70142
rect 25564 70196 25620 70206
rect 25564 70102 25620 70140
rect 25788 70194 25844 70206
rect 25788 70142 25790 70194
rect 25842 70142 25844 70194
rect 25116 70018 25172 70028
rect 25340 70082 25396 70094
rect 25340 70030 25342 70082
rect 25394 70030 25396 70082
rect 24008 69804 25208 69814
rect 24064 69802 24112 69804
rect 24168 69802 24216 69804
rect 24076 69750 24112 69802
rect 24200 69750 24216 69802
rect 24064 69748 24112 69750
rect 24168 69748 24216 69750
rect 24272 69802 24320 69804
rect 24376 69802 24424 69804
rect 24480 69802 24528 69804
rect 24376 69750 24396 69802
rect 24480 69750 24520 69802
rect 24272 69748 24320 69750
rect 24376 69748 24424 69750
rect 24480 69748 24528 69750
rect 24584 69748 24632 69804
rect 24688 69802 24736 69804
rect 24792 69802 24840 69804
rect 24896 69802 24944 69804
rect 24696 69750 24736 69802
rect 24820 69750 24840 69802
rect 24688 69748 24736 69750
rect 24792 69748 24840 69750
rect 24896 69748 24944 69750
rect 25000 69802 25048 69804
rect 25104 69802 25152 69804
rect 25000 69750 25016 69802
rect 25104 69750 25140 69802
rect 25000 69748 25048 69750
rect 25104 69748 25152 69750
rect 24008 69738 25208 69748
rect 23884 69358 23886 69410
rect 23938 69358 23940 69410
rect 23884 69346 23940 69358
rect 24556 69636 24612 69646
rect 24556 69410 24612 69580
rect 25340 69636 25396 70030
rect 25340 69570 25396 69580
rect 24556 69358 24558 69410
rect 24610 69358 24612 69410
rect 24556 69346 24612 69358
rect 25788 68964 25844 70142
rect 25452 68908 25844 68964
rect 25900 69524 25956 70476
rect 27020 70420 27076 70430
rect 23996 68628 24052 68638
rect 23772 68626 24052 68628
rect 23772 68574 23774 68626
rect 23826 68574 23998 68626
rect 24050 68574 24052 68626
rect 23772 68572 24052 68574
rect 23772 66948 23828 68572
rect 23996 68562 24052 68572
rect 24220 68628 24276 68638
rect 24220 68534 24276 68572
rect 24444 68626 24500 68638
rect 24444 68574 24446 68626
rect 24498 68574 24500 68626
rect 24444 68404 24500 68574
rect 24668 68626 24724 68638
rect 24668 68574 24670 68626
rect 24722 68574 24724 68626
rect 24668 68516 24724 68574
rect 24668 68450 24724 68460
rect 25340 68626 25396 68638
rect 25340 68574 25342 68626
rect 25394 68574 25396 68626
rect 24444 68338 24500 68348
rect 24008 68236 25208 68246
rect 24064 68234 24112 68236
rect 24168 68234 24216 68236
rect 24076 68182 24112 68234
rect 24200 68182 24216 68234
rect 24064 68180 24112 68182
rect 24168 68180 24216 68182
rect 24272 68234 24320 68236
rect 24376 68234 24424 68236
rect 24480 68234 24528 68236
rect 24376 68182 24396 68234
rect 24480 68182 24520 68234
rect 24272 68180 24320 68182
rect 24376 68180 24424 68182
rect 24480 68180 24528 68182
rect 24584 68180 24632 68236
rect 24688 68234 24736 68236
rect 24792 68234 24840 68236
rect 24896 68234 24944 68236
rect 24696 68182 24736 68234
rect 24820 68182 24840 68234
rect 24688 68180 24736 68182
rect 24792 68180 24840 68182
rect 24896 68180 24944 68182
rect 25000 68234 25048 68236
rect 25104 68234 25152 68236
rect 25000 68182 25016 68234
rect 25104 68182 25140 68234
rect 25000 68180 25048 68182
rect 25104 68180 25152 68182
rect 24008 68170 25208 68180
rect 24444 68068 24500 68078
rect 24444 67842 24500 68012
rect 24444 67790 24446 67842
rect 24498 67790 24500 67842
rect 24444 67778 24500 67790
rect 25116 67844 25172 67854
rect 25340 67844 25396 68574
rect 25116 67842 25396 67844
rect 25116 67790 25118 67842
rect 25170 67790 25396 67842
rect 25116 67788 25396 67790
rect 25116 67778 25172 67788
rect 23772 66882 23828 66892
rect 23884 67282 23940 67294
rect 23884 67230 23886 67282
rect 23938 67230 23940 67282
rect 22540 66836 22596 66846
rect 22540 66164 22596 66780
rect 22540 66070 22596 66108
rect 23884 66052 23940 67230
rect 25340 67284 25396 67788
rect 25452 67620 25508 68908
rect 25564 68740 25620 68750
rect 25564 67842 25620 68684
rect 25676 68628 25732 68638
rect 25676 68534 25732 68572
rect 25564 67790 25566 67842
rect 25618 67790 25620 67842
rect 25564 67778 25620 67790
rect 25452 67564 25620 67620
rect 25228 66948 25284 66958
rect 24444 66836 24500 66874
rect 25228 66854 25284 66892
rect 24444 66770 24500 66780
rect 24008 66668 25208 66678
rect 24064 66666 24112 66668
rect 24168 66666 24216 66668
rect 24076 66614 24112 66666
rect 24200 66614 24216 66666
rect 24064 66612 24112 66614
rect 24168 66612 24216 66614
rect 24272 66666 24320 66668
rect 24376 66666 24424 66668
rect 24480 66666 24528 66668
rect 24376 66614 24396 66666
rect 24480 66614 24520 66666
rect 24272 66612 24320 66614
rect 24376 66612 24424 66614
rect 24480 66612 24528 66614
rect 24584 66612 24632 66668
rect 24688 66666 24736 66668
rect 24792 66666 24840 66668
rect 24896 66666 24944 66668
rect 24696 66614 24736 66666
rect 24820 66614 24840 66666
rect 24688 66612 24736 66614
rect 24792 66612 24840 66614
rect 24896 66612 24944 66614
rect 25000 66666 25048 66668
rect 25104 66666 25152 66668
rect 25000 66614 25016 66666
rect 25104 66614 25140 66666
rect 25000 66612 25048 66614
rect 25104 66612 25152 66614
rect 24008 66602 25208 66612
rect 23436 63140 23492 63150
rect 23772 63140 23828 63150
rect 22316 62468 22372 62478
rect 22316 61458 22372 62412
rect 22316 61406 22318 61458
rect 22370 61406 22372 61458
rect 22316 61394 22372 61406
rect 22092 59378 22148 59388
rect 23436 59780 23492 63084
rect 21644 59332 21700 59342
rect 21644 59330 21812 59332
rect 21644 59278 21646 59330
rect 21698 59278 21812 59330
rect 21644 59276 21812 59278
rect 21644 59266 21700 59276
rect 21532 59126 21588 59164
rect 21756 59108 21812 59276
rect 21644 58996 21700 59006
rect 21308 58994 21700 58996
rect 21308 58942 21646 58994
rect 21698 58942 21700 58994
rect 21308 58940 21700 58942
rect 21644 58930 21700 58940
rect 21084 57598 21086 57650
rect 21138 57598 21140 57650
rect 20300 55122 20356 55132
rect 21084 55188 21140 57598
rect 21308 58434 21364 58446
rect 21308 58382 21310 58434
rect 21362 58382 21364 58434
rect 21308 56754 21364 58382
rect 21644 58436 21700 58474
rect 21644 58370 21700 58380
rect 21644 58210 21700 58222
rect 21644 58158 21646 58210
rect 21698 58158 21700 58210
rect 21532 57652 21588 57662
rect 21532 57092 21588 57596
rect 21644 57650 21700 58158
rect 21644 57598 21646 57650
rect 21698 57598 21700 57650
rect 21644 57586 21700 57598
rect 21532 57036 21700 57092
rect 21308 56702 21310 56754
rect 21362 56702 21364 56754
rect 21308 56084 21364 56702
rect 21532 56868 21588 56878
rect 21532 56642 21588 56812
rect 21644 56866 21700 57036
rect 21644 56814 21646 56866
rect 21698 56814 21700 56866
rect 21644 56802 21700 56814
rect 21532 56590 21534 56642
rect 21586 56590 21588 56642
rect 21532 56578 21588 56590
rect 21756 56196 21812 59052
rect 22204 59108 22260 59118
rect 22204 59014 22260 59052
rect 23436 58996 23492 59724
rect 23212 58940 23492 58996
rect 23548 63084 23772 63140
rect 21980 58322 22036 58334
rect 21980 58270 21982 58322
rect 22034 58270 22036 58322
rect 21532 56140 21812 56196
rect 21868 56754 21924 56766
rect 21868 56702 21870 56754
rect 21922 56702 21924 56754
rect 21420 56084 21476 56094
rect 21308 56028 21420 56084
rect 21420 55990 21476 56028
rect 21084 55122 21140 55132
rect 21196 54740 21252 54750
rect 21196 54646 21252 54684
rect 20188 53778 20244 53788
rect 21532 53956 21588 56140
rect 21644 55972 21700 55982
rect 21644 55410 21700 55916
rect 21868 55522 21924 56702
rect 21980 55970 22036 58270
rect 22540 58212 22596 58222
rect 22428 58210 22596 58212
rect 22428 58158 22542 58210
rect 22594 58158 22596 58210
rect 22428 58156 22596 58158
rect 22092 56644 22148 56654
rect 22092 56642 22260 56644
rect 22092 56590 22094 56642
rect 22146 56590 22260 56642
rect 22092 56588 22260 56590
rect 22092 56578 22148 56588
rect 21980 55918 21982 55970
rect 22034 55918 22036 55970
rect 21980 55906 22036 55918
rect 22092 56194 22148 56206
rect 22092 56142 22094 56194
rect 22146 56142 22148 56194
rect 22092 55972 22148 56142
rect 22204 56196 22260 56588
rect 22204 56130 22260 56140
rect 22428 56196 22484 58156
rect 22540 58146 22596 58156
rect 22876 56756 22932 56766
rect 23100 56756 23156 56766
rect 22876 56754 23100 56756
rect 22876 56702 22878 56754
rect 22930 56702 23100 56754
rect 22876 56700 23100 56702
rect 22764 56308 22820 56318
rect 22092 55906 22148 55916
rect 22316 56084 22372 56094
rect 22428 56084 22484 56140
rect 22372 56028 22484 56084
rect 22540 56252 22764 56308
rect 22316 55524 22372 56028
rect 21868 55470 21870 55522
rect 21922 55470 21924 55522
rect 21868 55458 21924 55470
rect 22092 55468 22372 55524
rect 21644 55358 21646 55410
rect 21698 55358 21700 55410
rect 21644 55346 21700 55358
rect 22092 55410 22148 55468
rect 22092 55358 22094 55410
rect 22146 55358 22148 55410
rect 22092 55346 22148 55358
rect 21756 55300 21812 55310
rect 21756 54738 21812 55244
rect 21756 54686 21758 54738
rect 21810 54686 21812 54738
rect 21756 54674 21812 54686
rect 22092 54740 22148 54750
rect 22092 54646 22148 54684
rect 21532 53900 21812 53956
rect 21532 53620 21588 53900
rect 21532 53554 21588 53564
rect 21644 53732 21700 53742
rect 21644 53170 21700 53676
rect 21644 53118 21646 53170
rect 21698 53118 21700 53170
rect 20972 52836 21028 52846
rect 20972 52834 21588 52836
rect 20972 52782 20974 52834
rect 21026 52782 21588 52834
rect 20972 52780 21588 52782
rect 20972 52770 21028 52780
rect 20412 52612 20468 52622
rect 19404 52052 19460 52062
rect 19404 51958 19460 51996
rect 19964 51378 20020 52108
rect 20300 52162 20356 52174
rect 20300 52110 20302 52162
rect 20354 52110 20356 52162
rect 19964 51326 19966 51378
rect 20018 51326 20020 51378
rect 19964 51314 20020 51326
rect 20188 52052 20244 52062
rect 19180 50708 19236 50718
rect 19068 50706 19236 50708
rect 19068 50654 19182 50706
rect 19234 50654 19236 50706
rect 19068 50652 19236 50654
rect 18620 50614 18676 50652
rect 19180 50642 19236 50652
rect 19852 50708 19908 50718
rect 19852 50614 19908 50652
rect 18172 49982 18174 50034
rect 18226 49982 18228 50034
rect 18172 49970 18228 49982
rect 18284 50372 18452 50428
rect 18844 50596 18900 50606
rect 18060 49870 18062 49922
rect 18114 49870 18116 49922
rect 18060 49858 18116 49870
rect 17948 49758 17950 49810
rect 18002 49758 18004 49810
rect 17948 49746 18004 49758
rect 16492 49086 16494 49138
rect 16546 49086 16548 49138
rect 16492 49074 16548 49086
rect 17500 49700 17556 49710
rect 17052 49028 17108 49038
rect 17500 49028 17556 49644
rect 17724 49028 17780 49038
rect 17500 49026 17780 49028
rect 17500 48974 17726 49026
rect 17778 48974 17780 49026
rect 17500 48972 17780 48974
rect 17052 48934 17108 48972
rect 16716 48804 16772 48814
rect 16716 48130 16772 48748
rect 17724 48804 17780 48972
rect 17948 48916 18004 48926
rect 17948 48822 18004 48860
rect 17724 48738 17780 48748
rect 18284 48356 18340 50372
rect 18844 49140 18900 50540
rect 19404 50594 19460 50606
rect 19404 50542 19406 50594
rect 19458 50542 19460 50594
rect 19292 50484 19348 50522
rect 19292 50418 19348 50428
rect 19404 50428 19460 50542
rect 19404 50372 19684 50428
rect 19516 49924 19572 49934
rect 19068 49922 19572 49924
rect 19068 49870 19518 49922
rect 19570 49870 19572 49922
rect 19068 49868 19572 49870
rect 18956 49812 19012 49822
rect 18956 49718 19012 49756
rect 18508 49084 18788 49140
rect 18396 49026 18452 49038
rect 18396 48974 18398 49026
rect 18450 48974 18452 49026
rect 18396 48804 18452 48974
rect 18508 49026 18564 49084
rect 18508 48974 18510 49026
rect 18562 48974 18564 49026
rect 18508 48962 18564 48974
rect 18620 48916 18676 48926
rect 18620 48822 18676 48860
rect 18396 48748 18564 48804
rect 18508 48692 18564 48748
rect 18508 48636 18676 48692
rect 18284 48300 18564 48356
rect 18508 48242 18564 48300
rect 18508 48190 18510 48242
rect 18562 48190 18564 48242
rect 16716 48078 16718 48130
rect 16770 48078 16772 48130
rect 16716 46564 16772 48078
rect 17836 48132 17892 48142
rect 18172 48132 18228 48142
rect 17836 48130 18228 48132
rect 17836 48078 17838 48130
rect 17890 48078 18174 48130
rect 18226 48078 18228 48130
rect 17836 48076 18228 48078
rect 17612 47460 17668 47470
rect 17612 47366 17668 47404
rect 17836 47068 17892 48076
rect 18172 48066 18228 48076
rect 16380 45826 16436 45836
rect 16492 46508 16772 46564
rect 17276 47012 17332 47022
rect 16492 45668 16548 46508
rect 17276 46114 17332 46956
rect 17612 47012 17892 47068
rect 18396 47012 18452 47022
rect 17500 46674 17556 46686
rect 17500 46622 17502 46674
rect 17554 46622 17556 46674
rect 17500 46564 17556 46622
rect 17612 46564 17668 47012
rect 17500 46508 17612 46564
rect 17612 46498 17668 46508
rect 18284 46788 18340 46798
rect 17276 46062 17278 46114
rect 17330 46062 17332 46114
rect 17276 46050 17332 46062
rect 16828 46004 16884 46014
rect 16716 46002 16884 46004
rect 16716 45950 16830 46002
rect 16882 45950 16884 46002
rect 16716 45948 16884 45950
rect 16604 45890 16660 45902
rect 16604 45838 16606 45890
rect 16658 45838 16660 45890
rect 16604 45780 16660 45838
rect 16604 45714 16660 45724
rect 16268 45612 16548 45668
rect 15932 45332 15988 45342
rect 15820 45220 15876 45230
rect 15820 44100 15876 45164
rect 15932 44994 15988 45276
rect 15932 44942 15934 44994
rect 15986 44942 15988 44994
rect 15932 44884 15988 44942
rect 15932 44818 15988 44828
rect 16268 44772 16324 45612
rect 16380 45332 16436 45342
rect 16604 45332 16660 45342
rect 16380 45238 16436 45276
rect 16492 45276 16604 45332
rect 16268 44716 16436 44772
rect 16268 44100 16324 44110
rect 15820 44098 16324 44100
rect 15820 44046 16270 44098
rect 16322 44046 16324 44098
rect 15820 44044 16324 44046
rect 15820 43762 15876 44044
rect 16268 44034 16324 44044
rect 16380 43876 16436 44716
rect 15820 43710 15822 43762
rect 15874 43710 15876 43762
rect 15820 39396 15876 43710
rect 16268 43820 16436 43876
rect 16156 43538 16212 43550
rect 16156 43486 16158 43538
rect 16210 43486 16212 43538
rect 16156 43316 16212 43486
rect 16044 43260 16156 43316
rect 16044 42866 16100 43260
rect 16156 43250 16212 43260
rect 16044 42814 16046 42866
rect 16098 42814 16100 42866
rect 16044 42802 16100 42814
rect 15932 40404 15988 40414
rect 15932 40310 15988 40348
rect 15820 39394 16100 39396
rect 15820 39342 15822 39394
rect 15874 39342 16100 39394
rect 15820 39340 16100 39342
rect 15820 39330 15876 39340
rect 15260 38612 15316 38622
rect 15708 38612 15876 38668
rect 13244 37202 13300 37212
rect 12908 36654 12910 36706
rect 12962 36654 12964 36706
rect 12572 36484 12628 36494
rect 12460 36260 12516 36270
rect 12572 36260 12628 36428
rect 12460 36258 12628 36260
rect 12460 36206 12462 36258
rect 12514 36206 12628 36258
rect 12460 36204 12628 36206
rect 12460 36194 12516 36204
rect 12460 35476 12516 35486
rect 12460 35138 12516 35420
rect 12460 35086 12462 35138
rect 12514 35086 12516 35138
rect 12460 35074 12516 35086
rect 12460 34804 12516 34814
rect 12460 34356 12516 34748
rect 12460 34290 12516 34300
rect 12460 30210 12516 30222
rect 12460 30158 12462 30210
rect 12514 30158 12516 30210
rect 12460 30100 12516 30158
rect 12460 30034 12516 30044
rect 12348 29586 12404 29596
rect 12460 29540 12516 29550
rect 12460 28418 12516 29484
rect 12460 28366 12462 28418
rect 12514 28366 12516 28418
rect 12460 28354 12516 28366
rect 12012 28030 12014 28082
rect 12066 28030 12068 28082
rect 12012 28018 12068 28030
rect 9772 27636 9828 27646
rect 9772 27542 9828 27580
rect 9772 27188 9828 27198
rect 9660 27186 9828 27188
rect 9660 27134 9774 27186
rect 9826 27134 9828 27186
rect 9660 27132 9828 27134
rect 9772 27122 9828 27132
rect 8876 25732 8932 27020
rect 9884 25732 9940 27692
rect 11564 27860 11620 27870
rect 11564 27746 11620 27804
rect 11564 27694 11566 27746
rect 11618 27694 11620 27746
rect 11564 27188 11620 27694
rect 12348 27748 12404 27758
rect 12348 27654 12404 27692
rect 12460 27524 12516 27534
rect 12572 27524 12628 36204
rect 12908 36260 12964 36654
rect 13580 36484 13636 38612
rect 15260 38050 15316 38556
rect 15260 37998 15262 38050
rect 15314 37998 15316 38050
rect 15260 37986 15316 37998
rect 15708 38050 15764 38062
rect 15708 37998 15710 38050
rect 15762 37998 15764 38050
rect 13692 37826 13748 37838
rect 13692 37774 13694 37826
rect 13746 37774 13748 37826
rect 13692 36932 13748 37774
rect 14008 37660 15208 37670
rect 14064 37658 14112 37660
rect 14168 37658 14216 37660
rect 14076 37606 14112 37658
rect 14200 37606 14216 37658
rect 14064 37604 14112 37606
rect 14168 37604 14216 37606
rect 14272 37658 14320 37660
rect 14376 37658 14424 37660
rect 14480 37658 14528 37660
rect 14376 37606 14396 37658
rect 14480 37606 14520 37658
rect 14272 37604 14320 37606
rect 14376 37604 14424 37606
rect 14480 37604 14528 37606
rect 14584 37604 14632 37660
rect 14688 37658 14736 37660
rect 14792 37658 14840 37660
rect 14896 37658 14944 37660
rect 14696 37606 14736 37658
rect 14820 37606 14840 37658
rect 14688 37604 14736 37606
rect 14792 37604 14840 37606
rect 14896 37604 14944 37606
rect 15000 37658 15048 37660
rect 15104 37658 15152 37660
rect 15000 37606 15016 37658
rect 15104 37606 15140 37658
rect 15000 37604 15048 37606
rect 15104 37604 15152 37606
rect 14008 37594 15208 37604
rect 14812 37492 14868 37502
rect 14812 37398 14868 37436
rect 15708 37492 15764 37998
rect 15708 37426 15764 37436
rect 14028 37380 14084 37390
rect 14028 37286 14084 37324
rect 13692 36866 13748 36876
rect 14252 37268 14308 37278
rect 14252 36594 14308 37212
rect 14252 36542 14254 36594
rect 14306 36542 14308 36594
rect 14252 36530 14308 36542
rect 15036 37266 15092 37278
rect 15036 37214 15038 37266
rect 15090 37214 15092 37266
rect 15036 36932 15092 37214
rect 13580 36390 13636 36428
rect 12908 36166 12964 36204
rect 13692 36370 13748 36382
rect 13692 36318 13694 36370
rect 13746 36318 13748 36370
rect 13692 36260 13748 36318
rect 14812 36372 14868 36382
rect 14812 36278 14868 36316
rect 15036 36260 15092 36876
rect 15036 36204 15428 36260
rect 13580 35812 13636 35822
rect 12796 35700 12852 35710
rect 12796 35138 12852 35644
rect 12796 35086 12798 35138
rect 12850 35086 12852 35138
rect 12796 35074 12852 35086
rect 13580 35138 13636 35756
rect 13580 35086 13582 35138
rect 13634 35086 13636 35138
rect 13580 35074 13636 35086
rect 13692 35028 13748 36204
rect 14008 36092 15208 36102
rect 14064 36090 14112 36092
rect 14168 36090 14216 36092
rect 14076 36038 14112 36090
rect 14200 36038 14216 36090
rect 14064 36036 14112 36038
rect 14168 36036 14216 36038
rect 14272 36090 14320 36092
rect 14376 36090 14424 36092
rect 14480 36090 14528 36092
rect 14376 36038 14396 36090
rect 14480 36038 14520 36090
rect 14272 36036 14320 36038
rect 14376 36036 14424 36038
rect 14480 36036 14528 36038
rect 14584 36036 14632 36092
rect 14688 36090 14736 36092
rect 14792 36090 14840 36092
rect 14896 36090 14944 36092
rect 14696 36038 14736 36090
rect 14820 36038 14840 36090
rect 14688 36036 14736 36038
rect 14792 36036 14840 36038
rect 14896 36036 14944 36038
rect 15000 36090 15048 36092
rect 15104 36090 15152 36092
rect 15000 36038 15016 36090
rect 15104 36038 15140 36090
rect 15000 36036 15048 36038
rect 15104 36036 15152 36038
rect 14008 36026 15208 36036
rect 14924 35812 14980 35822
rect 14924 35718 14980 35756
rect 14028 35700 14084 35710
rect 14028 35606 14084 35644
rect 14588 35700 14644 35710
rect 13692 34962 13748 34972
rect 14588 35140 14644 35644
rect 14700 35698 14756 35710
rect 14700 35646 14702 35698
rect 14754 35646 14756 35698
rect 14700 35252 14756 35646
rect 15148 35700 15204 35710
rect 15372 35700 15428 36204
rect 15204 35644 15428 35700
rect 15148 35606 15204 35644
rect 14700 35186 14756 35196
rect 15036 35252 15092 35262
rect 14588 35026 14644 35084
rect 14588 34974 14590 35026
rect 14642 34974 14644 35026
rect 14588 34962 14644 34974
rect 15036 35026 15092 35196
rect 15036 34974 15038 35026
rect 15090 34974 15092 35026
rect 15036 34962 15092 34974
rect 13468 34802 13524 34814
rect 13468 34750 13470 34802
rect 13522 34750 13524 34802
rect 13020 34580 13076 34590
rect 12908 34018 12964 34030
rect 12908 33966 12910 34018
rect 12962 33966 12964 34018
rect 12908 33908 12964 33966
rect 12908 33842 12964 33852
rect 12908 32564 12964 32574
rect 12908 32470 12964 32508
rect 12684 31892 12740 31902
rect 12684 31798 12740 31836
rect 13020 31780 13076 34524
rect 13468 33908 13524 34750
rect 13580 34690 13636 34702
rect 14140 34692 14196 34702
rect 13580 34638 13582 34690
rect 13634 34638 13636 34690
rect 13580 34580 13636 34638
rect 13580 34514 13636 34524
rect 13804 34690 14196 34692
rect 13804 34638 14142 34690
rect 14194 34638 14196 34690
rect 13804 34636 14196 34638
rect 13804 34580 13860 34636
rect 14140 34626 14196 34636
rect 13804 34514 13860 34524
rect 14008 34524 15208 34534
rect 14064 34522 14112 34524
rect 14168 34522 14216 34524
rect 14076 34470 14112 34522
rect 14200 34470 14216 34522
rect 14064 34468 14112 34470
rect 14168 34468 14216 34470
rect 14272 34522 14320 34524
rect 14376 34522 14424 34524
rect 14480 34522 14528 34524
rect 14376 34470 14396 34522
rect 14480 34470 14520 34522
rect 14272 34468 14320 34470
rect 14376 34468 14424 34470
rect 14480 34468 14528 34470
rect 14584 34468 14632 34524
rect 14688 34522 14736 34524
rect 14792 34522 14840 34524
rect 14896 34522 14944 34524
rect 14696 34470 14736 34522
rect 14820 34470 14840 34522
rect 14688 34468 14736 34470
rect 14792 34468 14840 34470
rect 14896 34468 14944 34470
rect 15000 34522 15048 34524
rect 15104 34522 15152 34524
rect 15000 34470 15016 34522
rect 15104 34470 15140 34522
rect 15000 34468 15048 34470
rect 15104 34468 15152 34470
rect 14008 34458 15208 34468
rect 15820 34356 15876 38612
rect 16044 37828 16100 39340
rect 16044 36596 16100 37772
rect 16156 38948 16212 38958
rect 16156 38834 16212 38892
rect 16156 38782 16158 38834
rect 16210 38782 16212 38834
rect 16156 37490 16212 38782
rect 16156 37438 16158 37490
rect 16210 37438 16212 37490
rect 16156 37426 16212 37438
rect 16044 36530 16100 36540
rect 15820 34262 15876 34300
rect 16268 34356 16324 43820
rect 16492 43650 16548 45276
rect 16604 45266 16660 45276
rect 16716 45220 16772 45948
rect 16828 45938 16884 45948
rect 18284 46002 18340 46732
rect 18284 45950 18286 46002
rect 18338 45950 18340 46002
rect 18284 45938 18340 45950
rect 17500 45892 17556 45902
rect 17500 45798 17556 45836
rect 17836 45780 17892 45790
rect 17724 45778 17892 45780
rect 17724 45726 17838 45778
rect 17890 45726 17892 45778
rect 17724 45724 17892 45726
rect 17724 45332 17780 45724
rect 17836 45714 17892 45724
rect 18060 45778 18116 45790
rect 18060 45726 18062 45778
rect 18114 45726 18116 45778
rect 18060 45332 18116 45726
rect 17724 45266 17780 45276
rect 17836 45276 18116 45332
rect 18284 45332 18340 45342
rect 17388 45220 17444 45230
rect 16716 45218 17108 45220
rect 16716 45166 16718 45218
rect 16770 45166 17108 45218
rect 16716 45164 17108 45166
rect 16716 43762 16772 45164
rect 16828 44996 16884 45006
rect 16828 44902 16884 44940
rect 17052 44546 17108 45164
rect 17388 44884 17444 45164
rect 17724 45106 17780 45118
rect 17724 45054 17726 45106
rect 17778 45054 17780 45106
rect 17388 44818 17444 44828
rect 17500 44994 17556 45006
rect 17500 44942 17502 44994
rect 17554 44942 17556 44994
rect 17052 44494 17054 44546
rect 17106 44494 17108 44546
rect 17052 44482 17108 44494
rect 16716 43710 16718 43762
rect 16770 43710 16772 43762
rect 16716 43698 16772 43710
rect 16492 43598 16494 43650
rect 16546 43598 16548 43650
rect 16492 43586 16548 43598
rect 17388 43652 17444 43662
rect 16380 43538 16436 43550
rect 16380 43486 16382 43538
rect 16434 43486 16436 43538
rect 16380 42980 16436 43486
rect 16604 43538 16660 43550
rect 16604 43486 16606 43538
rect 16658 43486 16660 43538
rect 16604 43428 16660 43486
rect 17388 43538 17444 43596
rect 17388 43486 17390 43538
rect 17442 43486 17444 43538
rect 17388 43474 17444 43486
rect 16604 43362 16660 43372
rect 16716 43204 16772 43214
rect 16380 42924 16548 42980
rect 16380 42754 16436 42766
rect 16380 42702 16382 42754
rect 16434 42702 16436 42754
rect 16380 38612 16436 42702
rect 16492 41412 16548 42924
rect 16716 42754 16772 43148
rect 17500 43204 17556 44942
rect 17612 44548 17668 44558
rect 17612 44434 17668 44492
rect 17612 44382 17614 44434
rect 17666 44382 17668 44434
rect 17612 44370 17668 44382
rect 17724 44436 17780 45054
rect 17724 44322 17780 44380
rect 17724 44270 17726 44322
rect 17778 44270 17780 44322
rect 17724 44258 17780 44270
rect 17612 44212 17668 44222
rect 17612 43762 17668 44156
rect 17612 43710 17614 43762
rect 17666 43710 17668 43762
rect 17612 43698 17668 43710
rect 17724 43764 17780 43774
rect 17836 43764 17892 45276
rect 17948 45106 18004 45118
rect 17948 45054 17950 45106
rect 18002 45054 18004 45106
rect 17948 44884 18004 45054
rect 18284 45106 18340 45276
rect 18284 45054 18286 45106
rect 18338 45054 18340 45106
rect 18284 45042 18340 45054
rect 18284 44884 18340 44894
rect 17948 44882 18340 44884
rect 17948 44830 18286 44882
rect 18338 44830 18340 44882
rect 17948 44828 18340 44830
rect 18284 44818 18340 44828
rect 18060 44322 18116 44334
rect 18060 44270 18062 44322
rect 18114 44270 18116 44322
rect 17724 43762 17892 43764
rect 17724 43710 17726 43762
rect 17778 43710 17892 43762
rect 17724 43708 17892 43710
rect 17948 44098 18004 44110
rect 17948 44046 17950 44098
rect 18002 44046 18004 44098
rect 17724 43698 17780 43708
rect 17500 43138 17556 43148
rect 17836 43538 17892 43550
rect 17836 43486 17838 43538
rect 17890 43486 17892 43538
rect 16716 42702 16718 42754
rect 16770 42702 16772 42754
rect 16716 42690 16772 42702
rect 17836 42420 17892 43486
rect 17612 42364 17892 42420
rect 16492 41346 16548 41356
rect 17500 41412 17556 41422
rect 16716 38948 16772 38958
rect 17500 38948 17556 41356
rect 17612 41074 17668 42364
rect 17836 42196 17892 42206
rect 17836 42102 17892 42140
rect 17724 42084 17780 42094
rect 17724 41990 17780 42028
rect 17612 41022 17614 41074
rect 17666 41022 17668 41074
rect 17612 40628 17668 41022
rect 17612 40562 17668 40572
rect 17948 40516 18004 44046
rect 18060 43652 18116 44270
rect 18060 43538 18116 43596
rect 18060 43486 18062 43538
rect 18114 43486 18116 43538
rect 18060 42196 18116 43486
rect 18060 42130 18116 42140
rect 18172 44212 18228 44222
rect 18172 41860 18228 44156
rect 18396 43764 18452 46956
rect 18508 44660 18564 48190
rect 18620 47068 18676 48636
rect 18620 47002 18676 47012
rect 18732 46564 18788 49084
rect 18844 49026 18900 49084
rect 18844 48974 18846 49026
rect 18898 48974 18900 49026
rect 18844 48962 18900 48974
rect 19068 48354 19124 49868
rect 19516 49858 19572 49868
rect 19292 49252 19348 49262
rect 19628 49252 19684 50372
rect 19292 49250 19684 49252
rect 19292 49198 19294 49250
rect 19346 49198 19684 49250
rect 19292 49196 19684 49198
rect 20188 49252 20244 51996
rect 20300 51378 20356 52110
rect 20412 52162 20468 52556
rect 20412 52110 20414 52162
rect 20466 52110 20468 52162
rect 20412 52098 20468 52110
rect 20860 52164 20916 52174
rect 21196 52164 21252 52174
rect 20860 52162 21252 52164
rect 20860 52110 20862 52162
rect 20914 52110 21198 52162
rect 21250 52110 21252 52162
rect 20860 52108 21252 52110
rect 20860 52098 20916 52108
rect 21196 52098 21252 52108
rect 21532 52162 21588 52780
rect 21644 52612 21700 53118
rect 21644 52546 21700 52556
rect 21532 52110 21534 52162
rect 21586 52110 21588 52162
rect 21532 52052 21588 52110
rect 21532 51986 21588 51996
rect 21420 51940 21476 51950
rect 21420 51846 21476 51884
rect 20300 51326 20302 51378
rect 20354 51326 20356 51378
rect 20300 51314 20356 51326
rect 19292 49186 19348 49196
rect 20076 49140 20132 49150
rect 20076 49046 20132 49084
rect 19628 48804 19684 48814
rect 19628 48710 19684 48748
rect 19068 48302 19070 48354
rect 19122 48302 19124 48354
rect 19068 48290 19124 48302
rect 19852 47236 19908 47246
rect 18956 46900 19012 46910
rect 19012 46844 19348 46900
rect 18956 46806 19012 46844
rect 19292 46674 19348 46844
rect 19292 46622 19294 46674
rect 19346 46622 19348 46674
rect 19292 46610 19348 46622
rect 18732 46508 19012 46564
rect 18732 45668 18788 45678
rect 18732 45574 18788 45612
rect 18620 44884 18676 44894
rect 18620 44790 18676 44828
rect 18508 44604 18676 44660
rect 18508 44436 18564 44446
rect 18508 44342 18564 44380
rect 18620 44434 18676 44604
rect 18956 44548 19012 46508
rect 19292 45666 19348 45678
rect 19292 45614 19294 45666
rect 19346 45614 19348 45666
rect 19292 45556 19348 45614
rect 18956 44482 19012 44492
rect 19068 45500 19292 45556
rect 18620 44382 18622 44434
rect 18674 44382 18676 44434
rect 18620 43988 18676 44382
rect 19068 44434 19124 45500
rect 19292 45490 19348 45500
rect 19628 45668 19684 45678
rect 19068 44382 19070 44434
rect 19122 44382 19124 44434
rect 19068 44212 19124 44382
rect 19068 44146 19124 44156
rect 19180 45332 19236 45342
rect 18620 43922 18676 43932
rect 18956 44098 19012 44110
rect 18956 44046 18958 44098
rect 19010 44046 19012 44098
rect 18844 43876 18900 43886
rect 18732 43764 18788 43774
rect 18396 43762 18788 43764
rect 18396 43710 18734 43762
rect 18786 43710 18788 43762
rect 18396 43708 18788 43710
rect 18732 43698 18788 43708
rect 18844 43762 18900 43820
rect 18844 43710 18846 43762
rect 18898 43710 18900 43762
rect 18844 43698 18900 43710
rect 18396 43538 18452 43550
rect 18620 43540 18676 43550
rect 18396 43486 18398 43538
rect 18450 43486 18452 43538
rect 18396 43316 18452 43486
rect 18396 42084 18452 43260
rect 18396 42018 18452 42028
rect 18508 43538 18676 43540
rect 18508 43486 18622 43538
rect 18674 43486 18676 43538
rect 18508 43484 18676 43486
rect 18396 41860 18452 41870
rect 18172 41858 18452 41860
rect 18172 41806 18398 41858
rect 18450 41806 18452 41858
rect 18172 41804 18452 41806
rect 18396 41298 18452 41804
rect 18396 41246 18398 41298
rect 18450 41246 18452 41298
rect 18396 41234 18452 41246
rect 17948 40460 18340 40516
rect 18172 39620 18228 39630
rect 17836 39618 18228 39620
rect 17836 39566 18174 39618
rect 18226 39566 18228 39618
rect 17836 39564 18228 39566
rect 17836 39058 17892 39564
rect 18172 39554 18228 39564
rect 17836 39006 17838 39058
rect 17890 39006 17892 39058
rect 17836 38994 17892 39006
rect 17612 38948 17668 38958
rect 17500 38946 17668 38948
rect 17500 38894 17614 38946
rect 17666 38894 17668 38946
rect 17500 38892 17668 38894
rect 16492 38724 16548 38762
rect 16492 38658 16548 38668
rect 16380 38546 16436 38556
rect 16716 37492 16772 38892
rect 17612 38882 17668 38892
rect 18284 38946 18340 40460
rect 18508 40404 18564 43484
rect 18620 43474 18676 43484
rect 18956 43538 19012 44046
rect 18956 43486 18958 43538
rect 19010 43486 19012 43538
rect 18956 43428 19012 43486
rect 18956 43362 19012 43372
rect 19068 42196 19124 42206
rect 19068 42102 19124 42140
rect 18732 41972 18788 41982
rect 18732 41298 18788 41916
rect 19180 41748 19236 45276
rect 19628 45330 19684 45612
rect 19628 45278 19630 45330
rect 19682 45278 19684 45330
rect 19628 45266 19684 45278
rect 19292 44996 19348 45006
rect 19516 44996 19572 45006
rect 19292 44994 19572 44996
rect 19292 44942 19294 44994
rect 19346 44942 19518 44994
rect 19570 44942 19572 44994
rect 19292 44940 19572 44942
rect 19292 44930 19348 44940
rect 19292 43540 19348 43550
rect 19292 43446 19348 43484
rect 19292 42756 19348 42766
rect 19404 42756 19460 44940
rect 19516 44930 19572 44940
rect 19852 44884 19908 47180
rect 20188 47068 20244 49196
rect 20972 48244 21028 48254
rect 20972 48150 21028 48188
rect 21420 48242 21476 48254
rect 21420 48190 21422 48242
rect 21474 48190 21476 48242
rect 21420 47572 21476 48190
rect 21420 47506 21476 47516
rect 21644 47236 21700 47246
rect 21644 47142 21700 47180
rect 20188 47012 20356 47068
rect 20300 46004 20356 47012
rect 20748 46004 20804 46014
rect 20300 46002 21364 46004
rect 20300 45950 20302 46002
rect 20354 45950 20750 46002
rect 20802 45950 21364 46002
rect 20300 45948 21364 45950
rect 20300 45938 20356 45948
rect 20748 45938 20804 45948
rect 21308 45892 21364 45948
rect 21308 45798 21364 45836
rect 21420 45666 21476 45678
rect 21420 45614 21422 45666
rect 21474 45614 21476 45666
rect 21420 45444 21476 45614
rect 21532 45668 21588 45678
rect 21532 45574 21588 45612
rect 20524 45388 21476 45444
rect 19852 44818 19908 44828
rect 20076 45106 20132 45118
rect 20076 45054 20078 45106
rect 20130 45054 20132 45106
rect 19964 44212 20020 44222
rect 19740 44100 19796 44110
rect 19964 44100 20020 44156
rect 19740 44098 20020 44100
rect 19740 44046 19742 44098
rect 19794 44046 20020 44098
rect 19740 44044 20020 44046
rect 19740 44034 19796 44044
rect 19516 43876 19572 43886
rect 19572 43820 19684 43876
rect 19516 43810 19572 43820
rect 19628 42980 19684 43820
rect 19964 43762 20020 44044
rect 19964 43710 19966 43762
rect 20018 43710 20020 43762
rect 19740 43652 19796 43662
rect 19740 43558 19796 43596
rect 19852 43428 19908 43438
rect 19852 43334 19908 43372
rect 19852 42980 19908 42990
rect 19628 42978 19908 42980
rect 19628 42926 19854 42978
rect 19906 42926 19908 42978
rect 19628 42924 19908 42926
rect 19852 42914 19908 42924
rect 19348 42700 19460 42756
rect 19292 42690 19348 42700
rect 19292 42530 19348 42542
rect 19292 42478 19294 42530
rect 19346 42478 19348 42530
rect 19292 41860 19348 42478
rect 19964 42196 20020 43710
rect 20076 42532 20132 45054
rect 20524 45106 20580 45388
rect 21756 45332 21812 53900
rect 22204 53284 22260 55468
rect 22540 55412 22596 56252
rect 22764 56214 22820 56252
rect 22652 55858 22708 55870
rect 22652 55806 22654 55858
rect 22706 55806 22708 55858
rect 22652 55522 22708 55806
rect 22652 55470 22654 55522
rect 22706 55470 22708 55522
rect 22652 55458 22708 55470
rect 22092 53172 22148 53182
rect 22204 53172 22260 53228
rect 22092 53170 22260 53172
rect 22092 53118 22094 53170
rect 22146 53118 22260 53170
rect 22092 53116 22260 53118
rect 22316 55410 22596 55412
rect 22316 55358 22542 55410
rect 22594 55358 22596 55410
rect 22316 55356 22596 55358
rect 21868 52164 21924 52174
rect 21868 52070 21924 52108
rect 21980 51940 22036 51950
rect 21980 49810 22036 51884
rect 21980 49758 21982 49810
rect 22034 49758 22036 49810
rect 21980 49746 22036 49758
rect 22092 47796 22148 53116
rect 22316 52948 22372 55356
rect 22540 55346 22596 55356
rect 22316 49028 22372 52892
rect 22540 55188 22596 55198
rect 22540 54402 22596 55132
rect 22876 54740 22932 56700
rect 23100 56690 23156 56700
rect 22988 56196 23044 56206
rect 22988 56102 23044 56140
rect 22876 54674 22932 54684
rect 22540 54350 22542 54402
rect 22594 54350 22596 54402
rect 22540 52500 22596 54350
rect 22876 53732 22932 53742
rect 22652 53284 22708 53294
rect 22652 53170 22708 53228
rect 22652 53118 22654 53170
rect 22706 53118 22708 53170
rect 22652 53106 22708 53118
rect 22876 53170 22932 53676
rect 22876 53118 22878 53170
rect 22930 53118 22932 53170
rect 22876 53106 22932 53118
rect 22764 52836 22820 52846
rect 22540 52434 22596 52444
rect 22652 52834 22820 52836
rect 22652 52782 22766 52834
rect 22818 52782 22820 52834
rect 22652 52780 22820 52782
rect 22652 52276 22708 52780
rect 22764 52770 22820 52780
rect 22428 52220 22708 52276
rect 22428 52162 22484 52220
rect 22428 52110 22430 52162
rect 22482 52110 22484 52162
rect 22428 52098 22484 52110
rect 22876 51604 22932 51614
rect 22876 51510 22932 51548
rect 22428 50708 22484 50718
rect 22428 49810 22484 50652
rect 23100 50708 23156 50718
rect 23100 50614 23156 50652
rect 23212 50428 23268 58940
rect 23548 54852 23604 63084
rect 23772 63046 23828 63084
rect 23884 62916 23940 65996
rect 24556 66052 24612 66062
rect 24556 65958 24612 65996
rect 25004 66050 25060 66062
rect 25004 65998 25006 66050
rect 25058 65998 25060 66050
rect 25004 65380 25060 65998
rect 25340 65490 25396 67228
rect 25452 67170 25508 67182
rect 25452 67118 25454 67170
rect 25506 67118 25508 67170
rect 25452 66276 25508 67118
rect 25564 66946 25620 67564
rect 25564 66894 25566 66946
rect 25618 66894 25620 66946
rect 25564 66882 25620 66894
rect 25900 66612 25956 69468
rect 26236 70196 26292 70206
rect 26348 70196 26404 70206
rect 26292 70194 26404 70196
rect 26292 70142 26350 70194
rect 26402 70142 26404 70194
rect 26292 70140 26404 70142
rect 26012 67844 26068 67854
rect 26236 67844 26292 70140
rect 26348 70130 26404 70140
rect 26460 70084 26516 70094
rect 26460 69990 26516 70028
rect 27020 69300 27076 70364
rect 27132 70196 27188 70206
rect 27132 70102 27188 70140
rect 27020 69186 27076 69244
rect 27020 69134 27022 69186
rect 27074 69134 27076 69186
rect 27020 69122 27076 69134
rect 26684 68628 26740 68638
rect 26012 67842 26292 67844
rect 26012 67790 26014 67842
rect 26066 67790 26292 67842
rect 26012 67788 26292 67790
rect 26348 68516 26404 68526
rect 26012 67778 26068 67788
rect 26124 67284 26180 67294
rect 26348 67284 26404 68460
rect 26460 68404 26516 68414
rect 26460 67844 26516 68348
rect 26684 68066 26740 68572
rect 26684 68014 26686 68066
rect 26738 68014 26740 68066
rect 26684 68002 26740 68014
rect 26460 67750 26516 67788
rect 26796 67954 26852 67966
rect 26796 67902 26798 67954
rect 26850 67902 26852 67954
rect 26124 67282 26404 67284
rect 26124 67230 26126 67282
rect 26178 67230 26404 67282
rect 26124 67228 26404 67230
rect 26124 67218 26180 67228
rect 25564 66556 25956 66612
rect 26012 67170 26068 67182
rect 26012 67118 26014 67170
rect 26066 67118 26068 67170
rect 25564 66386 25620 66556
rect 25564 66334 25566 66386
rect 25618 66334 25620 66386
rect 25564 66322 25620 66334
rect 25452 66052 25508 66220
rect 25900 66052 25956 66062
rect 25452 66050 25956 66052
rect 25452 65998 25902 66050
rect 25954 65998 25956 66050
rect 25452 65996 25956 65998
rect 26012 66052 26068 67118
rect 26236 66948 26292 66958
rect 26236 66854 26292 66892
rect 26684 66948 26740 66958
rect 26684 66854 26740 66892
rect 26348 66052 26404 66062
rect 26012 66050 26516 66052
rect 26012 65998 26350 66050
rect 26402 65998 26516 66050
rect 26012 65996 26516 65998
rect 25340 65438 25342 65490
rect 25394 65438 25396 65490
rect 25340 65426 25396 65438
rect 25004 65314 25060 65324
rect 24008 65100 25208 65110
rect 24064 65098 24112 65100
rect 24168 65098 24216 65100
rect 24076 65046 24112 65098
rect 24200 65046 24216 65098
rect 24064 65044 24112 65046
rect 24168 65044 24216 65046
rect 24272 65098 24320 65100
rect 24376 65098 24424 65100
rect 24480 65098 24528 65100
rect 24376 65046 24396 65098
rect 24480 65046 24520 65098
rect 24272 65044 24320 65046
rect 24376 65044 24424 65046
rect 24480 65044 24528 65046
rect 24584 65044 24632 65100
rect 24688 65098 24736 65100
rect 24792 65098 24840 65100
rect 24896 65098 24944 65100
rect 24696 65046 24736 65098
rect 24820 65046 24840 65098
rect 24688 65044 24736 65046
rect 24792 65044 24840 65046
rect 24896 65044 24944 65046
rect 25000 65098 25048 65100
rect 25104 65098 25152 65100
rect 25000 65046 25016 65098
rect 25104 65046 25140 65098
rect 25000 65044 25048 65046
rect 25104 65044 25152 65046
rect 24008 65034 25208 65044
rect 25340 63922 25396 63934
rect 25340 63870 25342 63922
rect 25394 63870 25396 63922
rect 24008 63532 25208 63542
rect 24064 63530 24112 63532
rect 24168 63530 24216 63532
rect 24076 63478 24112 63530
rect 24200 63478 24216 63530
rect 24064 63476 24112 63478
rect 24168 63476 24216 63478
rect 24272 63530 24320 63532
rect 24376 63530 24424 63532
rect 24480 63530 24528 63532
rect 24376 63478 24396 63530
rect 24480 63478 24520 63530
rect 24272 63476 24320 63478
rect 24376 63476 24424 63478
rect 24480 63476 24528 63478
rect 24584 63476 24632 63532
rect 24688 63530 24736 63532
rect 24792 63530 24840 63532
rect 24896 63530 24944 63532
rect 24696 63478 24736 63530
rect 24820 63478 24840 63530
rect 24688 63476 24736 63478
rect 24792 63476 24840 63478
rect 24896 63476 24944 63478
rect 25000 63530 25048 63532
rect 25104 63530 25152 63532
rect 25000 63478 25016 63530
rect 25104 63478 25140 63530
rect 25000 63476 25048 63478
rect 25104 63476 25152 63478
rect 24008 63466 25208 63476
rect 24780 63252 24836 63262
rect 24780 63158 24836 63196
rect 24892 63140 24948 63150
rect 24892 63046 24948 63084
rect 25228 63138 25284 63150
rect 25228 63086 25230 63138
rect 25282 63086 25284 63138
rect 24108 63028 24164 63038
rect 24108 62934 24164 62972
rect 24668 63028 24724 63038
rect 24668 62934 24724 62972
rect 23772 62860 23940 62916
rect 25228 62916 25284 63086
rect 23772 62188 23828 62860
rect 25228 62850 25284 62860
rect 24108 62580 24164 62590
rect 24108 62188 24164 62524
rect 24668 62468 24724 62478
rect 24668 62374 24724 62412
rect 25340 62356 25396 63870
rect 25676 63922 25732 63934
rect 25676 63870 25678 63922
rect 25730 63870 25732 63922
rect 25676 63252 25732 63870
rect 25676 63186 25732 63196
rect 25676 62914 25732 62926
rect 25676 62862 25678 62914
rect 25730 62862 25732 62914
rect 25676 62468 25732 62862
rect 25676 62402 25732 62412
rect 25340 62262 25396 62300
rect 25788 62354 25844 62366
rect 25788 62302 25790 62354
rect 25842 62302 25844 62354
rect 23660 62132 23828 62188
rect 23884 62132 24164 62188
rect 23660 58828 23716 62132
rect 23772 60002 23828 60014
rect 23772 59950 23774 60002
rect 23826 59950 23828 60002
rect 23772 59780 23828 59950
rect 23772 59714 23828 59724
rect 23884 59444 23940 62132
rect 24008 61964 25208 61974
rect 24064 61962 24112 61964
rect 24168 61962 24216 61964
rect 24076 61910 24112 61962
rect 24200 61910 24216 61962
rect 24064 61908 24112 61910
rect 24168 61908 24216 61910
rect 24272 61962 24320 61964
rect 24376 61962 24424 61964
rect 24480 61962 24528 61964
rect 24376 61910 24396 61962
rect 24480 61910 24520 61962
rect 24272 61908 24320 61910
rect 24376 61908 24424 61910
rect 24480 61908 24528 61910
rect 24584 61908 24632 61964
rect 24688 61962 24736 61964
rect 24792 61962 24840 61964
rect 24896 61962 24944 61964
rect 24696 61910 24736 61962
rect 24820 61910 24840 61962
rect 24688 61908 24736 61910
rect 24792 61908 24840 61910
rect 24896 61908 24944 61910
rect 25000 61962 25048 61964
rect 25104 61962 25152 61964
rect 25000 61910 25016 61962
rect 25104 61910 25140 61962
rect 25000 61908 25048 61910
rect 25104 61908 25152 61910
rect 24008 61898 25208 61908
rect 25788 61908 25844 62302
rect 25788 61842 25844 61852
rect 24220 61796 24276 61806
rect 24220 61682 24276 61740
rect 24220 61630 24222 61682
rect 24274 61630 24276 61682
rect 24220 61618 24276 61630
rect 25228 61796 25284 61806
rect 24556 61460 24612 61470
rect 24556 61366 24612 61404
rect 25228 61458 25284 61740
rect 25228 61406 25230 61458
rect 25282 61406 25284 61458
rect 25228 61394 25284 61406
rect 25788 61460 25844 61470
rect 25788 61366 25844 61404
rect 25900 60900 25956 65996
rect 26348 65986 26404 65996
rect 26012 65492 26068 65502
rect 26012 65398 26068 65436
rect 26012 62132 26068 62142
rect 26012 61794 26068 62076
rect 26124 61908 26180 61918
rect 26180 61852 26404 61908
rect 26124 61842 26180 61852
rect 26012 61742 26014 61794
rect 26066 61742 26068 61794
rect 26012 61730 26068 61742
rect 26348 61794 26404 61852
rect 26348 61742 26350 61794
rect 26402 61742 26404 61794
rect 26348 61730 26404 61742
rect 25900 60844 26180 60900
rect 25340 60676 25396 60686
rect 25340 60582 25396 60620
rect 26012 60676 26068 60686
rect 24008 60396 25208 60406
rect 24064 60394 24112 60396
rect 24168 60394 24216 60396
rect 24076 60342 24112 60394
rect 24200 60342 24216 60394
rect 24064 60340 24112 60342
rect 24168 60340 24216 60342
rect 24272 60394 24320 60396
rect 24376 60394 24424 60396
rect 24480 60394 24528 60396
rect 24376 60342 24396 60394
rect 24480 60342 24520 60394
rect 24272 60340 24320 60342
rect 24376 60340 24424 60342
rect 24480 60340 24528 60342
rect 24584 60340 24632 60396
rect 24688 60394 24736 60396
rect 24792 60394 24840 60396
rect 24896 60394 24944 60396
rect 24696 60342 24736 60394
rect 24820 60342 24840 60394
rect 24688 60340 24736 60342
rect 24792 60340 24840 60342
rect 24896 60340 24944 60342
rect 25000 60394 25048 60396
rect 25104 60394 25152 60396
rect 25000 60342 25016 60394
rect 25104 60342 25140 60394
rect 25000 60340 25048 60342
rect 25104 60340 25152 60342
rect 24008 60330 25208 60340
rect 26012 60114 26068 60620
rect 26012 60062 26014 60114
rect 26066 60062 26068 60114
rect 23660 58772 23828 58828
rect 23660 58212 23716 58222
rect 23660 57652 23716 58156
rect 23772 58100 23828 58772
rect 23884 58548 23940 59388
rect 25340 59444 25396 59454
rect 25340 59350 25396 59388
rect 26012 59218 26068 60062
rect 26012 59166 26014 59218
rect 26066 59166 26068 59218
rect 25788 59108 25844 59118
rect 26012 59108 26068 59166
rect 25788 59106 26068 59108
rect 25788 59054 25790 59106
rect 25842 59054 26068 59106
rect 25788 59052 26068 59054
rect 25788 59042 25844 59052
rect 24008 58828 25208 58838
rect 24064 58826 24112 58828
rect 24168 58826 24216 58828
rect 24076 58774 24112 58826
rect 24200 58774 24216 58826
rect 24064 58772 24112 58774
rect 24168 58772 24216 58774
rect 24272 58826 24320 58828
rect 24376 58826 24424 58828
rect 24480 58826 24528 58828
rect 24376 58774 24396 58826
rect 24480 58774 24520 58826
rect 24272 58772 24320 58774
rect 24376 58772 24424 58774
rect 24480 58772 24528 58774
rect 24584 58772 24632 58828
rect 24688 58826 24736 58828
rect 24792 58826 24840 58828
rect 24896 58826 24944 58828
rect 24696 58774 24736 58826
rect 24820 58774 24840 58826
rect 24688 58772 24736 58774
rect 24792 58772 24840 58774
rect 24896 58772 24944 58774
rect 25000 58826 25048 58828
rect 25104 58826 25152 58828
rect 25000 58774 25016 58826
rect 25104 58774 25140 58826
rect 25000 58772 25048 58774
rect 25104 58772 25152 58774
rect 24008 58762 25208 58772
rect 23884 58492 24388 58548
rect 24220 58210 24276 58222
rect 24220 58158 24222 58210
rect 24274 58158 24276 58210
rect 24220 58100 24276 58158
rect 23772 58044 24276 58100
rect 23660 57586 23716 57596
rect 23884 56644 23940 58044
rect 24220 57876 24276 57886
rect 24332 57876 24388 58492
rect 26012 58436 26068 59052
rect 26012 58370 26068 58380
rect 25676 58324 25732 58334
rect 24220 57874 24388 57876
rect 24220 57822 24222 57874
rect 24274 57822 24388 57874
rect 24220 57820 24388 57822
rect 25340 58268 25676 58324
rect 25340 57874 25396 58268
rect 25676 58258 25732 58268
rect 25340 57822 25342 57874
rect 25394 57822 25396 57874
rect 24220 57810 24276 57820
rect 25340 57810 25396 57822
rect 25452 57988 25508 57998
rect 26124 57988 26180 60844
rect 26236 57988 26292 57998
rect 26124 57932 26236 57988
rect 24780 57764 24836 57774
rect 24780 57670 24836 57708
rect 25340 57316 25396 57326
rect 24008 57260 25208 57270
rect 24064 57258 24112 57260
rect 24168 57258 24216 57260
rect 24076 57206 24112 57258
rect 24200 57206 24216 57258
rect 24064 57204 24112 57206
rect 24168 57204 24216 57206
rect 24272 57258 24320 57260
rect 24376 57258 24424 57260
rect 24480 57258 24528 57260
rect 24376 57206 24396 57258
rect 24480 57206 24520 57258
rect 24272 57204 24320 57206
rect 24376 57204 24424 57206
rect 24480 57204 24528 57206
rect 24584 57204 24632 57260
rect 24688 57258 24736 57260
rect 24792 57258 24840 57260
rect 24896 57258 24944 57260
rect 24696 57206 24736 57258
rect 24820 57206 24840 57258
rect 24688 57204 24736 57206
rect 24792 57204 24840 57206
rect 24896 57204 24944 57206
rect 25000 57258 25048 57260
rect 25104 57258 25152 57260
rect 25000 57206 25016 57258
rect 25104 57206 25140 57258
rect 25000 57204 25048 57206
rect 25104 57204 25152 57206
rect 24008 57194 25208 57204
rect 25340 57092 25396 57260
rect 24668 57036 25396 57092
rect 23996 56644 24052 56654
rect 23884 56588 23996 56644
rect 23996 56578 24052 56588
rect 24668 56306 24724 57036
rect 25116 56868 25172 56878
rect 25116 56774 25172 56812
rect 24668 56254 24670 56306
rect 24722 56254 24724 56306
rect 24668 56196 24724 56254
rect 25340 56308 25396 56318
rect 25452 56308 25508 57932
rect 25900 57762 25956 57774
rect 25900 57710 25902 57762
rect 25954 57710 25956 57762
rect 25676 57652 25732 57662
rect 25676 57558 25732 57596
rect 25900 57316 25956 57710
rect 26236 57762 26292 57932
rect 26236 57710 26238 57762
rect 26290 57710 26292 57762
rect 26236 57698 26292 57710
rect 26460 57316 26516 65996
rect 26796 64932 26852 67902
rect 26796 64866 26852 64876
rect 27020 63924 27076 63934
rect 26572 63028 26628 63038
rect 26572 62934 26628 62972
rect 27020 63026 27076 63868
rect 27020 62974 27022 63026
rect 27074 62974 27076 63026
rect 27020 62962 27076 62974
rect 27132 63028 27188 63038
rect 27132 62934 27188 62972
rect 26796 62916 26852 62926
rect 26796 62822 26852 62860
rect 26908 61460 26964 61470
rect 26684 61012 26740 61022
rect 26684 60674 26740 60956
rect 26684 60622 26686 60674
rect 26738 60622 26740 60674
rect 26684 59780 26740 60622
rect 26684 59714 26740 59724
rect 26684 59220 26740 59230
rect 26684 59218 26852 59220
rect 26684 59166 26686 59218
rect 26738 59166 26852 59218
rect 26684 59164 26852 59166
rect 26684 59154 26740 59164
rect 25900 57250 25956 57260
rect 26348 57260 26516 57316
rect 26572 58436 26628 58446
rect 25900 57090 25956 57102
rect 25900 57038 25902 57090
rect 25954 57038 25956 57090
rect 25340 56306 25508 56308
rect 25340 56254 25342 56306
rect 25394 56254 25508 56306
rect 25340 56252 25508 56254
rect 25340 56242 25396 56252
rect 24668 56130 24724 56140
rect 24008 55692 25208 55702
rect 24064 55690 24112 55692
rect 24168 55690 24216 55692
rect 24076 55638 24112 55690
rect 24200 55638 24216 55690
rect 24064 55636 24112 55638
rect 24168 55636 24216 55638
rect 24272 55690 24320 55692
rect 24376 55690 24424 55692
rect 24480 55690 24528 55692
rect 24376 55638 24396 55690
rect 24480 55638 24520 55690
rect 24272 55636 24320 55638
rect 24376 55636 24424 55638
rect 24480 55636 24528 55638
rect 24584 55636 24632 55692
rect 24688 55690 24736 55692
rect 24792 55690 24840 55692
rect 24896 55690 24944 55692
rect 24696 55638 24736 55690
rect 24820 55638 24840 55690
rect 24688 55636 24736 55638
rect 24792 55636 24840 55638
rect 24896 55636 24944 55638
rect 25000 55690 25048 55692
rect 25104 55690 25152 55692
rect 25000 55638 25016 55690
rect 25104 55638 25140 55690
rect 25000 55636 25048 55638
rect 25104 55636 25152 55638
rect 24008 55626 25208 55636
rect 23548 54796 23716 54852
rect 23548 54628 23604 54638
rect 23548 53844 23604 54572
rect 23548 53778 23604 53788
rect 23660 53732 23716 54796
rect 24008 54124 25208 54134
rect 24064 54122 24112 54124
rect 24168 54122 24216 54124
rect 24076 54070 24112 54122
rect 24200 54070 24216 54122
rect 24064 54068 24112 54070
rect 24168 54068 24216 54070
rect 24272 54122 24320 54124
rect 24376 54122 24424 54124
rect 24480 54122 24528 54124
rect 24376 54070 24396 54122
rect 24480 54070 24520 54122
rect 24272 54068 24320 54070
rect 24376 54068 24424 54070
rect 24480 54068 24528 54070
rect 24584 54068 24632 54124
rect 24688 54122 24736 54124
rect 24792 54122 24840 54124
rect 24896 54122 24944 54124
rect 24696 54070 24736 54122
rect 24820 54070 24840 54122
rect 24688 54068 24736 54070
rect 24792 54068 24840 54070
rect 24896 54068 24944 54070
rect 25000 54122 25048 54124
rect 25104 54122 25152 54124
rect 25000 54070 25016 54122
rect 25104 54070 25140 54122
rect 25000 54068 25048 54070
rect 25104 54068 25152 54070
rect 24008 54058 25208 54068
rect 23660 53666 23716 53676
rect 24668 53844 24724 53854
rect 24668 53730 24724 53788
rect 24668 53678 24670 53730
rect 24722 53678 24724 53730
rect 24668 53666 24724 53678
rect 25116 53508 25172 53518
rect 25116 53414 25172 53452
rect 23772 53284 23828 53294
rect 23436 53058 23492 53070
rect 23436 53006 23438 53058
rect 23490 53006 23492 53058
rect 23324 52948 23380 52958
rect 23436 52948 23492 53006
rect 23324 52946 23492 52948
rect 23324 52894 23326 52946
rect 23378 52894 23492 52946
rect 23324 52892 23492 52894
rect 23660 53060 23716 53070
rect 23324 52882 23380 52892
rect 23660 52388 23716 53004
rect 23772 53058 23828 53228
rect 24220 53284 24276 53294
rect 24220 53170 24276 53228
rect 24220 53118 24222 53170
rect 24274 53118 24276 53170
rect 24220 53106 24276 53118
rect 25340 53172 25396 53182
rect 25340 53078 25396 53116
rect 23772 53006 23774 53058
rect 23826 53006 23828 53058
rect 23772 52994 23828 53006
rect 24008 52556 25208 52566
rect 24064 52554 24112 52556
rect 24168 52554 24216 52556
rect 24076 52502 24112 52554
rect 24200 52502 24216 52554
rect 24064 52500 24112 52502
rect 24168 52500 24216 52502
rect 24272 52554 24320 52556
rect 24376 52554 24424 52556
rect 24480 52554 24528 52556
rect 24376 52502 24396 52554
rect 24480 52502 24520 52554
rect 24272 52500 24320 52502
rect 24376 52500 24424 52502
rect 24480 52500 24528 52502
rect 24584 52500 24632 52556
rect 24688 52554 24736 52556
rect 24792 52554 24840 52556
rect 24896 52554 24944 52556
rect 24696 52502 24736 52554
rect 24820 52502 24840 52554
rect 24688 52500 24736 52502
rect 24792 52500 24840 52502
rect 24896 52500 24944 52502
rect 25000 52554 25048 52556
rect 25104 52554 25152 52556
rect 25000 52502 25016 52554
rect 25104 52502 25140 52554
rect 25000 52500 25048 52502
rect 25104 52500 25152 52502
rect 25452 52500 25508 56252
rect 25788 56868 25844 56878
rect 25900 56868 25956 57038
rect 25788 56866 25956 56868
rect 25788 56814 25790 56866
rect 25842 56814 25956 56866
rect 25788 56812 25956 56814
rect 25788 55970 25844 56812
rect 26124 56644 26180 56654
rect 26124 56084 26180 56588
rect 26348 56308 26404 57260
rect 26572 57090 26628 58380
rect 26684 58434 26740 58446
rect 26684 58382 26686 58434
rect 26738 58382 26740 58434
rect 26684 58324 26740 58382
rect 26684 58258 26740 58268
rect 26796 57876 26852 59164
rect 26796 57810 26852 57820
rect 26908 57652 26964 61404
rect 27020 60788 27076 60798
rect 27356 60788 27412 70924
rect 27916 70196 27972 70206
rect 27916 70102 27972 70140
rect 28700 70196 28756 70206
rect 27580 70084 27636 70094
rect 27580 69634 27636 70028
rect 27580 69582 27582 69634
rect 27634 69582 27636 69634
rect 27580 69570 27636 69582
rect 27580 69300 27636 69310
rect 27580 67954 27636 69244
rect 27916 69298 27972 69310
rect 28364 69300 28420 69310
rect 27916 69246 27918 69298
rect 27970 69246 27972 69298
rect 27580 67902 27582 67954
rect 27634 67902 27636 67954
rect 27580 67890 27636 67902
rect 27804 69186 27860 69198
rect 27804 69134 27806 69186
rect 27858 69134 27860 69186
rect 27804 67844 27860 69134
rect 27916 68852 27972 69246
rect 27916 68786 27972 68796
rect 28252 69244 28364 69300
rect 28252 68850 28308 69244
rect 28364 69206 28420 69244
rect 28252 68798 28254 68850
rect 28306 68798 28308 68850
rect 28252 68786 28308 68798
rect 27804 67778 27860 67788
rect 28700 66836 28756 70140
rect 29148 69634 29204 69646
rect 29148 69582 29150 69634
rect 29202 69582 29204 69634
rect 29148 69300 29204 69582
rect 29260 69524 29316 69534
rect 29260 69430 29316 69468
rect 28812 68852 28868 68862
rect 28812 68758 28868 68796
rect 29148 68850 29204 69244
rect 29148 68798 29150 68850
rect 29202 68798 29204 68850
rect 29148 68786 29204 68798
rect 29596 68628 29652 78932
rect 34008 78428 35208 78438
rect 34064 78426 34112 78428
rect 34168 78426 34216 78428
rect 34076 78374 34112 78426
rect 34200 78374 34216 78426
rect 34064 78372 34112 78374
rect 34168 78372 34216 78374
rect 34272 78426 34320 78428
rect 34376 78426 34424 78428
rect 34480 78426 34528 78428
rect 34376 78374 34396 78426
rect 34480 78374 34520 78426
rect 34272 78372 34320 78374
rect 34376 78372 34424 78374
rect 34480 78372 34528 78374
rect 34584 78372 34632 78428
rect 34688 78426 34736 78428
rect 34792 78426 34840 78428
rect 34896 78426 34944 78428
rect 34696 78374 34736 78426
rect 34820 78374 34840 78426
rect 34688 78372 34736 78374
rect 34792 78372 34840 78374
rect 34896 78372 34944 78374
rect 35000 78426 35048 78428
rect 35104 78426 35152 78428
rect 35000 78374 35016 78426
rect 35104 78374 35140 78426
rect 35000 78372 35048 78374
rect 35104 78372 35152 78374
rect 34008 78362 35208 78372
rect 34008 76860 35208 76870
rect 34064 76858 34112 76860
rect 34168 76858 34216 76860
rect 34076 76806 34112 76858
rect 34200 76806 34216 76858
rect 34064 76804 34112 76806
rect 34168 76804 34216 76806
rect 34272 76858 34320 76860
rect 34376 76858 34424 76860
rect 34480 76858 34528 76860
rect 34376 76806 34396 76858
rect 34480 76806 34520 76858
rect 34272 76804 34320 76806
rect 34376 76804 34424 76806
rect 34480 76804 34528 76806
rect 34584 76804 34632 76860
rect 34688 76858 34736 76860
rect 34792 76858 34840 76860
rect 34896 76858 34944 76860
rect 34696 76806 34736 76858
rect 34820 76806 34840 76858
rect 34688 76804 34736 76806
rect 34792 76804 34840 76806
rect 34896 76804 34944 76806
rect 35000 76858 35048 76860
rect 35104 76858 35152 76860
rect 35000 76806 35016 76858
rect 35104 76806 35140 76858
rect 35000 76804 35048 76806
rect 35104 76804 35152 76806
rect 34008 76794 35208 76804
rect 34008 75292 35208 75302
rect 34064 75290 34112 75292
rect 34168 75290 34216 75292
rect 34076 75238 34112 75290
rect 34200 75238 34216 75290
rect 34064 75236 34112 75238
rect 34168 75236 34216 75238
rect 34272 75290 34320 75292
rect 34376 75290 34424 75292
rect 34480 75290 34528 75292
rect 34376 75238 34396 75290
rect 34480 75238 34520 75290
rect 34272 75236 34320 75238
rect 34376 75236 34424 75238
rect 34480 75236 34528 75238
rect 34584 75236 34632 75292
rect 34688 75290 34736 75292
rect 34792 75290 34840 75292
rect 34896 75290 34944 75292
rect 34696 75238 34736 75290
rect 34820 75238 34840 75290
rect 34688 75236 34736 75238
rect 34792 75236 34840 75238
rect 34896 75236 34944 75238
rect 35000 75290 35048 75292
rect 35104 75290 35152 75292
rect 35000 75238 35016 75290
rect 35104 75238 35140 75290
rect 35000 75236 35048 75238
rect 35104 75236 35152 75238
rect 34008 75226 35208 75236
rect 34008 73724 35208 73734
rect 34064 73722 34112 73724
rect 34168 73722 34216 73724
rect 34076 73670 34112 73722
rect 34200 73670 34216 73722
rect 34064 73668 34112 73670
rect 34168 73668 34216 73670
rect 34272 73722 34320 73724
rect 34376 73722 34424 73724
rect 34480 73722 34528 73724
rect 34376 73670 34396 73722
rect 34480 73670 34520 73722
rect 34272 73668 34320 73670
rect 34376 73668 34424 73670
rect 34480 73668 34528 73670
rect 34584 73668 34632 73724
rect 34688 73722 34736 73724
rect 34792 73722 34840 73724
rect 34896 73722 34944 73724
rect 34696 73670 34736 73722
rect 34820 73670 34840 73722
rect 34688 73668 34736 73670
rect 34792 73668 34840 73670
rect 34896 73668 34944 73670
rect 35000 73722 35048 73724
rect 35104 73722 35152 73724
rect 35000 73670 35016 73722
rect 35104 73670 35140 73722
rect 35000 73668 35048 73670
rect 35104 73668 35152 73670
rect 34008 73658 35208 73668
rect 34008 72156 35208 72166
rect 34064 72154 34112 72156
rect 34168 72154 34216 72156
rect 34076 72102 34112 72154
rect 34200 72102 34216 72154
rect 34064 72100 34112 72102
rect 34168 72100 34216 72102
rect 34272 72154 34320 72156
rect 34376 72154 34424 72156
rect 34480 72154 34528 72156
rect 34376 72102 34396 72154
rect 34480 72102 34520 72154
rect 34272 72100 34320 72102
rect 34376 72100 34424 72102
rect 34480 72100 34528 72102
rect 34584 72100 34632 72156
rect 34688 72154 34736 72156
rect 34792 72154 34840 72156
rect 34896 72154 34944 72156
rect 34696 72102 34736 72154
rect 34820 72102 34840 72154
rect 34688 72100 34736 72102
rect 34792 72100 34840 72102
rect 34896 72100 34944 72102
rect 35000 72154 35048 72156
rect 35104 72154 35152 72156
rect 35000 72102 35016 72154
rect 35104 72102 35140 72154
rect 35000 72100 35048 72102
rect 35104 72100 35152 72102
rect 34008 72090 35208 72100
rect 35532 71988 35588 71998
rect 35532 71986 36260 71988
rect 35532 71934 35534 71986
rect 35586 71934 36260 71986
rect 35532 71932 36260 71934
rect 35532 71922 35588 71932
rect 35868 71762 35924 71774
rect 35868 71710 35870 71762
rect 35922 71710 35924 71762
rect 30156 71650 30212 71662
rect 30156 71598 30158 71650
rect 30210 71598 30212 71650
rect 30156 70980 30212 71598
rect 35084 71650 35140 71662
rect 35084 71598 35086 71650
rect 35138 71598 35140 71650
rect 34972 71540 35028 71550
rect 34972 71446 35028 71484
rect 29820 70084 29876 70094
rect 29820 69634 29876 70028
rect 29820 69582 29822 69634
rect 29874 69582 29876 69634
rect 29820 69522 29876 69582
rect 29820 69470 29822 69522
rect 29874 69470 29876 69522
rect 29820 69458 29876 69470
rect 29596 68562 29652 68572
rect 30156 69410 30212 70924
rect 32396 70978 32452 70990
rect 32396 70926 32398 70978
rect 32450 70926 32452 70978
rect 31836 70756 31892 70766
rect 32060 70756 32116 70766
rect 31612 70196 31668 70206
rect 31388 70194 31668 70196
rect 31388 70142 31614 70194
rect 31666 70142 31668 70194
rect 31388 70140 31668 70142
rect 31164 70084 31220 70094
rect 31388 70084 31444 70140
rect 31612 70130 31668 70140
rect 31836 70196 31892 70700
rect 31836 70130 31892 70140
rect 31948 70754 32116 70756
rect 31948 70702 32062 70754
rect 32114 70702 32116 70754
rect 31948 70700 32116 70702
rect 31164 70082 31444 70084
rect 31164 70030 31166 70082
rect 31218 70030 31444 70082
rect 31164 70028 31444 70030
rect 31164 69860 31220 70028
rect 31500 69972 31556 69982
rect 30156 69358 30158 69410
rect 30210 69358 30212 69410
rect 29036 68404 29092 68414
rect 29036 67284 29092 68348
rect 30156 68404 30212 69358
rect 30604 69804 31220 69860
rect 31276 69970 31556 69972
rect 31276 69918 31502 69970
rect 31554 69918 31556 69970
rect 31276 69916 31556 69918
rect 30604 68852 30660 69804
rect 31276 69748 31332 69916
rect 31500 69906 31556 69916
rect 31836 69972 31892 69982
rect 31948 69972 32004 70700
rect 32060 70690 32116 70700
rect 32396 70532 32452 70926
rect 32620 70980 32676 70990
rect 33068 70980 33124 70990
rect 32620 70978 33012 70980
rect 32620 70926 32622 70978
rect 32674 70926 33012 70978
rect 32620 70924 33012 70926
rect 32620 70914 32676 70924
rect 32396 70466 32452 70476
rect 32956 70420 33012 70924
rect 33068 70886 33124 70924
rect 33516 70978 33572 70990
rect 33516 70926 33518 70978
rect 33570 70926 33572 70978
rect 33404 70532 33460 70542
rect 33180 70420 33236 70430
rect 32956 70364 33180 70420
rect 33180 70326 33236 70364
rect 33292 70308 33348 70318
rect 32060 70252 32676 70308
rect 32060 70194 32116 70252
rect 32060 70142 32062 70194
rect 32114 70142 32116 70194
rect 32060 70130 32116 70142
rect 32508 70084 32564 70094
rect 32620 70084 32676 70252
rect 33068 70084 33124 70094
rect 32620 70082 33124 70084
rect 32620 70030 33070 70082
rect 33122 70030 33124 70082
rect 32620 70028 33124 70030
rect 32508 69990 32564 70028
rect 33068 70018 33124 70028
rect 31836 69970 32004 69972
rect 31836 69918 31838 69970
rect 31890 69918 32004 69970
rect 31836 69916 32004 69918
rect 31836 69906 31892 69916
rect 30716 69692 31332 69748
rect 30716 69410 30772 69692
rect 30716 69358 30718 69410
rect 30770 69358 30772 69410
rect 30716 69346 30772 69358
rect 30156 68338 30212 68348
rect 30380 68516 30436 68526
rect 30604 68516 30660 68796
rect 30828 68852 30884 68862
rect 30828 68850 31332 68852
rect 30828 68798 30830 68850
rect 30882 68798 31332 68850
rect 30828 68796 31332 68798
rect 30828 68786 30884 68796
rect 30380 68514 30660 68516
rect 30380 68462 30382 68514
rect 30434 68462 30660 68514
rect 30380 68460 30660 68462
rect 31052 68626 31108 68638
rect 31052 68574 31054 68626
rect 31106 68574 31108 68626
rect 29820 67956 29876 67966
rect 30380 67956 30436 68460
rect 28924 67060 28980 67070
rect 29036 67060 29092 67228
rect 28924 67058 29092 67060
rect 28924 67006 28926 67058
rect 28978 67006 29092 67058
rect 28924 67004 29092 67006
rect 28924 66994 28980 67004
rect 28700 66780 28980 66836
rect 28588 66052 28644 66062
rect 28588 65958 28644 65996
rect 28364 65716 28420 65726
rect 28252 65660 28364 65716
rect 28252 64146 28308 65660
rect 28364 65622 28420 65660
rect 28252 64094 28254 64146
rect 28306 64094 28308 64146
rect 28252 62580 28308 64094
rect 28812 63924 28868 63934
rect 28812 63830 28868 63868
rect 28588 62914 28644 62926
rect 28588 62862 28590 62914
rect 28642 62862 28644 62914
rect 28588 62804 28644 62862
rect 28588 62738 28644 62748
rect 28252 62486 28308 62524
rect 28812 62244 28868 62282
rect 28812 62178 28868 62188
rect 28476 61460 28532 61470
rect 28476 61366 28532 61404
rect 28588 61348 28644 61358
rect 28588 61254 28644 61292
rect 27076 60732 27412 60788
rect 28588 61012 28644 61022
rect 27020 60694 27076 60732
rect 28588 60226 28644 60956
rect 28588 60174 28590 60226
rect 28642 60174 28644 60226
rect 28028 59780 28084 59790
rect 28364 59780 28420 59790
rect 28028 59778 28364 59780
rect 28028 59726 28030 59778
rect 28082 59726 28364 59778
rect 28028 59724 28364 59726
rect 28028 59714 28084 59724
rect 28364 59686 28420 59724
rect 28476 59778 28532 59790
rect 28476 59726 28478 59778
rect 28530 59726 28532 59778
rect 27244 59108 27300 59118
rect 27244 57764 27300 59052
rect 27804 58884 27860 58894
rect 27356 58436 27412 58446
rect 27356 58342 27412 58380
rect 27692 58210 27748 58222
rect 27692 58158 27694 58210
rect 27746 58158 27748 58210
rect 27244 57762 27524 57764
rect 27244 57710 27246 57762
rect 27298 57710 27524 57762
rect 27244 57708 27524 57710
rect 27244 57698 27300 57708
rect 27132 57652 27188 57662
rect 26908 57650 27188 57652
rect 26908 57598 27134 57650
rect 27186 57598 27188 57650
rect 26908 57596 27188 57598
rect 26572 57038 26574 57090
rect 26626 57038 26628 57090
rect 26572 56978 26628 57038
rect 26572 56926 26574 56978
rect 26626 56926 26628 56978
rect 26572 56914 26628 56926
rect 27020 56644 27076 56654
rect 27132 56644 27188 57596
rect 27468 56978 27524 57708
rect 27468 56926 27470 56978
rect 27522 56926 27524 56978
rect 27468 56914 27524 56926
rect 27020 56642 27188 56644
rect 27020 56590 27022 56642
rect 27074 56590 27188 56642
rect 27020 56588 27188 56590
rect 27020 56578 27076 56588
rect 26348 56242 26404 56252
rect 26460 56196 26516 56206
rect 26460 56084 26516 56140
rect 26124 56028 26516 56084
rect 25788 55918 25790 55970
rect 25842 55918 25844 55970
rect 25676 53620 25732 53630
rect 24008 52490 25208 52500
rect 25340 52444 25508 52500
rect 25564 53564 25676 53620
rect 23660 52332 23940 52388
rect 23884 52276 23940 52332
rect 23772 52164 23828 52174
rect 23660 52108 23772 52164
rect 22428 49758 22430 49810
rect 22482 49758 22484 49810
rect 22428 49746 22484 49758
rect 22764 50372 23268 50428
rect 23324 52052 23380 52062
rect 22316 48972 22484 49028
rect 22316 48802 22372 48814
rect 22316 48750 22318 48802
rect 22370 48750 22372 48802
rect 22316 48692 22372 48750
rect 22316 48626 22372 48636
rect 21980 47740 22148 47796
rect 21980 47236 22036 47740
rect 22092 47572 22148 47582
rect 22092 47478 22148 47516
rect 21980 47142 22036 47180
rect 22204 47234 22260 47246
rect 22204 47182 22206 47234
rect 22258 47182 22260 47234
rect 22204 46228 22260 47182
rect 21868 46172 22260 46228
rect 21868 45668 21924 46172
rect 22316 46116 22372 46126
rect 21980 46114 22372 46116
rect 21980 46062 22318 46114
rect 22370 46062 22372 46114
rect 21980 46060 22372 46062
rect 21980 45890 22036 46060
rect 22316 46050 22372 46060
rect 21980 45838 21982 45890
rect 22034 45838 22036 45890
rect 21980 45826 22036 45838
rect 22204 45892 22260 45902
rect 22204 45798 22260 45836
rect 21868 45602 21924 45612
rect 22316 45666 22372 45678
rect 22316 45614 22318 45666
rect 22370 45614 22372 45666
rect 20524 45054 20526 45106
rect 20578 45054 20580 45106
rect 20524 45042 20580 45054
rect 21420 45276 21812 45332
rect 22316 45332 22372 45614
rect 20300 44436 20356 44446
rect 20300 44434 21364 44436
rect 20300 44382 20302 44434
rect 20354 44382 21364 44434
rect 20300 44380 21364 44382
rect 20300 44370 20356 44380
rect 21308 44322 21364 44380
rect 21308 44270 21310 44322
rect 21362 44270 21364 44322
rect 21308 44258 21364 44270
rect 20412 44212 20468 44222
rect 20188 44098 20244 44110
rect 20188 44046 20190 44098
rect 20242 44046 20244 44098
rect 20188 43540 20244 44046
rect 20412 43762 20468 44156
rect 21420 44100 21476 45276
rect 22316 45266 22372 45276
rect 21756 45108 21812 45118
rect 21756 44434 21812 45052
rect 21756 44382 21758 44434
rect 21810 44382 21812 44434
rect 21756 44370 21812 44382
rect 22316 44996 22372 45006
rect 21980 44324 22036 44334
rect 21980 44230 22036 44268
rect 21308 44044 21476 44100
rect 21532 44210 21588 44222
rect 21532 44158 21534 44210
rect 21586 44158 21588 44210
rect 20412 43710 20414 43762
rect 20466 43710 20468 43762
rect 20412 43698 20468 43710
rect 20972 43764 21028 43774
rect 20972 43670 21028 43708
rect 20188 43474 20244 43484
rect 20748 42756 20804 42766
rect 20748 42662 20804 42700
rect 20188 42532 20244 42542
rect 20076 42476 20188 42532
rect 20188 42438 20244 42476
rect 20972 42532 21028 42542
rect 19964 42130 20020 42140
rect 20748 42196 20804 42206
rect 19964 41860 20020 41870
rect 19292 41858 20020 41860
rect 19292 41806 19966 41858
rect 20018 41806 20020 41858
rect 19292 41804 20020 41806
rect 19180 41692 19460 41748
rect 18732 41246 18734 41298
rect 18786 41246 18788 41298
rect 18732 41234 18788 41246
rect 18284 38894 18286 38946
rect 18338 38894 18340 38946
rect 16828 38836 16884 38846
rect 16828 38722 16884 38780
rect 17388 38836 17444 38846
rect 17388 38742 17444 38780
rect 17948 38834 18004 38846
rect 17948 38782 17950 38834
rect 18002 38782 18004 38834
rect 16828 38670 16830 38722
rect 16882 38670 16884 38722
rect 16828 38658 16884 38670
rect 17948 38724 18004 38782
rect 17948 38658 18004 38668
rect 17612 38500 17668 38510
rect 16716 37490 16884 37492
rect 16716 37438 16718 37490
rect 16770 37438 16884 37490
rect 16716 37436 16884 37438
rect 16716 37426 16772 37436
rect 16828 37380 16884 37436
rect 16828 37314 16884 37324
rect 16492 37268 16548 37278
rect 16492 37174 16548 37212
rect 17500 37266 17556 37278
rect 17500 37214 17502 37266
rect 17554 37214 17556 37266
rect 16828 37156 16884 37166
rect 16828 37062 16884 37100
rect 17500 37156 17556 37214
rect 17500 37090 17556 37100
rect 16380 35812 16436 35822
rect 16380 35718 16436 35756
rect 17052 35364 17108 35374
rect 16940 34804 16996 34814
rect 16716 34692 16772 34702
rect 16772 34636 16884 34692
rect 16716 34598 16772 34636
rect 16716 34356 16772 34366
rect 16268 34354 16660 34356
rect 16268 34302 16270 34354
rect 16322 34302 16660 34354
rect 16268 34300 16660 34302
rect 16268 34290 16324 34300
rect 16604 34242 16660 34300
rect 16716 34262 16772 34300
rect 16604 34190 16606 34242
rect 16658 34190 16660 34242
rect 16492 34132 16548 34142
rect 13468 33842 13524 33852
rect 16380 33908 16436 33918
rect 16380 33570 16436 33852
rect 16380 33518 16382 33570
rect 16434 33518 16436 33570
rect 16380 33506 16436 33518
rect 15372 33460 15428 33470
rect 13916 33348 13972 33358
rect 13916 33254 13972 33292
rect 14140 33234 14196 33246
rect 14140 33182 14142 33234
rect 14194 33182 14196 33234
rect 13580 33122 13636 33134
rect 14140 33124 14196 33182
rect 13580 33070 13582 33122
rect 13634 33070 13636 33122
rect 13580 32564 13636 33070
rect 13580 32498 13636 32508
rect 13804 33068 14196 33124
rect 14476 33234 14532 33246
rect 14476 33182 14478 33234
rect 14530 33182 14532 33234
rect 14476 33124 14532 33182
rect 13804 32002 13860 33068
rect 14476 33058 14532 33068
rect 14008 32956 15208 32966
rect 14064 32954 14112 32956
rect 14168 32954 14216 32956
rect 14076 32902 14112 32954
rect 14200 32902 14216 32954
rect 14064 32900 14112 32902
rect 14168 32900 14216 32902
rect 14272 32954 14320 32956
rect 14376 32954 14424 32956
rect 14480 32954 14528 32956
rect 14376 32902 14396 32954
rect 14480 32902 14520 32954
rect 14272 32900 14320 32902
rect 14376 32900 14424 32902
rect 14480 32900 14528 32902
rect 14584 32900 14632 32956
rect 14688 32954 14736 32956
rect 14792 32954 14840 32956
rect 14896 32954 14944 32956
rect 14696 32902 14736 32954
rect 14820 32902 14840 32954
rect 14688 32900 14736 32902
rect 14792 32900 14840 32902
rect 14896 32900 14944 32902
rect 15000 32954 15048 32956
rect 15104 32954 15152 32956
rect 15000 32902 15016 32954
rect 15104 32902 15140 32954
rect 15000 32900 15048 32902
rect 15104 32900 15152 32902
rect 14008 32890 15208 32900
rect 13804 31950 13806 32002
rect 13858 31950 13860 32002
rect 13804 31938 13860 31950
rect 14476 32788 14532 32798
rect 14476 32004 14532 32732
rect 15372 32788 15428 33404
rect 16268 33348 16324 33358
rect 16044 33292 16268 33348
rect 15932 33122 15988 33134
rect 15932 33070 15934 33122
rect 15986 33070 15988 33122
rect 15932 33012 15988 33070
rect 15372 32694 15428 32732
rect 15820 32956 15932 33012
rect 15820 32452 15876 32956
rect 15932 32946 15988 32956
rect 15932 32788 15988 32798
rect 16044 32788 16100 33292
rect 16268 33254 16324 33292
rect 16380 33122 16436 33134
rect 16380 33070 16382 33122
rect 16434 33070 16436 33122
rect 16380 33012 16436 33070
rect 15932 32786 16100 32788
rect 15932 32734 15934 32786
rect 15986 32734 16100 32786
rect 15932 32732 16100 32734
rect 16268 32788 16324 32798
rect 15932 32722 15988 32732
rect 16268 32694 16324 32732
rect 15820 32386 15876 32396
rect 14588 32004 14644 32014
rect 14476 32002 14644 32004
rect 14476 31950 14590 32002
rect 14642 31950 14644 32002
rect 14476 31948 14644 31950
rect 14588 31938 14644 31948
rect 16268 32002 16324 32014
rect 16268 31950 16270 32002
rect 16322 31950 16324 32002
rect 16268 31890 16324 31950
rect 16268 31838 16270 31890
rect 16322 31838 16324 31890
rect 16268 31826 16324 31838
rect 13020 31714 13076 31724
rect 14924 31778 14980 31790
rect 14924 31726 14926 31778
rect 14978 31726 14980 31778
rect 13468 31666 13524 31678
rect 13468 31614 13470 31666
rect 13522 31614 13524 31666
rect 13356 30884 13412 30894
rect 13020 30212 13076 30222
rect 13020 28868 13076 30156
rect 13356 30212 13412 30828
rect 13356 30146 13412 30156
rect 13468 30100 13524 31614
rect 13692 31668 13748 31678
rect 13692 31574 13748 31612
rect 14140 31668 14196 31678
rect 14140 31556 14196 31612
rect 14924 31668 14980 31726
rect 15708 31780 15764 31790
rect 15708 31778 15876 31780
rect 15708 31726 15710 31778
rect 15762 31726 15876 31778
rect 15708 31724 15876 31726
rect 15708 31714 15764 31724
rect 15596 31668 15652 31678
rect 14924 31602 14980 31612
rect 15372 31612 15596 31668
rect 13804 31554 14196 31556
rect 13804 31502 14142 31554
rect 14194 31502 14196 31554
rect 13804 31500 14196 31502
rect 13692 31108 13748 31118
rect 13804 31108 13860 31500
rect 14140 31490 14196 31500
rect 14008 31388 15208 31398
rect 14064 31386 14112 31388
rect 14168 31386 14216 31388
rect 14076 31334 14112 31386
rect 14200 31334 14216 31386
rect 14064 31332 14112 31334
rect 14168 31332 14216 31334
rect 14272 31386 14320 31388
rect 14376 31386 14424 31388
rect 14480 31386 14528 31388
rect 14376 31334 14396 31386
rect 14480 31334 14520 31386
rect 14272 31332 14320 31334
rect 14376 31332 14424 31334
rect 14480 31332 14528 31334
rect 14584 31332 14632 31388
rect 14688 31386 14736 31388
rect 14792 31386 14840 31388
rect 14896 31386 14944 31388
rect 14696 31334 14736 31386
rect 14820 31334 14840 31386
rect 14688 31332 14736 31334
rect 14792 31332 14840 31334
rect 14896 31332 14944 31334
rect 15000 31386 15048 31388
rect 15104 31386 15152 31388
rect 15000 31334 15016 31386
rect 15104 31334 15140 31386
rect 15000 31332 15048 31334
rect 15104 31332 15152 31334
rect 14008 31322 15208 31332
rect 15260 31220 15316 31230
rect 15372 31220 15428 31612
rect 15596 31574 15652 31612
rect 15260 31218 15428 31220
rect 15260 31166 15262 31218
rect 15314 31166 15428 31218
rect 15260 31164 15428 31166
rect 15820 31556 15876 31724
rect 15260 31154 15316 31164
rect 13748 31052 13860 31108
rect 15596 31108 15652 31118
rect 15596 31106 15764 31108
rect 15596 31054 15598 31106
rect 15650 31054 15764 31106
rect 15596 31052 15764 31054
rect 13692 31042 13748 31052
rect 15596 31042 15652 31052
rect 15484 30996 15540 31006
rect 15372 30994 15540 30996
rect 15372 30942 15486 30994
rect 15538 30942 15540 30994
rect 15372 30940 15540 30942
rect 14364 30882 14420 30894
rect 14364 30830 14366 30882
rect 14418 30830 14420 30882
rect 14364 30772 14420 30830
rect 14252 30212 14308 30222
rect 14252 30118 14308 30156
rect 13468 28980 13524 30044
rect 14364 29988 14420 30716
rect 14700 30882 14756 30894
rect 14700 30830 14702 30882
rect 14754 30830 14756 30882
rect 14700 30324 14756 30830
rect 14700 30258 14756 30268
rect 14364 29922 14420 29932
rect 14008 29820 15208 29830
rect 14064 29818 14112 29820
rect 14168 29818 14216 29820
rect 14076 29766 14112 29818
rect 14200 29766 14216 29818
rect 14064 29764 14112 29766
rect 14168 29764 14216 29766
rect 14272 29818 14320 29820
rect 14376 29818 14424 29820
rect 14480 29818 14528 29820
rect 14376 29766 14396 29818
rect 14480 29766 14520 29818
rect 14272 29764 14320 29766
rect 14376 29764 14424 29766
rect 14480 29764 14528 29766
rect 14584 29764 14632 29820
rect 14688 29818 14736 29820
rect 14792 29818 14840 29820
rect 14896 29818 14944 29820
rect 14696 29766 14736 29818
rect 14820 29766 14840 29818
rect 14688 29764 14736 29766
rect 14792 29764 14840 29766
rect 14896 29764 14944 29766
rect 15000 29818 15048 29820
rect 15104 29818 15152 29820
rect 15000 29766 15016 29818
rect 15104 29766 15140 29818
rect 15000 29764 15048 29766
rect 15104 29764 15152 29766
rect 14008 29754 15208 29764
rect 14476 29652 14532 29662
rect 15372 29652 15428 30940
rect 15484 30930 15540 30940
rect 15596 30772 15652 30782
rect 15596 30678 15652 30716
rect 15596 30324 15652 30334
rect 15708 30324 15764 31052
rect 15652 30268 15764 30324
rect 15596 30258 15652 30268
rect 15708 29988 15764 29998
rect 14476 29558 14532 29596
rect 15036 29596 15428 29652
rect 15596 29652 15652 29662
rect 13804 29540 13860 29550
rect 13468 28914 13524 28924
rect 13580 29428 13636 29438
rect 13020 28866 13412 28868
rect 13020 28814 13022 28866
rect 13074 28814 13412 28866
rect 13020 28812 13412 28814
rect 13020 28802 13076 28812
rect 13356 28644 13412 28812
rect 13580 28866 13636 29372
rect 13580 28814 13582 28866
rect 13634 28814 13636 28866
rect 13580 28802 13636 28814
rect 13356 28588 13636 28644
rect 13132 28420 13188 28430
rect 12684 27970 12740 27982
rect 12684 27918 12686 27970
rect 12738 27918 12740 27970
rect 12684 27860 12740 27918
rect 12684 27794 12740 27804
rect 13132 27970 13188 28364
rect 13132 27918 13134 27970
rect 13186 27918 13188 27970
rect 12516 27468 12628 27524
rect 12460 27458 12516 27468
rect 11564 27122 11620 27132
rect 13020 27188 13076 27198
rect 13132 27188 13188 27918
rect 13020 27186 13188 27188
rect 13020 27134 13022 27186
rect 13074 27134 13188 27186
rect 13020 27132 13188 27134
rect 13468 28308 13524 28318
rect 13020 27122 13076 27132
rect 12236 26964 12292 26974
rect 9996 25732 10052 25742
rect 9884 25730 10052 25732
rect 9884 25678 9998 25730
rect 10050 25678 10052 25730
rect 9884 25676 10052 25678
rect 8876 25666 8932 25676
rect 9996 25666 10052 25676
rect 10220 25394 10276 25406
rect 10556 25396 10612 25406
rect 10220 25342 10222 25394
rect 10274 25342 10276 25394
rect 9212 25284 9268 25294
rect 9212 25190 9268 25228
rect 9660 25284 9716 25294
rect 10220 25284 10276 25342
rect 9660 25282 10052 25284
rect 9660 25230 9662 25282
rect 9714 25230 10052 25282
rect 9660 25228 10052 25230
rect 9660 25218 9716 25228
rect 8540 24894 8542 24946
rect 8594 24894 8596 24946
rect 7756 22978 7812 22988
rect 7308 22418 7364 22428
rect 6748 21812 6804 21822
rect 6748 20914 6804 21756
rect 6972 21700 7028 21710
rect 6972 21606 7028 21644
rect 6860 21588 6916 21598
rect 6860 21494 6916 21532
rect 7532 21588 7588 21598
rect 7532 21494 7588 21532
rect 6748 20862 6750 20914
rect 6802 20862 6804 20914
rect 6748 20692 6804 20862
rect 6748 20626 6804 20636
rect 6636 20580 6692 20590
rect 6636 14868 6692 20524
rect 7420 18788 7476 18798
rect 7084 17556 7140 17566
rect 6972 16884 7028 16894
rect 6972 16790 7028 16828
rect 6860 16772 6916 16782
rect 6860 16678 6916 16716
rect 7084 16098 7140 17500
rect 7420 17106 7476 18732
rect 7420 17054 7422 17106
rect 7474 17054 7476 17106
rect 7420 17042 7476 17054
rect 7196 16884 7252 16894
rect 7196 16882 7588 16884
rect 7196 16830 7198 16882
rect 7250 16830 7588 16882
rect 7196 16828 7588 16830
rect 7196 16818 7252 16828
rect 7420 16436 7476 16446
rect 7084 16046 7086 16098
rect 7138 16046 7140 16098
rect 7084 16034 7140 16046
rect 7196 16380 7420 16436
rect 7196 15652 7252 16380
rect 7420 16370 7476 16380
rect 7084 15596 7252 15652
rect 7420 16210 7476 16222
rect 7420 16158 7422 16210
rect 7474 16158 7476 16210
rect 6860 15316 6916 15326
rect 7084 15316 7140 15596
rect 7308 15540 7364 15550
rect 7196 15428 7252 15438
rect 7196 15334 7252 15372
rect 6860 15314 7140 15316
rect 6860 15262 6862 15314
rect 6914 15262 7140 15314
rect 6860 15260 7140 15262
rect 6860 15250 6916 15260
rect 7084 15148 7140 15260
rect 6972 15092 7028 15102
rect 7084 15092 7252 15148
rect 6972 14998 7028 15036
rect 6636 14812 7140 14868
rect 6524 14690 6580 14700
rect 6972 14642 7028 14654
rect 6972 14590 6974 14642
rect 7026 14590 7028 14642
rect 6972 14532 7028 14590
rect 6412 14476 7028 14532
rect 6412 14420 6468 14476
rect 6412 14354 6468 14364
rect 6972 13972 7028 14476
rect 7084 14530 7140 14812
rect 7084 14478 7086 14530
rect 7138 14478 7140 14530
rect 7084 14084 7140 14478
rect 7196 14420 7252 15092
rect 7196 14354 7252 14364
rect 7084 14028 7252 14084
rect 6972 13916 7140 13972
rect 6972 13748 7028 13758
rect 6524 13076 6580 13086
rect 6300 13020 6524 13076
rect 4060 12114 4116 12124
rect 5292 12180 5348 12190
rect 4008 11788 5208 11798
rect 4064 11786 4112 11788
rect 4168 11786 4216 11788
rect 4076 11734 4112 11786
rect 4200 11734 4216 11786
rect 4064 11732 4112 11734
rect 4168 11732 4216 11734
rect 4272 11786 4320 11788
rect 4376 11786 4424 11788
rect 4480 11786 4528 11788
rect 4376 11734 4396 11786
rect 4480 11734 4520 11786
rect 4272 11732 4320 11734
rect 4376 11732 4424 11734
rect 4480 11732 4528 11734
rect 4584 11732 4632 11788
rect 4688 11786 4736 11788
rect 4792 11786 4840 11788
rect 4896 11786 4944 11788
rect 4696 11734 4736 11786
rect 4820 11734 4840 11786
rect 4688 11732 4736 11734
rect 4792 11732 4840 11734
rect 4896 11732 4944 11734
rect 5000 11786 5048 11788
rect 5104 11786 5152 11788
rect 5000 11734 5016 11786
rect 5104 11734 5140 11786
rect 5000 11732 5048 11734
rect 5104 11732 5152 11734
rect 4008 11722 5208 11732
rect 3724 11618 3892 11620
rect 3724 11566 3726 11618
rect 3778 11566 3892 11618
rect 3724 11564 3892 11566
rect 3724 11554 3780 11564
rect 4396 11508 4452 11518
rect 4396 11394 4452 11452
rect 5068 11508 5124 11518
rect 5068 11414 5124 11452
rect 4396 11342 4398 11394
rect 4450 11342 4452 11394
rect 4396 11330 4452 11342
rect 4508 11396 4564 11406
rect 4508 11282 4564 11340
rect 4508 11230 4510 11282
rect 4562 11230 4564 11282
rect 4508 11218 4564 11230
rect 4732 10836 4788 10846
rect 4732 10742 4788 10780
rect 5292 10834 5348 12124
rect 5516 12068 5572 12078
rect 5404 11954 5460 11966
rect 5404 11902 5406 11954
rect 5458 11902 5460 11954
rect 5404 11396 5460 11902
rect 5404 11330 5460 11340
rect 5292 10782 5294 10834
rect 5346 10782 5348 10834
rect 5292 10770 5348 10782
rect 5404 10836 5460 10846
rect 5516 10836 5572 12012
rect 5740 11788 5796 12348
rect 6076 12404 6132 12414
rect 6076 12310 6132 12348
rect 6524 12178 6580 13020
rect 6972 12964 7028 13692
rect 6524 12126 6526 12178
rect 6578 12126 6580 12178
rect 6524 12114 6580 12126
rect 6748 12962 7028 12964
rect 6748 12910 6974 12962
rect 7026 12910 7028 12962
rect 6748 12908 7028 12910
rect 6748 12404 6804 12908
rect 6972 12898 7028 12908
rect 7084 13636 7140 13916
rect 7196 13748 7252 14028
rect 7196 13682 7252 13692
rect 6748 12178 6804 12348
rect 7084 12850 7140 13580
rect 7196 13076 7252 13086
rect 7196 12962 7252 13020
rect 7196 12910 7198 12962
rect 7250 12910 7252 12962
rect 7196 12898 7252 12910
rect 7084 12798 7086 12850
rect 7138 12798 7140 12850
rect 6860 12292 6916 12302
rect 6860 12198 6916 12236
rect 6748 12126 6750 12178
rect 6802 12126 6804 12178
rect 6748 12114 6804 12126
rect 7084 12178 7140 12798
rect 7084 12126 7086 12178
rect 7138 12126 7140 12178
rect 7084 12068 7140 12126
rect 7084 12002 7140 12012
rect 7308 12068 7364 15484
rect 7420 13188 7476 16158
rect 7532 15540 7588 16828
rect 7980 16772 8036 24892
rect 8092 24724 8148 24734
rect 8540 24724 8596 24894
rect 8092 24722 8596 24724
rect 8092 24670 8094 24722
rect 8146 24670 8596 24722
rect 8092 24668 8596 24670
rect 8988 24724 9044 24734
rect 8092 23042 8148 24668
rect 8988 24630 9044 24668
rect 9996 24722 10052 25228
rect 10220 25218 10276 25228
rect 10332 25394 10612 25396
rect 10332 25342 10558 25394
rect 10610 25342 10612 25394
rect 10332 25340 10612 25342
rect 9996 24670 9998 24722
rect 10050 24670 10052 24722
rect 9996 24658 10052 24670
rect 8316 24500 8372 24510
rect 8316 23938 8372 24444
rect 9660 24500 9716 24510
rect 9660 24406 9716 24444
rect 8316 23886 8318 23938
rect 8370 23886 8372 23938
rect 8316 23874 8372 23886
rect 8092 22990 8094 23042
rect 8146 22990 8148 23042
rect 8092 22978 8148 22990
rect 9660 23156 9716 23166
rect 8540 22146 8596 22158
rect 9212 22148 9268 22158
rect 8540 22094 8542 22146
rect 8594 22094 8596 22146
rect 8428 21812 8484 21822
rect 8428 21718 8484 21756
rect 8428 20804 8484 20814
rect 8428 20710 8484 20748
rect 8540 17668 8596 22094
rect 8764 22146 9268 22148
rect 8764 22094 9214 22146
rect 9266 22094 9268 22146
rect 8764 22092 9268 22094
rect 8764 21700 8820 22092
rect 9212 22082 9268 22092
rect 9548 22146 9604 22158
rect 9548 22094 9550 22146
rect 9602 22094 9604 22146
rect 8876 21812 8932 21822
rect 8876 21718 8932 21756
rect 8764 21606 8820 21644
rect 8876 21362 8932 21374
rect 8876 21310 8878 21362
rect 8930 21310 8932 21362
rect 8540 17442 8596 17612
rect 8764 20580 8820 20590
rect 8540 17390 8542 17442
rect 8594 17390 8596 17442
rect 8540 17378 8596 17390
rect 8652 17444 8708 17454
rect 8652 17108 8708 17388
rect 8540 17106 8708 17108
rect 8540 17054 8654 17106
rect 8706 17054 8708 17106
rect 8540 17052 8708 17054
rect 8428 16996 8484 17006
rect 8204 16882 8260 16894
rect 8204 16830 8206 16882
rect 8258 16830 8260 16882
rect 8092 16772 8148 16782
rect 7980 16716 8092 16772
rect 8092 16706 8148 16716
rect 7756 16660 7812 16670
rect 7756 16566 7812 16604
rect 7868 16658 7924 16670
rect 7868 16606 7870 16658
rect 7922 16606 7924 16658
rect 7868 16436 7924 16606
rect 8204 16548 8260 16830
rect 8316 16660 8372 16670
rect 8316 16566 8372 16604
rect 7868 16370 7924 16380
rect 7980 16492 8260 16548
rect 7756 16212 7812 16222
rect 7980 16212 8036 16492
rect 7756 16210 8036 16212
rect 7756 16158 7758 16210
rect 7810 16158 8036 16210
rect 7756 16156 8036 16158
rect 7756 16146 7812 16156
rect 7532 15426 7588 15484
rect 7532 15374 7534 15426
rect 7586 15374 7588 15426
rect 7532 15362 7588 15374
rect 8092 15484 8372 15540
rect 7756 15314 7812 15326
rect 7756 15262 7758 15314
rect 7810 15262 7812 15314
rect 7756 15148 7812 15262
rect 7644 15092 7812 15148
rect 7868 15204 7924 15214
rect 8092 15204 8148 15484
rect 7868 15202 8148 15204
rect 7868 15150 7870 15202
rect 7922 15150 8148 15202
rect 7868 15148 8148 15150
rect 8204 15314 8260 15326
rect 8204 15262 8206 15314
rect 8258 15262 8260 15314
rect 7868 15138 7924 15148
rect 7644 14308 7700 15092
rect 7756 14644 7812 14654
rect 8204 14644 8260 15262
rect 7756 14642 8260 14644
rect 7756 14590 7758 14642
rect 7810 14590 8260 14642
rect 7756 14588 8260 14590
rect 7756 14578 7812 14588
rect 8204 14420 8260 14430
rect 8204 14326 8260 14364
rect 7644 14252 8148 14308
rect 8092 13970 8148 14252
rect 8092 13918 8094 13970
rect 8146 13918 8148 13970
rect 8092 13906 8148 13918
rect 7756 13748 7812 13758
rect 7756 13654 7812 13692
rect 8204 13636 8260 13646
rect 8204 13542 8260 13580
rect 8316 13524 8372 15484
rect 8428 15538 8484 16940
rect 8428 15486 8430 15538
rect 8482 15486 8484 15538
rect 8428 15148 8484 15486
rect 8540 15540 8596 17052
rect 8652 17042 8708 17052
rect 8764 16884 8820 20524
rect 8876 20020 8932 21310
rect 9100 20804 9156 20814
rect 9548 20804 9604 22094
rect 9660 21586 9716 23100
rect 9660 21534 9662 21586
rect 9714 21534 9716 21586
rect 9660 21522 9716 21534
rect 9996 22146 10052 22158
rect 9996 22094 9998 22146
rect 10050 22094 10052 22146
rect 9100 20710 9156 20748
rect 9436 20748 9604 20804
rect 9772 20804 9828 20814
rect 9324 20692 9380 20702
rect 9324 20598 9380 20636
rect 8876 19954 8932 19964
rect 9436 17780 9492 20748
rect 9548 20580 9604 20590
rect 9548 20486 9604 20524
rect 9660 20578 9716 20590
rect 9660 20526 9662 20578
rect 9714 20526 9716 20578
rect 9660 20132 9716 20526
rect 9660 20066 9716 20076
rect 9548 17780 9604 17790
rect 9436 17778 9604 17780
rect 9436 17726 9550 17778
rect 9602 17726 9604 17778
rect 9436 17724 9604 17726
rect 9212 17556 9268 17566
rect 9212 17462 9268 17500
rect 8876 16884 8932 16894
rect 8764 16882 9156 16884
rect 8764 16830 8878 16882
rect 8930 16830 9156 16882
rect 8764 16828 9156 16830
rect 8876 16818 8932 16828
rect 8652 16212 8708 16222
rect 8652 16098 8708 16156
rect 8652 16046 8654 16098
rect 8706 16046 8708 16098
rect 8652 16034 8708 16046
rect 8652 15540 8708 15550
rect 8540 15538 9044 15540
rect 8540 15486 8654 15538
rect 8706 15486 9044 15538
rect 8540 15484 9044 15486
rect 8652 15474 8708 15484
rect 8876 15314 8932 15326
rect 8876 15262 8878 15314
rect 8930 15262 8932 15314
rect 8428 15092 8708 15148
rect 8428 14532 8484 14542
rect 8428 14438 8484 14476
rect 8652 14420 8708 15092
rect 8764 15092 8820 15102
rect 8764 14998 8820 15036
rect 8876 14980 8932 15262
rect 8764 14420 8820 14430
rect 8652 14364 8764 14420
rect 8764 14326 8820 14364
rect 8876 13860 8932 14924
rect 8988 14420 9044 15484
rect 9100 14980 9156 16828
rect 9100 14914 9156 14924
rect 9436 16210 9492 17724
rect 9548 17714 9604 17724
rect 9660 17556 9716 17566
rect 9660 16994 9716 17500
rect 9660 16942 9662 16994
rect 9714 16942 9716 16994
rect 9660 16930 9716 16942
rect 9548 16884 9604 16894
rect 9548 16790 9604 16828
rect 9436 16158 9438 16210
rect 9490 16158 9492 16210
rect 9212 14530 9268 14542
rect 9212 14478 9214 14530
rect 9266 14478 9268 14530
rect 9100 14420 9156 14430
rect 8988 14418 9156 14420
rect 8988 14366 9102 14418
rect 9154 14366 9156 14418
rect 8988 14364 9156 14366
rect 9100 13972 9156 14364
rect 9100 13906 9156 13916
rect 8876 13804 9044 13860
rect 8988 13748 9044 13804
rect 9100 13748 9156 13758
rect 8988 13746 9156 13748
rect 8988 13694 9102 13746
rect 9154 13694 9156 13746
rect 8988 13692 9156 13694
rect 9100 13682 9156 13692
rect 8540 13636 8596 13646
rect 8316 13468 8484 13524
rect 7644 13188 7700 13198
rect 7420 13186 7812 13188
rect 7420 13134 7646 13186
rect 7698 13134 7812 13186
rect 7420 13132 7812 13134
rect 7644 13122 7700 13132
rect 7420 12292 7476 12302
rect 7476 12236 7588 12292
rect 7420 12226 7476 12236
rect 7532 12178 7588 12236
rect 7532 12126 7534 12178
rect 7586 12126 7588 12178
rect 7532 12114 7588 12126
rect 7756 12178 7812 13132
rect 8316 12962 8372 12974
rect 8316 12910 8318 12962
rect 8370 12910 8372 12962
rect 8204 12740 8260 12750
rect 8204 12402 8260 12684
rect 8204 12350 8206 12402
rect 8258 12350 8260 12402
rect 8204 12338 8260 12350
rect 7756 12126 7758 12178
rect 7810 12126 7812 12178
rect 7756 12114 7812 12126
rect 7364 12012 7476 12068
rect 7308 11974 7364 12012
rect 6972 11956 7028 11966
rect 5740 11732 6020 11788
rect 5404 10834 5572 10836
rect 5404 10782 5406 10834
rect 5458 10782 5572 10834
rect 5404 10780 5572 10782
rect 5740 11172 5796 11182
rect 5404 10770 5460 10780
rect 4008 10220 5208 10230
rect 4064 10218 4112 10220
rect 4168 10218 4216 10220
rect 4076 10166 4112 10218
rect 4200 10166 4216 10218
rect 4064 10164 4112 10166
rect 4168 10164 4216 10166
rect 4272 10218 4320 10220
rect 4376 10218 4424 10220
rect 4480 10218 4528 10220
rect 4376 10166 4396 10218
rect 4480 10166 4520 10218
rect 4272 10164 4320 10166
rect 4376 10164 4424 10166
rect 4480 10164 4528 10166
rect 4584 10164 4632 10220
rect 4688 10218 4736 10220
rect 4792 10218 4840 10220
rect 4896 10218 4944 10220
rect 4696 10166 4736 10218
rect 4820 10166 4840 10218
rect 4688 10164 4736 10166
rect 4792 10164 4840 10166
rect 4896 10164 4944 10166
rect 5000 10218 5048 10220
rect 5104 10218 5152 10220
rect 5000 10166 5016 10218
rect 5104 10166 5140 10218
rect 5000 10164 5048 10166
rect 5104 10164 5152 10166
rect 4008 10154 5208 10164
rect 5740 9602 5796 11116
rect 5964 10836 6020 11732
rect 6972 11618 7028 11900
rect 6972 11566 6974 11618
rect 7026 11566 7028 11618
rect 6972 11554 7028 11566
rect 7420 11508 7476 12012
rect 8316 11956 8372 12910
rect 8316 11890 8372 11900
rect 7532 11508 7588 11518
rect 7084 11506 7588 11508
rect 7084 11454 7534 11506
rect 7586 11454 7588 11506
rect 7084 11452 7588 11454
rect 6860 11396 6916 11406
rect 6860 11302 6916 11340
rect 6972 11284 7028 11294
rect 7084 11284 7140 11452
rect 7532 11442 7588 11452
rect 6972 11282 7140 11284
rect 6972 11230 6974 11282
rect 7026 11230 7140 11282
rect 6972 11228 7140 11230
rect 7980 11394 8036 11406
rect 7980 11342 7982 11394
rect 8034 11342 8036 11394
rect 6972 11218 7028 11228
rect 7980 11172 8036 11342
rect 7980 11106 8036 11116
rect 6020 10780 6244 10836
rect 5964 10742 6020 10780
rect 6188 9940 6244 10780
rect 8428 10610 8484 13468
rect 8540 12402 8596 13580
rect 9212 13636 9268 14478
rect 9212 13570 9268 13580
rect 9324 13188 9380 13198
rect 8876 13186 9380 13188
rect 8876 13134 9326 13186
rect 9378 13134 9380 13186
rect 8876 13132 9380 13134
rect 8764 13076 8820 13086
rect 8540 12350 8542 12402
rect 8594 12350 8596 12402
rect 8540 12338 8596 12350
rect 8652 13074 8820 13076
rect 8652 13022 8766 13074
rect 8818 13022 8820 13074
rect 8652 13020 8820 13022
rect 8652 11394 8708 13020
rect 8764 13010 8820 13020
rect 8764 12852 8820 12862
rect 8764 12758 8820 12796
rect 8876 12850 8932 13132
rect 9324 13122 9380 13132
rect 8876 12798 8878 12850
rect 8930 12798 8932 12850
rect 8876 12786 8932 12798
rect 9100 12740 9156 12750
rect 9100 12646 9156 12684
rect 8988 12404 9044 12414
rect 8988 12068 9044 12348
rect 8988 12002 9044 12012
rect 8652 11342 8654 11394
rect 8706 11342 8708 11394
rect 8652 11330 8708 11342
rect 8428 10558 8430 10610
rect 8482 10558 8484 10610
rect 8428 10546 8484 10558
rect 8876 11172 8932 11182
rect 9436 11172 9492 16158
rect 9660 15540 9716 15550
rect 9660 15446 9716 15484
rect 9772 15538 9828 20748
rect 9884 20020 9940 20030
rect 9884 19926 9940 19964
rect 9996 17668 10052 22094
rect 10108 21586 10164 21598
rect 10108 21534 10110 21586
rect 10162 21534 10164 21586
rect 10108 19908 10164 21534
rect 10332 21364 10388 25340
rect 10556 25330 10612 25340
rect 10780 24836 10836 24846
rect 10780 24834 11396 24836
rect 10780 24782 10782 24834
rect 10834 24782 11396 24834
rect 10780 24780 11396 24782
rect 10780 24770 10836 24780
rect 10556 24724 10612 24734
rect 10556 22596 10612 24668
rect 10780 24388 10836 24398
rect 10780 23714 10836 24332
rect 11340 24164 11396 24780
rect 11564 24610 11620 24622
rect 11564 24558 11566 24610
rect 11618 24558 11620 24610
rect 11564 24388 11620 24558
rect 11564 24322 11620 24332
rect 11340 24162 11620 24164
rect 11340 24110 11342 24162
rect 11394 24110 11620 24162
rect 11340 24108 11620 24110
rect 11340 24098 11396 24108
rect 11564 23938 11620 24108
rect 11564 23886 11566 23938
rect 11618 23886 11620 23938
rect 11564 23874 11620 23886
rect 11676 23828 11732 23838
rect 11676 23734 11732 23772
rect 12236 23828 12292 26908
rect 12572 25284 12628 25294
rect 12572 24946 12628 25228
rect 13468 25172 13524 28252
rect 13580 27972 13636 28588
rect 13580 27906 13636 27916
rect 13692 28532 13748 28542
rect 13692 27748 13748 28476
rect 13692 27186 13748 27692
rect 13692 27134 13694 27186
rect 13746 27134 13748 27186
rect 13692 27122 13748 27134
rect 13804 27188 13860 29484
rect 14700 29204 14756 29214
rect 13916 29092 13972 29102
rect 13916 28866 13972 29036
rect 13916 28814 13918 28866
rect 13970 28814 13972 28866
rect 13916 28802 13972 28814
rect 14364 28644 14420 28654
rect 14364 28550 14420 28588
rect 14700 28530 14756 29148
rect 15036 29202 15092 29596
rect 15036 29150 15038 29202
rect 15090 29150 15092 29202
rect 14924 29092 14980 29102
rect 15036 29092 15092 29150
rect 15372 29204 15428 29214
rect 15372 29110 15428 29148
rect 14980 29036 15092 29092
rect 14924 29026 14980 29036
rect 14700 28478 14702 28530
rect 14754 28478 14756 28530
rect 14700 28466 14756 28478
rect 15484 28644 15540 28654
rect 15260 28420 15316 28458
rect 15260 28354 15316 28364
rect 14008 28252 15208 28262
rect 14064 28250 14112 28252
rect 14168 28250 14216 28252
rect 14076 28198 14112 28250
rect 14200 28198 14216 28250
rect 14064 28196 14112 28198
rect 14168 28196 14216 28198
rect 14272 28250 14320 28252
rect 14376 28250 14424 28252
rect 14480 28250 14528 28252
rect 14376 28198 14396 28250
rect 14480 28198 14520 28250
rect 14272 28196 14320 28198
rect 14376 28196 14424 28198
rect 14480 28196 14528 28198
rect 14584 28196 14632 28252
rect 14688 28250 14736 28252
rect 14792 28250 14840 28252
rect 14896 28250 14944 28252
rect 14696 28198 14736 28250
rect 14820 28198 14840 28250
rect 14688 28196 14736 28198
rect 14792 28196 14840 28198
rect 14896 28196 14944 28198
rect 15000 28250 15048 28252
rect 15104 28250 15152 28252
rect 15000 28198 15016 28250
rect 15104 28198 15140 28250
rect 15000 28196 15048 28198
rect 15104 28196 15152 28198
rect 14008 28186 15208 28196
rect 15484 28082 15540 28588
rect 15596 28420 15652 29596
rect 15708 29426 15764 29932
rect 15820 29540 15876 31500
rect 16268 31220 16324 31230
rect 16380 31220 16436 32956
rect 16268 31218 16380 31220
rect 16268 31166 16270 31218
rect 16322 31166 16380 31218
rect 16268 31164 16380 31166
rect 16268 31154 16324 31164
rect 16380 31126 16436 31164
rect 16044 30324 16100 30334
rect 15932 29540 15988 29550
rect 15820 29538 15988 29540
rect 15820 29486 15934 29538
rect 15986 29486 15988 29538
rect 15820 29484 15988 29486
rect 15932 29474 15988 29484
rect 15708 29374 15710 29426
rect 15762 29374 15764 29426
rect 15708 29362 15764 29374
rect 16044 29428 16100 30268
rect 16492 29764 16548 34076
rect 15820 28420 15876 28430
rect 15596 28418 15876 28420
rect 15596 28366 15822 28418
rect 15874 28366 15876 28418
rect 15596 28364 15876 28366
rect 15820 28354 15876 28364
rect 15484 28030 15486 28082
rect 15538 28030 15540 28082
rect 15484 28018 15540 28030
rect 14028 27972 14084 27982
rect 14252 27972 14308 27982
rect 14084 27970 14308 27972
rect 14084 27918 14254 27970
rect 14306 27918 14308 27970
rect 14084 27916 14308 27918
rect 14028 27906 14084 27916
rect 14252 27906 14308 27916
rect 14364 27970 14420 27982
rect 14364 27918 14366 27970
rect 14418 27918 14420 27970
rect 13916 27860 13972 27870
rect 13916 27766 13972 27804
rect 14028 27188 14084 27198
rect 13804 27132 14028 27188
rect 14028 27094 14084 27132
rect 14364 26964 14420 27918
rect 14588 27972 14644 27982
rect 14588 27878 14644 27916
rect 15708 27972 15764 27982
rect 15708 27878 15764 27916
rect 15820 27860 15876 27870
rect 15820 27766 15876 27804
rect 15260 27748 15316 27758
rect 16044 27748 16100 29372
rect 16380 29708 16548 29764
rect 16604 32788 16660 34190
rect 16828 33460 16884 34636
rect 16940 34354 16996 34748
rect 16940 34302 16942 34354
rect 16994 34302 16996 34354
rect 16940 34290 16996 34302
rect 16940 33460 16996 33470
rect 16828 33458 16996 33460
rect 16828 33406 16942 33458
rect 16994 33406 16996 33458
rect 16828 33404 16996 33406
rect 16716 32788 16772 32798
rect 16604 32786 16772 32788
rect 16604 32734 16718 32786
rect 16770 32734 16772 32786
rect 16604 32732 16772 32734
rect 16604 32002 16660 32732
rect 16716 32722 16772 32732
rect 16828 32004 16884 33404
rect 16940 33394 16996 33404
rect 17052 33124 17108 35308
rect 17500 35252 17556 35262
rect 17612 35252 17668 38444
rect 18284 38276 18340 38894
rect 18284 38210 18340 38220
rect 18396 40348 18564 40404
rect 18396 39058 18452 40348
rect 18956 39842 19012 39854
rect 18956 39790 18958 39842
rect 19010 39790 19012 39842
rect 18396 39006 18398 39058
rect 18450 39006 18452 39058
rect 18396 38052 18452 39006
rect 17724 37996 18452 38052
rect 18620 39618 18676 39630
rect 18620 39566 18622 39618
rect 18674 39566 18676 39618
rect 18620 38612 18676 39566
rect 17724 37266 17780 37996
rect 17948 37828 18004 37838
rect 17948 37734 18004 37772
rect 17836 37492 17892 37502
rect 17836 37398 17892 37436
rect 17724 37214 17726 37266
rect 17778 37214 17780 37266
rect 17724 37202 17780 37214
rect 18060 37268 18116 37278
rect 18060 37174 18116 37212
rect 18620 37266 18676 38556
rect 18732 38276 18788 38286
rect 18732 38182 18788 38220
rect 18956 37828 19012 39790
rect 19180 39732 19236 39742
rect 19068 39060 19124 39070
rect 19180 39060 19236 39676
rect 19068 39058 19236 39060
rect 19068 39006 19070 39058
rect 19122 39006 19236 39058
rect 19068 39004 19236 39006
rect 19068 38612 19124 39004
rect 19068 38546 19124 38556
rect 19292 37828 19348 37838
rect 18956 37762 19012 37772
rect 19068 37826 19348 37828
rect 19068 37774 19294 37826
rect 19346 37774 19348 37826
rect 19068 37772 19348 37774
rect 18620 37214 18622 37266
rect 18674 37214 18676 37266
rect 18620 35588 18676 37214
rect 18620 35252 18676 35532
rect 17612 35196 18116 35252
rect 17164 35140 17220 35150
rect 17164 35138 17444 35140
rect 17164 35086 17166 35138
rect 17218 35086 17444 35138
rect 17164 35084 17444 35086
rect 17164 35074 17220 35084
rect 17276 34802 17332 34814
rect 17276 34750 17278 34802
rect 17330 34750 17332 34802
rect 17164 34690 17220 34702
rect 17164 34638 17166 34690
rect 17218 34638 17220 34690
rect 17164 33908 17220 34638
rect 17164 33842 17220 33852
rect 17276 33458 17332 34750
rect 17388 33908 17444 35084
rect 17500 34130 17556 35196
rect 17948 35026 18004 35038
rect 17948 34974 17950 35026
rect 18002 34974 18004 35026
rect 17612 34804 17668 34814
rect 17612 34710 17668 34748
rect 17836 34692 17892 34702
rect 17836 34356 17892 34636
rect 17836 34290 17892 34300
rect 17500 34078 17502 34130
rect 17554 34078 17556 34130
rect 17500 34066 17556 34078
rect 17836 34130 17892 34142
rect 17836 34078 17838 34130
rect 17890 34078 17892 34130
rect 17836 33908 17892 34078
rect 17388 33852 17892 33908
rect 17948 33796 18004 34974
rect 17276 33406 17278 33458
rect 17330 33406 17332 33458
rect 17276 33394 17332 33406
rect 17724 33740 18004 33796
rect 18060 34804 18116 35196
rect 18620 35186 18676 35196
rect 18732 37380 18788 37390
rect 18508 34804 18564 34814
rect 18060 34802 18564 34804
rect 18060 34750 18062 34802
rect 18114 34750 18510 34802
rect 18562 34750 18564 34802
rect 18060 34748 18564 34750
rect 17052 33058 17108 33068
rect 17612 33234 17668 33246
rect 17612 33182 17614 33234
rect 17666 33182 17668 33234
rect 17612 33124 17668 33182
rect 17724 33234 17780 33740
rect 18060 33684 18116 34748
rect 18508 34738 18564 34748
rect 18060 33348 18116 33628
rect 17724 33182 17726 33234
rect 17778 33182 17780 33234
rect 17724 33170 17780 33182
rect 17836 33292 18116 33348
rect 18172 34356 18228 34366
rect 17836 33234 17892 33292
rect 17836 33182 17838 33234
rect 17890 33182 17892 33234
rect 17612 33058 17668 33068
rect 17612 32788 17668 32798
rect 17836 32788 17892 33182
rect 18060 33124 18116 33134
rect 18172 33124 18228 34300
rect 18060 33122 18228 33124
rect 18060 33070 18062 33122
rect 18114 33070 18228 33122
rect 18060 33068 18228 33070
rect 18508 33124 18564 33134
rect 18060 33058 18116 33068
rect 18508 33030 18564 33068
rect 18732 32900 18788 37324
rect 19068 37266 19124 37772
rect 19292 37762 19348 37772
rect 19068 37214 19070 37266
rect 19122 37214 19124 37266
rect 19068 37202 19124 37214
rect 18844 36260 18900 36270
rect 18844 36166 18900 36204
rect 19404 35924 19460 41692
rect 19628 39844 19684 39854
rect 19964 39844 20020 41804
rect 20748 41298 20804 42140
rect 20748 41246 20750 41298
rect 20802 41246 20804 41298
rect 20748 41188 20804 41246
rect 20748 41122 20804 41132
rect 20972 41970 21028 42476
rect 20972 41918 20974 41970
rect 21026 41918 21028 41970
rect 19628 39842 20020 39844
rect 19628 39790 19630 39842
rect 19682 39790 20020 39842
rect 19628 39788 20020 39790
rect 19628 39730 19684 39788
rect 19628 39678 19630 39730
rect 19682 39678 19684 39730
rect 19628 39666 19684 39678
rect 20972 39732 21028 41918
rect 20972 39666 21028 39676
rect 19292 35868 19460 35924
rect 19516 39396 19572 39406
rect 19516 38948 19572 39340
rect 19516 38892 20132 38948
rect 19516 38834 19572 38892
rect 19516 38782 19518 38834
rect 19570 38782 19572 38834
rect 19068 34804 19124 34814
rect 19068 34710 19124 34748
rect 18956 33684 19012 33694
rect 18956 33458 19012 33628
rect 18956 33406 18958 33458
rect 19010 33406 19012 33458
rect 18956 33394 19012 33406
rect 19292 33460 19348 35868
rect 19404 35698 19460 35710
rect 19404 35646 19406 35698
rect 19458 35646 19460 35698
rect 19404 35588 19460 35646
rect 19404 35522 19460 35532
rect 19516 34804 19572 38782
rect 19852 38724 19908 38734
rect 19628 38052 19684 38062
rect 19628 37958 19684 37996
rect 19852 37938 19908 38668
rect 20076 38668 20132 38892
rect 21308 38668 21364 44044
rect 21532 43764 21588 44158
rect 21532 43698 21588 43708
rect 21420 43426 21476 43438
rect 21420 43374 21422 43426
rect 21474 43374 21476 43426
rect 21420 43316 21476 43374
rect 21420 43250 21476 43260
rect 21756 43428 21812 43438
rect 21756 42978 21812 43372
rect 21756 42926 21758 42978
rect 21810 42926 21812 42978
rect 21756 42914 21812 42926
rect 22316 42756 22372 44940
rect 22428 42868 22484 48972
rect 22540 47460 22596 47470
rect 22540 47366 22596 47404
rect 22764 46900 22820 50372
rect 22876 49700 22932 49710
rect 22876 49698 23044 49700
rect 22876 49646 22878 49698
rect 22930 49646 23044 49698
rect 22876 49644 23044 49646
rect 22876 49634 22932 49644
rect 22876 49026 22932 49038
rect 22876 48974 22878 49026
rect 22930 48974 22932 49026
rect 22876 48468 22932 48974
rect 22876 48402 22932 48412
rect 22988 47682 23044 49644
rect 23324 49026 23380 51996
rect 23436 51940 23492 51950
rect 23436 51602 23492 51884
rect 23436 51550 23438 51602
rect 23490 51550 23492 51602
rect 23436 51538 23492 51550
rect 23436 50482 23492 50494
rect 23436 50430 23438 50482
rect 23490 50430 23492 50482
rect 23436 50428 23492 50430
rect 23660 50428 23716 52108
rect 23772 52098 23828 52108
rect 23772 51604 23828 51614
rect 23772 51510 23828 51548
rect 23884 50594 23940 52220
rect 24220 52164 24276 52174
rect 24220 51602 24276 52108
rect 24220 51550 24222 51602
rect 24274 51550 24276 51602
rect 24220 51538 24276 51550
rect 24892 51938 24948 51950
rect 24892 51886 24894 51938
rect 24946 51886 24948 51938
rect 24892 51604 24948 51886
rect 24892 51538 24948 51548
rect 25340 51492 25396 52444
rect 25452 52276 25508 52286
rect 25452 52182 25508 52220
rect 25340 51436 25508 51492
rect 25340 51266 25396 51278
rect 25340 51214 25342 51266
rect 25394 51214 25396 51266
rect 25340 51154 25396 51214
rect 25340 51102 25342 51154
rect 25394 51102 25396 51154
rect 24008 50988 25208 50998
rect 24064 50986 24112 50988
rect 24168 50986 24216 50988
rect 24076 50934 24112 50986
rect 24200 50934 24216 50986
rect 24064 50932 24112 50934
rect 24168 50932 24216 50934
rect 24272 50986 24320 50988
rect 24376 50986 24424 50988
rect 24480 50986 24528 50988
rect 24376 50934 24396 50986
rect 24480 50934 24520 50986
rect 24272 50932 24320 50934
rect 24376 50932 24424 50934
rect 24480 50932 24528 50934
rect 24584 50932 24632 50988
rect 24688 50986 24736 50988
rect 24792 50986 24840 50988
rect 24896 50986 24944 50988
rect 24696 50934 24736 50986
rect 24820 50934 24840 50986
rect 24688 50932 24736 50934
rect 24792 50932 24840 50934
rect 24896 50932 24944 50934
rect 25000 50986 25048 50988
rect 25104 50986 25152 50988
rect 25000 50934 25016 50986
rect 25104 50934 25140 50986
rect 25000 50932 25048 50934
rect 25104 50932 25152 50934
rect 24008 50922 25208 50932
rect 24332 50708 24388 50718
rect 24332 50614 24388 50652
rect 24892 50708 24948 50718
rect 24892 50614 24948 50652
rect 23884 50542 23886 50594
rect 23938 50542 23940 50594
rect 23884 50530 23940 50542
rect 23996 50484 24052 50494
rect 23436 50372 23604 50428
rect 23660 50372 23940 50428
rect 23548 50148 23604 50372
rect 23548 50092 23828 50148
rect 23548 49810 23604 49822
rect 23548 49758 23550 49810
rect 23602 49758 23604 49810
rect 23324 48974 23326 49026
rect 23378 48974 23380 49026
rect 23324 48692 23380 48974
rect 23436 49698 23492 49710
rect 23436 49646 23438 49698
rect 23490 49646 23492 49698
rect 23436 48916 23492 49646
rect 23548 49138 23604 49758
rect 23772 49810 23828 50092
rect 23772 49758 23774 49810
rect 23826 49758 23828 49810
rect 23772 49746 23828 49758
rect 23884 49588 23940 50372
rect 23996 50034 24052 50428
rect 23996 49982 23998 50034
rect 24050 49982 24052 50034
rect 23996 49970 24052 49982
rect 23548 49086 23550 49138
rect 23602 49086 23604 49138
rect 23548 49074 23604 49086
rect 23772 49532 23940 49588
rect 23436 48860 23604 48916
rect 23380 48636 23492 48692
rect 23324 48598 23380 48636
rect 22988 47630 22990 47682
rect 23042 47630 23044 47682
rect 22988 47618 23044 47630
rect 23212 47460 23268 47470
rect 22988 47458 23268 47460
rect 22988 47406 23214 47458
rect 23266 47406 23268 47458
rect 22988 47404 23268 47406
rect 22764 46834 22820 46844
rect 22876 47346 22932 47358
rect 22876 47294 22878 47346
rect 22930 47294 22932 47346
rect 22876 46788 22932 47294
rect 22876 46722 22932 46732
rect 22988 46564 23044 47404
rect 23212 47394 23268 47404
rect 23324 47458 23380 47470
rect 23324 47406 23326 47458
rect 23378 47406 23380 47458
rect 22764 46508 23044 46564
rect 22764 46002 22820 46508
rect 22764 45950 22766 46002
rect 22818 45950 22820 46002
rect 22764 45938 22820 45950
rect 22988 45330 23044 45342
rect 22988 45278 22990 45330
rect 23042 45278 23044 45330
rect 22988 44100 23044 45278
rect 22988 44034 23044 44044
rect 23324 43092 23380 47406
rect 23436 45890 23492 48636
rect 23548 46228 23604 48860
rect 23660 48356 23716 48366
rect 23660 48262 23716 48300
rect 23772 48244 23828 49532
rect 24008 49420 25208 49430
rect 24064 49418 24112 49420
rect 24168 49418 24216 49420
rect 24076 49366 24112 49418
rect 24200 49366 24216 49418
rect 24064 49364 24112 49366
rect 24168 49364 24216 49366
rect 24272 49418 24320 49420
rect 24376 49418 24424 49420
rect 24480 49418 24528 49420
rect 24376 49366 24396 49418
rect 24480 49366 24520 49418
rect 24272 49364 24320 49366
rect 24376 49364 24424 49366
rect 24480 49364 24528 49366
rect 24584 49364 24632 49420
rect 24688 49418 24736 49420
rect 24792 49418 24840 49420
rect 24896 49418 24944 49420
rect 24696 49366 24736 49418
rect 24820 49366 24840 49418
rect 24688 49364 24736 49366
rect 24792 49364 24840 49366
rect 24896 49364 24944 49366
rect 25000 49418 25048 49420
rect 25104 49418 25152 49420
rect 25000 49366 25016 49418
rect 25104 49366 25140 49418
rect 25000 49364 25048 49366
rect 25104 49364 25152 49366
rect 24008 49354 25208 49364
rect 24332 49028 24388 49038
rect 24332 48934 24388 48972
rect 25340 48916 25396 51102
rect 25452 50428 25508 51436
rect 25564 50708 25620 53564
rect 25676 53526 25732 53564
rect 25788 52836 25844 55918
rect 26460 54740 26516 56028
rect 26348 54738 26516 54740
rect 26348 54686 26462 54738
rect 26514 54686 26516 54738
rect 26348 54684 26516 54686
rect 25676 52834 25844 52836
rect 25676 52782 25790 52834
rect 25842 52782 25844 52834
rect 25676 52780 25844 52782
rect 25676 52164 25732 52780
rect 25788 52770 25844 52780
rect 25900 53730 25956 53742
rect 25900 53678 25902 53730
rect 25954 53678 25956 53730
rect 25900 53508 25956 53678
rect 25676 52098 25732 52108
rect 25900 52162 25956 53452
rect 26348 53172 26404 54684
rect 26460 54674 26516 54684
rect 27020 54402 27076 54414
rect 27020 54350 27022 54402
rect 27074 54350 27076 54402
rect 26460 53956 26516 53966
rect 26460 53862 26516 53900
rect 26796 53956 26852 53966
rect 26572 53844 26628 53854
rect 25900 52110 25902 52162
rect 25954 52110 25956 52162
rect 25788 52052 25844 52062
rect 25788 51958 25844 51996
rect 25788 51604 25844 51614
rect 25788 51510 25844 51548
rect 25900 51154 25956 52110
rect 25900 51102 25902 51154
rect 25954 51102 25956 51154
rect 25900 51090 25956 51102
rect 26236 53170 26404 53172
rect 26236 53118 26350 53170
rect 26402 53118 26404 53170
rect 26236 53116 26404 53118
rect 26236 51604 26292 53116
rect 26348 53106 26404 53116
rect 26460 53172 26516 53182
rect 26460 52388 26516 53116
rect 26572 52946 26628 53788
rect 26796 53730 26852 53900
rect 26796 53678 26798 53730
rect 26850 53678 26852 53730
rect 26796 53666 26852 53678
rect 26572 52894 26574 52946
rect 26626 52894 26628 52946
rect 26572 52882 26628 52894
rect 26572 52388 26628 52398
rect 26460 52386 26628 52388
rect 26460 52334 26574 52386
rect 26626 52334 26628 52386
rect 26460 52332 26628 52334
rect 26572 52322 26628 52332
rect 25564 50642 25620 50652
rect 25452 50372 25620 50428
rect 25340 48850 25396 48860
rect 25452 49252 25508 49262
rect 23772 47572 23828 48188
rect 23772 47506 23828 47516
rect 23884 48468 23940 48478
rect 23660 47460 23716 47470
rect 23660 47366 23716 47404
rect 23884 47346 23940 48412
rect 24444 48468 24500 48478
rect 24444 48374 24500 48412
rect 25340 48468 25396 48478
rect 25452 48468 25508 49196
rect 25340 48466 25508 48468
rect 25340 48414 25342 48466
rect 25394 48414 25508 48466
rect 25340 48412 25508 48414
rect 25340 48356 25396 48412
rect 25340 48290 25396 48300
rect 24008 47852 25208 47862
rect 24064 47850 24112 47852
rect 24168 47850 24216 47852
rect 24076 47798 24112 47850
rect 24200 47798 24216 47850
rect 24064 47796 24112 47798
rect 24168 47796 24216 47798
rect 24272 47850 24320 47852
rect 24376 47850 24424 47852
rect 24480 47850 24528 47852
rect 24376 47798 24396 47850
rect 24480 47798 24520 47850
rect 24272 47796 24320 47798
rect 24376 47796 24424 47798
rect 24480 47796 24528 47798
rect 24584 47796 24632 47852
rect 24688 47850 24736 47852
rect 24792 47850 24840 47852
rect 24896 47850 24944 47852
rect 24696 47798 24736 47850
rect 24820 47798 24840 47850
rect 24688 47796 24736 47798
rect 24792 47796 24840 47798
rect 24896 47796 24944 47798
rect 25000 47850 25048 47852
rect 25104 47850 25152 47852
rect 25000 47798 25016 47850
rect 25104 47798 25140 47850
rect 25000 47796 25048 47798
rect 25104 47796 25152 47798
rect 24008 47786 25208 47796
rect 24444 47572 24500 47582
rect 24444 47458 24500 47516
rect 24444 47406 24446 47458
rect 24498 47406 24500 47458
rect 24444 47394 24500 47406
rect 24780 47458 24836 47470
rect 24780 47406 24782 47458
rect 24834 47406 24836 47458
rect 23884 47294 23886 47346
rect 23938 47294 23940 47346
rect 23884 47282 23940 47294
rect 23996 47346 24052 47358
rect 23996 47294 23998 47346
rect 24050 47294 24052 47346
rect 23996 47236 24052 47294
rect 23996 47170 24052 47180
rect 23772 46900 23828 46910
rect 23772 46562 23828 46844
rect 23772 46510 23774 46562
rect 23826 46510 23828 46562
rect 23548 46172 23716 46228
rect 23436 45838 23438 45890
rect 23490 45838 23492 45890
rect 23436 45220 23492 45838
rect 23548 46002 23604 46014
rect 23548 45950 23550 46002
rect 23602 45950 23604 46002
rect 23548 45332 23604 45950
rect 23548 45238 23604 45276
rect 23436 45154 23492 45164
rect 23660 44324 23716 46172
rect 22764 43036 23380 43092
rect 23548 44268 23716 44324
rect 22540 42868 22596 42878
rect 22428 42812 22540 42868
rect 22540 42802 22596 42812
rect 22204 42700 22316 42756
rect 21420 42530 21476 42542
rect 21420 42478 21422 42530
rect 21474 42478 21476 42530
rect 21420 41970 21476 42478
rect 21420 41918 21422 41970
rect 21474 41918 21476 41970
rect 21420 41906 21476 41918
rect 21532 41300 21588 41310
rect 21532 41206 21588 41244
rect 21868 41188 21924 41198
rect 21532 40404 21588 40414
rect 20076 38612 20244 38668
rect 21308 38612 21476 38668
rect 19852 37886 19854 37938
rect 19906 37886 19908 37938
rect 19852 37874 19908 37886
rect 20188 37938 20244 38612
rect 20188 37886 20190 37938
rect 20242 37886 20244 37938
rect 20188 37874 20244 37886
rect 21084 37380 21140 37390
rect 19628 37268 19684 37278
rect 19628 34914 19684 37212
rect 20188 36260 20244 36270
rect 19852 35698 19908 35710
rect 19852 35646 19854 35698
rect 19906 35646 19908 35698
rect 19852 35140 19908 35646
rect 20188 35308 20244 36204
rect 19852 35074 19908 35084
rect 20076 35252 20244 35308
rect 20300 35924 20356 35934
rect 19628 34862 19630 34914
rect 19682 34862 19684 34914
rect 19628 34850 19684 34862
rect 19516 34710 19572 34748
rect 19292 33394 19348 33404
rect 20076 34130 20132 35252
rect 20300 35138 20356 35868
rect 20300 35086 20302 35138
rect 20354 35086 20356 35138
rect 20300 35074 20356 35086
rect 20636 35140 20692 35150
rect 20636 35046 20692 35084
rect 20076 34078 20078 34130
rect 20130 34078 20132 34130
rect 20076 34020 20132 34078
rect 18732 32844 18900 32900
rect 18060 32788 18116 32798
rect 16604 31950 16606 32002
rect 16658 31950 16660 32002
rect 16604 31780 16660 31950
rect 16604 30210 16660 31724
rect 16716 31948 16884 32004
rect 17276 32786 18452 32788
rect 17276 32734 17614 32786
rect 17666 32734 18062 32786
rect 18114 32734 18452 32786
rect 17276 32732 18452 32734
rect 16716 31890 16772 31948
rect 16716 31838 16718 31890
rect 16770 31838 16772 31890
rect 16716 31220 16772 31838
rect 17052 31780 17108 31790
rect 17052 31686 17108 31724
rect 17276 31778 17332 32732
rect 17612 32722 17668 32732
rect 18060 32722 18116 32732
rect 17276 31726 17278 31778
rect 17330 31726 17332 31778
rect 17276 31668 17332 31726
rect 18172 31780 18228 31790
rect 18172 31686 18228 31724
rect 18396 31778 18452 32732
rect 18396 31726 18398 31778
rect 18450 31726 18452 31778
rect 18396 31714 18452 31726
rect 17276 31602 17332 31612
rect 17388 31666 17444 31678
rect 17388 31614 17390 31666
rect 17442 31614 17444 31666
rect 17388 31556 17444 31614
rect 18732 31666 18788 31678
rect 18732 31614 18734 31666
rect 18786 31614 18788 31666
rect 16828 31220 16884 31230
rect 17388 31220 17444 31500
rect 17836 31554 17892 31566
rect 17836 31502 17838 31554
rect 17890 31502 17892 31554
rect 16716 31218 17444 31220
rect 16716 31166 16830 31218
rect 16882 31166 17444 31218
rect 16716 31164 17444 31166
rect 17500 31220 17556 31230
rect 16828 31154 16884 31164
rect 17500 30994 17556 31164
rect 17500 30942 17502 30994
rect 17554 30942 17556 30994
rect 17500 30930 17556 30942
rect 17724 30882 17780 30894
rect 17724 30830 17726 30882
rect 17778 30830 17780 30882
rect 17388 30772 17444 30782
rect 17388 30678 17444 30716
rect 16604 30158 16606 30210
rect 16658 30158 16660 30210
rect 16380 28532 16436 29708
rect 16492 29540 16548 29550
rect 16604 29540 16660 30158
rect 17164 30212 17220 30222
rect 17724 30212 17780 30830
rect 17836 30772 17892 31502
rect 18508 31554 18564 31566
rect 18508 31502 18510 31554
rect 18562 31502 18564 31554
rect 18508 31220 18564 31502
rect 18732 31556 18788 31614
rect 18732 31490 18788 31500
rect 17948 31164 18564 31220
rect 17948 30994 18004 31164
rect 17948 30942 17950 30994
rect 18002 30942 18004 30994
rect 17948 30930 18004 30942
rect 18172 30772 18228 30782
rect 17836 30770 18228 30772
rect 17836 30718 18174 30770
rect 18226 30718 18228 30770
rect 17836 30716 18228 30718
rect 17836 30212 17892 30222
rect 17724 30156 17836 30212
rect 16492 29538 16996 29540
rect 16492 29486 16494 29538
rect 16546 29486 16996 29538
rect 16492 29484 16996 29486
rect 16492 29474 16548 29484
rect 16380 28466 16436 28476
rect 16828 28532 16884 28542
rect 16828 28082 16884 28476
rect 16828 28030 16830 28082
rect 16882 28030 16884 28082
rect 16828 28018 16884 28030
rect 16380 27748 16436 27758
rect 16044 27746 16436 27748
rect 16044 27694 16382 27746
rect 16434 27694 16436 27746
rect 16044 27692 16436 27694
rect 15260 27654 15316 27692
rect 15148 27188 15204 27198
rect 15148 27094 15204 27132
rect 15484 27076 15540 27086
rect 14364 26898 14420 26908
rect 14700 26964 14756 27002
rect 14700 26898 14756 26908
rect 14008 26684 15208 26694
rect 14064 26682 14112 26684
rect 14168 26682 14216 26684
rect 14076 26630 14112 26682
rect 14200 26630 14216 26682
rect 14064 26628 14112 26630
rect 14168 26628 14216 26630
rect 14272 26682 14320 26684
rect 14376 26682 14424 26684
rect 14480 26682 14528 26684
rect 14376 26630 14396 26682
rect 14480 26630 14520 26682
rect 14272 26628 14320 26630
rect 14376 26628 14424 26630
rect 14480 26628 14528 26630
rect 14584 26628 14632 26684
rect 14688 26682 14736 26684
rect 14792 26682 14840 26684
rect 14896 26682 14944 26684
rect 14696 26630 14736 26682
rect 14820 26630 14840 26682
rect 14688 26628 14736 26630
rect 14792 26628 14840 26630
rect 14896 26628 14944 26630
rect 15000 26682 15048 26684
rect 15104 26682 15152 26684
rect 15000 26630 15016 26682
rect 15104 26630 15140 26682
rect 15000 26628 15048 26630
rect 15104 26628 15152 26630
rect 14008 26618 15208 26628
rect 14028 25620 14084 25630
rect 14028 25526 14084 25564
rect 14476 25620 14532 25630
rect 14364 25394 14420 25406
rect 14364 25342 14366 25394
rect 14418 25342 14420 25394
rect 13580 25284 13636 25294
rect 14364 25284 14420 25342
rect 14476 25394 14532 25564
rect 14700 25508 14756 25518
rect 14700 25506 15204 25508
rect 14700 25454 14702 25506
rect 14754 25454 15204 25506
rect 14700 25452 15204 25454
rect 14700 25442 14756 25452
rect 14476 25342 14478 25394
rect 14530 25342 14532 25394
rect 14476 25330 14532 25342
rect 13636 25228 14420 25284
rect 15036 25284 15092 25322
rect 15148 25284 15204 25452
rect 15484 25284 15540 27020
rect 16380 26964 16436 27692
rect 16940 27186 16996 29484
rect 16940 27134 16942 27186
rect 16994 27134 16996 27186
rect 16940 27122 16996 27134
rect 16380 26898 16436 26908
rect 15148 25228 15428 25284
rect 13580 25190 13636 25228
rect 15036 25218 15092 25228
rect 12572 24894 12574 24946
rect 12626 24894 12628 24946
rect 12572 24836 12628 24894
rect 13020 25116 13524 25172
rect 13020 24946 13076 25116
rect 13468 25060 13524 25116
rect 14008 25116 15208 25126
rect 14064 25114 14112 25116
rect 14168 25114 14216 25116
rect 14076 25062 14112 25114
rect 14200 25062 14216 25114
rect 14064 25060 14112 25062
rect 14168 25060 14216 25062
rect 14272 25114 14320 25116
rect 14376 25114 14424 25116
rect 14480 25114 14528 25116
rect 14376 25062 14396 25114
rect 14480 25062 14520 25114
rect 14272 25060 14320 25062
rect 14376 25060 14424 25062
rect 14480 25060 14528 25062
rect 14584 25060 14632 25116
rect 14688 25114 14736 25116
rect 14792 25114 14840 25116
rect 14896 25114 14944 25116
rect 14696 25062 14736 25114
rect 14820 25062 14840 25114
rect 14688 25060 14736 25062
rect 14792 25060 14840 25062
rect 14896 25060 14944 25062
rect 15000 25114 15048 25116
rect 15104 25114 15152 25116
rect 15000 25062 15016 25114
rect 15104 25062 15140 25114
rect 15000 25060 15048 25062
rect 15104 25060 15152 25062
rect 13468 25004 13860 25060
rect 14008 25050 15208 25060
rect 13020 24894 13022 24946
rect 13074 24894 13076 24946
rect 13020 24882 13076 24894
rect 12572 24770 12628 24780
rect 13804 24722 13860 25004
rect 14028 24836 14084 24846
rect 14028 24742 14084 24780
rect 14364 24834 14420 24846
rect 14364 24782 14366 24834
rect 14418 24782 14420 24834
rect 13804 24670 13806 24722
rect 13858 24670 13860 24722
rect 13804 24658 13860 24670
rect 13468 24500 13524 24510
rect 13468 24498 13860 24500
rect 13468 24446 13470 24498
rect 13522 24446 13860 24498
rect 13468 24444 13860 24446
rect 13468 24434 13524 24444
rect 10780 23662 10782 23714
rect 10834 23662 10836 23714
rect 10780 23650 10836 23662
rect 11228 23716 11284 23726
rect 11116 23156 11172 23166
rect 11116 23062 11172 23100
rect 10556 22530 10612 22540
rect 11228 22370 11284 23660
rect 11900 23716 11956 23726
rect 11900 23622 11956 23660
rect 12236 23714 12292 23772
rect 12236 23662 12238 23714
rect 12290 23662 12292 23714
rect 12236 23604 12292 23662
rect 13468 23938 13524 23950
rect 13468 23886 13470 23938
rect 13522 23886 13524 23938
rect 12236 23548 12628 23604
rect 11564 23154 11620 23166
rect 11564 23102 11566 23154
rect 11618 23102 11620 23154
rect 11564 22482 11620 23102
rect 11564 22430 11566 22482
rect 11618 22430 11620 22482
rect 11564 22418 11620 22430
rect 12460 23044 12516 23054
rect 11228 22318 11230 22370
rect 11282 22318 11284 22370
rect 11228 22306 11284 22318
rect 11788 22372 11844 22382
rect 11564 22260 11620 22270
rect 11564 22166 11620 22204
rect 10332 20802 10388 21308
rect 11676 22146 11732 22158
rect 11676 22094 11678 22146
rect 11730 22094 11732 22146
rect 11676 21140 11732 22094
rect 10332 20750 10334 20802
rect 10386 20750 10388 20802
rect 10332 20692 10388 20750
rect 10332 20626 10388 20636
rect 10444 21084 11732 21140
rect 10332 20132 10388 20170
rect 10332 20066 10388 20076
rect 10444 20130 10500 21084
rect 10444 20078 10446 20130
rect 10498 20078 10500 20130
rect 10332 19908 10388 19918
rect 10108 19906 10388 19908
rect 10108 19854 10334 19906
rect 10386 19854 10388 19906
rect 10108 19852 10388 19854
rect 10332 19842 10388 19852
rect 10444 17890 10500 20078
rect 10556 20914 10612 20926
rect 10556 20862 10558 20914
rect 10610 20862 10612 20914
rect 10556 20132 10612 20862
rect 11788 20804 11844 22316
rect 12460 22372 12516 22988
rect 12460 22278 12516 22316
rect 12124 22260 12180 22270
rect 12124 22166 12180 22204
rect 11900 22148 11956 22158
rect 12236 22148 12292 22158
rect 11900 22146 12068 22148
rect 11900 22094 11902 22146
rect 11954 22094 12068 22146
rect 11900 22092 12068 22094
rect 11900 22082 11956 22092
rect 12012 21364 12068 22092
rect 12236 22054 12292 22092
rect 12348 21698 12404 21710
rect 12348 21646 12350 21698
rect 12402 21646 12404 21698
rect 12012 21308 12292 21364
rect 12236 20914 12292 21308
rect 12236 20862 12238 20914
rect 12290 20862 12292 20914
rect 12236 20850 12292 20862
rect 11788 20802 12068 20804
rect 11788 20750 11790 20802
rect 11842 20750 12068 20802
rect 11788 20748 12068 20750
rect 11788 20738 11844 20748
rect 10892 20692 10948 20702
rect 10780 20690 10948 20692
rect 10780 20638 10894 20690
rect 10946 20638 10948 20690
rect 10780 20636 10948 20638
rect 10668 20244 10724 20254
rect 10780 20244 10836 20636
rect 10892 20626 10948 20636
rect 10668 20242 10836 20244
rect 10668 20190 10670 20242
rect 10722 20190 10836 20242
rect 10668 20188 10836 20190
rect 11564 20242 11620 20254
rect 11564 20190 11566 20242
rect 11618 20190 11620 20242
rect 10668 20178 10724 20188
rect 10556 20066 10612 20076
rect 11564 20132 11620 20190
rect 11676 20242 11732 20254
rect 11676 20190 11678 20242
rect 11730 20190 11732 20242
rect 11676 20132 11732 20190
rect 11788 20132 11844 20142
rect 11676 20076 11788 20132
rect 12012 20132 12068 20748
rect 12124 20802 12180 20814
rect 12124 20750 12126 20802
rect 12178 20750 12180 20802
rect 12124 20468 12180 20750
rect 12348 20580 12404 21646
rect 12572 21476 12628 23548
rect 13356 23268 13412 23278
rect 12796 22372 12852 22382
rect 12796 22370 12964 22372
rect 12796 22318 12798 22370
rect 12850 22318 12964 22370
rect 12796 22316 12964 22318
rect 12796 22306 12852 22316
rect 12572 21410 12628 21420
rect 12908 20914 12964 22316
rect 12908 20862 12910 20914
rect 12962 20862 12964 20914
rect 12908 20804 12964 20862
rect 12908 20738 12964 20748
rect 13132 21364 13188 21374
rect 12348 20514 12404 20524
rect 12124 20412 12292 20468
rect 12124 20132 12180 20142
rect 12012 20130 12180 20132
rect 12012 20078 12126 20130
rect 12178 20078 12180 20130
rect 12012 20076 12180 20078
rect 12236 20132 12292 20412
rect 13132 20244 13188 21308
rect 13020 20188 13132 20244
rect 12348 20132 12404 20142
rect 12236 20130 12404 20132
rect 12236 20078 12350 20130
rect 12402 20078 12404 20130
rect 12236 20076 12404 20078
rect 11564 20066 11620 20076
rect 10444 17838 10446 17890
rect 10498 17838 10500 17890
rect 10444 17826 10500 17838
rect 9996 17574 10052 17612
rect 10892 17668 10948 17678
rect 10556 17442 10612 17454
rect 10556 17390 10558 17442
rect 10610 17390 10612 17442
rect 10556 17220 10612 17390
rect 10780 17444 10836 17454
rect 10780 17350 10836 17388
rect 10108 17164 10612 17220
rect 10108 17106 10164 17164
rect 10108 17054 10110 17106
rect 10162 17054 10164 17106
rect 10108 17042 10164 17054
rect 10444 16996 10500 17006
rect 10444 16902 10500 16940
rect 9772 15486 9774 15538
rect 9826 15486 9828 15538
rect 9548 15428 9604 15438
rect 9548 15148 9604 15372
rect 9772 15148 9828 15486
rect 10556 15538 10612 17164
rect 10892 16994 10948 17612
rect 11116 17666 11172 17678
rect 11116 17614 11118 17666
rect 11170 17614 11172 17666
rect 11116 17444 11172 17614
rect 11116 17378 11172 17388
rect 11452 17442 11508 17454
rect 11452 17390 11454 17442
rect 11506 17390 11508 17442
rect 11228 17332 11284 17342
rect 10892 16942 10894 16994
rect 10946 16942 10948 16994
rect 10892 16930 10948 16942
rect 11004 16996 11060 17006
rect 11004 16902 11060 16940
rect 11116 16996 11172 17006
rect 11228 16996 11284 17276
rect 11116 16994 11284 16996
rect 11116 16942 11118 16994
rect 11170 16942 11284 16994
rect 11116 16940 11284 16942
rect 11116 16930 11172 16940
rect 11228 16772 11284 16782
rect 11228 16212 11284 16716
rect 11228 16118 11284 16156
rect 10556 15486 10558 15538
rect 10610 15486 10612 15538
rect 10220 15314 10276 15326
rect 10220 15262 10222 15314
rect 10274 15262 10276 15314
rect 10220 15148 10276 15262
rect 10556 15148 10612 15486
rect 9548 15092 9716 15148
rect 9772 15092 10052 15148
rect 9660 14532 9716 15092
rect 9772 14532 9828 14542
rect 9660 14530 9828 14532
rect 9660 14478 9774 14530
rect 9826 14478 9828 14530
rect 9660 14476 9828 14478
rect 9772 14466 9828 14476
rect 9996 14532 10052 15092
rect 9548 14420 9604 14430
rect 9548 13860 9604 14364
rect 9996 14418 10052 14476
rect 9996 14366 9998 14418
rect 10050 14366 10052 14418
rect 9996 14354 10052 14366
rect 10108 15092 10612 15148
rect 11004 15202 11060 15214
rect 11004 15150 11006 15202
rect 11058 15150 11060 15202
rect 11004 15148 11060 15150
rect 11004 15092 11172 15148
rect 10108 14418 10164 15092
rect 10556 14980 10612 15092
rect 10556 14914 10612 14924
rect 10556 14532 10612 14542
rect 10108 14366 10110 14418
rect 10162 14366 10164 14418
rect 10108 14354 10164 14366
rect 10332 14418 10388 14430
rect 10332 14366 10334 14418
rect 10386 14366 10388 14418
rect 9884 14308 9940 14318
rect 9548 13766 9604 13804
rect 9772 14306 9940 14308
rect 9772 14254 9886 14306
rect 9938 14254 9940 14306
rect 9772 14252 9940 14254
rect 9548 13636 9604 13646
rect 9548 13074 9604 13580
rect 9660 13634 9716 13646
rect 9660 13582 9662 13634
rect 9714 13582 9716 13634
rect 9660 13186 9716 13582
rect 9660 13134 9662 13186
rect 9714 13134 9716 13186
rect 9660 13122 9716 13134
rect 9548 13022 9550 13074
rect 9602 13022 9604 13074
rect 9548 13010 9604 13022
rect 9772 12852 9828 14252
rect 9884 14242 9940 14252
rect 9884 13972 9940 13982
rect 9884 13858 9940 13916
rect 9884 13806 9886 13858
rect 9938 13806 9940 13858
rect 9884 13794 9940 13806
rect 10108 13746 10164 13758
rect 10108 13694 10110 13746
rect 10162 13694 10164 13746
rect 10108 13524 10164 13694
rect 10164 13468 10276 13524
rect 10108 13458 10164 13468
rect 10220 12852 10276 13468
rect 10332 13076 10388 14366
rect 10556 13970 10612 14476
rect 11116 14532 11172 15092
rect 11452 14980 11508 17390
rect 11564 17444 11620 17454
rect 11564 15428 11620 17388
rect 11788 17444 11844 20076
rect 11900 20020 11956 20030
rect 11900 20018 12068 20020
rect 11900 19966 11902 20018
rect 11954 19966 12068 20018
rect 11900 19964 12068 19966
rect 11900 19954 11956 19964
rect 12012 18562 12068 19964
rect 12012 18510 12014 18562
rect 12066 18510 12068 18562
rect 11900 18226 11956 18238
rect 11900 18174 11902 18226
rect 11954 18174 11956 18226
rect 11900 17668 11956 18174
rect 12012 18004 12068 18510
rect 12124 18564 12180 20076
rect 12348 20066 12404 20076
rect 12572 20132 12628 20142
rect 12572 20038 12628 20076
rect 12684 20018 12740 20030
rect 12684 19966 12686 20018
rect 12738 19966 12740 20018
rect 12236 18564 12292 18574
rect 12124 18508 12236 18564
rect 12236 18470 12292 18508
rect 12012 17938 12068 17948
rect 12572 18340 12628 18350
rect 11900 17574 11956 17612
rect 12012 17554 12068 17566
rect 12012 17502 12014 17554
rect 12066 17502 12068 17554
rect 12012 17444 12068 17502
rect 12572 17554 12628 18284
rect 12572 17502 12574 17554
rect 12626 17502 12628 17554
rect 11788 17388 12068 17444
rect 12348 17444 12404 17454
rect 11788 16996 11844 17388
rect 12348 17350 12404 17388
rect 12572 17332 12628 17502
rect 12572 17266 12628 17276
rect 12684 18004 12740 19966
rect 13020 18340 13076 20188
rect 13132 20178 13188 20188
rect 13020 18274 13076 18284
rect 13132 18562 13188 18574
rect 13132 18510 13134 18562
rect 13186 18510 13188 18562
rect 13132 18004 13188 18510
rect 12740 17948 13188 18004
rect 13244 18450 13300 18462
rect 13244 18398 13246 18450
rect 13298 18398 13300 18450
rect 11788 16930 11844 16940
rect 12348 16996 12404 17006
rect 12124 16882 12180 16894
rect 12124 16830 12126 16882
rect 12178 16830 12180 16882
rect 12124 16772 12180 16830
rect 12124 16706 12180 16716
rect 12348 16100 12404 16940
rect 12684 16660 12740 17948
rect 12908 17444 12964 17454
rect 12964 17388 13076 17444
rect 12908 17378 12964 17388
rect 12348 16098 12516 16100
rect 12348 16046 12350 16098
rect 12402 16046 12516 16098
rect 12348 16044 12516 16046
rect 12348 16034 12404 16044
rect 11564 15314 11620 15372
rect 11564 15262 11566 15314
rect 11618 15262 11620 15314
rect 11564 15250 11620 15262
rect 12236 15876 12292 15886
rect 12236 15314 12292 15820
rect 12236 15262 12238 15314
rect 12290 15262 12292 15314
rect 12236 15250 12292 15262
rect 12012 15202 12068 15214
rect 12012 15150 12014 15202
rect 12066 15150 12068 15202
rect 11788 15092 11844 15102
rect 11788 15090 11956 15092
rect 11788 15038 11790 15090
rect 11842 15038 11956 15090
rect 11788 15036 11956 15038
rect 11788 15026 11844 15036
rect 11452 14914 11508 14924
rect 11452 14644 11508 14654
rect 11116 14438 11172 14476
rect 11228 14588 11452 14644
rect 10556 13918 10558 13970
rect 10610 13918 10612 13970
rect 10556 13906 10612 13918
rect 11116 13970 11172 13982
rect 11116 13918 11118 13970
rect 11170 13918 11172 13970
rect 10780 13860 10836 13870
rect 10780 13746 10836 13804
rect 10780 13694 10782 13746
rect 10834 13694 10836 13746
rect 10780 13682 10836 13694
rect 10444 13076 10500 13086
rect 10332 13020 10444 13076
rect 10444 13010 10500 13020
rect 10780 12964 10836 12974
rect 10556 12962 10836 12964
rect 10556 12910 10782 12962
rect 10834 12910 10836 12962
rect 10556 12908 10836 12910
rect 11116 12964 11172 13918
rect 11228 13972 11284 14588
rect 11452 14550 11508 14588
rect 11900 14532 11956 15036
rect 11900 14438 11956 14476
rect 11228 13858 11284 13916
rect 12012 13860 12068 15150
rect 12348 15090 12404 15102
rect 12348 15038 12350 15090
rect 12402 15038 12404 15090
rect 12348 14980 12404 15038
rect 11228 13806 11230 13858
rect 11282 13806 11284 13858
rect 11228 13794 11284 13806
rect 11564 13804 12068 13860
rect 12124 14924 12348 14980
rect 11452 13746 11508 13758
rect 11452 13694 11454 13746
rect 11506 13694 11508 13746
rect 11452 13636 11508 13694
rect 11452 13570 11508 13580
rect 11228 12964 11284 12974
rect 11116 12962 11284 12964
rect 11116 12910 11230 12962
rect 11282 12910 11284 12962
rect 11116 12908 11284 12910
rect 10332 12852 10388 12862
rect 10220 12850 10388 12852
rect 10220 12798 10334 12850
rect 10386 12798 10388 12850
rect 10220 12796 10388 12798
rect 9772 12786 9828 12796
rect 10332 12404 10388 12796
rect 10332 12310 10388 12348
rect 10556 12402 10612 12908
rect 10780 12898 10836 12908
rect 11228 12898 11284 12908
rect 11452 12964 11508 12974
rect 11564 12964 11620 13804
rect 12012 13636 12068 13646
rect 12124 13636 12180 14924
rect 12348 14914 12404 14924
rect 12348 14532 12404 14542
rect 12348 14438 12404 14476
rect 12348 13972 12404 13982
rect 12348 13878 12404 13916
rect 12460 13748 12516 16044
rect 12684 16098 12740 16604
rect 12684 16046 12686 16098
rect 12738 16046 12740 16098
rect 12684 16034 12740 16046
rect 12908 15988 12964 15998
rect 12796 15986 12964 15988
rect 12796 15934 12910 15986
rect 12962 15934 12964 15986
rect 12796 15932 12964 15934
rect 12796 15314 12852 15932
rect 12908 15922 12964 15932
rect 12908 15540 12964 15550
rect 13020 15540 13076 17388
rect 13244 17332 13300 18398
rect 13132 17276 13300 17332
rect 13132 15876 13188 17276
rect 13356 17220 13412 23212
rect 13244 17164 13412 17220
rect 13468 23156 13524 23886
rect 13468 20468 13524 23100
rect 13580 23716 13636 23726
rect 13580 22594 13636 23660
rect 13804 23604 13860 24444
rect 13916 23938 13972 23950
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13916 23716 13972 23886
rect 14364 23828 14420 24782
rect 15372 24834 15428 25228
rect 15372 24782 15374 24834
rect 15426 24782 15428 24834
rect 15372 24770 15428 24782
rect 15484 24722 15540 25228
rect 15484 24670 15486 24722
rect 15538 24670 15540 24722
rect 15484 24658 15540 24670
rect 16604 24610 16660 24622
rect 16604 24558 16606 24610
rect 16658 24558 16660 24610
rect 14364 23762 14420 23772
rect 15372 24500 15428 24510
rect 13916 23650 13972 23660
rect 13692 23548 13860 23604
rect 15372 23604 15428 24444
rect 16492 24388 16548 24398
rect 16492 23716 16548 24332
rect 16492 23622 16548 23660
rect 16604 23828 16660 24558
rect 15484 23604 15540 23614
rect 14008 23548 15208 23558
rect 13692 23492 13748 23548
rect 14064 23546 14112 23548
rect 14168 23546 14216 23548
rect 14076 23494 14112 23546
rect 14200 23494 14216 23546
rect 14064 23492 14112 23494
rect 14168 23492 14216 23494
rect 14272 23546 14320 23548
rect 14376 23546 14424 23548
rect 14480 23546 14528 23548
rect 14376 23494 14396 23546
rect 14480 23494 14520 23546
rect 14272 23492 14320 23494
rect 14376 23492 14424 23494
rect 14480 23492 14528 23494
rect 14584 23492 14632 23548
rect 14688 23546 14736 23548
rect 14792 23546 14840 23548
rect 14896 23546 14944 23548
rect 14696 23494 14736 23546
rect 14820 23494 14840 23546
rect 14688 23492 14736 23494
rect 14792 23492 14840 23494
rect 14896 23492 14944 23494
rect 15000 23546 15048 23548
rect 15104 23546 15152 23548
rect 15000 23494 15016 23546
rect 15104 23494 15140 23546
rect 15000 23492 15048 23494
rect 15104 23492 15152 23494
rect 14008 23482 15208 23492
rect 15372 23548 15484 23604
rect 13692 23426 13748 23436
rect 15148 23380 15204 23390
rect 15372 23380 15428 23548
rect 15484 23538 15540 23548
rect 16268 23604 16324 23614
rect 15148 23378 15428 23380
rect 15148 23326 15150 23378
rect 15202 23326 15428 23378
rect 15148 23324 15428 23326
rect 15932 23380 15988 23390
rect 15148 23314 15204 23324
rect 13804 23266 13860 23278
rect 13804 23214 13806 23266
rect 13858 23214 13860 23266
rect 13804 22708 13860 23214
rect 14588 23156 14644 23166
rect 14588 23062 14644 23100
rect 15932 23154 15988 23324
rect 15932 23102 15934 23154
rect 15986 23102 15988 23154
rect 15932 23090 15988 23102
rect 16268 23266 16324 23548
rect 16268 23214 16270 23266
rect 16322 23214 16324 23266
rect 13804 22642 13860 22652
rect 13916 22932 13972 22942
rect 15596 22932 15652 22942
rect 13580 22542 13582 22594
rect 13634 22542 13636 22594
rect 13580 22530 13636 22542
rect 13916 22594 13972 22876
rect 13916 22542 13918 22594
rect 13970 22542 13972 22594
rect 13916 22530 13972 22542
rect 15484 22930 15652 22932
rect 15484 22878 15598 22930
rect 15650 22878 15652 22930
rect 15484 22876 15652 22878
rect 15372 22372 15428 22382
rect 14140 22260 14196 22270
rect 14140 22166 14196 22204
rect 14700 22260 14756 22270
rect 14700 22166 14756 22204
rect 13692 22148 13748 22158
rect 13692 21810 13748 22092
rect 14008 21980 15208 21990
rect 14064 21978 14112 21980
rect 14168 21978 14216 21980
rect 14076 21926 14112 21978
rect 14200 21926 14216 21978
rect 14064 21924 14112 21926
rect 14168 21924 14216 21926
rect 14272 21978 14320 21980
rect 14376 21978 14424 21980
rect 14480 21978 14528 21980
rect 14376 21926 14396 21978
rect 14480 21926 14520 21978
rect 14272 21924 14320 21926
rect 14376 21924 14424 21926
rect 14480 21924 14528 21926
rect 14584 21924 14632 21980
rect 14688 21978 14736 21980
rect 14792 21978 14840 21980
rect 14896 21978 14944 21980
rect 14696 21926 14736 21978
rect 14820 21926 14840 21978
rect 14688 21924 14736 21926
rect 14792 21924 14840 21926
rect 14896 21924 14944 21926
rect 15000 21978 15048 21980
rect 15104 21978 15152 21980
rect 15000 21926 15016 21978
rect 15104 21926 15140 21978
rect 15000 21924 15048 21926
rect 15104 21924 15152 21926
rect 14008 21914 15208 21924
rect 15260 21812 15316 21822
rect 13692 21758 13694 21810
rect 13746 21758 13748 21810
rect 13692 21252 13748 21758
rect 15148 21756 15260 21812
rect 15148 21754 15204 21756
rect 15036 21698 15092 21710
rect 15036 21646 15038 21698
rect 15090 21646 15092 21698
rect 15148 21702 15150 21754
rect 15202 21702 15204 21754
rect 15260 21746 15316 21756
rect 15148 21690 15204 21702
rect 15036 21588 15092 21646
rect 15036 21532 15204 21588
rect 13692 21186 13748 21196
rect 14140 21474 14196 21486
rect 14140 21422 14142 21474
rect 14194 21422 14196 21474
rect 14140 21028 14196 21422
rect 14140 20962 14196 20972
rect 14588 21474 14644 21486
rect 14588 21422 14590 21474
rect 14642 21422 14644 21474
rect 13692 20916 13748 20926
rect 13692 20578 13748 20860
rect 13692 20526 13694 20578
rect 13746 20526 13748 20578
rect 13692 20468 13748 20526
rect 14140 20580 14196 20618
rect 14140 20514 14196 20524
rect 14588 20580 14644 21422
rect 15036 21362 15092 21374
rect 15036 21310 15038 21362
rect 15090 21310 15092 21362
rect 15036 20580 15092 21310
rect 15148 21364 15204 21532
rect 15148 21298 15204 21308
rect 15148 20916 15204 20926
rect 15372 20916 15428 22316
rect 15484 21588 15540 22876
rect 15596 22866 15652 22876
rect 15932 22372 15988 22382
rect 15596 22370 15988 22372
rect 15596 22318 15934 22370
rect 15986 22318 15988 22370
rect 15596 22316 15988 22318
rect 15596 21810 15652 22316
rect 15932 22306 15988 22316
rect 15596 21758 15598 21810
rect 15650 21758 15652 21810
rect 15596 21746 15652 21758
rect 15932 21588 15988 21598
rect 15484 21586 15988 21588
rect 15484 21534 15934 21586
rect 15986 21534 15988 21586
rect 15484 21532 15988 21534
rect 15932 21522 15988 21532
rect 15204 20860 15428 20916
rect 15596 21364 15652 21374
rect 15596 20914 15652 21308
rect 15596 20862 15598 20914
rect 15650 20862 15652 20914
rect 15148 20822 15204 20860
rect 15036 20524 15428 20580
rect 14588 20514 14644 20524
rect 13468 20412 13748 20468
rect 14008 20412 15208 20422
rect 13244 16772 13300 17164
rect 13356 16996 13412 17006
rect 13468 16996 13524 20412
rect 14064 20410 14112 20412
rect 14168 20410 14216 20412
rect 14076 20358 14112 20410
rect 14200 20358 14216 20410
rect 14064 20356 14112 20358
rect 14168 20356 14216 20358
rect 14272 20410 14320 20412
rect 14376 20410 14424 20412
rect 14480 20410 14528 20412
rect 14376 20358 14396 20410
rect 14480 20358 14520 20410
rect 14272 20356 14320 20358
rect 14376 20356 14424 20358
rect 14480 20356 14528 20358
rect 14584 20356 14632 20412
rect 14688 20410 14736 20412
rect 14792 20410 14840 20412
rect 14896 20410 14944 20412
rect 14696 20358 14736 20410
rect 14820 20358 14840 20410
rect 14688 20356 14736 20358
rect 14792 20356 14840 20358
rect 14896 20356 14944 20358
rect 15000 20410 15048 20412
rect 15104 20410 15152 20412
rect 15000 20358 15016 20410
rect 15104 20358 15140 20410
rect 15000 20356 15048 20358
rect 15104 20356 15152 20358
rect 14008 20346 15208 20356
rect 14028 20244 14084 20254
rect 15372 20244 15428 20524
rect 14084 20188 14196 20244
rect 14028 20178 14084 20188
rect 13692 20132 13748 20142
rect 13692 19348 13748 20076
rect 13916 20130 13972 20142
rect 13916 20078 13918 20130
rect 13970 20078 13972 20130
rect 13916 20020 13972 20078
rect 14140 20130 14196 20188
rect 14140 20078 14142 20130
rect 14194 20078 14196 20130
rect 14140 20066 14196 20078
rect 15036 20188 15428 20244
rect 13916 19954 13972 19964
rect 14364 20018 14420 20030
rect 14364 19966 14366 20018
rect 14418 19966 14420 20018
rect 14252 19908 14308 19918
rect 14252 19814 14308 19852
rect 13692 19292 13860 19348
rect 13692 19124 13748 19134
rect 13692 18228 13748 19068
rect 13804 18562 13860 19292
rect 14364 19124 14420 19966
rect 14812 20020 14868 20030
rect 14812 19926 14868 19964
rect 14588 19348 14644 19386
rect 14588 19282 14644 19292
rect 14700 19236 14756 19246
rect 14700 19142 14756 19180
rect 15036 19234 15092 20188
rect 15596 20132 15652 20862
rect 15596 20066 15652 20076
rect 16044 20132 16100 20142
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 15036 19170 15092 19182
rect 15708 19908 15764 19918
rect 14420 19068 14532 19124
rect 14364 19058 14420 19068
rect 14252 19012 14308 19050
rect 14252 18946 14308 18956
rect 14476 19010 14532 19068
rect 14476 18958 14478 19010
rect 14530 18958 14532 19010
rect 14476 18946 14532 18958
rect 14008 18844 15208 18854
rect 14064 18842 14112 18844
rect 14168 18842 14216 18844
rect 14076 18790 14112 18842
rect 14200 18790 14216 18842
rect 14064 18788 14112 18790
rect 14168 18788 14216 18790
rect 14272 18842 14320 18844
rect 14376 18842 14424 18844
rect 14480 18842 14528 18844
rect 14376 18790 14396 18842
rect 14480 18790 14520 18842
rect 14272 18788 14320 18790
rect 14376 18788 14424 18790
rect 14480 18788 14528 18790
rect 14584 18788 14632 18844
rect 14688 18842 14736 18844
rect 14792 18842 14840 18844
rect 14896 18842 14944 18844
rect 14696 18790 14736 18842
rect 14820 18790 14840 18842
rect 14688 18788 14736 18790
rect 14792 18788 14840 18790
rect 14896 18788 14944 18790
rect 15000 18842 15048 18844
rect 15104 18842 15152 18844
rect 15000 18790 15016 18842
rect 15104 18790 15140 18842
rect 15000 18788 15048 18790
rect 15104 18788 15152 18790
rect 14008 18778 15208 18788
rect 15372 18674 15428 18686
rect 15372 18622 15374 18674
rect 15426 18622 15428 18674
rect 13804 18510 13806 18562
rect 13858 18510 13860 18562
rect 13804 18498 13860 18510
rect 13916 18564 13972 18574
rect 13916 18450 13972 18508
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13916 18386 13972 18398
rect 14812 18450 14868 18462
rect 14812 18398 14814 18450
rect 14866 18398 14868 18450
rect 14812 18340 14868 18398
rect 15372 18452 15428 18622
rect 15708 18562 15764 19852
rect 15708 18510 15710 18562
rect 15762 18510 15764 18562
rect 15708 18498 15764 18510
rect 15820 19348 15876 19358
rect 15596 18452 15652 18462
rect 15372 18450 15652 18452
rect 15372 18398 15598 18450
rect 15650 18398 15652 18450
rect 15372 18396 15652 18398
rect 15596 18386 15652 18396
rect 14812 18274 14868 18284
rect 15820 18340 15876 19292
rect 15820 18274 15876 18284
rect 13692 18172 13972 18228
rect 13804 18004 13860 18014
rect 13580 17892 13636 17902
rect 13804 17892 13860 17948
rect 13580 17890 13860 17892
rect 13580 17838 13582 17890
rect 13634 17838 13860 17890
rect 13580 17836 13860 17838
rect 13580 17826 13636 17836
rect 13916 17780 13972 18172
rect 13356 16994 13524 16996
rect 13356 16942 13358 16994
rect 13410 16942 13524 16994
rect 13356 16940 13524 16942
rect 13692 17724 13972 17780
rect 13356 16930 13412 16940
rect 13244 16212 13300 16716
rect 13580 16660 13636 16670
rect 13244 16146 13300 16156
rect 13356 16436 13412 16446
rect 13132 15810 13188 15820
rect 12908 15538 13076 15540
rect 12908 15486 12910 15538
rect 12962 15486 13076 15538
rect 12908 15484 13076 15486
rect 13356 15538 13412 16380
rect 13580 16210 13636 16604
rect 13692 16322 13748 17724
rect 14364 17444 14420 17482
rect 14364 17378 14420 17388
rect 14008 17276 15208 17286
rect 14064 17274 14112 17276
rect 14168 17274 14216 17276
rect 14076 17222 14112 17274
rect 14200 17222 14216 17274
rect 14064 17220 14112 17222
rect 14168 17220 14216 17222
rect 14272 17274 14320 17276
rect 14376 17274 14424 17276
rect 14480 17274 14528 17276
rect 14376 17222 14396 17274
rect 14480 17222 14520 17274
rect 14272 17220 14320 17222
rect 14376 17220 14424 17222
rect 14480 17220 14528 17222
rect 14584 17220 14632 17276
rect 14688 17274 14736 17276
rect 14792 17274 14840 17276
rect 14896 17274 14944 17276
rect 14696 17222 14736 17274
rect 14820 17222 14840 17274
rect 14688 17220 14736 17222
rect 14792 17220 14840 17222
rect 14896 17220 14944 17222
rect 15000 17274 15048 17276
rect 15104 17274 15152 17276
rect 15000 17222 15016 17274
rect 15104 17222 15140 17274
rect 15000 17220 15048 17222
rect 15104 17220 15152 17222
rect 14008 17210 15208 17220
rect 15372 17220 15428 17230
rect 14924 17108 14980 17118
rect 15372 17108 15428 17164
rect 14924 16882 14980 17052
rect 14924 16830 14926 16882
rect 14978 16830 14980 16882
rect 14588 16658 14644 16670
rect 14588 16606 14590 16658
rect 14642 16606 14644 16658
rect 13692 16270 13694 16322
rect 13746 16270 13748 16322
rect 13692 16258 13748 16270
rect 14028 16324 14084 16334
rect 13580 16158 13582 16210
rect 13634 16158 13636 16210
rect 13580 16146 13636 16158
rect 14028 16210 14084 16268
rect 14028 16158 14030 16210
rect 14082 16158 14084 16210
rect 14028 16146 14084 16158
rect 14028 15988 14084 15998
rect 14028 15876 14084 15932
rect 14588 15988 14644 16606
rect 14700 16212 14756 16222
rect 14924 16212 14980 16830
rect 15260 17052 15428 17108
rect 15260 16436 15316 17052
rect 15484 16996 15540 17006
rect 15484 16902 15540 16940
rect 15708 16996 15764 17006
rect 15596 16884 15652 16894
rect 15260 16380 15428 16436
rect 15036 16212 15092 16222
rect 14924 16210 15092 16212
rect 14924 16158 15038 16210
rect 15090 16158 15092 16210
rect 14924 16156 15092 16158
rect 14700 16118 14756 16156
rect 15036 16146 15092 16156
rect 14588 15922 14644 15932
rect 13356 15486 13358 15538
rect 13410 15486 13412 15538
rect 12908 15474 12964 15484
rect 13356 15474 13412 15486
rect 13804 15820 14084 15876
rect 14140 15876 14196 15914
rect 12796 15262 12798 15314
rect 12850 15262 12852 15314
rect 12796 15250 12852 15262
rect 13132 15314 13188 15326
rect 13132 15262 13134 15314
rect 13186 15262 13188 15314
rect 12796 14980 12852 14990
rect 12796 14642 12852 14924
rect 12796 14590 12798 14642
rect 12850 14590 12852 14642
rect 12796 14578 12852 14590
rect 13132 14644 13188 15262
rect 13356 15314 13412 15326
rect 13356 15262 13358 15314
rect 13410 15262 13412 15314
rect 13356 14980 13412 15262
rect 13412 14924 13636 14980
rect 13356 14914 13412 14924
rect 13132 14578 13188 14588
rect 13580 14642 13636 14924
rect 13580 14590 13582 14642
rect 13634 14590 13636 14642
rect 13580 14578 13636 14590
rect 13468 13972 13524 13982
rect 12460 13682 12516 13692
rect 13244 13748 13300 13758
rect 12012 13634 12180 13636
rect 12012 13582 12014 13634
rect 12066 13582 12180 13634
rect 12012 13580 12180 13582
rect 12012 13570 12068 13580
rect 11452 12962 11620 12964
rect 11452 12910 11454 12962
rect 11506 12910 11620 12962
rect 11452 12908 11620 12910
rect 11676 13076 11732 13086
rect 11452 12898 11508 12908
rect 11340 12740 11396 12750
rect 11004 12738 11396 12740
rect 11004 12686 11342 12738
rect 11394 12686 11396 12738
rect 11004 12684 11396 12686
rect 10556 12350 10558 12402
rect 10610 12350 10612 12402
rect 10556 12338 10612 12350
rect 10892 12404 10948 12414
rect 10892 12310 10948 12348
rect 10220 12180 10276 12190
rect 10220 12086 10276 12124
rect 9660 11172 9716 11182
rect 9436 11116 9660 11172
rect 8876 10610 8932 11116
rect 9660 10836 9716 11116
rect 10892 11170 10948 11182
rect 10892 11118 10894 11170
rect 10946 11118 10948 11170
rect 10892 11060 10948 11118
rect 10108 10836 10164 10846
rect 9660 10834 10388 10836
rect 9660 10782 9662 10834
rect 9714 10782 10110 10834
rect 10162 10782 10388 10834
rect 9660 10780 10388 10782
rect 9660 10770 9716 10780
rect 10108 10770 10164 10780
rect 8876 10558 8878 10610
rect 8930 10558 8932 10610
rect 8876 10546 8932 10558
rect 10332 10610 10388 10780
rect 10332 10558 10334 10610
rect 10386 10558 10388 10610
rect 10332 10546 10388 10558
rect 5740 9550 5742 9602
rect 5794 9550 5796 9602
rect 4008 8652 5208 8662
rect 4064 8650 4112 8652
rect 4168 8650 4216 8652
rect 4076 8598 4112 8650
rect 4200 8598 4216 8650
rect 4064 8596 4112 8598
rect 4168 8596 4216 8598
rect 4272 8650 4320 8652
rect 4376 8650 4424 8652
rect 4480 8650 4528 8652
rect 4376 8598 4396 8650
rect 4480 8598 4520 8650
rect 4272 8596 4320 8598
rect 4376 8596 4424 8598
rect 4480 8596 4528 8598
rect 4584 8596 4632 8652
rect 4688 8650 4736 8652
rect 4792 8650 4840 8652
rect 4896 8650 4944 8652
rect 4696 8598 4736 8650
rect 4820 8598 4840 8650
rect 4688 8596 4736 8598
rect 4792 8596 4840 8598
rect 4896 8596 4944 8598
rect 5000 8650 5048 8652
rect 5104 8650 5152 8652
rect 5000 8598 5016 8650
rect 5104 8598 5140 8650
rect 5000 8596 5048 8598
rect 5104 8596 5152 8598
rect 4008 8586 5208 8596
rect 5404 8036 5460 8046
rect 4732 7700 4788 7710
rect 4732 7606 4788 7644
rect 5292 7250 5348 7262
rect 5292 7198 5294 7250
rect 5346 7198 5348 7250
rect 4008 7084 5208 7094
rect 4064 7082 4112 7084
rect 4168 7082 4216 7084
rect 4076 7030 4112 7082
rect 4200 7030 4216 7082
rect 4064 7028 4112 7030
rect 4168 7028 4216 7030
rect 4272 7082 4320 7084
rect 4376 7082 4424 7084
rect 4480 7082 4528 7084
rect 4376 7030 4396 7082
rect 4480 7030 4520 7082
rect 4272 7028 4320 7030
rect 4376 7028 4424 7030
rect 4480 7028 4528 7030
rect 4584 7028 4632 7084
rect 4688 7082 4736 7084
rect 4792 7082 4840 7084
rect 4896 7082 4944 7084
rect 4696 7030 4736 7082
rect 4820 7030 4840 7082
rect 4688 7028 4736 7030
rect 4792 7028 4840 7030
rect 4896 7028 4944 7030
rect 5000 7082 5048 7084
rect 5104 7082 5152 7084
rect 5000 7030 5016 7082
rect 5104 7030 5140 7082
rect 5000 7028 5048 7030
rect 5104 7028 5152 7030
rect 4008 7018 5208 7028
rect 3612 6738 3668 6748
rect 4172 6916 4228 6926
rect 2268 6692 2324 6702
rect 2492 6692 2548 6702
rect 2268 6690 2492 6692
rect 2268 6638 2270 6690
rect 2322 6638 2492 6690
rect 2268 6636 2492 6638
rect 2268 6626 2324 6636
rect 2492 6598 2548 6636
rect 4060 6692 4116 6702
rect 4060 6598 4116 6636
rect 2604 6580 2660 6590
rect 2940 6580 2996 6590
rect 2604 6578 2996 6580
rect 2604 6526 2606 6578
rect 2658 6526 2942 6578
rect 2994 6526 2996 6578
rect 2604 6524 2996 6526
rect 2604 6514 2660 6524
rect 2940 6514 2996 6524
rect 3612 6578 3668 6590
rect 3612 6526 3614 6578
rect 3666 6526 3668 6578
rect 3052 6468 3108 6478
rect 3276 6468 3332 6478
rect 3612 6468 3668 6526
rect 3052 6374 3108 6412
rect 3164 6466 3332 6468
rect 3164 6414 3278 6466
rect 3330 6414 3332 6466
rect 3164 6412 3332 6414
rect 3164 6244 3220 6412
rect 3276 6402 3332 6412
rect 3388 6412 3668 6468
rect 3388 6244 3444 6412
rect 2156 5954 2212 5964
rect 2492 6188 3220 6244
rect 3276 6188 3444 6244
rect 2492 6018 2548 6188
rect 2492 5966 2494 6018
rect 2546 5966 2548 6018
rect 2492 5954 2548 5966
rect 3164 6020 3220 6030
rect 3276 6020 3332 6188
rect 3164 6018 3332 6020
rect 3164 5966 3166 6018
rect 3218 5966 3332 6018
rect 3164 5964 3332 5966
rect 3500 6020 3556 6030
rect 3164 5954 3220 5964
rect 3500 5926 3556 5964
rect 2828 5906 2884 5918
rect 2828 5854 2830 5906
rect 2882 5854 2884 5906
rect 2044 5794 2100 5806
rect 2044 5742 2046 5794
rect 2098 5742 2100 5794
rect 2044 5684 2100 5742
rect 2380 5684 2436 5694
rect 2044 5618 2100 5628
rect 2268 5682 2436 5684
rect 2268 5630 2382 5682
rect 2434 5630 2436 5682
rect 2268 5628 2436 5630
rect 1932 4340 1988 4350
rect 1708 4338 1932 4340
rect 1708 4286 1710 4338
rect 1762 4286 1932 4338
rect 1708 4284 1932 4286
rect 1708 4274 1764 4284
rect 1932 4274 1988 4284
rect 2268 4338 2324 5628
rect 2380 5618 2436 5628
rect 2828 5684 2884 5854
rect 4172 5906 4228 6860
rect 4508 6804 4564 6814
rect 4508 6710 4564 6748
rect 4732 6804 4788 6814
rect 4172 5854 4174 5906
rect 4226 5854 4228 5906
rect 3612 5796 3668 5806
rect 4172 5796 4228 5854
rect 4732 5906 4788 6748
rect 4732 5854 4734 5906
rect 4786 5854 4788 5906
rect 4732 5842 4788 5854
rect 5292 6692 5348 7198
rect 3612 5702 3668 5740
rect 3836 5740 4228 5796
rect 2828 5618 2884 5628
rect 2268 4286 2270 4338
rect 2322 4286 2324 4338
rect 2268 4274 2324 4286
rect 3836 4340 3892 5740
rect 4008 5516 5208 5526
rect 4064 5514 4112 5516
rect 4168 5514 4216 5516
rect 4076 5462 4112 5514
rect 4200 5462 4216 5514
rect 4064 5460 4112 5462
rect 4168 5460 4216 5462
rect 4272 5514 4320 5516
rect 4376 5514 4424 5516
rect 4480 5514 4528 5516
rect 4376 5462 4396 5514
rect 4480 5462 4520 5514
rect 4272 5460 4320 5462
rect 4376 5460 4424 5462
rect 4480 5460 4528 5462
rect 4584 5460 4632 5516
rect 4688 5514 4736 5516
rect 4792 5514 4840 5516
rect 4896 5514 4944 5516
rect 4696 5462 4736 5514
rect 4820 5462 4840 5514
rect 4688 5460 4736 5462
rect 4792 5460 4840 5462
rect 4896 5460 4944 5462
rect 5000 5514 5048 5516
rect 5104 5514 5152 5516
rect 5000 5462 5016 5514
rect 5104 5462 5140 5514
rect 5000 5460 5048 5462
rect 5104 5460 5152 5462
rect 4008 5450 5208 5460
rect 5292 5124 5348 6636
rect 5292 5058 5348 5068
rect 4732 5012 4788 5022
rect 4732 4562 4788 4956
rect 4732 4510 4734 4562
rect 4786 4510 4788 4562
rect 4732 4498 4788 4510
rect 5404 4564 5460 7980
rect 5516 7364 5572 7374
rect 5516 6692 5572 7308
rect 5628 7364 5684 7374
rect 5740 7364 5796 9550
rect 6076 9938 6244 9940
rect 6076 9886 6190 9938
rect 6242 9886 6244 9938
rect 6076 9884 6244 9886
rect 6076 8372 6132 9884
rect 6188 9874 6244 9884
rect 9212 10164 9268 10174
rect 9212 9602 9268 10108
rect 10892 10164 10948 11004
rect 11004 10610 11060 12684
rect 11340 12674 11396 12684
rect 11676 11618 11732 13020
rect 12908 12852 12964 12862
rect 12908 12758 12964 12796
rect 13244 12402 13300 13692
rect 13468 12516 13524 13916
rect 13804 13188 13860 15820
rect 14140 15810 14196 15820
rect 14008 15708 15208 15718
rect 14064 15706 14112 15708
rect 14168 15706 14216 15708
rect 14076 15654 14112 15706
rect 14200 15654 14216 15706
rect 14064 15652 14112 15654
rect 14168 15652 14216 15654
rect 14272 15706 14320 15708
rect 14376 15706 14424 15708
rect 14480 15706 14528 15708
rect 14376 15654 14396 15706
rect 14480 15654 14520 15706
rect 14272 15652 14320 15654
rect 14376 15652 14424 15654
rect 14480 15652 14528 15654
rect 14584 15652 14632 15708
rect 14688 15706 14736 15708
rect 14792 15706 14840 15708
rect 14896 15706 14944 15708
rect 14696 15654 14736 15706
rect 14820 15654 14840 15706
rect 14688 15652 14736 15654
rect 14792 15652 14840 15654
rect 14896 15652 14944 15654
rect 15000 15706 15048 15708
rect 15104 15706 15152 15708
rect 15000 15654 15016 15706
rect 15104 15654 15140 15706
rect 15000 15652 15048 15654
rect 15104 15652 15152 15654
rect 14008 15642 15208 15652
rect 13916 15428 13972 15438
rect 13916 15334 13972 15372
rect 14364 15204 14420 15214
rect 14364 15110 14420 15148
rect 15372 14532 15428 16380
rect 15148 14420 15204 14430
rect 15372 14420 15428 14476
rect 15148 14418 15428 14420
rect 15148 14366 15150 14418
rect 15202 14366 15428 14418
rect 15148 14364 15428 14366
rect 15148 14354 15204 14364
rect 14008 14140 15208 14150
rect 14064 14138 14112 14140
rect 14168 14138 14216 14140
rect 14076 14086 14112 14138
rect 14200 14086 14216 14138
rect 14064 14084 14112 14086
rect 14168 14084 14216 14086
rect 14272 14138 14320 14140
rect 14376 14138 14424 14140
rect 14480 14138 14528 14140
rect 14376 14086 14396 14138
rect 14480 14086 14520 14138
rect 14272 14084 14320 14086
rect 14376 14084 14424 14086
rect 14480 14084 14528 14086
rect 14584 14084 14632 14140
rect 14688 14138 14736 14140
rect 14792 14138 14840 14140
rect 14896 14138 14944 14140
rect 14696 14086 14736 14138
rect 14820 14086 14840 14138
rect 14688 14084 14736 14086
rect 14792 14084 14840 14086
rect 14896 14084 14944 14086
rect 15000 14138 15048 14140
rect 15104 14138 15152 14140
rect 15000 14086 15016 14138
rect 15104 14086 15140 14138
rect 15000 14084 15048 14086
rect 15104 14084 15152 14086
rect 14008 14074 15208 14084
rect 14252 13748 14308 13758
rect 14252 13654 14308 13692
rect 14812 13748 14868 13758
rect 14812 13654 14868 13692
rect 15372 13748 15428 14364
rect 15372 13682 15428 13692
rect 15596 13970 15652 16828
rect 15708 16882 15764 16940
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 15428 15764 16830
rect 15708 15362 15764 15372
rect 15596 13918 15598 13970
rect 15650 13918 15652 13970
rect 14924 13634 14980 13646
rect 14924 13582 14926 13634
rect 14978 13582 14980 13634
rect 14028 13188 14084 13198
rect 13804 13186 14084 13188
rect 13804 13134 14030 13186
rect 14082 13134 14084 13186
rect 13804 13132 14084 13134
rect 14028 13122 14084 13132
rect 14924 13188 14980 13582
rect 14924 13122 14980 13132
rect 15260 13524 15316 13534
rect 14364 12852 14420 12862
rect 14364 12758 14420 12796
rect 14588 12850 14644 12862
rect 14588 12798 14590 12850
rect 14642 12798 14644 12850
rect 13692 12740 13748 12750
rect 14588 12740 14644 12798
rect 13692 12738 13860 12740
rect 13692 12686 13694 12738
rect 13746 12686 13860 12738
rect 13692 12684 13860 12686
rect 13692 12674 13748 12684
rect 13468 12460 13748 12516
rect 13244 12350 13246 12402
rect 13298 12350 13300 12402
rect 13244 12338 13300 12350
rect 13580 11844 13636 11854
rect 11676 11566 11678 11618
rect 11730 11566 11732 11618
rect 11676 11554 11732 11566
rect 13244 11620 13300 11630
rect 12012 11172 12068 11182
rect 12012 11078 12068 11116
rect 12460 11170 12516 11182
rect 12460 11118 12462 11170
rect 12514 11118 12516 11170
rect 12460 11060 12516 11118
rect 12460 10994 12516 11004
rect 13244 11060 13300 11564
rect 13244 10836 13300 11004
rect 13244 10742 13300 10780
rect 13580 11394 13636 11788
rect 13580 11342 13582 11394
rect 13634 11342 13636 11394
rect 11004 10558 11006 10610
rect 11058 10558 11060 10610
rect 11004 10546 11060 10558
rect 10892 10098 10948 10108
rect 9212 9550 9214 9602
rect 9266 9550 9268 9602
rect 5852 8036 5908 8046
rect 5852 7942 5908 7980
rect 6076 7700 6132 8316
rect 7308 8372 7364 8382
rect 6636 8036 6692 8046
rect 6692 7980 6804 8036
rect 6636 7970 6692 7980
rect 6076 7606 6132 7644
rect 6748 7476 6804 7980
rect 5628 7362 5796 7364
rect 5628 7310 5630 7362
rect 5682 7310 5796 7362
rect 5628 7308 5796 7310
rect 6636 7364 6692 7374
rect 5628 6916 5684 7308
rect 6636 7270 6692 7308
rect 6524 7250 6580 7262
rect 6524 7198 6526 7250
rect 6578 7198 6580 7250
rect 5628 6850 5684 6860
rect 5740 6972 6132 7028
rect 5740 6914 5796 6972
rect 5740 6862 5742 6914
rect 5794 6862 5796 6914
rect 5740 6850 5796 6862
rect 6076 6916 6132 6972
rect 6188 6916 6244 6926
rect 6076 6914 6244 6916
rect 6076 6862 6190 6914
rect 6242 6862 6244 6914
rect 6076 6860 6244 6862
rect 6188 6850 6244 6860
rect 6300 6914 6356 6926
rect 6300 6862 6302 6914
rect 6354 6862 6356 6914
rect 6300 6804 6356 6862
rect 6524 6916 6580 7198
rect 6748 7140 6804 7420
rect 6860 7474 6916 7486
rect 6860 7422 6862 7474
rect 6914 7422 6916 7474
rect 6860 7364 6916 7422
rect 6860 7298 6916 7308
rect 6748 7084 7028 7140
rect 6748 6916 6804 6926
rect 6524 6914 6804 6916
rect 6524 6862 6750 6914
rect 6802 6862 6804 6914
rect 6524 6860 6804 6862
rect 6300 6738 6356 6748
rect 5852 6692 5908 6702
rect 5516 6690 5908 6692
rect 5516 6638 5854 6690
rect 5906 6638 5908 6690
rect 5516 6636 5908 6638
rect 5740 6468 5796 6478
rect 5740 5122 5796 6412
rect 5740 5070 5742 5122
rect 5794 5070 5796 5122
rect 5740 5058 5796 5070
rect 5852 5122 5908 6636
rect 6748 6692 6804 6860
rect 6972 6914 7028 7084
rect 6972 6862 6974 6914
rect 7026 6862 7028 6914
rect 6972 6850 7028 6862
rect 6412 6580 6468 6590
rect 6412 6486 6468 6524
rect 6748 5908 6804 6636
rect 5964 5796 6020 5806
rect 5964 5234 6020 5740
rect 6748 5348 6804 5852
rect 7308 6130 7364 8316
rect 7980 8372 8036 8382
rect 7980 8278 8036 8316
rect 9212 8372 9268 9550
rect 9212 8306 9268 8316
rect 7980 7586 8036 7598
rect 7980 7534 7982 7586
rect 8034 7534 8036 7586
rect 7532 7476 7588 7486
rect 7532 7382 7588 7420
rect 7980 7476 8036 7534
rect 8540 7586 8596 7598
rect 8540 7534 8542 7586
rect 8594 7534 8596 7586
rect 7980 7410 8036 7420
rect 8092 7476 8148 7486
rect 8092 7474 8372 7476
rect 8092 7422 8094 7474
rect 8146 7422 8372 7474
rect 8092 7420 8372 7422
rect 8092 7410 8148 7420
rect 7644 7364 7700 7374
rect 7700 7308 7924 7364
rect 7644 7298 7700 7308
rect 7756 6692 7812 6702
rect 7756 6598 7812 6636
rect 7308 6078 7310 6130
rect 7362 6078 7364 6130
rect 6860 5348 6916 5358
rect 5964 5182 5966 5234
rect 6018 5182 6020 5234
rect 5964 5170 6020 5182
rect 6524 5346 6916 5348
rect 6524 5294 6862 5346
rect 6914 5294 6916 5346
rect 6524 5292 6916 5294
rect 5852 5070 5854 5122
rect 5906 5070 5908 5122
rect 5852 5058 5908 5070
rect 6076 5124 6132 5134
rect 6076 5030 6132 5068
rect 6300 5124 6356 5134
rect 6300 5122 6468 5124
rect 6300 5070 6302 5122
rect 6354 5070 6468 5122
rect 6300 5068 6468 5070
rect 6300 5058 6356 5068
rect 6076 4564 6132 4574
rect 6300 4564 6356 4574
rect 5404 4562 6356 4564
rect 5404 4510 6078 4562
rect 6130 4510 6302 4562
rect 6354 4510 6356 4562
rect 5404 4508 6356 4510
rect 5404 4450 5460 4508
rect 6076 4498 6132 4508
rect 6300 4498 6356 4508
rect 6412 4562 6468 5068
rect 6412 4510 6414 4562
rect 6466 4510 6468 4562
rect 6412 4498 6468 4510
rect 6524 4562 6580 5292
rect 6860 5282 6916 5292
rect 6524 4510 6526 4562
rect 6578 4510 6580 4562
rect 6524 4498 6580 4510
rect 6636 5012 6692 5022
rect 5404 4398 5406 4450
rect 5458 4398 5460 4450
rect 5404 4386 5460 4398
rect 3836 4274 3892 4284
rect 5964 4340 6020 4350
rect 6636 4340 6692 4956
rect 7308 5012 7364 6078
rect 7532 6578 7588 6590
rect 7532 6526 7534 6578
rect 7586 6526 7588 6578
rect 7532 6468 7588 6526
rect 7532 5796 7588 6412
rect 7868 6132 7924 7308
rect 7980 7252 8036 7262
rect 7980 7158 8036 7196
rect 8092 6916 8148 6926
rect 8092 6822 8148 6860
rect 8316 6804 8372 7420
rect 8204 6748 8372 6804
rect 8428 7474 8484 7486
rect 8428 7422 8430 7474
rect 8482 7422 8484 7474
rect 8428 7252 8484 7422
rect 7980 6580 8036 6590
rect 8036 6524 8148 6580
rect 7980 6486 8036 6524
rect 7532 5730 7588 5740
rect 7644 6130 7924 6132
rect 7644 6078 7870 6130
rect 7922 6078 7924 6130
rect 7644 6076 7924 6078
rect 7308 4946 7364 4956
rect 7532 5012 7588 5022
rect 7532 4898 7588 4956
rect 7532 4846 7534 4898
rect 7586 4846 7588 4898
rect 7532 4834 7588 4846
rect 7644 4676 7700 6076
rect 7868 6066 7924 6076
rect 7420 4620 7700 4676
rect 7420 4452 7476 4620
rect 4008 3948 5208 3958
rect 4064 3946 4112 3948
rect 4168 3946 4216 3948
rect 4076 3894 4112 3946
rect 4200 3894 4216 3946
rect 4064 3892 4112 3894
rect 4168 3892 4216 3894
rect 4272 3946 4320 3948
rect 4376 3946 4424 3948
rect 4480 3946 4528 3948
rect 4376 3894 4396 3946
rect 4480 3894 4520 3946
rect 4272 3892 4320 3894
rect 4376 3892 4424 3894
rect 4480 3892 4528 3894
rect 4584 3892 4632 3948
rect 4688 3946 4736 3948
rect 4792 3946 4840 3948
rect 4896 3946 4944 3948
rect 4696 3894 4736 3946
rect 4820 3894 4840 3946
rect 4688 3892 4736 3894
rect 4792 3892 4840 3894
rect 4896 3892 4944 3894
rect 5000 3946 5048 3948
rect 5104 3946 5152 3948
rect 5000 3894 5016 3946
rect 5104 3894 5140 3946
rect 5000 3892 5048 3894
rect 5104 3892 5152 3894
rect 4008 3882 5208 3892
rect 5964 3668 6020 4284
rect 5964 3574 6020 3612
rect 6412 4284 6692 4340
rect 6972 4450 7476 4452
rect 6972 4398 7422 4450
rect 7474 4398 7476 4450
rect 6972 4396 7476 4398
rect 6972 4338 7028 4396
rect 7420 4386 7476 4396
rect 8092 4340 8148 6524
rect 8204 5684 8260 6748
rect 8316 6580 8372 6590
rect 8316 6018 8372 6524
rect 8428 6132 8484 7196
rect 8540 6916 8596 7534
rect 11900 7586 11956 7598
rect 11900 7534 11902 7586
rect 11954 7534 11956 7586
rect 8540 6850 8596 6860
rect 8764 7474 8820 7486
rect 8764 7422 8766 7474
rect 8818 7422 8820 7474
rect 8764 6916 8820 7422
rect 8764 6850 8820 6860
rect 9660 7364 9716 7374
rect 10108 7364 10164 7374
rect 9660 7362 10164 7364
rect 9660 7310 9662 7362
rect 9714 7310 10110 7362
rect 10162 7310 10164 7362
rect 9660 7308 10164 7310
rect 8540 6692 8596 6702
rect 8540 6690 8932 6692
rect 8540 6638 8542 6690
rect 8594 6638 8932 6690
rect 8540 6636 8932 6638
rect 8540 6626 8596 6636
rect 8652 6466 8708 6478
rect 8652 6414 8654 6466
rect 8706 6414 8708 6466
rect 8540 6132 8596 6142
rect 8428 6076 8540 6132
rect 8540 6066 8596 6076
rect 8316 5966 8318 6018
rect 8370 5966 8372 6018
rect 8316 5954 8372 5966
rect 8428 5908 8484 5918
rect 8316 5684 8372 5694
rect 8204 5628 8316 5684
rect 8316 4562 8372 5628
rect 8316 4510 8318 4562
rect 8370 4510 8372 4562
rect 8316 4498 8372 4510
rect 8428 4450 8484 5852
rect 8540 5906 8596 5918
rect 8540 5854 8542 5906
rect 8594 5854 8596 5906
rect 8540 5796 8596 5854
rect 8540 5730 8596 5740
rect 8428 4398 8430 4450
rect 8482 4398 8484 4450
rect 8428 4386 8484 4398
rect 8652 4452 8708 6414
rect 8764 6466 8820 6478
rect 8764 6414 8766 6466
rect 8818 6414 8820 6466
rect 8764 5684 8820 6414
rect 8876 6132 8932 6636
rect 9212 6690 9268 6702
rect 9212 6638 9214 6690
rect 9266 6638 9268 6690
rect 8988 6132 9044 6142
rect 8876 6130 9044 6132
rect 8876 6078 8990 6130
rect 9042 6078 9044 6130
rect 8876 6076 9044 6078
rect 8988 6066 9044 6076
rect 8764 5618 8820 5628
rect 8876 5908 8932 5918
rect 8876 4562 8932 5852
rect 8876 4510 8878 4562
rect 8930 4510 8932 4562
rect 8876 4498 8932 4510
rect 9100 5908 9156 5918
rect 9100 4562 9156 5852
rect 9212 5684 9268 6638
rect 9212 5618 9268 5628
rect 9324 6692 9380 6702
rect 9660 6692 9716 7308
rect 10108 7298 10164 7308
rect 11116 7250 11172 7262
rect 11116 7198 11118 7250
rect 11170 7198 11172 7250
rect 9324 6690 9716 6692
rect 9324 6638 9326 6690
rect 9378 6638 9716 6690
rect 9324 6636 9716 6638
rect 9772 6916 9828 6926
rect 9324 5908 9380 6636
rect 9436 5908 9492 5918
rect 9324 5906 9492 5908
rect 9324 5854 9438 5906
rect 9490 5854 9492 5906
rect 9324 5852 9492 5854
rect 9100 4510 9102 4562
rect 9154 4510 9156 4562
rect 9100 4498 9156 4510
rect 9324 5124 9380 5852
rect 9436 5842 9492 5852
rect 9772 5124 9828 6860
rect 9996 6692 10052 6702
rect 9996 6598 10052 6636
rect 9996 5908 10052 5918
rect 9996 5814 10052 5852
rect 11116 5796 11172 7198
rect 11116 5730 11172 5740
rect 11900 6580 11956 7534
rect 13580 7476 13636 11342
rect 13692 10836 13748 12460
rect 13804 11396 13860 12684
rect 14588 12674 14644 12684
rect 15260 12740 15316 13468
rect 15596 12964 15652 13918
rect 16044 13970 16100 20076
rect 16268 16996 16324 23214
rect 16492 23266 16548 23278
rect 16492 23214 16494 23266
rect 16546 23214 16548 23266
rect 16380 21252 16436 21262
rect 16380 19796 16436 21196
rect 16492 20020 16548 23214
rect 16604 21588 16660 23772
rect 17052 23714 17108 23726
rect 17052 23662 17054 23714
rect 17106 23662 17108 23714
rect 17052 22260 17108 23662
rect 17052 22194 17108 22204
rect 17164 21868 17220 30156
rect 17836 30146 17892 30156
rect 17276 29986 17332 29998
rect 17276 29934 17278 29986
rect 17330 29934 17332 29986
rect 17276 29652 17332 29934
rect 17724 29652 17780 29662
rect 17276 29586 17332 29596
rect 17500 29650 17780 29652
rect 17500 29598 17726 29650
rect 17778 29598 17780 29650
rect 17500 29596 17780 29598
rect 17388 29428 17444 29438
rect 17388 29334 17444 29372
rect 17500 28082 17556 29596
rect 17724 29586 17780 29596
rect 17948 29538 18004 30716
rect 18172 30706 18228 30716
rect 17948 29486 17950 29538
rect 18002 29486 18004 29538
rect 17612 29426 17668 29438
rect 17612 29374 17614 29426
rect 17666 29374 17668 29426
rect 17612 28532 17668 29374
rect 17668 28476 17780 28532
rect 17612 28466 17668 28476
rect 17724 28084 17780 28476
rect 17500 28030 17502 28082
rect 17554 28030 17556 28082
rect 17500 28018 17556 28030
rect 17612 28082 17780 28084
rect 17612 28030 17726 28082
rect 17778 28030 17780 28082
rect 17612 28028 17780 28030
rect 17388 27188 17444 27198
rect 17612 27188 17668 28028
rect 17724 28018 17780 28028
rect 17948 28082 18004 29486
rect 18732 29428 18788 29438
rect 18732 29334 18788 29372
rect 18844 28868 18900 32844
rect 19740 30212 19796 30222
rect 19740 30118 19796 30156
rect 20076 30212 20132 33964
rect 20860 32564 20916 32574
rect 20076 29988 20132 30156
rect 20412 30212 20468 30222
rect 20860 30212 20916 32508
rect 20412 30210 20916 30212
rect 20412 30158 20414 30210
rect 20466 30158 20862 30210
rect 20914 30158 20916 30210
rect 20412 30156 20916 30158
rect 20412 30146 20468 30156
rect 20860 30146 20916 30156
rect 19740 29932 20132 29988
rect 19292 29652 19348 29662
rect 19292 29558 19348 29596
rect 19740 29652 19796 29932
rect 18844 28812 19684 28868
rect 18284 28644 18340 28654
rect 18284 28550 18340 28588
rect 17948 28030 17950 28082
rect 18002 28030 18004 28082
rect 17948 28018 18004 28030
rect 18396 28084 18452 28094
rect 17836 27860 17892 27870
rect 17836 27766 17892 27804
rect 17388 27186 17668 27188
rect 17388 27134 17390 27186
rect 17442 27134 17668 27186
rect 17388 27132 17668 27134
rect 17388 27122 17444 27132
rect 18396 26908 18452 28028
rect 18844 28082 18900 28812
rect 18956 28644 19012 28654
rect 19292 28644 19348 28654
rect 18956 28642 19348 28644
rect 18956 28590 18958 28642
rect 19010 28590 19294 28642
rect 19346 28590 19348 28642
rect 18956 28588 19348 28590
rect 18956 28578 19012 28588
rect 18844 28030 18846 28082
rect 18898 28030 18900 28082
rect 18844 28018 18900 28030
rect 19292 27860 19348 28588
rect 19292 27794 19348 27804
rect 19628 27858 19684 28812
rect 19740 28754 19796 29596
rect 21084 29652 21140 37324
rect 21196 33906 21252 33918
rect 21196 33854 21198 33906
rect 21250 33854 21252 33906
rect 21196 33684 21252 33854
rect 21196 33618 21252 33628
rect 21308 33572 21364 33582
rect 21308 32564 21364 33516
rect 21308 32470 21364 32508
rect 21420 31668 21476 38612
rect 21532 37490 21588 40348
rect 21756 39732 21812 39742
rect 21756 39618 21812 39676
rect 21756 39566 21758 39618
rect 21810 39566 21812 39618
rect 21756 39554 21812 39566
rect 21532 37438 21534 37490
rect 21586 37438 21588 37490
rect 21532 37380 21588 37438
rect 21868 37492 21924 41132
rect 22092 41188 22148 41198
rect 22092 41074 22148 41132
rect 22092 41022 22094 41074
rect 22146 41022 22148 41074
rect 21980 40628 22036 40638
rect 21980 38948 22036 40572
rect 22092 39396 22148 41022
rect 22204 40628 22260 42700
rect 22316 42662 22372 42700
rect 22540 42642 22596 42654
rect 22540 42590 22542 42642
rect 22594 42590 22596 42642
rect 22540 41972 22596 42590
rect 22540 41906 22596 41916
rect 22652 41300 22708 41310
rect 22652 41206 22708 41244
rect 22204 40534 22260 40572
rect 22652 40180 22708 40190
rect 22316 40178 22708 40180
rect 22316 40126 22654 40178
rect 22706 40126 22708 40178
rect 22316 40124 22708 40126
rect 22316 39618 22372 40124
rect 22652 40114 22708 40124
rect 22316 39566 22318 39618
rect 22370 39566 22372 39618
rect 22316 39554 22372 39566
rect 22092 39340 22372 39396
rect 21980 38892 22148 38948
rect 21980 38722 22036 38734
rect 21980 38670 21982 38722
rect 22034 38670 22036 38722
rect 21980 38052 22036 38670
rect 22092 38668 22148 38892
rect 22316 38836 22372 39340
rect 22764 38946 22820 43036
rect 23324 42868 23380 42878
rect 22988 40962 23044 40974
rect 22988 40910 22990 40962
rect 23042 40910 23044 40962
rect 22988 40402 23044 40910
rect 23100 40628 23156 40638
rect 23156 40572 23268 40628
rect 23100 40562 23156 40572
rect 23212 40514 23268 40572
rect 23212 40462 23214 40514
rect 23266 40462 23268 40514
rect 23212 40450 23268 40462
rect 22988 40350 22990 40402
rect 23042 40350 23044 40402
rect 22988 40338 23044 40350
rect 22764 38894 22766 38946
rect 22818 38894 22820 38946
rect 22764 38882 22820 38894
rect 22316 38834 22708 38836
rect 22316 38782 22318 38834
rect 22370 38782 22708 38834
rect 22316 38780 22708 38782
rect 22316 38770 22372 38780
rect 22652 38724 22708 38780
rect 23212 38724 23268 38734
rect 22652 38722 23268 38724
rect 22652 38670 23214 38722
rect 23266 38670 23268 38722
rect 22652 38668 23268 38670
rect 22092 38612 22260 38668
rect 23212 38658 23268 38668
rect 23324 38668 23380 42812
rect 23548 39844 23604 44268
rect 23660 44100 23716 44110
rect 23660 42644 23716 44044
rect 23660 42194 23716 42588
rect 23660 42142 23662 42194
rect 23714 42142 23716 42194
rect 23660 40740 23716 42142
rect 23660 40674 23716 40684
rect 23660 40514 23716 40526
rect 23660 40462 23662 40514
rect 23714 40462 23716 40514
rect 23660 40292 23716 40462
rect 23660 40226 23716 40236
rect 23548 39778 23604 39788
rect 23548 38834 23604 38846
rect 23548 38782 23550 38834
rect 23602 38782 23604 38834
rect 23324 38612 23492 38668
rect 22092 38052 22148 38062
rect 21980 37996 22092 38052
rect 21868 37426 21924 37436
rect 22092 37490 22148 37996
rect 22204 37716 22260 38612
rect 22204 37650 22260 37660
rect 22092 37438 22094 37490
rect 22146 37438 22148 37490
rect 22092 37426 22148 37438
rect 21532 37314 21588 37324
rect 22428 37380 22484 37390
rect 22428 37286 22484 37324
rect 22876 37154 22932 37166
rect 22876 37102 22878 37154
rect 22930 37102 22932 37154
rect 22876 36596 22932 37102
rect 23324 36596 23380 36606
rect 22876 36594 23380 36596
rect 22876 36542 23326 36594
rect 23378 36542 23380 36594
rect 22876 36540 23380 36542
rect 21532 36482 21588 36494
rect 21532 36430 21534 36482
rect 21586 36430 21588 36482
rect 21532 35700 21588 36430
rect 23100 36260 23156 36270
rect 23100 36148 23156 36204
rect 22316 36092 23156 36148
rect 22316 35922 22372 36092
rect 22316 35870 22318 35922
rect 22370 35870 22372 35922
rect 22316 35858 22372 35870
rect 22876 35924 22932 35934
rect 23100 35924 23156 36092
rect 23212 35924 23268 35934
rect 23100 35922 23268 35924
rect 23100 35870 23214 35922
rect 23266 35870 23268 35922
rect 23100 35868 23268 35870
rect 22876 35830 22932 35868
rect 21532 31892 21588 35644
rect 23100 34916 23156 34926
rect 23100 34822 23156 34860
rect 21532 31826 21588 31836
rect 21644 34804 21700 34814
rect 21420 31602 21476 31612
rect 21420 30212 21476 30222
rect 21420 30118 21476 30156
rect 21308 29652 21364 29662
rect 21084 29650 21364 29652
rect 21084 29598 21310 29650
rect 21362 29598 21364 29650
rect 21084 29596 21364 29598
rect 19740 28702 19742 28754
rect 19794 28702 19796 28754
rect 19740 28690 19796 28702
rect 19852 29540 19908 29550
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19628 27794 19684 27806
rect 19292 27636 19348 27646
rect 19292 27634 19572 27636
rect 19292 27582 19294 27634
rect 19346 27582 19572 27634
rect 19292 27580 19572 27582
rect 19292 27570 19348 27580
rect 19516 27300 19572 27580
rect 19628 27300 19684 27310
rect 19516 27298 19684 27300
rect 19516 27246 19630 27298
rect 19682 27246 19684 27298
rect 19516 27244 19684 27246
rect 19628 27234 19684 27244
rect 18844 27076 18900 27086
rect 19852 27076 19908 29484
rect 21084 29428 21140 29596
rect 21308 29586 21364 29596
rect 21084 29362 21140 29372
rect 21644 28868 21700 34748
rect 23212 34804 23268 35868
rect 23324 35588 23380 36540
rect 23436 36372 23492 38612
rect 23436 36306 23492 36316
rect 23548 35924 23604 38782
rect 23548 35858 23604 35868
rect 23660 37380 23716 37390
rect 23772 37380 23828 46510
rect 24780 46452 24836 47406
rect 25340 47236 25396 47246
rect 25340 46898 25396 47180
rect 25340 46846 25342 46898
rect 25394 46846 25396 46898
rect 25340 46834 25396 46846
rect 23884 46396 24836 46452
rect 23884 46116 23940 46396
rect 24008 46284 25208 46294
rect 24064 46282 24112 46284
rect 24168 46282 24216 46284
rect 24076 46230 24112 46282
rect 24200 46230 24216 46282
rect 24064 46228 24112 46230
rect 24168 46228 24216 46230
rect 24272 46282 24320 46284
rect 24376 46282 24424 46284
rect 24480 46282 24528 46284
rect 24376 46230 24396 46282
rect 24480 46230 24520 46282
rect 24272 46228 24320 46230
rect 24376 46228 24424 46230
rect 24480 46228 24528 46230
rect 24584 46228 24632 46284
rect 24688 46282 24736 46284
rect 24792 46282 24840 46284
rect 24896 46282 24944 46284
rect 24696 46230 24736 46282
rect 24820 46230 24840 46282
rect 24688 46228 24736 46230
rect 24792 46228 24840 46230
rect 24896 46228 24944 46230
rect 25000 46282 25048 46284
rect 25104 46282 25152 46284
rect 25000 46230 25016 46282
rect 25104 46230 25140 46282
rect 25000 46228 25048 46230
rect 25104 46228 25152 46230
rect 24008 46218 25208 46228
rect 25564 46116 25620 50372
rect 26236 49252 26292 51548
rect 26908 51938 26964 51950
rect 26908 51886 26910 51938
rect 26962 51886 26964 51938
rect 26908 51492 26964 51886
rect 27020 51604 27076 54350
rect 27132 52724 27188 56588
rect 27692 56196 27748 58158
rect 27804 57650 27860 58828
rect 28140 58436 28196 58446
rect 28140 58342 28196 58380
rect 28476 58436 28532 59726
rect 28476 58370 28532 58380
rect 28140 57876 28196 57886
rect 28140 57782 28196 57820
rect 28588 57876 28644 60174
rect 28588 57810 28644 57820
rect 28700 60674 28756 60686
rect 28700 60622 28702 60674
rect 28754 60622 28756 60674
rect 28700 60452 28756 60622
rect 27804 57598 27806 57650
rect 27858 57598 27860 57650
rect 27804 57586 27860 57598
rect 28588 56868 28644 56878
rect 28700 56868 28756 60396
rect 28924 59556 28980 66780
rect 29036 66274 29092 67004
rect 29260 67954 29876 67956
rect 29260 67902 29822 67954
rect 29874 67902 29876 67954
rect 29260 67900 29876 67902
rect 29260 67058 29316 67900
rect 29820 67890 29876 67900
rect 30044 67900 30436 67956
rect 30716 68402 30772 68414
rect 30716 68350 30718 68402
rect 30770 68350 30772 68402
rect 29372 67732 29428 67742
rect 29372 67638 29428 67676
rect 29484 67620 29540 67630
rect 29932 67620 29988 67630
rect 30044 67620 30100 67900
rect 30156 67732 30212 67742
rect 30492 67732 30548 67742
rect 30156 67730 30548 67732
rect 30156 67678 30158 67730
rect 30210 67678 30494 67730
rect 30546 67678 30548 67730
rect 30156 67676 30548 67678
rect 30156 67666 30212 67676
rect 30492 67666 30548 67676
rect 30716 67732 30772 68350
rect 31052 68068 31108 68574
rect 31276 68180 31332 68796
rect 31388 68628 31444 68638
rect 31388 68626 31892 68628
rect 31388 68574 31390 68626
rect 31442 68574 31892 68626
rect 31388 68572 31892 68574
rect 31388 68562 31444 68572
rect 31276 68124 31556 68180
rect 31052 68012 31332 68068
rect 30716 67666 30772 67676
rect 31164 67842 31220 67854
rect 31164 67790 31166 67842
rect 31218 67790 31220 67842
rect 29484 67618 29652 67620
rect 29484 67566 29486 67618
rect 29538 67566 29652 67618
rect 29484 67564 29652 67566
rect 29484 67554 29540 67564
rect 29260 67006 29262 67058
rect 29314 67006 29316 67058
rect 29260 66994 29316 67006
rect 29036 66222 29038 66274
rect 29090 66222 29092 66274
rect 29036 66210 29092 66222
rect 29372 66276 29428 66286
rect 29372 65716 29428 66220
rect 29596 66274 29652 67564
rect 29932 67618 30100 67620
rect 29932 67566 29934 67618
rect 29986 67566 30100 67618
rect 29932 67564 30100 67566
rect 29932 67554 29988 67564
rect 29596 66222 29598 66274
rect 29650 66222 29652 66274
rect 29596 66210 29652 66222
rect 29372 65492 29428 65660
rect 29260 65490 29428 65492
rect 29260 65438 29374 65490
rect 29426 65438 29428 65490
rect 29260 65436 29428 65438
rect 29036 65268 29092 65278
rect 29036 65266 29204 65268
rect 29036 65214 29038 65266
rect 29090 65214 29204 65266
rect 29036 65212 29204 65214
rect 29036 65202 29092 65212
rect 29148 64034 29204 65212
rect 29260 64818 29316 65436
rect 29372 65426 29428 65436
rect 29260 64766 29262 64818
rect 29314 64766 29316 64818
rect 29260 64754 29316 64766
rect 29148 63982 29150 64034
rect 29202 63982 29204 64034
rect 29148 63970 29204 63982
rect 29820 64482 29876 64494
rect 29820 64430 29822 64482
rect 29874 64430 29876 64482
rect 29260 63924 29316 63934
rect 29260 63830 29316 63868
rect 29260 62914 29316 62926
rect 29260 62862 29262 62914
rect 29314 62862 29316 62914
rect 29148 62356 29204 62366
rect 29148 62188 29204 62300
rect 29260 62188 29316 62862
rect 29596 62580 29652 62590
rect 29596 62486 29652 62524
rect 29820 62356 29876 64430
rect 29932 63812 29988 63822
rect 29932 63718 29988 63756
rect 30044 62916 30100 67564
rect 31164 66836 31220 67790
rect 31276 67844 31332 68012
rect 31388 67844 31444 67854
rect 31276 67842 31444 67844
rect 31276 67790 31390 67842
rect 31442 67790 31444 67842
rect 31276 67788 31444 67790
rect 31164 66770 31220 66780
rect 31276 67172 31332 67182
rect 30828 65492 30884 65502
rect 30828 65398 30884 65436
rect 31276 65490 31332 67116
rect 31388 66948 31444 67788
rect 31388 66882 31444 66892
rect 31276 65438 31278 65490
rect 31330 65438 31332 65490
rect 31276 65426 31332 65438
rect 31500 65490 31556 68124
rect 31836 68066 31892 68572
rect 31836 68014 31838 68066
rect 31890 68014 31892 68066
rect 31836 68002 31892 68014
rect 31948 67844 32004 69916
rect 33180 69188 33236 69198
rect 33292 69188 33348 70252
rect 33404 70306 33460 70476
rect 33404 70254 33406 70306
rect 33458 70254 33460 70306
rect 33404 69860 33460 70254
rect 33404 69794 33460 69804
rect 33516 69636 33572 70926
rect 33852 70980 33908 70990
rect 33516 69570 33572 69580
rect 33740 70420 33796 70430
rect 33740 69634 33796 70364
rect 33740 69582 33742 69634
rect 33794 69582 33796 69634
rect 33740 69570 33796 69582
rect 33852 70194 33908 70924
rect 35084 70756 35140 71598
rect 35756 70756 35812 70766
rect 35084 70700 35364 70756
rect 34008 70588 35208 70598
rect 34064 70586 34112 70588
rect 34168 70586 34216 70588
rect 34076 70534 34112 70586
rect 34200 70534 34216 70586
rect 34064 70532 34112 70534
rect 34168 70532 34216 70534
rect 34272 70586 34320 70588
rect 34376 70586 34424 70588
rect 34480 70586 34528 70588
rect 34376 70534 34396 70586
rect 34480 70534 34520 70586
rect 34272 70532 34320 70534
rect 34376 70532 34424 70534
rect 34480 70532 34528 70534
rect 34584 70532 34632 70588
rect 34688 70586 34736 70588
rect 34792 70586 34840 70588
rect 34896 70586 34944 70588
rect 34696 70534 34736 70586
rect 34820 70534 34840 70586
rect 34688 70532 34736 70534
rect 34792 70532 34840 70534
rect 34896 70532 34944 70534
rect 35000 70586 35048 70588
rect 35104 70586 35152 70588
rect 35000 70534 35016 70586
rect 35104 70534 35140 70586
rect 35000 70532 35048 70534
rect 35104 70532 35152 70534
rect 34008 70522 35208 70532
rect 35308 70532 35364 70700
rect 35756 70662 35812 70700
rect 35308 70466 35364 70476
rect 35644 70532 35700 70542
rect 33852 70142 33854 70194
rect 33906 70142 33908 70194
rect 33180 69186 33348 69188
rect 33180 69134 33182 69186
rect 33234 69134 33348 69186
rect 33180 69132 33348 69134
rect 33180 69122 33236 69132
rect 32172 67844 32228 67854
rect 31948 67842 32228 67844
rect 31948 67790 32174 67842
rect 32226 67790 32228 67842
rect 31948 67788 32228 67790
rect 32060 67620 32116 67630
rect 31948 67564 32060 67620
rect 31836 67284 31892 67294
rect 31948 67284 32004 67564
rect 32060 67554 32116 67564
rect 31836 67282 32004 67284
rect 31836 67230 31838 67282
rect 31890 67230 32004 67282
rect 31836 67228 32004 67230
rect 31500 65438 31502 65490
rect 31554 65438 31556 65490
rect 30268 64596 30324 64606
rect 30268 64146 30324 64540
rect 30268 64094 30270 64146
rect 30322 64094 30324 64146
rect 30268 64082 30324 64094
rect 31276 63810 31332 63822
rect 31276 63758 31278 63810
rect 31330 63758 31332 63810
rect 30492 63140 30548 63150
rect 30156 62916 30212 62926
rect 30044 62914 30212 62916
rect 30044 62862 30158 62914
rect 30210 62862 30212 62914
rect 30044 62860 30212 62862
rect 30044 62356 30100 62366
rect 29820 62300 30044 62356
rect 30044 62262 30100 62300
rect 29148 62132 29428 62188
rect 29372 61570 29428 62132
rect 29932 61572 29988 61582
rect 29372 61518 29374 61570
rect 29426 61518 29428 61570
rect 29372 60452 29428 61518
rect 29820 61570 29988 61572
rect 29820 61518 29934 61570
rect 29986 61518 29988 61570
rect 29820 61516 29988 61518
rect 29596 61348 29652 61358
rect 29652 61292 29764 61348
rect 29596 61282 29652 61292
rect 29372 60386 29428 60396
rect 29596 60564 29652 60574
rect 29596 59890 29652 60508
rect 29596 59838 29598 59890
rect 29650 59838 29652 59890
rect 29596 59826 29652 59838
rect 29708 59892 29764 61292
rect 29820 60116 29876 61516
rect 29932 61506 29988 61516
rect 30156 61124 30212 62860
rect 30492 62244 30548 63084
rect 31052 63140 31108 63150
rect 31052 63046 31108 63084
rect 31276 63138 31332 63758
rect 31276 63086 31278 63138
rect 31330 63086 31332 63138
rect 30716 63026 30772 63038
rect 30716 62974 30718 63026
rect 30770 62974 30772 63026
rect 30716 62804 30772 62974
rect 30716 62738 30772 62748
rect 31052 62916 31108 62926
rect 30492 62178 30548 62188
rect 30604 62524 30996 62580
rect 30604 61684 30660 62524
rect 30940 62466 30996 62524
rect 30940 62414 30942 62466
rect 30994 62414 30996 62466
rect 30940 62402 30996 62414
rect 31052 62466 31108 62860
rect 31052 62414 31054 62466
rect 31106 62414 31108 62466
rect 31052 62402 31108 62414
rect 31276 62804 31332 63086
rect 31500 63364 31556 65438
rect 31612 66836 31668 66846
rect 31612 65490 31668 66780
rect 31836 66276 31892 67228
rect 32172 67172 32228 67788
rect 32396 67730 32452 67742
rect 32396 67678 32398 67730
rect 32450 67678 32452 67730
rect 32396 67172 32452 67678
rect 32956 67620 33012 67630
rect 32956 67526 33012 67564
rect 33180 67172 33236 67182
rect 32396 67170 33236 67172
rect 32396 67118 33182 67170
rect 33234 67118 33236 67170
rect 32396 67116 33236 67118
rect 32172 67106 32228 67116
rect 32396 66836 32452 66846
rect 32396 66742 32452 66780
rect 31836 66210 31892 66220
rect 31948 66164 32004 66174
rect 31948 66070 32004 66108
rect 31612 65438 31614 65490
rect 31666 65438 31668 65490
rect 31612 65426 31668 65438
rect 31836 66052 31892 66062
rect 31836 65490 31892 65996
rect 32732 66052 32788 66062
rect 33068 66052 33124 67116
rect 33180 67106 33236 67116
rect 33292 67172 33348 67182
rect 33292 67078 33348 67116
rect 33852 67060 33908 70142
rect 34412 70420 34468 70430
rect 34412 70194 34468 70364
rect 34412 70142 34414 70194
rect 34466 70142 34468 70194
rect 34412 70130 34468 70142
rect 35196 70084 35252 70094
rect 34972 69860 35028 69870
rect 34636 69636 34692 69646
rect 34636 69542 34692 69580
rect 34972 69634 35028 69804
rect 34972 69582 34974 69634
rect 35026 69582 35028 69634
rect 34972 69570 35028 69582
rect 34748 69410 34804 69422
rect 34748 69358 34750 69410
rect 34802 69358 34804 69410
rect 33964 69188 34020 69198
rect 34300 69188 34356 69198
rect 34748 69188 34804 69358
rect 35196 69410 35252 70028
rect 35532 69860 35588 69870
rect 35532 69634 35588 69804
rect 35532 69582 35534 69634
rect 35586 69582 35588 69634
rect 35532 69570 35588 69582
rect 35196 69358 35198 69410
rect 35250 69358 35252 69410
rect 35196 69346 35252 69358
rect 34020 69186 34804 69188
rect 34020 69134 34302 69186
rect 34354 69134 34804 69186
rect 34020 69132 34804 69134
rect 35532 69300 35588 69310
rect 33964 69122 34020 69132
rect 34300 69122 34356 69132
rect 34008 69020 35208 69030
rect 34064 69018 34112 69020
rect 34168 69018 34216 69020
rect 34076 68966 34112 69018
rect 34200 68966 34216 69018
rect 34064 68964 34112 68966
rect 34168 68964 34216 68966
rect 34272 69018 34320 69020
rect 34376 69018 34424 69020
rect 34480 69018 34528 69020
rect 34376 68966 34396 69018
rect 34480 68966 34520 69018
rect 34272 68964 34320 68966
rect 34376 68964 34424 68966
rect 34480 68964 34528 68966
rect 34584 68964 34632 69020
rect 34688 69018 34736 69020
rect 34792 69018 34840 69020
rect 34896 69018 34944 69020
rect 34696 68966 34736 69018
rect 34820 68966 34840 69018
rect 34688 68964 34736 68966
rect 34792 68964 34840 68966
rect 34896 68964 34944 68966
rect 35000 69018 35048 69020
rect 35104 69018 35152 69020
rect 35000 68966 35016 69018
rect 35104 68966 35140 69018
rect 35000 68964 35048 68966
rect 35104 68964 35152 68966
rect 34008 68954 35208 68964
rect 34972 68852 35028 68862
rect 34972 67956 35028 68796
rect 35532 68626 35588 69244
rect 35644 68850 35700 70476
rect 35868 69636 35924 71710
rect 36092 71762 36148 71774
rect 36092 71710 36094 71762
rect 36146 71710 36148 71762
rect 35756 69580 35924 69636
rect 35980 71650 36036 71662
rect 35980 71598 35982 71650
rect 36034 71598 36036 71650
rect 35756 69300 35812 69580
rect 35980 69524 36036 71598
rect 35756 69234 35812 69244
rect 35868 69468 36036 69524
rect 36092 69972 36148 71710
rect 35644 68798 35646 68850
rect 35698 68798 35700 68850
rect 35644 68786 35700 68798
rect 35868 68852 35924 69468
rect 36092 69410 36148 69916
rect 36092 69358 36094 69410
rect 36146 69358 36148 69410
rect 35980 69300 36036 69310
rect 35980 69206 36036 69244
rect 35980 68852 36036 68862
rect 35868 68850 36036 68852
rect 35868 68798 35982 68850
rect 36034 68798 36036 68850
rect 35868 68796 36036 68798
rect 35980 68786 36036 68796
rect 35532 68574 35534 68626
rect 35586 68574 35588 68626
rect 35420 67956 35476 67966
rect 34972 67954 35476 67956
rect 34972 67902 34974 67954
rect 35026 67902 35422 67954
rect 35474 67902 35476 67954
rect 34972 67900 35476 67902
rect 34972 67890 35028 67900
rect 35308 67730 35364 67742
rect 35308 67678 35310 67730
rect 35362 67678 35364 67730
rect 34008 67452 35208 67462
rect 34064 67450 34112 67452
rect 34168 67450 34216 67452
rect 34076 67398 34112 67450
rect 34200 67398 34216 67450
rect 34064 67396 34112 67398
rect 34168 67396 34216 67398
rect 34272 67450 34320 67452
rect 34376 67450 34424 67452
rect 34480 67450 34528 67452
rect 34376 67398 34396 67450
rect 34480 67398 34520 67450
rect 34272 67396 34320 67398
rect 34376 67396 34424 67398
rect 34480 67396 34528 67398
rect 34584 67396 34632 67452
rect 34688 67450 34736 67452
rect 34792 67450 34840 67452
rect 34896 67450 34944 67452
rect 34696 67398 34736 67450
rect 34820 67398 34840 67450
rect 34688 67396 34736 67398
rect 34792 67396 34840 67398
rect 34896 67396 34944 67398
rect 35000 67450 35048 67452
rect 35104 67450 35152 67452
rect 35000 67398 35016 67450
rect 35104 67398 35140 67450
rect 35000 67396 35048 67398
rect 35104 67396 35152 67398
rect 34008 67386 35208 67396
rect 34524 67284 34580 67294
rect 33964 67060 34020 67070
rect 33852 67058 34020 67060
rect 33852 67006 33966 67058
rect 34018 67006 34020 67058
rect 33852 67004 34020 67006
rect 33180 66948 33236 66958
rect 33180 66834 33236 66892
rect 33180 66782 33182 66834
rect 33234 66782 33236 66834
rect 33180 66770 33236 66782
rect 33740 66946 33796 66958
rect 33740 66894 33742 66946
rect 33794 66894 33796 66946
rect 32788 65996 33124 66052
rect 33740 66164 33796 66894
rect 32732 65958 32788 65996
rect 33740 65714 33796 66108
rect 33740 65662 33742 65714
rect 33794 65662 33796 65714
rect 33740 65650 33796 65662
rect 31836 65438 31838 65490
rect 31890 65438 31892 65490
rect 31836 65426 31892 65438
rect 33852 65492 33908 67004
rect 33964 66994 34020 67004
rect 34524 67058 34580 67228
rect 35308 67284 35364 67678
rect 35308 67218 35364 67228
rect 35420 67060 35476 67900
rect 35532 67844 35588 68574
rect 35756 68628 35812 68638
rect 36092 68628 36148 69358
rect 36204 71764 36260 71932
rect 36316 71764 36372 71774
rect 36204 71762 36372 71764
rect 36204 71710 36318 71762
rect 36370 71710 36372 71762
rect 36204 71708 36372 71710
rect 36204 68852 36260 71708
rect 36316 71698 36372 71708
rect 36540 70756 36596 70766
rect 36316 70754 36596 70756
rect 36316 70702 36542 70754
rect 36594 70702 36596 70754
rect 36316 70700 36596 70702
rect 36316 70196 36372 70700
rect 36540 70690 36596 70700
rect 36652 70308 36708 70318
rect 36652 70214 36708 70252
rect 36316 69410 36372 70140
rect 37548 70194 37604 70206
rect 37548 70142 37550 70194
rect 37602 70142 37604 70194
rect 37436 69972 37492 69982
rect 37436 69878 37492 69916
rect 36316 69358 36318 69410
rect 36370 69358 36372 69410
rect 36316 69346 36372 69358
rect 37548 69300 37604 70142
rect 37884 70194 37940 70206
rect 37884 70142 37886 70194
rect 37938 70142 37940 70194
rect 37772 70084 37828 70094
rect 37772 69990 37828 70028
rect 37884 69972 37940 70142
rect 38108 70196 38164 70206
rect 38108 70102 38164 70140
rect 37884 69906 37940 69916
rect 37548 69234 37604 69244
rect 36204 68786 36260 68796
rect 35756 68626 36148 68628
rect 35756 68574 35758 68626
rect 35810 68574 36148 68626
rect 35756 68572 36148 68574
rect 35756 68562 35812 68572
rect 35644 67844 35700 67854
rect 35532 67842 35700 67844
rect 35532 67790 35646 67842
rect 35698 67790 35700 67842
rect 35532 67788 35700 67790
rect 34524 67006 34526 67058
rect 34578 67006 34580 67058
rect 34524 66994 34580 67006
rect 35196 67004 35476 67060
rect 35196 66052 35252 67004
rect 35644 66388 35700 67788
rect 35868 67844 35924 67854
rect 35868 67750 35924 67788
rect 37100 67844 37156 67854
rect 37100 67750 37156 67788
rect 37324 67844 37380 67854
rect 37324 67842 37716 67844
rect 37324 67790 37326 67842
rect 37378 67790 37716 67842
rect 37324 67788 37716 67790
rect 37324 67778 37380 67788
rect 36988 67730 37044 67742
rect 36988 67678 36990 67730
rect 37042 67678 37044 67730
rect 35644 66322 35700 66332
rect 36876 67170 36932 67182
rect 36876 67118 36878 67170
rect 36930 67118 36932 67170
rect 36092 66162 36148 66174
rect 36092 66110 36094 66162
rect 36146 66110 36148 66162
rect 35196 65996 35364 66052
rect 34008 65884 35208 65894
rect 34064 65882 34112 65884
rect 34168 65882 34216 65884
rect 34076 65830 34112 65882
rect 34200 65830 34216 65882
rect 34064 65828 34112 65830
rect 34168 65828 34216 65830
rect 34272 65882 34320 65884
rect 34376 65882 34424 65884
rect 34480 65882 34528 65884
rect 34376 65830 34396 65882
rect 34480 65830 34520 65882
rect 34272 65828 34320 65830
rect 34376 65828 34424 65830
rect 34480 65828 34528 65830
rect 34584 65828 34632 65884
rect 34688 65882 34736 65884
rect 34792 65882 34840 65884
rect 34896 65882 34944 65884
rect 34696 65830 34736 65882
rect 34820 65830 34840 65882
rect 34688 65828 34736 65830
rect 34792 65828 34840 65830
rect 34896 65828 34944 65830
rect 35000 65882 35048 65884
rect 35104 65882 35152 65884
rect 35000 65830 35016 65882
rect 35104 65830 35140 65882
rect 35000 65828 35048 65830
rect 35104 65828 35152 65830
rect 34008 65818 35208 65828
rect 35308 65716 35364 65996
rect 35196 65660 35364 65716
rect 33964 65492 34020 65502
rect 33852 65490 34020 65492
rect 33852 65438 33966 65490
rect 34018 65438 34020 65490
rect 33852 65436 34020 65438
rect 33964 65426 34020 65436
rect 34636 65490 34692 65502
rect 34636 65438 34638 65490
rect 34690 65438 34692 65490
rect 34636 64932 34692 65438
rect 34636 64866 34692 64876
rect 35196 64820 35252 65660
rect 36092 65044 36148 66110
rect 36876 66164 36932 67118
rect 36988 66612 37044 67678
rect 37660 67284 37716 67788
rect 37548 67282 37716 67284
rect 37548 67230 37662 67282
rect 37714 67230 37716 67282
rect 37548 67228 37716 67230
rect 36988 66556 37380 66612
rect 36988 66388 37044 66398
rect 36988 66294 37044 66332
rect 36092 64978 36148 64988
rect 36204 66050 36260 66062
rect 36204 65998 36206 66050
rect 36258 65998 36260 66050
rect 35532 64932 35588 64942
rect 35532 64838 35588 64876
rect 35868 64932 35924 64942
rect 35868 64838 35924 64876
rect 35196 64818 35476 64820
rect 35196 64766 35198 64818
rect 35250 64766 35476 64818
rect 35196 64764 35476 64766
rect 35196 64754 35252 64764
rect 35420 64708 35476 64764
rect 35644 64708 35700 64718
rect 35420 64706 35700 64708
rect 35420 64654 35646 64706
rect 35698 64654 35700 64706
rect 35420 64652 35700 64654
rect 34008 64316 35208 64326
rect 34064 64314 34112 64316
rect 34168 64314 34216 64316
rect 34076 64262 34112 64314
rect 34200 64262 34216 64314
rect 34064 64260 34112 64262
rect 34168 64260 34216 64262
rect 34272 64314 34320 64316
rect 34376 64314 34424 64316
rect 34480 64314 34528 64316
rect 34376 64262 34396 64314
rect 34480 64262 34520 64314
rect 34272 64260 34320 64262
rect 34376 64260 34424 64262
rect 34480 64260 34528 64262
rect 34584 64260 34632 64316
rect 34688 64314 34736 64316
rect 34792 64314 34840 64316
rect 34896 64314 34944 64316
rect 34696 64262 34736 64314
rect 34820 64262 34840 64314
rect 34688 64260 34736 64262
rect 34792 64260 34840 64262
rect 34896 64260 34944 64262
rect 35000 64314 35048 64316
rect 35104 64314 35152 64316
rect 35000 64262 35016 64314
rect 35104 64262 35140 64314
rect 35000 64260 35048 64262
rect 35104 64260 35152 64262
rect 34008 64250 35208 64260
rect 31836 63922 31892 63934
rect 31836 63870 31838 63922
rect 31890 63870 31892 63922
rect 31836 63812 31892 63870
rect 31724 63364 31780 63374
rect 31500 63362 31780 63364
rect 31500 63310 31726 63362
rect 31778 63310 31780 63362
rect 31500 63308 31780 63310
rect 31500 62916 31556 63308
rect 31724 63298 31780 63308
rect 31500 62850 31556 62860
rect 30156 61058 30212 61068
rect 30380 61628 30660 61684
rect 30716 62354 30772 62366
rect 30716 62302 30718 62354
rect 30770 62302 30772 62354
rect 29932 61012 29988 61022
rect 29932 60898 29988 60956
rect 29932 60846 29934 60898
rect 29986 60846 29988 60898
rect 29932 60834 29988 60846
rect 30044 60900 30100 60910
rect 30044 60898 30212 60900
rect 30044 60846 30046 60898
rect 30098 60846 30212 60898
rect 30044 60844 30212 60846
rect 30044 60834 30100 60844
rect 30044 60562 30100 60574
rect 30044 60510 30046 60562
rect 30098 60510 30100 60562
rect 29932 60116 29988 60126
rect 29820 60114 29988 60116
rect 29820 60062 29934 60114
rect 29986 60062 29988 60114
rect 29820 60060 29988 60062
rect 29932 60050 29988 60060
rect 30044 60116 30100 60510
rect 30044 60050 30100 60060
rect 29820 59892 29876 59902
rect 29708 59890 29876 59892
rect 29708 59838 29822 59890
rect 29874 59838 29876 59890
rect 29708 59836 29876 59838
rect 29820 59826 29876 59836
rect 30044 59892 30100 59902
rect 30044 59798 30100 59836
rect 28924 59500 29204 59556
rect 28812 59444 28868 59454
rect 28868 59388 28980 59444
rect 28812 59378 28868 59388
rect 28924 59330 28980 59388
rect 28924 59278 28926 59330
rect 28978 59278 28980 59330
rect 28924 59266 28980 59278
rect 29148 59220 29204 59500
rect 29932 59444 29988 59454
rect 29988 59388 30100 59444
rect 29932 59378 29988 59388
rect 29932 59220 29988 59230
rect 29148 59218 29988 59220
rect 29148 59166 29934 59218
rect 29986 59166 29988 59218
rect 29148 59164 29988 59166
rect 29708 58994 29764 59006
rect 29708 58942 29710 58994
rect 29762 58942 29764 58994
rect 29708 58884 29764 58942
rect 29708 58818 29764 58828
rect 29596 58212 29652 58222
rect 29820 58212 29876 59164
rect 29932 59154 29988 59164
rect 29932 58436 29988 58446
rect 29932 58342 29988 58380
rect 29596 58210 29876 58212
rect 29596 58158 29598 58210
rect 29650 58158 29876 58210
rect 29596 58156 29876 58158
rect 29036 56868 29092 56878
rect 28588 56866 29092 56868
rect 28588 56814 28590 56866
rect 28642 56814 29038 56866
rect 29090 56814 29092 56866
rect 28588 56812 29092 56814
rect 28588 56802 28644 56812
rect 29036 56802 29092 56812
rect 27692 56130 27748 56140
rect 28140 56642 28196 56654
rect 28140 56590 28142 56642
rect 28194 56590 28196 56642
rect 28140 56196 28196 56590
rect 28140 56130 28196 56140
rect 27356 54516 27412 54526
rect 27692 54516 27748 54526
rect 27356 53844 27412 54460
rect 27356 53778 27412 53788
rect 27468 54514 27748 54516
rect 27468 54462 27694 54514
rect 27746 54462 27748 54514
rect 27468 54460 27748 54462
rect 27356 53508 27412 53518
rect 27244 53506 27412 53508
rect 27244 53454 27358 53506
rect 27410 53454 27412 53506
rect 27244 53452 27412 53454
rect 27244 52946 27300 53452
rect 27356 53442 27412 53452
rect 27244 52894 27246 52946
rect 27298 52894 27300 52946
rect 27244 52882 27300 52894
rect 27132 52668 27300 52724
rect 27020 51602 27188 51604
rect 27020 51550 27022 51602
rect 27074 51550 27188 51602
rect 27020 51548 27188 51550
rect 27020 51538 27076 51548
rect 26908 51426 26964 51436
rect 27132 50372 27188 51548
rect 27244 50428 27300 52668
rect 27468 51602 27524 54460
rect 27692 54450 27748 54460
rect 27692 53956 27748 53966
rect 27692 53862 27748 53900
rect 28028 53618 28084 53630
rect 28028 53566 28030 53618
rect 28082 53566 28084 53618
rect 27580 52052 27636 52062
rect 27580 51958 27636 51996
rect 27468 51550 27470 51602
rect 27522 51550 27524 51602
rect 27468 51538 27524 51550
rect 27580 51492 27636 51502
rect 27636 51436 27860 51492
rect 27580 51426 27636 51436
rect 27804 51378 27860 51436
rect 27804 51326 27806 51378
rect 27858 51326 27860 51378
rect 27804 51314 27860 51326
rect 28028 51490 28084 53566
rect 28476 53620 28532 53630
rect 28476 53526 28532 53564
rect 29372 53508 29428 53518
rect 28028 51438 28030 51490
rect 28082 51438 28084 51490
rect 27244 50372 27524 50428
rect 26460 49924 26516 49934
rect 26460 49830 26516 49868
rect 26236 49158 26292 49196
rect 27132 49698 27188 50316
rect 27132 49646 27134 49698
rect 27186 49646 27188 49698
rect 25676 49028 25732 49038
rect 25676 47348 25732 48972
rect 26684 49028 26740 49038
rect 26236 48916 26292 48926
rect 26236 48468 26292 48860
rect 26124 48466 26292 48468
rect 26124 48414 26238 48466
rect 26290 48414 26292 48466
rect 26124 48412 26292 48414
rect 25788 48130 25844 48142
rect 25788 48078 25790 48130
rect 25842 48078 25844 48130
rect 25788 47572 25844 48078
rect 25788 47506 25844 47516
rect 25676 47292 25844 47348
rect 23884 46060 24276 46116
rect 24220 46002 24276 46060
rect 24220 45950 24222 46002
rect 24274 45950 24276 46002
rect 24220 45938 24276 45950
rect 25340 46060 25620 46116
rect 24780 45892 24836 45902
rect 24780 45798 24836 45836
rect 25116 45890 25172 45902
rect 25116 45838 25118 45890
rect 25170 45838 25172 45890
rect 24108 45780 24164 45790
rect 24108 45666 24164 45724
rect 24108 45614 24110 45666
rect 24162 45614 24164 45666
rect 23884 44996 23940 45006
rect 24108 44996 24164 45614
rect 24332 45668 24388 45678
rect 24332 45574 24388 45612
rect 24332 45332 24388 45342
rect 24332 45238 24388 45276
rect 23884 44994 24164 44996
rect 23884 44942 23886 44994
rect 23938 44942 24164 44994
rect 23884 44940 24164 44942
rect 23884 44436 23940 44940
rect 25116 44884 25172 45838
rect 25116 44818 25172 44828
rect 24008 44716 25208 44726
rect 24064 44714 24112 44716
rect 24168 44714 24216 44716
rect 24076 44662 24112 44714
rect 24200 44662 24216 44714
rect 24064 44660 24112 44662
rect 24168 44660 24216 44662
rect 24272 44714 24320 44716
rect 24376 44714 24424 44716
rect 24480 44714 24528 44716
rect 24376 44662 24396 44714
rect 24480 44662 24520 44714
rect 24272 44660 24320 44662
rect 24376 44660 24424 44662
rect 24480 44660 24528 44662
rect 24584 44660 24632 44716
rect 24688 44714 24736 44716
rect 24792 44714 24840 44716
rect 24896 44714 24944 44716
rect 24696 44662 24736 44714
rect 24820 44662 24840 44714
rect 24688 44660 24736 44662
rect 24792 44660 24840 44662
rect 24896 44660 24944 44662
rect 25000 44714 25048 44716
rect 25104 44714 25152 44716
rect 25000 44662 25016 44714
rect 25104 44662 25140 44714
rect 25000 44660 25048 44662
rect 25104 44660 25152 44662
rect 24008 44650 25208 44660
rect 25340 44548 25396 46060
rect 25788 46004 25844 47292
rect 25788 45938 25844 45948
rect 26012 46564 26068 46574
rect 25676 45890 25732 45902
rect 25676 45838 25678 45890
rect 25730 45838 25732 45890
rect 25676 45780 25732 45838
rect 26012 45780 26068 46508
rect 25676 45724 25956 45780
rect 25900 45330 25956 45724
rect 26012 45714 26068 45724
rect 26124 45332 26180 48412
rect 26236 48402 26292 48412
rect 26684 48466 26740 48972
rect 27020 49028 27076 49038
rect 27020 48934 27076 48972
rect 26908 48914 26964 48926
rect 26908 48862 26910 48914
rect 26962 48862 26964 48914
rect 26908 48804 26964 48862
rect 26908 48738 26964 48748
rect 26684 48414 26686 48466
rect 26738 48414 26740 48466
rect 26684 48402 26740 48414
rect 27020 48356 27076 48366
rect 26460 46900 26516 46910
rect 27020 46900 27076 48300
rect 27132 47908 27188 49646
rect 27356 48244 27412 48254
rect 27356 48150 27412 48188
rect 27132 47852 27412 47908
rect 27132 47234 27188 47246
rect 27132 47182 27134 47234
rect 27186 47182 27188 47234
rect 27132 47124 27188 47182
rect 27132 47058 27188 47068
rect 27132 46900 27188 46910
rect 27020 46898 27188 46900
rect 27020 46846 27134 46898
rect 27186 46846 27188 46898
rect 27020 46844 27188 46846
rect 26460 46806 26516 46844
rect 27132 46834 27188 46844
rect 26572 46788 26628 46798
rect 26236 46674 26292 46686
rect 26236 46622 26238 46674
rect 26290 46622 26292 46674
rect 26236 45892 26292 46622
rect 26572 46674 26628 46732
rect 26572 46622 26574 46674
rect 26626 46622 26628 46674
rect 26572 46564 26628 46622
rect 26572 46498 26628 46508
rect 26236 45826 26292 45836
rect 25900 45278 25902 45330
rect 25954 45278 25956 45330
rect 25900 45266 25956 45278
rect 26012 45276 26180 45332
rect 25788 45108 25844 45118
rect 25788 45014 25844 45052
rect 25452 44996 25508 45006
rect 25452 44902 25508 44940
rect 25340 44492 25620 44548
rect 23884 44370 23940 44380
rect 24108 44100 24164 44110
rect 23884 44098 24164 44100
rect 23884 44046 24110 44098
rect 24162 44046 24164 44098
rect 23884 44044 24164 44046
rect 23884 42868 23940 44044
rect 24108 44034 24164 44044
rect 24008 43148 25208 43158
rect 24064 43146 24112 43148
rect 24168 43146 24216 43148
rect 24076 43094 24112 43146
rect 24200 43094 24216 43146
rect 24064 43092 24112 43094
rect 24168 43092 24216 43094
rect 24272 43146 24320 43148
rect 24376 43146 24424 43148
rect 24480 43146 24528 43148
rect 24376 43094 24396 43146
rect 24480 43094 24520 43146
rect 24272 43092 24320 43094
rect 24376 43092 24424 43094
rect 24480 43092 24528 43094
rect 24584 43092 24632 43148
rect 24688 43146 24736 43148
rect 24792 43146 24840 43148
rect 24896 43146 24944 43148
rect 24696 43094 24736 43146
rect 24820 43094 24840 43146
rect 24688 43092 24736 43094
rect 24792 43092 24840 43094
rect 24896 43092 24944 43094
rect 25000 43146 25048 43148
rect 25104 43146 25152 43148
rect 25000 43094 25016 43146
rect 25104 43094 25140 43146
rect 25000 43092 25048 43094
rect 25104 43092 25152 43094
rect 24008 43082 25208 43092
rect 23884 42802 23940 42812
rect 25004 42868 25060 42878
rect 25004 42774 25060 42812
rect 24556 42644 24612 42654
rect 24556 42550 24612 42588
rect 24444 41972 24500 41982
rect 24444 41878 24500 41916
rect 25340 41972 25396 41982
rect 25340 41878 25396 41916
rect 25452 41748 25508 41758
rect 25452 41654 25508 41692
rect 24008 41580 25208 41590
rect 24064 41578 24112 41580
rect 24168 41578 24216 41580
rect 24076 41526 24112 41578
rect 24200 41526 24216 41578
rect 24064 41524 24112 41526
rect 24168 41524 24216 41526
rect 24272 41578 24320 41580
rect 24376 41578 24424 41580
rect 24480 41578 24528 41580
rect 24376 41526 24396 41578
rect 24480 41526 24520 41578
rect 24272 41524 24320 41526
rect 24376 41524 24424 41526
rect 24480 41524 24528 41526
rect 24584 41524 24632 41580
rect 24688 41578 24736 41580
rect 24792 41578 24840 41580
rect 24896 41578 24944 41580
rect 24696 41526 24736 41578
rect 24820 41526 24840 41578
rect 24688 41524 24736 41526
rect 24792 41524 24840 41526
rect 24896 41524 24944 41526
rect 25000 41578 25048 41580
rect 25104 41578 25152 41580
rect 25000 41526 25016 41578
rect 25104 41526 25140 41578
rect 25000 41524 25048 41526
rect 25104 41524 25152 41526
rect 24008 41514 25208 41524
rect 25452 41412 25508 41422
rect 24668 41300 24724 41310
rect 24668 41186 24724 41244
rect 24668 41134 24670 41186
rect 24722 41134 24724 41186
rect 24668 41122 24724 41134
rect 24780 41188 24836 41198
rect 24780 41094 24836 41132
rect 25452 41188 25508 41356
rect 24556 41076 24612 41086
rect 24556 40982 24612 41020
rect 25228 41076 25284 41086
rect 25228 40982 25284 41020
rect 23884 40964 23940 40974
rect 23884 40870 23940 40908
rect 24332 40962 24388 40974
rect 24332 40910 24334 40962
rect 24386 40910 24388 40962
rect 24332 40292 24388 40910
rect 24444 40964 24500 40974
rect 24444 40870 24500 40908
rect 25452 40628 25508 41132
rect 25452 40562 25508 40572
rect 24332 40226 24388 40236
rect 25452 40292 25508 40302
rect 24008 40012 25208 40022
rect 24064 40010 24112 40012
rect 24168 40010 24216 40012
rect 24076 39958 24112 40010
rect 24200 39958 24216 40010
rect 24064 39956 24112 39958
rect 24168 39956 24216 39958
rect 24272 40010 24320 40012
rect 24376 40010 24424 40012
rect 24480 40010 24528 40012
rect 24376 39958 24396 40010
rect 24480 39958 24520 40010
rect 24272 39956 24320 39958
rect 24376 39956 24424 39958
rect 24480 39956 24528 39958
rect 24584 39956 24632 40012
rect 24688 40010 24736 40012
rect 24792 40010 24840 40012
rect 24896 40010 24944 40012
rect 24696 39958 24736 40010
rect 24820 39958 24840 40010
rect 24688 39956 24736 39958
rect 24792 39956 24840 39958
rect 24896 39956 24944 39958
rect 25000 40010 25048 40012
rect 25104 40010 25152 40012
rect 25000 39958 25016 40010
rect 25104 39958 25140 40010
rect 25000 39956 25048 39958
rect 25104 39956 25152 39958
rect 24008 39946 25208 39956
rect 24108 39844 24164 39854
rect 24108 38946 24164 39788
rect 24556 39620 24612 39630
rect 24556 39506 24612 39564
rect 24556 39454 24558 39506
rect 24610 39454 24612 39506
rect 24556 39442 24612 39454
rect 25340 39508 25396 39518
rect 25452 39508 25508 40236
rect 25340 39506 25508 39508
rect 25340 39454 25342 39506
rect 25394 39454 25508 39506
rect 25340 39452 25508 39454
rect 25340 39442 25396 39452
rect 24108 38894 24110 38946
rect 24162 38894 24164 38946
rect 24108 38882 24164 38894
rect 24008 38444 25208 38454
rect 24064 38442 24112 38444
rect 24168 38442 24216 38444
rect 24076 38390 24112 38442
rect 24200 38390 24216 38442
rect 24064 38388 24112 38390
rect 24168 38388 24216 38390
rect 24272 38442 24320 38444
rect 24376 38442 24424 38444
rect 24480 38442 24528 38444
rect 24376 38390 24396 38442
rect 24480 38390 24520 38442
rect 24272 38388 24320 38390
rect 24376 38388 24424 38390
rect 24480 38388 24528 38390
rect 24584 38388 24632 38444
rect 24688 38442 24736 38444
rect 24792 38442 24840 38444
rect 24896 38442 24944 38444
rect 24696 38390 24736 38442
rect 24820 38390 24840 38442
rect 24688 38388 24736 38390
rect 24792 38388 24840 38390
rect 24896 38388 24944 38390
rect 25000 38442 25048 38444
rect 25104 38442 25152 38444
rect 25000 38390 25016 38442
rect 25104 38390 25140 38442
rect 25000 38388 25048 38390
rect 25104 38388 25152 38390
rect 24008 38378 25208 38388
rect 24892 38164 24948 38174
rect 24892 38070 24948 38108
rect 25564 38164 25620 44492
rect 26012 44324 26068 45276
rect 26124 45106 26180 45118
rect 26124 45054 26126 45106
rect 26178 45054 26180 45106
rect 26124 44996 26180 45054
rect 26348 45108 26404 45118
rect 26348 45014 26404 45052
rect 26124 44930 26180 44940
rect 27244 44996 27300 45006
rect 27356 44996 27412 47852
rect 27468 46788 27524 50372
rect 28028 50372 28084 51438
rect 28476 53172 28532 53182
rect 28476 51490 28532 53116
rect 28476 51438 28478 51490
rect 28530 51438 28532 51490
rect 28476 51426 28532 51438
rect 29372 51380 29428 53452
rect 29372 51314 29428 51324
rect 28084 50316 28196 50372
rect 28028 50306 28084 50316
rect 27692 49924 27748 49934
rect 27580 49586 27636 49598
rect 27580 49534 27582 49586
rect 27634 49534 27636 49586
rect 27580 48244 27636 49534
rect 27692 49250 27748 49868
rect 28140 49922 28196 50316
rect 28140 49870 28142 49922
rect 28194 49870 28196 49922
rect 28140 49858 28196 49870
rect 28700 49922 28756 49934
rect 28700 49870 28702 49922
rect 28754 49870 28756 49922
rect 27916 49588 27972 49598
rect 27916 49586 28084 49588
rect 27916 49534 27918 49586
rect 27970 49534 28084 49586
rect 27916 49532 28084 49534
rect 27916 49522 27972 49532
rect 27692 49198 27694 49250
rect 27746 49198 27748 49250
rect 27692 49186 27748 49198
rect 28028 49250 28084 49532
rect 28028 49198 28030 49250
rect 28082 49198 28084 49250
rect 28028 49186 28084 49198
rect 28588 48804 28644 48814
rect 28588 48710 28644 48748
rect 28700 48468 28756 49870
rect 29596 49252 29652 58156
rect 29932 57876 29988 57886
rect 30044 57876 30100 59388
rect 30156 59332 30212 60844
rect 30268 60452 30324 60462
rect 30268 60002 30324 60396
rect 30268 59950 30270 60002
rect 30322 59950 30324 60002
rect 30268 59938 30324 59950
rect 30156 59266 30212 59276
rect 30380 58884 30436 61628
rect 30604 61460 30660 61470
rect 30604 60900 30660 61404
rect 30604 60786 30660 60844
rect 30604 60734 30606 60786
rect 30658 60734 30660 60786
rect 30604 60722 30660 60734
rect 30716 59892 30772 62302
rect 31276 62188 31332 62748
rect 31836 62188 31892 63756
rect 34860 63924 34916 63934
rect 34748 63252 34804 63262
rect 34748 63158 34804 63196
rect 34860 63026 34916 63868
rect 34860 62974 34862 63026
rect 34914 62974 34916 63026
rect 34860 62962 34916 62974
rect 35084 63028 35140 63038
rect 35084 62934 35140 62972
rect 33628 62914 33684 62926
rect 33628 62862 33630 62914
rect 33682 62862 33684 62914
rect 33628 62580 33684 62862
rect 34008 62748 35208 62758
rect 34064 62746 34112 62748
rect 34168 62746 34216 62748
rect 34076 62694 34112 62746
rect 34200 62694 34216 62746
rect 34064 62692 34112 62694
rect 34168 62692 34216 62694
rect 34272 62746 34320 62748
rect 34376 62746 34424 62748
rect 34480 62746 34528 62748
rect 34376 62694 34396 62746
rect 34480 62694 34520 62746
rect 34272 62692 34320 62694
rect 34376 62692 34424 62694
rect 34480 62692 34528 62694
rect 34584 62692 34632 62748
rect 34688 62746 34736 62748
rect 34792 62746 34840 62748
rect 34896 62746 34944 62748
rect 34696 62694 34736 62746
rect 34820 62694 34840 62746
rect 34688 62692 34736 62694
rect 34792 62692 34840 62694
rect 34896 62692 34944 62694
rect 35000 62746 35048 62748
rect 35104 62746 35152 62748
rect 35000 62694 35016 62746
rect 35104 62694 35140 62746
rect 35000 62692 35048 62694
rect 35104 62692 35152 62694
rect 34008 62682 35208 62692
rect 33404 62356 33460 62366
rect 33404 62262 33460 62300
rect 31276 62132 31444 62188
rect 31836 62132 32116 62188
rect 30828 61124 30884 61134
rect 30884 61068 30996 61124
rect 30828 61058 30884 61068
rect 30940 60228 30996 61068
rect 30604 59836 30716 59892
rect 30492 59444 30548 59454
rect 30492 59350 30548 59388
rect 30380 58818 30436 58828
rect 30268 58436 30324 58446
rect 30268 58434 30436 58436
rect 30268 58382 30270 58434
rect 30322 58382 30436 58434
rect 30268 58380 30436 58382
rect 30268 58370 30324 58380
rect 29932 57874 30100 57876
rect 29932 57822 29934 57874
rect 29986 57822 30100 57874
rect 29932 57820 30100 57822
rect 30268 58210 30324 58222
rect 30268 58158 30270 58210
rect 30322 58158 30324 58210
rect 29932 57810 29988 57820
rect 30268 57316 30324 58158
rect 30380 58212 30436 58380
rect 30604 58434 30660 59836
rect 30716 59826 30772 59836
rect 30828 60172 30996 60228
rect 31052 60786 31108 60798
rect 31052 60734 31054 60786
rect 31106 60734 31108 60786
rect 31052 60676 31108 60734
rect 30604 58382 30606 58434
rect 30658 58382 30660 58434
rect 30604 58370 30660 58382
rect 30380 58146 30436 58156
rect 30828 58100 30884 60172
rect 30940 60004 30996 60014
rect 30940 59910 30996 59948
rect 31052 59780 31108 60620
rect 31052 59108 31108 59724
rect 30940 59052 31108 59108
rect 31276 59332 31332 59342
rect 30940 58212 30996 59052
rect 30940 58118 30996 58156
rect 31052 58884 31108 58894
rect 30492 58044 30884 58100
rect 30492 57874 30548 58044
rect 30492 57822 30494 57874
rect 30546 57822 30548 57874
rect 30492 57810 30548 57822
rect 29708 57260 30324 57316
rect 30716 57316 30772 58044
rect 30828 57876 30884 57886
rect 30828 57538 30884 57820
rect 30940 57876 30996 57886
rect 31052 57876 31108 58828
rect 31276 58658 31332 59276
rect 31276 58606 31278 58658
rect 31330 58606 31332 58658
rect 31276 58594 31332 58606
rect 31388 58436 31444 62132
rect 31724 60900 31780 60910
rect 31500 60788 31556 60798
rect 31724 60788 31780 60844
rect 31500 60694 31556 60732
rect 31612 60786 31780 60788
rect 31612 60734 31726 60786
rect 31778 60734 31780 60786
rect 31612 60732 31780 60734
rect 31612 60004 31668 60732
rect 31724 60722 31780 60732
rect 32060 60786 32116 62132
rect 32508 61348 32564 61358
rect 32060 60734 32062 60786
rect 32114 60734 32116 60786
rect 31948 60674 32004 60686
rect 31948 60622 31950 60674
rect 32002 60622 32004 60674
rect 31500 59948 31668 60004
rect 31724 60004 31780 60014
rect 31500 58772 31556 59948
rect 31612 59780 31668 59790
rect 31612 59442 31668 59724
rect 31612 59390 31614 59442
rect 31666 59390 31668 59442
rect 31612 59378 31668 59390
rect 31724 59442 31780 59948
rect 31724 59390 31726 59442
rect 31778 59390 31780 59442
rect 31724 59378 31780 59390
rect 31836 59330 31892 59342
rect 31836 59278 31838 59330
rect 31890 59278 31892 59330
rect 31836 58772 31892 59278
rect 31948 59218 32004 60622
rect 32060 60676 32116 60734
rect 32060 60610 32116 60620
rect 32396 60786 32452 60798
rect 32396 60734 32398 60786
rect 32450 60734 32452 60786
rect 32396 60228 32452 60734
rect 31948 59166 31950 59218
rect 32002 59166 32004 59218
rect 31948 59154 32004 59166
rect 32284 60116 32340 60126
rect 32284 59218 32340 60060
rect 32284 59166 32286 59218
rect 32338 59166 32340 59218
rect 32284 59154 32340 59166
rect 31500 58716 31780 58772
rect 31836 58716 32228 58772
rect 31612 58548 31668 58558
rect 31388 58380 31556 58436
rect 31388 58212 31444 58222
rect 31388 58118 31444 58156
rect 30940 57874 31108 57876
rect 30940 57822 30942 57874
rect 30994 57822 31108 57874
rect 30940 57820 31108 57822
rect 30940 57810 30996 57820
rect 30828 57486 30830 57538
rect 30882 57486 30884 57538
rect 30828 57474 30884 57486
rect 31164 57426 31220 57438
rect 31164 57374 31166 57426
rect 31218 57374 31220 57426
rect 31164 57316 31220 57374
rect 30716 57260 31220 57316
rect 29708 56866 29764 57260
rect 29708 56814 29710 56866
rect 29762 56814 29764 56866
rect 29708 56802 29764 56814
rect 31164 56644 31220 57260
rect 31164 56578 31220 56588
rect 30268 56196 30324 56206
rect 30268 54740 30324 56140
rect 31164 56084 31220 56094
rect 31164 54740 31220 56028
rect 29708 54738 30324 54740
rect 29708 54686 30270 54738
rect 30322 54686 30324 54738
rect 29708 54684 30324 54686
rect 29708 53170 29764 54684
rect 30268 54674 30324 54684
rect 31052 54738 31220 54740
rect 31052 54686 31166 54738
rect 31218 54686 31220 54738
rect 31052 54684 31220 54686
rect 30380 54516 30436 54526
rect 30380 53954 30436 54460
rect 30828 54292 30884 54302
rect 30828 54290 30996 54292
rect 30828 54238 30830 54290
rect 30882 54238 30996 54290
rect 30828 54236 30996 54238
rect 30828 54226 30884 54236
rect 30380 53902 30382 53954
rect 30434 53902 30436 53954
rect 30380 53842 30436 53902
rect 30380 53790 30382 53842
rect 30434 53790 30436 53842
rect 30380 53778 30436 53790
rect 30940 53732 30996 54236
rect 30940 53666 30996 53676
rect 31052 53954 31108 54684
rect 31164 54674 31220 54684
rect 31052 53902 31054 53954
rect 31106 53902 31108 53954
rect 29708 53118 29710 53170
rect 29762 53118 29764 53170
rect 29708 53106 29764 53118
rect 30268 53620 30324 53630
rect 30268 53170 30324 53564
rect 30828 53620 30884 53630
rect 30828 53172 30884 53564
rect 30268 53118 30270 53170
rect 30322 53118 30324 53170
rect 30268 52948 30324 53118
rect 30268 52882 30324 52892
rect 30492 53116 30996 53172
rect 30044 52276 30100 52286
rect 30044 52182 30100 52220
rect 30268 52164 30324 52174
rect 30268 52070 30324 52108
rect 29596 49186 29652 49196
rect 30156 50708 30212 50718
rect 28700 48402 28756 48412
rect 30156 48466 30212 50652
rect 30156 48414 30158 48466
rect 30210 48414 30212 48466
rect 30156 48402 30212 48414
rect 30380 48580 30436 48590
rect 27692 48244 27748 48254
rect 27580 48242 27748 48244
rect 27580 48190 27694 48242
rect 27746 48190 27748 48242
rect 27580 48188 27748 48190
rect 27692 48178 27748 48188
rect 29260 47572 29316 47582
rect 29260 47478 29316 47516
rect 29484 47348 29540 47358
rect 27468 46722 27524 46732
rect 27916 47234 27972 47246
rect 27916 47182 27918 47234
rect 27970 47182 27972 47234
rect 27916 46900 27972 47182
rect 27916 46674 27972 46844
rect 28364 47234 28420 47246
rect 28364 47182 28366 47234
rect 28418 47182 28420 47234
rect 28364 47012 28420 47182
rect 27916 46622 27918 46674
rect 27970 46622 27972 46674
rect 27916 46610 27972 46622
rect 28028 46786 28084 46798
rect 28028 46734 28030 46786
rect 28082 46734 28084 46786
rect 27300 44940 27412 44996
rect 27468 46562 27524 46574
rect 27468 46510 27470 46562
rect 27522 46510 27524 46562
rect 27468 46452 27524 46510
rect 28028 46452 28084 46734
rect 27468 46396 28084 46452
rect 27244 44902 27300 44940
rect 26012 44258 26068 44268
rect 26236 44884 26292 44894
rect 26012 43316 26068 43326
rect 26012 42082 26068 43260
rect 26012 42030 26014 42082
rect 26066 42030 26068 42082
rect 26012 42018 26068 42030
rect 26124 42868 26180 42878
rect 26124 42082 26180 42812
rect 26124 42030 26126 42082
rect 26178 42030 26180 42082
rect 26124 42018 26180 42030
rect 26236 42866 26292 44828
rect 26796 43426 26852 43438
rect 26796 43374 26798 43426
rect 26850 43374 26852 43426
rect 26796 43316 26852 43374
rect 26852 43260 27076 43316
rect 26796 43222 26852 43260
rect 26236 42814 26238 42866
rect 26290 42814 26292 42866
rect 25788 41970 25844 41982
rect 25788 41918 25790 41970
rect 25842 41918 25844 41970
rect 25788 41412 25844 41918
rect 26236 41972 26292 42814
rect 26572 42868 26628 42878
rect 26572 42754 26628 42812
rect 26572 42702 26574 42754
rect 26626 42702 26628 42754
rect 26572 42690 26628 42702
rect 26796 42754 26852 42766
rect 26796 42702 26798 42754
rect 26850 42702 26852 42754
rect 26684 42530 26740 42542
rect 26684 42478 26686 42530
rect 26738 42478 26740 42530
rect 26684 41972 26740 42478
rect 26236 41860 26292 41916
rect 25788 41346 25844 41356
rect 25900 41804 26292 41860
rect 26460 41916 26740 41972
rect 25788 41188 25844 41198
rect 25788 41094 25844 41132
rect 25900 40402 25956 41804
rect 26460 41410 26516 41916
rect 26460 41358 26462 41410
rect 26514 41358 26516 41410
rect 26460 41346 26516 41358
rect 26572 41746 26628 41758
rect 26572 41694 26574 41746
rect 26626 41694 26628 41746
rect 26572 41412 26628 41694
rect 26684 41412 26740 41422
rect 26572 41410 26740 41412
rect 26572 41358 26686 41410
rect 26738 41358 26740 41410
rect 26572 41356 26740 41358
rect 26684 41346 26740 41356
rect 26012 41300 26068 41310
rect 26012 41206 26068 41244
rect 26124 40964 26180 40974
rect 26124 40962 26516 40964
rect 26124 40910 26126 40962
rect 26178 40910 26516 40962
rect 26124 40908 26516 40910
rect 26124 40898 26180 40908
rect 25900 40350 25902 40402
rect 25954 40350 25956 40402
rect 25900 40338 25956 40350
rect 26460 40402 26516 40908
rect 26796 40628 26852 42702
rect 27020 42756 27076 43260
rect 27020 42662 27076 42700
rect 27020 41972 27076 41982
rect 27356 41972 27412 41982
rect 26908 41188 26964 41198
rect 26908 41094 26964 41132
rect 26796 40562 26852 40572
rect 26460 40350 26462 40402
rect 26514 40350 26516 40402
rect 26460 40338 26516 40350
rect 27020 40404 27076 41916
rect 27244 41970 27412 41972
rect 27244 41918 27358 41970
rect 27410 41918 27412 41970
rect 27244 41916 27412 41918
rect 27132 41748 27188 41758
rect 27132 41186 27188 41692
rect 27244 41298 27300 41916
rect 27356 41906 27412 41916
rect 27244 41246 27246 41298
rect 27298 41246 27300 41298
rect 27244 41234 27300 41246
rect 27356 41412 27412 41422
rect 27132 41134 27134 41186
rect 27186 41134 27188 41186
rect 27132 41122 27188 41134
rect 27356 41186 27412 41356
rect 27356 41134 27358 41186
rect 27410 41134 27412 41186
rect 27356 41122 27412 41134
rect 27020 40338 27076 40348
rect 26124 39732 26180 39742
rect 26124 39638 26180 39676
rect 25676 39620 25732 39630
rect 25676 39526 25732 39564
rect 27468 38668 27524 46396
rect 27804 45780 27860 45790
rect 27804 45330 27860 45724
rect 28140 45668 28196 45678
rect 28364 45668 28420 46956
rect 28700 47012 28756 47022
rect 28700 46674 28756 46956
rect 28700 46622 28702 46674
rect 28754 46622 28756 46674
rect 28700 46610 28756 46622
rect 29036 46452 29092 46462
rect 29484 46452 29540 47292
rect 30380 47348 30436 48524
rect 30492 48356 30548 53116
rect 30940 53058 30996 53116
rect 30940 53006 30942 53058
rect 30994 53006 30996 53058
rect 30940 52994 30996 53006
rect 30828 52948 30884 52958
rect 30828 52854 30884 52892
rect 31052 52276 31108 53902
rect 31276 53732 31332 53742
rect 31276 53618 31332 53676
rect 31276 53566 31278 53618
rect 31330 53566 31332 53618
rect 31276 53172 31332 53566
rect 31388 53620 31444 53630
rect 31500 53620 31556 58380
rect 31612 58434 31668 58492
rect 31612 58382 31614 58434
rect 31666 58382 31668 58434
rect 31612 58370 31668 58382
rect 31724 58436 31780 58716
rect 32172 58658 32228 58716
rect 32172 58606 32174 58658
rect 32226 58606 32228 58658
rect 32172 58594 32228 58606
rect 32284 58548 32340 58558
rect 32396 58548 32452 60172
rect 32508 59444 32564 61292
rect 33068 61346 33124 61358
rect 33068 61294 33070 61346
rect 33122 61294 33124 61346
rect 33068 60900 33124 61294
rect 33404 61346 33460 61358
rect 33404 61294 33406 61346
rect 33458 61294 33460 61346
rect 33180 61012 33236 61022
rect 33180 60918 33236 60956
rect 33068 60834 33124 60844
rect 33292 60788 33348 60798
rect 33292 60694 33348 60732
rect 33404 60676 33460 61294
rect 33628 61348 33684 62524
rect 34412 62468 34468 62478
rect 33628 61282 33684 61292
rect 33740 62356 33796 62366
rect 33852 62356 33908 62366
rect 33796 62354 33908 62356
rect 33796 62302 33854 62354
rect 33906 62302 33908 62354
rect 33796 62300 33908 62302
rect 33740 61012 33796 62300
rect 33852 62290 33908 62300
rect 34412 62354 34468 62412
rect 34412 62302 34414 62354
rect 34466 62302 34468 62354
rect 34412 62290 34468 62302
rect 35420 62188 35476 64652
rect 35644 64642 35700 64652
rect 36092 64708 36148 64718
rect 36204 64708 36260 65998
rect 36316 66050 36372 66062
rect 36316 65998 36318 66050
rect 36370 65998 36372 66050
rect 36316 65492 36372 65998
rect 36876 65714 36932 66108
rect 36876 65662 36878 65714
rect 36930 65662 36932 65714
rect 36876 65650 36932 65662
rect 36316 65426 36372 65436
rect 36988 64932 37044 64942
rect 37100 64932 37156 66556
rect 37324 66498 37380 66556
rect 37324 66446 37326 66498
rect 37378 66446 37380 66498
rect 37324 66434 37380 66446
rect 37548 66386 37604 67228
rect 37660 67218 37716 67228
rect 37548 66334 37550 66386
rect 37602 66334 37604 66386
rect 37548 66322 37604 66334
rect 37660 65492 37716 65502
rect 37548 65436 37660 65492
rect 37044 64876 37156 64932
rect 37324 65044 37380 65054
rect 37324 64930 37380 64988
rect 37324 64878 37326 64930
rect 37378 64878 37380 64930
rect 36988 64838 37044 64876
rect 36092 64706 36260 64708
rect 36092 64654 36094 64706
rect 36146 64654 36260 64706
rect 36092 64652 36260 64654
rect 36092 64642 36148 64652
rect 37324 63924 37380 64878
rect 37548 64818 37604 65436
rect 37660 65398 37716 65436
rect 37548 64766 37550 64818
rect 37602 64766 37604 64818
rect 37548 64754 37604 64766
rect 35868 63028 35924 63038
rect 35868 62934 35924 62972
rect 35532 62916 35588 62926
rect 35532 62822 35588 62860
rect 35756 62916 35812 62926
rect 35756 62822 35812 62860
rect 35980 62914 36036 62926
rect 35980 62862 35982 62914
rect 36034 62862 36036 62914
rect 35980 62188 36036 62862
rect 36764 62580 36820 62590
rect 35420 62132 35588 62188
rect 35980 62132 36260 62188
rect 35532 61684 35588 62132
rect 35980 61684 36036 61694
rect 35532 61682 36036 61684
rect 35532 61630 35534 61682
rect 35586 61630 35982 61682
rect 36034 61630 36036 61682
rect 35532 61628 36036 61630
rect 35532 61618 35588 61628
rect 35980 61618 36036 61628
rect 36204 61572 36260 62132
rect 36764 62132 36820 62524
rect 37324 62188 37380 63868
rect 36764 62066 36820 62076
rect 36988 62132 37380 62188
rect 37548 62916 37604 62926
rect 37548 62578 37604 62860
rect 37548 62526 37550 62578
rect 37602 62526 37604 62578
rect 36988 61794 37044 62132
rect 36988 61742 36990 61794
rect 37042 61742 37044 61794
rect 36988 61730 37044 61742
rect 37548 61682 37604 62526
rect 37548 61630 37550 61682
rect 37602 61630 37604 61682
rect 37548 61618 37604 61630
rect 37772 62132 37828 62142
rect 36204 61478 36260 61516
rect 36316 61570 36372 61582
rect 36316 61518 36318 61570
rect 36370 61518 36372 61570
rect 35868 61460 35924 61470
rect 35644 61458 35924 61460
rect 35644 61406 35870 61458
rect 35922 61406 35924 61458
rect 35644 61404 35924 61406
rect 33852 61348 33908 61358
rect 33852 61254 33908 61292
rect 34412 61348 34468 61386
rect 34412 61282 34468 61292
rect 34008 61180 35208 61190
rect 34064 61178 34112 61180
rect 34168 61178 34216 61180
rect 34076 61126 34112 61178
rect 34200 61126 34216 61178
rect 34064 61124 34112 61126
rect 34168 61124 34216 61126
rect 34272 61178 34320 61180
rect 34376 61178 34424 61180
rect 34480 61178 34528 61180
rect 34376 61126 34396 61178
rect 34480 61126 34520 61178
rect 34272 61124 34320 61126
rect 34376 61124 34424 61126
rect 34480 61124 34528 61126
rect 34584 61124 34632 61180
rect 34688 61178 34736 61180
rect 34792 61178 34840 61180
rect 34896 61178 34944 61180
rect 34696 61126 34736 61178
rect 34820 61126 34840 61178
rect 34688 61124 34736 61126
rect 34792 61124 34840 61126
rect 34896 61124 34944 61126
rect 35000 61178 35048 61180
rect 35104 61178 35152 61180
rect 35000 61126 35016 61178
rect 35104 61126 35140 61178
rect 35000 61124 35048 61126
rect 35104 61124 35152 61126
rect 34008 61114 35208 61124
rect 34188 61012 34244 61022
rect 33740 61010 34692 61012
rect 33740 60958 34190 61010
rect 34242 60958 34692 61010
rect 33740 60956 34692 60958
rect 33404 60610 33460 60620
rect 33740 60676 33796 60686
rect 33740 60582 33796 60620
rect 33180 60564 33236 60574
rect 33180 60470 33236 60508
rect 32508 59378 32564 59388
rect 33180 59780 33236 59790
rect 33180 59444 33236 59724
rect 33180 59378 33236 59388
rect 33068 59332 33124 59342
rect 33068 59238 33124 59276
rect 33292 59330 33348 59342
rect 33292 59278 33294 59330
rect 33346 59278 33348 59330
rect 33292 58884 33348 59278
rect 33292 58818 33348 58828
rect 33404 58994 33460 59006
rect 33404 58942 33406 58994
rect 33458 58942 33460 58994
rect 32340 58492 32452 58548
rect 32284 58454 32340 58492
rect 31836 58436 31892 58446
rect 31724 58434 31892 58436
rect 31724 58382 31838 58434
rect 31890 58382 31892 58434
rect 31724 58380 31892 58382
rect 31836 58370 31892 58380
rect 33404 58436 33460 58942
rect 32732 58212 32788 58222
rect 32060 56642 32116 56654
rect 32060 56590 32062 56642
rect 32114 56590 32116 56642
rect 32060 56196 32116 56590
rect 32060 56102 32116 56140
rect 32732 56642 32788 58156
rect 33404 57652 33460 58380
rect 33740 57876 33796 57886
rect 33852 57876 33908 60956
rect 34188 60946 34244 60956
rect 34636 60786 34692 60956
rect 34636 60734 34638 60786
rect 34690 60734 34692 60786
rect 34636 60722 34692 60734
rect 35308 60788 35364 60798
rect 35644 60788 35700 61404
rect 35868 61394 35924 61404
rect 35308 60786 35700 60788
rect 35308 60734 35310 60786
rect 35362 60734 35700 60786
rect 35308 60732 35700 60734
rect 35308 60722 35364 60732
rect 33964 60228 34020 60238
rect 33964 60134 34020 60172
rect 36204 60228 36260 60238
rect 36204 59890 36260 60172
rect 36316 60114 36372 61518
rect 37324 61572 37380 61582
rect 36988 60228 37044 60238
rect 37324 60228 37380 61516
rect 37772 61010 37828 62076
rect 37772 60958 37774 61010
rect 37826 60958 37828 61010
rect 37772 60946 37828 60958
rect 38332 60562 38388 60574
rect 38332 60510 38334 60562
rect 38386 60510 38388 60562
rect 36988 60226 37380 60228
rect 36988 60174 36990 60226
rect 37042 60174 37380 60226
rect 36988 60172 37380 60174
rect 37548 60228 37604 60238
rect 36988 60162 37044 60172
rect 36316 60062 36318 60114
rect 36370 60062 36372 60114
rect 36316 60050 36372 60062
rect 37548 60114 37604 60172
rect 38332 60228 38388 60510
rect 38332 60162 38388 60172
rect 37548 60062 37550 60114
rect 37602 60062 37604 60114
rect 37548 60050 37604 60062
rect 36428 60004 36484 60014
rect 37324 60004 37380 60014
rect 36428 59910 36484 59948
rect 37212 59948 37324 60004
rect 36204 59838 36206 59890
rect 36258 59838 36260 59890
rect 36204 59826 36260 59838
rect 34300 59780 34356 59818
rect 34300 59714 34356 59724
rect 34008 59612 35208 59622
rect 34064 59610 34112 59612
rect 34168 59610 34216 59612
rect 34076 59558 34112 59610
rect 34200 59558 34216 59610
rect 34064 59556 34112 59558
rect 34168 59556 34216 59558
rect 34272 59610 34320 59612
rect 34376 59610 34424 59612
rect 34480 59610 34528 59612
rect 34376 59558 34396 59610
rect 34480 59558 34520 59610
rect 34272 59556 34320 59558
rect 34376 59556 34424 59558
rect 34480 59556 34528 59558
rect 34584 59556 34632 59612
rect 34688 59610 34736 59612
rect 34792 59610 34840 59612
rect 34896 59610 34944 59612
rect 34696 59558 34736 59610
rect 34820 59558 34840 59610
rect 34688 59556 34736 59558
rect 34792 59556 34840 59558
rect 34896 59556 34944 59558
rect 35000 59610 35048 59612
rect 35104 59610 35152 59612
rect 35000 59558 35016 59610
rect 35104 59558 35140 59610
rect 35000 59556 35048 59558
rect 35104 59556 35152 59558
rect 34008 59546 35208 59556
rect 34972 58434 35028 58446
rect 34972 58382 34974 58434
rect 35026 58382 35028 58434
rect 34412 58324 34468 58334
rect 34412 58210 34468 58268
rect 34412 58158 34414 58210
rect 34466 58158 34468 58210
rect 34412 58146 34468 58158
rect 34972 58212 35028 58382
rect 35196 58436 35252 58446
rect 35196 58342 35252 58380
rect 36876 58434 36932 58446
rect 36876 58382 36878 58434
rect 36930 58382 36932 58434
rect 35084 58324 35140 58334
rect 35084 58212 35140 58268
rect 35532 58324 35588 58334
rect 35084 58156 35364 58212
rect 34972 58146 35028 58156
rect 34008 58044 35208 58054
rect 34064 58042 34112 58044
rect 34168 58042 34216 58044
rect 34076 57990 34112 58042
rect 34200 57990 34216 58042
rect 34064 57988 34112 57990
rect 34168 57988 34216 57990
rect 34272 58042 34320 58044
rect 34376 58042 34424 58044
rect 34480 58042 34528 58044
rect 34376 57990 34396 58042
rect 34480 57990 34520 58042
rect 34272 57988 34320 57990
rect 34376 57988 34424 57990
rect 34480 57988 34528 57990
rect 34584 57988 34632 58044
rect 34688 58042 34736 58044
rect 34792 58042 34840 58044
rect 34896 58042 34944 58044
rect 34696 57990 34736 58042
rect 34820 57990 34840 58042
rect 34688 57988 34736 57990
rect 34792 57988 34840 57990
rect 34896 57988 34944 57990
rect 35000 58042 35048 58044
rect 35104 58042 35152 58044
rect 35000 57990 35016 58042
rect 35104 57990 35140 58042
rect 35000 57988 35048 57990
rect 35104 57988 35152 57990
rect 34008 57978 35208 57988
rect 34300 57876 34356 57886
rect 35308 57876 35364 58156
rect 33404 57586 33460 57596
rect 33628 57874 34244 57876
rect 33628 57822 33742 57874
rect 33794 57822 34244 57874
rect 33628 57820 34244 57822
rect 32732 56590 32734 56642
rect 32786 56590 32788 56642
rect 32508 56084 32564 56094
rect 32508 55990 32564 56028
rect 31444 53564 31556 53620
rect 31948 53620 32004 53630
rect 31388 53526 31444 53564
rect 31948 53526 32004 53564
rect 31276 53106 31332 53116
rect 31612 53506 31668 53518
rect 31612 53454 31614 53506
rect 31666 53454 31668 53506
rect 31164 52948 31220 52958
rect 31500 52948 31556 52958
rect 31164 52946 31556 52948
rect 31164 52894 31166 52946
rect 31218 52894 31502 52946
rect 31554 52894 31556 52946
rect 31164 52892 31556 52894
rect 31164 52882 31220 52892
rect 31500 52882 31556 52892
rect 31052 52164 31108 52220
rect 31164 52164 31220 52174
rect 31052 52162 31220 52164
rect 31052 52110 31166 52162
rect 31218 52110 31220 52162
rect 31052 52108 31220 52110
rect 30716 52052 30772 52062
rect 30716 51958 30772 51996
rect 30828 51940 30884 51950
rect 30828 51846 30884 51884
rect 30940 51940 30996 51950
rect 30940 51938 31108 51940
rect 30940 51886 30942 51938
rect 30994 51886 31108 51938
rect 30940 51884 31108 51886
rect 30940 51874 30996 51884
rect 30940 51604 30996 51614
rect 30716 51548 30940 51604
rect 30716 50708 30772 51548
rect 30940 51510 30996 51548
rect 30716 50614 30772 50652
rect 31052 49140 31108 51884
rect 31052 49074 31108 49084
rect 31164 50706 31220 52108
rect 31612 52164 31668 53454
rect 31948 52946 32004 52958
rect 31948 52894 31950 52946
rect 32002 52894 32004 52946
rect 31948 52388 32004 52894
rect 32172 52948 32228 52958
rect 32172 52946 32452 52948
rect 32172 52894 32174 52946
rect 32226 52894 32452 52946
rect 32172 52892 32452 52894
rect 32172 52882 32228 52892
rect 31612 52098 31668 52108
rect 31724 52332 32004 52388
rect 32060 52834 32116 52846
rect 32060 52782 32062 52834
rect 32114 52782 32116 52834
rect 31724 52052 31780 52332
rect 31836 52164 31892 52174
rect 32060 52164 32116 52782
rect 31836 52162 32116 52164
rect 31836 52110 31838 52162
rect 31890 52110 32116 52162
rect 31836 52108 32116 52110
rect 31836 52098 31892 52108
rect 31724 51716 31780 51996
rect 32172 51940 32228 51950
rect 31724 51660 31892 51716
rect 31612 51266 31668 51278
rect 31612 51214 31614 51266
rect 31666 51214 31668 51266
rect 31612 50820 31668 51214
rect 31612 50764 31780 50820
rect 31164 50654 31166 50706
rect 31218 50654 31220 50706
rect 31164 50596 31220 50654
rect 31612 50596 31668 50606
rect 31164 50594 31668 50596
rect 31164 50542 31614 50594
rect 31666 50542 31668 50594
rect 31164 50540 31668 50542
rect 31164 49700 31220 50540
rect 31612 50530 31668 50540
rect 30828 48468 30884 48478
rect 30884 48412 31108 48468
rect 30828 48374 30884 48412
rect 30492 48290 30548 48300
rect 30716 47570 30772 47582
rect 30716 47518 30718 47570
rect 30770 47518 30772 47570
rect 30716 47460 30772 47518
rect 30716 47394 30772 47404
rect 31052 47458 31108 48412
rect 31164 48244 31220 49644
rect 31724 49252 31780 50764
rect 31612 49140 31668 49150
rect 31724 49140 31780 49196
rect 31612 49138 31780 49140
rect 31612 49086 31614 49138
rect 31666 49086 31780 49138
rect 31612 49084 31780 49086
rect 31612 49074 31668 49084
rect 31276 49026 31332 49038
rect 31836 49028 31892 51660
rect 31948 51380 32004 51390
rect 31948 51286 32004 51324
rect 32172 50594 32228 51884
rect 32396 51490 32452 52892
rect 32396 51438 32398 51490
rect 32450 51438 32452 51490
rect 32396 51426 32452 51438
rect 32172 50542 32174 50594
rect 32226 50542 32228 50594
rect 32172 50530 32228 50542
rect 32620 51380 32676 51390
rect 32172 49700 32228 49710
rect 32172 49698 32340 49700
rect 32172 49646 32174 49698
rect 32226 49646 32340 49698
rect 32172 49644 32340 49646
rect 32172 49634 32228 49644
rect 31276 48974 31278 49026
rect 31330 48974 31332 49026
rect 31276 48580 31332 48974
rect 31724 48972 31892 49028
rect 31948 49586 32004 49598
rect 31948 49534 31950 49586
rect 32002 49534 32004 49586
rect 31612 48916 31668 48926
rect 31612 48822 31668 48860
rect 31276 48514 31332 48524
rect 31164 48150 31220 48188
rect 31276 48356 31332 48366
rect 31052 47406 31054 47458
rect 31106 47406 31108 47458
rect 31052 47394 31108 47406
rect 31276 47458 31332 48300
rect 31724 48244 31780 48972
rect 31836 48804 31892 48814
rect 31948 48804 32004 49534
rect 32172 49140 32228 49150
rect 32172 49046 32228 49084
rect 31892 48748 32004 48804
rect 31836 48710 31892 48748
rect 31836 48244 31892 48254
rect 31724 48188 31836 48244
rect 31836 48150 31892 48188
rect 31612 48018 31668 48030
rect 31612 47966 31614 48018
rect 31666 47966 31668 48018
rect 31612 47796 31668 47966
rect 31388 47740 31668 47796
rect 31388 47570 31444 47740
rect 31388 47518 31390 47570
rect 31442 47518 31444 47570
rect 31388 47506 31444 47518
rect 31276 47406 31278 47458
rect 31330 47406 31332 47458
rect 30380 47254 30436 47292
rect 30156 47234 30212 47246
rect 30156 47182 30158 47234
rect 30210 47182 30212 47234
rect 30156 47124 30212 47182
rect 30604 47234 30660 47246
rect 30604 47182 30606 47234
rect 30658 47182 30660 47234
rect 30604 47124 30660 47182
rect 31276 47236 31332 47406
rect 31276 47170 31332 47180
rect 31500 47460 31556 47470
rect 30156 47068 30660 47124
rect 29596 47012 29652 47022
rect 29596 46898 29652 46956
rect 29596 46846 29598 46898
rect 29650 46846 29652 46898
rect 29596 46834 29652 46846
rect 30604 46900 30660 47068
rect 31164 46900 31220 46910
rect 30604 46898 31220 46900
rect 30604 46846 30606 46898
rect 30658 46846 31166 46898
rect 31218 46846 31220 46898
rect 30604 46844 31220 46846
rect 30604 46834 30660 46844
rect 30156 46562 30212 46574
rect 30156 46510 30158 46562
rect 30210 46510 30212 46562
rect 30156 46452 30212 46510
rect 29036 46450 29540 46452
rect 29036 46398 29038 46450
rect 29090 46398 29540 46450
rect 29036 46396 29540 46398
rect 29036 46386 29092 46396
rect 28700 45780 28756 45790
rect 28700 45686 28756 45724
rect 28196 45612 28420 45668
rect 29260 45668 29316 45678
rect 28140 45574 28196 45612
rect 27804 45278 27806 45330
rect 27858 45278 27860 45330
rect 27804 45266 27860 45278
rect 27692 45108 27748 45118
rect 27692 45014 27748 45052
rect 27580 44996 27636 45006
rect 27580 44902 27636 44940
rect 29148 43652 29204 43662
rect 28140 42868 28196 42878
rect 27580 42756 27636 42766
rect 27580 42662 27636 42700
rect 28140 41410 28196 42812
rect 29036 41412 29092 41422
rect 28140 41358 28142 41410
rect 28194 41358 28196 41410
rect 28140 41346 28196 41358
rect 28588 41410 29092 41412
rect 28588 41358 29038 41410
rect 29090 41358 29092 41410
rect 28588 41356 29092 41358
rect 27804 41300 27860 41310
rect 27804 41206 27860 41244
rect 28588 41298 28644 41356
rect 29036 41346 29092 41356
rect 28588 41246 28590 41298
rect 28642 41246 28644 41298
rect 28588 41234 28644 41246
rect 29148 41300 29204 43596
rect 29260 41972 29316 45612
rect 29372 45556 29428 45566
rect 29372 43428 29428 45500
rect 29484 43540 29540 46396
rect 29932 46396 30212 46452
rect 29708 45666 29764 45678
rect 29708 45614 29710 45666
rect 29762 45614 29764 45666
rect 29708 44996 29764 45614
rect 29820 45668 29876 45678
rect 29932 45668 29988 46396
rect 30156 46116 30212 46126
rect 30156 46022 30212 46060
rect 30380 45890 30436 45902
rect 30380 45838 30382 45890
rect 30434 45838 30436 45890
rect 30044 45780 30100 45790
rect 30044 45686 30100 45724
rect 29876 45612 29988 45668
rect 29820 45602 29876 45612
rect 30380 45444 30436 45838
rect 30156 45388 30436 45444
rect 29932 44996 29988 45006
rect 30156 44996 30212 45388
rect 30604 44996 30660 45006
rect 29708 44994 30212 44996
rect 29708 44942 29934 44994
rect 29986 44942 30212 44994
rect 29708 44940 30212 44942
rect 30268 44994 30660 44996
rect 30268 44942 30606 44994
rect 30658 44942 30660 44994
rect 30268 44940 30660 44942
rect 29932 44930 29988 44940
rect 29484 43474 29540 43484
rect 29820 43650 29876 43662
rect 29820 43598 29822 43650
rect 29874 43598 29876 43650
rect 29372 43316 29428 43372
rect 29484 43316 29540 43326
rect 29372 43314 29540 43316
rect 29372 43262 29486 43314
rect 29538 43262 29540 43314
rect 29372 43260 29540 43262
rect 29484 43250 29540 43260
rect 29596 43314 29652 43326
rect 29596 43262 29598 43314
rect 29650 43262 29652 43314
rect 29596 42868 29652 43262
rect 29596 42802 29652 42812
rect 29260 41906 29316 41916
rect 29820 41410 29876 43598
rect 29820 41358 29822 41410
rect 29874 41358 29876 41410
rect 29260 41300 29316 41310
rect 29708 41300 29764 41310
rect 29148 41298 29540 41300
rect 29148 41246 29262 41298
rect 29314 41246 29540 41298
rect 29148 41244 29540 41246
rect 28476 41188 28532 41198
rect 28476 41094 28532 41132
rect 27916 40964 27972 40974
rect 27916 40870 27972 40908
rect 29148 40964 29204 41244
rect 29260 41234 29316 41244
rect 29148 40898 29204 40908
rect 29036 40740 29092 40750
rect 29036 40626 29092 40684
rect 29036 40574 29038 40626
rect 29090 40574 29092 40626
rect 29036 40562 29092 40574
rect 24668 37492 24724 37502
rect 24668 37398 24724 37436
rect 23772 37324 24052 37380
rect 23436 35588 23492 35598
rect 23324 35532 23436 35588
rect 21756 34020 21812 34030
rect 21756 33926 21812 33964
rect 22204 34018 22260 34030
rect 22204 33966 22206 34018
rect 22258 33966 22260 34018
rect 22204 33572 22260 33966
rect 23212 33684 23268 34748
rect 23212 33618 23268 33628
rect 22204 33506 22260 33516
rect 23436 33572 23492 35532
rect 23548 35476 23604 35486
rect 23548 34914 23604 35420
rect 23660 35252 23716 37324
rect 23996 37044 24052 37324
rect 25564 37268 25620 38108
rect 27132 38612 27524 38668
rect 27804 40404 27860 40414
rect 26684 37826 26740 37838
rect 26684 37774 26686 37826
rect 26738 37774 26740 37826
rect 26460 37604 26516 37614
rect 25900 37492 25956 37502
rect 25900 37378 25956 37436
rect 25900 37326 25902 37378
rect 25954 37326 25956 37378
rect 25900 37314 25956 37326
rect 26460 37378 26516 37548
rect 26684 37492 26740 37774
rect 26684 37426 26740 37436
rect 26460 37326 26462 37378
rect 26514 37326 26516 37378
rect 26460 37314 26516 37326
rect 27020 37380 27076 37390
rect 27020 37286 27076 37324
rect 25676 37268 25732 37278
rect 25564 37266 25732 37268
rect 25564 37214 25678 37266
rect 25730 37214 25732 37266
rect 25564 37212 25732 37214
rect 25676 37202 25732 37212
rect 26684 37268 26740 37278
rect 24108 37154 24164 37166
rect 24108 37102 24110 37154
rect 24162 37102 24164 37154
rect 24108 37044 24164 37102
rect 23884 36988 24164 37044
rect 25340 37044 25396 37054
rect 26460 37044 26516 37054
rect 25340 37042 25620 37044
rect 25340 36990 25342 37042
rect 25394 36990 25620 37042
rect 25340 36988 25620 36990
rect 23884 35700 23940 36988
rect 25340 36978 25396 36988
rect 24008 36876 25208 36886
rect 24064 36874 24112 36876
rect 24168 36874 24216 36876
rect 24076 36822 24112 36874
rect 24200 36822 24216 36874
rect 24064 36820 24112 36822
rect 24168 36820 24216 36822
rect 24272 36874 24320 36876
rect 24376 36874 24424 36876
rect 24480 36874 24528 36876
rect 24376 36822 24396 36874
rect 24480 36822 24520 36874
rect 24272 36820 24320 36822
rect 24376 36820 24424 36822
rect 24480 36820 24528 36822
rect 24584 36820 24632 36876
rect 24688 36874 24736 36876
rect 24792 36874 24840 36876
rect 24896 36874 24944 36876
rect 24696 36822 24736 36874
rect 24820 36822 24840 36874
rect 24688 36820 24736 36822
rect 24792 36820 24840 36822
rect 24896 36820 24944 36822
rect 25000 36874 25048 36876
rect 25104 36874 25152 36876
rect 25000 36822 25016 36874
rect 25104 36822 25140 36874
rect 25000 36820 25048 36822
rect 25104 36820 25152 36822
rect 24008 36810 25208 36820
rect 24332 36482 24388 36494
rect 24332 36430 24334 36482
rect 24386 36430 24388 36482
rect 23996 35700 24052 35710
rect 24332 35700 24388 36430
rect 25340 35812 25396 35822
rect 25396 35756 25508 35812
rect 25340 35746 25396 35756
rect 23660 35186 23716 35196
rect 23772 35644 23996 35700
rect 24052 35644 24388 35700
rect 23548 34862 23550 34914
rect 23602 34862 23604 34914
rect 23548 34850 23604 34862
rect 22540 33460 22596 33470
rect 22540 33366 22596 33404
rect 22428 33124 22484 33134
rect 21756 32562 21812 32574
rect 21756 32510 21758 32562
rect 21810 32510 21812 32562
rect 21756 31892 21812 32510
rect 21756 31826 21812 31836
rect 22316 29540 22372 29550
rect 22316 29446 22372 29484
rect 20076 28756 20132 28766
rect 20076 28084 20132 28700
rect 21644 28754 21700 28812
rect 21644 28702 21646 28754
rect 21698 28702 21700 28754
rect 21644 28690 21700 28702
rect 21980 28756 22036 28766
rect 21980 28662 22036 28700
rect 20076 27858 20132 28028
rect 20076 27806 20078 27858
rect 20130 27806 20132 27858
rect 20076 27794 20132 27806
rect 20300 27970 20356 27982
rect 20300 27918 20302 27970
rect 20354 27918 20356 27970
rect 18844 27074 19908 27076
rect 18844 27022 18846 27074
rect 18898 27022 19908 27074
rect 18844 27020 19908 27022
rect 18844 27010 18900 27020
rect 18284 26852 18452 26908
rect 19852 26962 19908 27020
rect 19852 26910 19854 26962
rect 19906 26910 19908 26962
rect 18172 26290 18228 26302
rect 18172 26238 18174 26290
rect 18226 26238 18228 26290
rect 17388 23714 17444 23726
rect 17388 23662 17390 23714
rect 17442 23662 17444 23714
rect 17388 23044 17444 23662
rect 17836 23716 17892 23726
rect 17836 23622 17892 23660
rect 18172 23156 18228 26238
rect 18284 24612 18340 26852
rect 19292 26850 19348 26862
rect 19292 26798 19294 26850
rect 19346 26798 19348 26850
rect 18732 26292 18788 26302
rect 19292 26292 19348 26798
rect 18732 26290 19348 26292
rect 18732 26238 18734 26290
rect 18786 26238 19348 26290
rect 18732 26236 19348 26238
rect 18732 26226 18788 26236
rect 18732 24948 18788 24958
rect 18732 24854 18788 24892
rect 19516 24948 19572 24958
rect 19516 24722 19572 24892
rect 19516 24670 19518 24722
rect 19570 24670 19572 24722
rect 19516 24658 19572 24670
rect 19740 24834 19796 24846
rect 19740 24782 19742 24834
rect 19794 24782 19796 24834
rect 18284 23604 18340 24556
rect 19740 24612 19796 24782
rect 19740 24546 19796 24556
rect 19180 24500 19236 24510
rect 19180 24498 19460 24500
rect 19180 24446 19182 24498
rect 19234 24446 19460 24498
rect 19180 24444 19460 24446
rect 19180 24434 19236 24444
rect 19404 24276 19460 24444
rect 19404 24220 19684 24276
rect 19628 24162 19684 24220
rect 19628 24110 19630 24162
rect 19682 24110 19684 24162
rect 19628 24098 19684 24110
rect 18844 23828 18900 23838
rect 18844 23734 18900 23772
rect 19852 23828 19908 26910
rect 20300 25732 20356 27918
rect 20972 27860 21028 27870
rect 20972 27300 21028 27804
rect 20972 27234 21028 27244
rect 21420 27858 21476 27870
rect 21420 27806 21422 27858
rect 21474 27806 21476 27858
rect 20412 26962 20468 26974
rect 20412 26910 20414 26962
rect 20466 26910 20468 26962
rect 20412 26516 20468 26910
rect 20412 26450 20468 26460
rect 21196 26740 21252 26750
rect 21196 26514 21252 26684
rect 21420 26628 21476 27806
rect 22316 27300 22372 27310
rect 22204 27076 22260 27086
rect 22316 27076 22372 27244
rect 22204 27074 22372 27076
rect 22204 27022 22206 27074
rect 22258 27022 22372 27074
rect 22204 27020 22372 27022
rect 22204 27010 22260 27020
rect 21420 26562 21476 26572
rect 21980 26740 22036 26750
rect 21196 26462 21198 26514
rect 21250 26462 21252 26514
rect 21196 26450 21252 26462
rect 21756 26516 21812 26526
rect 21756 26422 21812 26460
rect 20300 25666 20356 25676
rect 20748 25732 20804 25742
rect 20300 24834 20356 24846
rect 20300 24782 20302 24834
rect 20354 24782 20356 24834
rect 19852 23734 19908 23772
rect 20188 24612 20244 24622
rect 19292 23716 19348 23726
rect 18284 23538 18340 23548
rect 18956 23714 19348 23716
rect 18956 23662 19294 23714
rect 19346 23662 19348 23714
rect 18956 23660 19348 23662
rect 18284 23156 18340 23166
rect 18172 23154 18340 23156
rect 18172 23102 18286 23154
rect 18338 23102 18340 23154
rect 18172 23100 18340 23102
rect 17500 23044 17556 23054
rect 17388 23042 17556 23044
rect 17388 22990 17502 23042
rect 17554 22990 17556 23042
rect 17388 22988 17556 22990
rect 18284 23044 18340 23100
rect 18732 23156 18788 23166
rect 18956 23156 19012 23660
rect 19292 23650 19348 23660
rect 18732 23154 19012 23156
rect 18732 23102 18734 23154
rect 18786 23102 19012 23154
rect 18732 23100 19012 23102
rect 18732 23090 18788 23100
rect 18396 23044 18452 23054
rect 18284 22988 18396 23044
rect 17500 22372 17556 22988
rect 18396 22978 18452 22988
rect 17500 22306 17556 22316
rect 20188 22260 20244 24556
rect 20300 22372 20356 24782
rect 20412 23828 20468 23838
rect 20412 23734 20468 23772
rect 20636 23716 20692 23726
rect 20412 22372 20468 22382
rect 20300 22316 20412 22372
rect 18508 22148 18564 22158
rect 19068 22148 19124 22158
rect 18508 22054 18564 22092
rect 18620 22146 19124 22148
rect 18620 22094 19070 22146
rect 19122 22094 19124 22146
rect 18620 22092 19124 22094
rect 17164 21812 17444 21868
rect 16716 21700 16772 21710
rect 16716 21606 16772 21644
rect 16604 20132 16660 21532
rect 16716 20916 16772 20926
rect 16716 20244 16772 20860
rect 16716 20188 16884 20244
rect 16604 20076 16772 20132
rect 16492 19954 16548 19964
rect 16604 19908 16660 19918
rect 16380 19740 16548 19796
rect 16268 16930 16324 16940
rect 16380 19012 16436 19022
rect 16380 16660 16436 18956
rect 16492 17444 16548 19740
rect 16604 18674 16660 19852
rect 16716 18900 16772 20076
rect 16828 19012 16884 20188
rect 17164 19012 17220 19022
rect 16828 19010 17220 19012
rect 16828 18958 17166 19010
rect 17218 18958 17220 19010
rect 16828 18956 17220 18958
rect 16716 18844 16884 18900
rect 16604 18622 16606 18674
rect 16658 18622 16660 18674
rect 16604 18610 16660 18622
rect 16716 18452 16772 18462
rect 16716 18358 16772 18396
rect 16604 18340 16660 18350
rect 16604 17666 16660 18284
rect 16604 17614 16606 17666
rect 16658 17614 16660 17666
rect 16604 17602 16660 17614
rect 16492 17388 16660 17444
rect 16492 17220 16548 17230
rect 16492 16994 16548 17164
rect 16492 16942 16494 16994
rect 16546 16942 16548 16994
rect 16492 16930 16548 16942
rect 16604 16996 16660 17388
rect 16604 16994 16772 16996
rect 16604 16942 16606 16994
rect 16658 16942 16772 16994
rect 16604 16940 16772 16942
rect 16604 16930 16660 16940
rect 16604 16660 16660 16670
rect 16380 16658 16660 16660
rect 16380 16606 16606 16658
rect 16658 16606 16660 16658
rect 16380 16604 16660 16606
rect 16604 16594 16660 16604
rect 16716 16100 16772 16940
rect 16716 14980 16772 16044
rect 16716 14914 16772 14924
rect 16044 13918 16046 13970
rect 16098 13918 16100 13970
rect 16044 13524 16100 13918
rect 16828 13970 16884 18844
rect 17164 18452 17220 18956
rect 17388 18676 17444 21812
rect 18620 21700 18676 22092
rect 19068 22082 19124 22092
rect 19404 22148 19460 22158
rect 20188 22148 20244 22204
rect 20300 22148 20356 22158
rect 20188 22146 20356 22148
rect 20188 22094 20302 22146
rect 20354 22094 20356 22146
rect 20188 22092 20356 22094
rect 19404 22054 19460 22092
rect 20300 22082 20356 22092
rect 17500 21588 17556 21598
rect 17500 21494 17556 21532
rect 18284 20132 18340 20142
rect 18340 20076 18452 20132
rect 18284 20038 18340 20076
rect 18060 19012 18116 19022
rect 17388 18620 17556 18676
rect 17388 18452 17444 18462
rect 17164 18450 17444 18452
rect 17164 18398 17390 18450
rect 17442 18398 17444 18450
rect 17164 18396 17444 18398
rect 17052 17668 17108 17678
rect 17388 17668 17444 18396
rect 17052 17666 17444 17668
rect 17052 17614 17054 17666
rect 17106 17614 17444 17666
rect 17052 17612 17444 17614
rect 17052 16884 17108 17612
rect 17052 16818 17108 16828
rect 17164 15874 17220 15886
rect 17164 15822 17166 15874
rect 17218 15822 17220 15874
rect 17164 14756 17220 15822
rect 17164 14690 17220 14700
rect 17500 14644 17556 18620
rect 18060 18450 18116 18956
rect 18396 18564 18452 20076
rect 18620 20130 18676 21644
rect 20412 21026 20468 22316
rect 20412 20974 20414 21026
rect 20466 20974 20468 21026
rect 20412 20962 20468 20974
rect 20524 20578 20580 20590
rect 20524 20526 20526 20578
rect 20578 20526 20580 20578
rect 18620 20078 18622 20130
rect 18674 20078 18676 20130
rect 18620 20066 18676 20078
rect 18732 20132 18788 20142
rect 18732 20038 18788 20076
rect 20300 20132 20356 20142
rect 18956 20020 19012 20030
rect 18956 20018 19236 20020
rect 18956 19966 18958 20018
rect 19010 19966 19236 20018
rect 18956 19964 19236 19966
rect 18956 19954 19012 19964
rect 18844 19234 18900 19246
rect 18844 19182 18846 19234
rect 18898 19182 18900 19234
rect 18508 19124 18564 19134
rect 18844 19124 18900 19182
rect 18956 19236 19012 19246
rect 18956 19142 19012 19180
rect 18564 19068 18900 19124
rect 18508 19058 18564 19068
rect 18396 18508 18564 18564
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 18060 18386 18116 18398
rect 17948 17780 18004 17790
rect 17948 17686 18004 17724
rect 18172 17554 18228 17566
rect 18172 17502 18174 17554
rect 18226 17502 18228 17554
rect 17612 17444 17668 17454
rect 18060 17444 18116 17454
rect 17612 17442 17892 17444
rect 17612 17390 17614 17442
rect 17666 17390 17892 17442
rect 17612 17388 17892 17390
rect 17612 17378 17668 17388
rect 17612 16884 17668 16894
rect 17612 16790 17668 16828
rect 17612 16100 17668 16110
rect 17612 16006 17668 16044
rect 17612 14644 17668 14654
rect 17500 14642 17668 14644
rect 17500 14590 17614 14642
rect 17666 14590 17668 14642
rect 17500 14588 17668 14590
rect 17612 14420 17668 14588
rect 17612 14354 17668 14364
rect 16828 13918 16830 13970
rect 16882 13918 16884 13970
rect 16828 13860 16884 13918
rect 16828 13794 16884 13804
rect 17836 13746 17892 17388
rect 18060 16770 18116 17388
rect 18060 16718 18062 16770
rect 18114 16718 18116 16770
rect 18060 15988 18116 16718
rect 18060 15922 18116 15932
rect 18172 16996 18228 17502
rect 18508 17444 18564 18508
rect 18620 17556 18676 17566
rect 18620 17462 18676 17500
rect 18508 17378 18564 17388
rect 18844 17332 18900 19068
rect 19180 19122 19236 19964
rect 19180 19070 19182 19122
rect 19234 19070 19236 19122
rect 19180 19058 19236 19070
rect 19516 19124 19572 19134
rect 19516 19030 19572 19068
rect 19740 19122 19796 19134
rect 20188 19124 20244 19134
rect 19740 19070 19742 19122
rect 19794 19070 19796 19122
rect 19628 19012 19684 19022
rect 19628 18918 19684 18956
rect 19740 18452 19796 19070
rect 19628 18396 19796 18452
rect 19852 19122 20244 19124
rect 19852 19070 20190 19122
rect 20242 19070 20244 19122
rect 19852 19068 20244 19070
rect 19292 18228 19348 18238
rect 19292 17666 19348 18172
rect 19292 17614 19294 17666
rect 19346 17614 19348 17666
rect 19292 17556 19348 17614
rect 19404 17668 19460 17678
rect 19628 17668 19684 18396
rect 19852 18340 19908 19068
rect 20188 19058 20244 19068
rect 20300 19124 20356 20076
rect 20524 19460 20580 20526
rect 20524 19394 20580 19404
rect 20524 19236 20580 19246
rect 20524 19142 20580 19180
rect 20300 18788 20356 19068
rect 19740 18284 19908 18340
rect 20076 18732 20356 18788
rect 19740 17778 19796 18284
rect 19740 17726 19742 17778
rect 19794 17726 19796 17778
rect 19740 17714 19796 17726
rect 19460 17612 19684 17668
rect 19404 17574 19460 17612
rect 19292 17490 19348 17500
rect 18844 17276 19460 17332
rect 18508 17220 18564 17230
rect 18508 17106 18564 17164
rect 18508 17054 18510 17106
rect 18562 17054 18564 17106
rect 18508 17042 18564 17054
rect 18172 14756 18228 16940
rect 19292 16772 19348 16782
rect 19180 16716 19292 16772
rect 18732 15316 18788 15326
rect 18732 15222 18788 15260
rect 19180 15314 19236 16716
rect 19292 16706 19348 16716
rect 19404 16770 19460 17276
rect 20076 17108 20132 18732
rect 20524 18676 20580 18686
rect 20636 18676 20692 23660
rect 20748 20916 20804 25676
rect 21980 25618 22036 26684
rect 22092 26516 22148 26526
rect 22092 26402 22148 26460
rect 22092 26350 22094 26402
rect 22146 26350 22148 26402
rect 22092 26338 22148 26350
rect 21980 25566 21982 25618
rect 22034 25566 22036 25618
rect 21980 25554 22036 25566
rect 21420 25284 21476 25294
rect 21420 23716 21476 25228
rect 22316 25284 22372 27020
rect 22428 26908 22484 33068
rect 22988 33122 23044 33134
rect 22988 33070 22990 33122
rect 23042 33070 23044 33122
rect 22988 32676 23044 33070
rect 23436 32788 23492 33516
rect 23436 32722 23492 32732
rect 23548 33122 23604 33134
rect 23548 33070 23550 33122
rect 23602 33070 23604 33122
rect 22988 32610 23044 32620
rect 23548 32452 23604 33070
rect 23324 32396 23604 32452
rect 23660 32676 23716 32686
rect 22988 31892 23044 31902
rect 22988 31798 23044 31836
rect 23324 31890 23380 32396
rect 23660 31948 23716 32620
rect 23324 31838 23326 31890
rect 23378 31838 23380 31890
rect 23324 31826 23380 31838
rect 23436 31892 23716 31948
rect 22540 31780 22596 31790
rect 22540 31686 22596 31724
rect 23212 30324 23268 30334
rect 23100 29428 23156 29438
rect 22652 29426 23156 29428
rect 22652 29374 23102 29426
rect 23154 29374 23156 29426
rect 22652 29372 23156 29374
rect 22652 28866 22708 29372
rect 23100 29362 23156 29372
rect 22652 28814 22654 28866
rect 22706 28814 22708 28866
rect 22652 28802 22708 28814
rect 22764 29202 22820 29214
rect 22764 29150 22766 29202
rect 22818 29150 22820 29202
rect 22652 27076 22708 27086
rect 22764 27076 22820 29150
rect 22988 28868 23044 28878
rect 22988 28774 23044 28812
rect 23212 27972 23268 30268
rect 23324 29540 23380 29550
rect 23324 29446 23380 29484
rect 23436 28756 23492 31892
rect 23436 28642 23492 28700
rect 23436 28590 23438 28642
rect 23490 28590 23492 28642
rect 23436 28578 23492 28590
rect 22652 27074 22820 27076
rect 22652 27022 22654 27074
rect 22706 27022 22820 27074
rect 22652 27020 22820 27022
rect 22988 27916 23268 27972
rect 23548 28530 23604 28542
rect 23548 28478 23550 28530
rect 23602 28478 23604 28530
rect 22652 27010 22708 27020
rect 22428 26852 22708 26908
rect 22652 26402 22708 26852
rect 22652 26350 22654 26402
rect 22706 26350 22708 26402
rect 22652 26180 22708 26350
rect 22652 26114 22708 26124
rect 22316 25190 22372 25228
rect 22876 26066 22932 26078
rect 22876 26014 22878 26066
rect 22930 26014 22932 26066
rect 22876 24052 22932 26014
rect 22876 23986 22932 23996
rect 21308 23714 21476 23716
rect 21308 23662 21422 23714
rect 21474 23662 21476 23714
rect 21308 23660 21476 23662
rect 20972 23380 21028 23390
rect 20972 23266 21028 23324
rect 20972 23214 20974 23266
rect 21026 23214 21028 23266
rect 20860 22484 20916 22494
rect 20860 22390 20916 22428
rect 20972 22148 21028 23214
rect 20972 22082 21028 22092
rect 21308 23044 21364 23660
rect 21420 23650 21476 23660
rect 21756 23828 21812 23838
rect 21756 23378 21812 23772
rect 22764 23828 22820 23838
rect 22764 23734 22820 23772
rect 21756 23326 21758 23378
rect 21810 23326 21812 23378
rect 21756 23314 21812 23326
rect 21868 23714 21924 23726
rect 21868 23662 21870 23714
rect 21922 23662 21924 23714
rect 21868 23380 21924 23662
rect 22428 23714 22484 23726
rect 22428 23662 22430 23714
rect 22482 23662 22484 23714
rect 22428 23604 22484 23662
rect 22876 23716 22932 23726
rect 22988 23716 23044 27916
rect 23548 27748 23604 28478
rect 23212 26628 23268 26638
rect 23212 26514 23268 26572
rect 23212 26462 23214 26514
rect 23266 26462 23268 26514
rect 23212 26450 23268 26462
rect 23436 25284 23492 25294
rect 23100 24500 23156 24510
rect 23100 23938 23156 24444
rect 23100 23886 23102 23938
rect 23154 23886 23156 23938
rect 23100 23874 23156 23886
rect 22876 23714 23044 23716
rect 22876 23662 22878 23714
rect 22930 23662 23044 23714
rect 22876 23660 23044 23662
rect 22876 23604 22932 23660
rect 22428 23548 22932 23604
rect 21868 23314 21924 23324
rect 23436 23380 23492 25228
rect 23436 23314 23492 23324
rect 21980 23268 22036 23278
rect 21980 23154 22036 23212
rect 21980 23102 21982 23154
rect 22034 23102 22036 23154
rect 21980 23090 22036 23102
rect 20748 20802 20804 20860
rect 20748 20750 20750 20802
rect 20802 20750 20804 20802
rect 20748 20738 20804 20750
rect 21308 21586 21364 22988
rect 21756 22484 21812 22494
rect 21756 22390 21812 22428
rect 23100 22372 23156 22382
rect 23100 22278 23156 22316
rect 21980 22260 22036 22270
rect 21980 22166 22036 22204
rect 22540 22258 22596 22270
rect 22540 22206 22542 22258
rect 22594 22206 22596 22258
rect 21308 21534 21310 21586
rect 21362 21534 21364 21586
rect 21308 20580 21364 21534
rect 21420 22146 21476 22158
rect 21420 22094 21422 22146
rect 21474 22094 21476 22146
rect 21420 21028 21476 22094
rect 21420 20962 21476 20972
rect 21532 21588 21588 21598
rect 21420 20804 21476 20814
rect 21532 20804 21588 21532
rect 21756 21588 21812 21598
rect 21756 21586 21924 21588
rect 21756 21534 21758 21586
rect 21810 21534 21924 21586
rect 21756 21532 21924 21534
rect 21756 21522 21812 21532
rect 21868 21026 21924 21532
rect 21868 20974 21870 21026
rect 21922 20974 21924 21026
rect 21868 20962 21924 20974
rect 22204 21028 22260 21038
rect 22204 20934 22260 20972
rect 21420 20802 21532 20804
rect 21420 20750 21422 20802
rect 21474 20750 21532 20802
rect 21420 20748 21532 20750
rect 21420 20738 21476 20748
rect 21532 20710 21588 20748
rect 22428 20804 22484 20814
rect 22428 20690 22484 20748
rect 22428 20638 22430 20690
rect 22482 20638 22484 20690
rect 22428 20626 22484 20638
rect 21308 20524 21476 20580
rect 21420 19796 21476 20524
rect 22540 20020 22596 22206
rect 23212 22146 23268 22158
rect 23212 22094 23214 22146
rect 23266 22094 23268 22146
rect 22988 21364 23044 21374
rect 22988 20690 23044 21308
rect 23212 20804 23268 22094
rect 23324 22148 23380 22158
rect 23324 21588 23380 22092
rect 23436 22146 23492 22158
rect 23436 22094 23438 22146
rect 23490 22094 23492 22146
rect 23436 22036 23492 22094
rect 23436 21970 23492 21980
rect 23548 21812 23604 27692
rect 23660 28084 23716 28094
rect 23660 26740 23716 28028
rect 23772 26908 23828 35644
rect 23996 35606 24052 35644
rect 24444 35588 24500 35598
rect 24444 35494 24500 35532
rect 25340 35476 25396 35486
rect 25340 35382 25396 35420
rect 24008 35308 25208 35318
rect 24064 35306 24112 35308
rect 24168 35306 24216 35308
rect 24076 35254 24112 35306
rect 24200 35254 24216 35306
rect 24064 35252 24112 35254
rect 24168 35252 24216 35254
rect 24272 35306 24320 35308
rect 24376 35306 24424 35308
rect 24480 35306 24528 35308
rect 24376 35254 24396 35306
rect 24480 35254 24520 35306
rect 24272 35252 24320 35254
rect 24376 35252 24424 35254
rect 24480 35252 24528 35254
rect 24584 35252 24632 35308
rect 24688 35306 24736 35308
rect 24792 35306 24840 35308
rect 24896 35306 24944 35308
rect 24696 35254 24736 35306
rect 24820 35254 24840 35306
rect 24688 35252 24736 35254
rect 24792 35252 24840 35254
rect 24896 35252 24944 35254
rect 25000 35306 25048 35308
rect 25104 35306 25152 35308
rect 25000 35254 25016 35306
rect 25104 35254 25140 35306
rect 25000 35252 25048 35254
rect 25104 35252 25152 35254
rect 24008 35242 25208 35252
rect 25452 34804 25508 35756
rect 25564 35700 25620 36988
rect 25900 35812 25956 35822
rect 25900 35718 25956 35756
rect 26460 35812 26516 36988
rect 26684 36594 26740 37212
rect 26684 36542 26686 36594
rect 26738 36542 26740 36594
rect 26684 36530 26740 36542
rect 26908 37268 26964 37278
rect 26460 35810 26628 35812
rect 26460 35758 26462 35810
rect 26514 35758 26628 35810
rect 26460 35756 26628 35758
rect 26460 35746 26516 35756
rect 25676 35700 25732 35710
rect 25564 35698 25732 35700
rect 25564 35646 25678 35698
rect 25730 35646 25732 35698
rect 25564 35644 25732 35646
rect 25676 35634 25732 35644
rect 26572 35138 26628 35756
rect 26572 35086 26574 35138
rect 26626 35086 26628 35138
rect 26572 35074 26628 35086
rect 26684 35476 26740 35486
rect 26012 34916 26068 34926
rect 25340 34748 25508 34804
rect 25788 34804 25844 34814
rect 25340 34354 25396 34748
rect 25788 34710 25844 34748
rect 25340 34302 25342 34354
rect 25394 34302 25396 34354
rect 24008 33740 25208 33750
rect 24064 33738 24112 33740
rect 24168 33738 24216 33740
rect 24076 33686 24112 33738
rect 24200 33686 24216 33738
rect 24064 33684 24112 33686
rect 24168 33684 24216 33686
rect 24272 33738 24320 33740
rect 24376 33738 24424 33740
rect 24480 33738 24528 33740
rect 24376 33686 24396 33738
rect 24480 33686 24520 33738
rect 24272 33684 24320 33686
rect 24376 33684 24424 33686
rect 24480 33684 24528 33686
rect 24584 33684 24632 33740
rect 24688 33738 24736 33740
rect 24792 33738 24840 33740
rect 24896 33738 24944 33740
rect 24696 33686 24736 33738
rect 24820 33686 24840 33738
rect 24688 33684 24736 33686
rect 24792 33684 24840 33686
rect 24896 33684 24944 33686
rect 25000 33738 25048 33740
rect 25104 33738 25152 33740
rect 25000 33686 25016 33738
rect 25104 33686 25140 33738
rect 25000 33684 25048 33686
rect 25104 33684 25152 33686
rect 24008 33674 25208 33684
rect 23996 33572 24052 33582
rect 23884 33460 23940 33470
rect 23884 33366 23940 33404
rect 23996 32900 24052 33516
rect 23996 32786 24052 32844
rect 23996 32734 23998 32786
rect 24050 32734 24052 32786
rect 23996 32722 24052 32734
rect 24444 33346 24500 33358
rect 24444 33294 24446 33346
rect 24498 33294 24500 33346
rect 24444 32676 24500 33294
rect 24668 33234 24724 33246
rect 24668 33182 24670 33234
rect 24722 33182 24724 33234
rect 24668 33124 24724 33182
rect 24668 33058 24724 33068
rect 25228 33124 25284 33134
rect 25340 33124 25396 34302
rect 25452 34580 25508 34590
rect 25452 33460 25508 34524
rect 26012 34132 26068 34860
rect 25452 33394 25508 33404
rect 25676 34130 26068 34132
rect 25676 34078 26014 34130
rect 26066 34078 26068 34130
rect 25676 34076 26068 34078
rect 25340 33068 25508 33124
rect 25228 33030 25284 33068
rect 24444 32610 24500 32620
rect 25340 32900 25396 32910
rect 25340 32786 25396 32844
rect 25340 32734 25342 32786
rect 25394 32734 25396 32786
rect 23884 32340 23940 32350
rect 23884 31666 23940 32284
rect 24780 32340 24836 32378
rect 24780 32274 24836 32284
rect 24008 32172 25208 32182
rect 24064 32170 24112 32172
rect 24168 32170 24216 32172
rect 24076 32118 24112 32170
rect 24200 32118 24216 32170
rect 24064 32116 24112 32118
rect 24168 32116 24216 32118
rect 24272 32170 24320 32172
rect 24376 32170 24424 32172
rect 24480 32170 24528 32172
rect 24376 32118 24396 32170
rect 24480 32118 24520 32170
rect 24272 32116 24320 32118
rect 24376 32116 24424 32118
rect 24480 32116 24528 32118
rect 24584 32116 24632 32172
rect 24688 32170 24736 32172
rect 24792 32170 24840 32172
rect 24896 32170 24944 32172
rect 24696 32118 24736 32170
rect 24820 32118 24840 32170
rect 24688 32116 24736 32118
rect 24792 32116 24840 32118
rect 24896 32116 24944 32118
rect 25000 32170 25048 32172
rect 25104 32170 25152 32172
rect 25000 32118 25016 32170
rect 25104 32118 25140 32170
rect 25000 32116 25048 32118
rect 25104 32116 25152 32118
rect 24008 32106 25208 32116
rect 23996 31892 24052 31902
rect 23996 31778 24052 31836
rect 23996 31726 23998 31778
rect 24050 31726 24052 31778
rect 23996 31714 24052 31726
rect 23884 31614 23886 31666
rect 23938 31614 23940 31666
rect 23884 31602 23940 31614
rect 24008 30604 25208 30614
rect 24064 30602 24112 30604
rect 24168 30602 24216 30604
rect 24076 30550 24112 30602
rect 24200 30550 24216 30602
rect 24064 30548 24112 30550
rect 24168 30548 24216 30550
rect 24272 30602 24320 30604
rect 24376 30602 24424 30604
rect 24480 30602 24528 30604
rect 24376 30550 24396 30602
rect 24480 30550 24520 30602
rect 24272 30548 24320 30550
rect 24376 30548 24424 30550
rect 24480 30548 24528 30550
rect 24584 30548 24632 30604
rect 24688 30602 24736 30604
rect 24792 30602 24840 30604
rect 24896 30602 24944 30604
rect 24696 30550 24736 30602
rect 24820 30550 24840 30602
rect 24688 30548 24736 30550
rect 24792 30548 24840 30550
rect 24896 30548 24944 30550
rect 25000 30602 25048 30604
rect 25104 30602 25152 30604
rect 25000 30550 25016 30602
rect 25104 30550 25140 30602
rect 25000 30548 25048 30550
rect 25104 30548 25152 30550
rect 24008 30538 25208 30548
rect 25340 30212 25396 32734
rect 23884 29538 23940 29550
rect 23884 29486 23886 29538
rect 23938 29486 23940 29538
rect 23884 27860 23940 29486
rect 24008 29036 25208 29046
rect 24064 29034 24112 29036
rect 24168 29034 24216 29036
rect 24076 28982 24112 29034
rect 24200 28982 24216 29034
rect 24064 28980 24112 28982
rect 24168 28980 24216 28982
rect 24272 29034 24320 29036
rect 24376 29034 24424 29036
rect 24480 29034 24528 29036
rect 24376 28982 24396 29034
rect 24480 28982 24520 29034
rect 24272 28980 24320 28982
rect 24376 28980 24424 28982
rect 24480 28980 24528 28982
rect 24584 28980 24632 29036
rect 24688 29034 24736 29036
rect 24792 29034 24840 29036
rect 24896 29034 24944 29036
rect 24696 28982 24736 29034
rect 24820 28982 24840 29034
rect 24688 28980 24736 28982
rect 24792 28980 24840 28982
rect 24896 28980 24944 28982
rect 25000 29034 25048 29036
rect 25104 29034 25152 29036
rect 25000 28982 25016 29034
rect 25104 28982 25140 29034
rect 25000 28980 25048 28982
rect 25104 28980 25152 28982
rect 24008 28970 25208 28980
rect 23884 27794 23940 27804
rect 25340 28084 25396 30156
rect 25452 31892 25508 33068
rect 25452 29988 25508 31836
rect 25564 31668 25620 31678
rect 25564 31574 25620 31612
rect 25564 30996 25620 31006
rect 25676 30996 25732 34076
rect 26012 34066 26068 34076
rect 26684 34130 26740 35420
rect 26908 34916 26964 37212
rect 27020 36484 27076 36494
rect 27020 35026 27076 36428
rect 27020 34974 27022 35026
rect 27074 34974 27076 35026
rect 27020 34962 27076 34974
rect 26908 34850 26964 34860
rect 27132 34692 27188 38612
rect 27580 37828 27636 37838
rect 27580 37380 27636 37772
rect 27804 37828 27860 40348
rect 29484 39732 29540 41244
rect 29708 41206 29764 41244
rect 29484 39638 29540 39676
rect 29820 39730 29876 41358
rect 29932 42530 29988 42542
rect 29932 42478 29934 42530
rect 29986 42478 29988 42530
rect 29932 42194 29988 42478
rect 29932 42142 29934 42194
rect 29986 42142 29988 42194
rect 29932 41972 29988 42142
rect 29932 40740 29988 41916
rect 29932 40674 29988 40684
rect 29932 40404 29988 40414
rect 30044 40404 30100 44940
rect 30268 43762 30324 44940
rect 30604 44930 30660 44940
rect 30716 43764 30772 46844
rect 31164 46834 31220 46844
rect 31388 46900 31444 46910
rect 31500 46900 31556 47404
rect 31724 47460 31780 47470
rect 31948 47460 32004 48748
rect 32284 48916 32340 49644
rect 32508 49698 32564 49710
rect 32508 49646 32510 49698
rect 32562 49646 32564 49698
rect 32508 49586 32564 49646
rect 32508 49534 32510 49586
rect 32562 49534 32564 49586
rect 32508 49522 32564 49534
rect 31724 47458 32004 47460
rect 31724 47406 31726 47458
rect 31778 47406 32004 47458
rect 31724 47404 32004 47406
rect 31724 47394 31780 47404
rect 31388 46898 31556 46900
rect 31388 46846 31390 46898
rect 31442 46846 31556 46898
rect 31388 46844 31556 46846
rect 31612 46900 31668 46910
rect 31388 46834 31444 46844
rect 31612 46786 31668 46844
rect 31612 46734 31614 46786
rect 31666 46734 31668 46786
rect 31612 46722 31668 46734
rect 30940 46674 30996 46686
rect 30940 46622 30942 46674
rect 30994 46622 30996 46674
rect 30940 46116 30996 46622
rect 30940 46050 30996 46060
rect 31276 46562 31332 46574
rect 31276 46510 31278 46562
rect 31330 46510 31332 46562
rect 31052 45892 31108 45902
rect 31052 45890 31220 45892
rect 31052 45838 31054 45890
rect 31106 45838 31220 45890
rect 31052 45836 31220 45838
rect 31052 45826 31108 45836
rect 31164 45330 31220 45836
rect 31164 45278 31166 45330
rect 31218 45278 31220 45330
rect 31164 45266 31220 45278
rect 30828 45108 30884 45118
rect 31276 45108 31332 46510
rect 31948 46564 32004 47404
rect 31948 46498 32004 46508
rect 32060 48244 32116 48254
rect 30828 45106 31332 45108
rect 30828 45054 30830 45106
rect 30882 45054 31332 45106
rect 30828 45052 31332 45054
rect 30828 45042 30884 45052
rect 30268 43710 30270 43762
rect 30322 43710 30324 43762
rect 30268 43698 30324 43710
rect 30492 43708 30772 43764
rect 30492 43652 30548 43708
rect 30156 43540 30212 43550
rect 30156 42532 30212 43484
rect 30492 43538 30548 43596
rect 30492 43486 30494 43538
rect 30546 43486 30548 43538
rect 30492 43474 30548 43486
rect 30940 43428 30996 43438
rect 30940 43334 30996 43372
rect 31724 43426 31780 43438
rect 31724 43374 31726 43426
rect 31778 43374 31780 43426
rect 30268 42868 30324 42878
rect 30268 42774 30324 42812
rect 30156 42466 30212 42476
rect 30492 42756 30548 42766
rect 30492 42196 30548 42700
rect 30828 42754 30884 42766
rect 30828 42702 30830 42754
rect 30882 42702 30884 42754
rect 30828 42196 30884 42702
rect 31052 42756 31108 42766
rect 31388 42756 31444 42766
rect 31052 42754 31444 42756
rect 31052 42702 31054 42754
rect 31106 42702 31390 42754
rect 31442 42702 31444 42754
rect 31052 42700 31444 42702
rect 31052 42690 31108 42700
rect 30492 42194 30772 42196
rect 30492 42142 30494 42194
rect 30546 42142 30772 42194
rect 30492 42140 30772 42142
rect 30492 42130 30548 42140
rect 30268 41972 30324 41982
rect 30268 41300 30324 41916
rect 30716 41636 30772 42140
rect 30828 42130 30884 42140
rect 31276 42532 31332 42542
rect 31052 41972 31108 41982
rect 31052 41878 31108 41916
rect 30716 41580 31108 41636
rect 30828 41412 30884 41422
rect 30604 41300 30660 41310
rect 30324 41244 30436 41300
rect 30268 41206 30324 41244
rect 30268 40628 30324 40638
rect 29988 40348 30100 40404
rect 30156 40516 30212 40526
rect 29932 40338 29988 40348
rect 30044 40180 30100 40190
rect 30156 40180 30212 40460
rect 30044 40178 30212 40180
rect 30044 40126 30046 40178
rect 30098 40126 30212 40178
rect 30044 40124 30212 40126
rect 30044 40114 30100 40124
rect 29820 39678 29822 39730
rect 29874 39678 29876 39730
rect 28252 39620 28308 39630
rect 27804 37826 27972 37828
rect 27804 37774 27806 37826
rect 27858 37774 27972 37826
rect 27804 37772 27972 37774
rect 27804 37762 27860 37772
rect 27580 37286 27636 37324
rect 27356 37266 27412 37278
rect 27356 37214 27358 37266
rect 27410 37214 27412 37266
rect 27356 37044 27412 37214
rect 27804 37266 27860 37278
rect 27804 37214 27806 37266
rect 27858 37214 27860 37266
rect 27356 36978 27412 36988
rect 27692 37154 27748 37166
rect 27692 37102 27694 37154
rect 27746 37102 27748 37154
rect 27692 36708 27748 37102
rect 27804 37044 27860 37214
rect 27916 37268 27972 37772
rect 28252 37826 28308 39564
rect 28252 37774 28254 37826
rect 28306 37774 28308 37826
rect 28028 37604 28084 37614
rect 28028 37378 28084 37548
rect 28252 37492 28308 37774
rect 28252 37426 28308 37436
rect 28028 37326 28030 37378
rect 28082 37326 28084 37378
rect 28028 37314 28084 37326
rect 27916 37202 27972 37212
rect 28252 37268 28308 37278
rect 28252 37174 28308 37212
rect 28924 37268 28980 37278
rect 28924 37266 29652 37268
rect 28924 37214 28926 37266
rect 28978 37214 29652 37266
rect 28924 37212 29652 37214
rect 28924 37202 28980 37212
rect 27804 36978 27860 36988
rect 28028 37156 28084 37166
rect 27692 36642 27748 36652
rect 27692 36484 27748 36494
rect 27692 36390 27748 36428
rect 28028 36370 28084 37100
rect 29484 37044 29540 37054
rect 29036 36708 29092 36718
rect 29036 36482 29092 36652
rect 29036 36430 29038 36482
rect 29090 36430 29092 36482
rect 29036 36418 29092 36430
rect 29484 36482 29540 36988
rect 29596 36594 29652 37212
rect 29820 37044 29876 39678
rect 30156 39732 30212 39742
rect 30156 39618 30212 39676
rect 30268 39730 30324 40572
rect 30268 39678 30270 39730
rect 30322 39678 30324 39730
rect 30268 39666 30324 39678
rect 30156 39566 30158 39618
rect 30210 39566 30212 39618
rect 30156 39554 30212 39566
rect 30380 39508 30436 41244
rect 30604 41206 30660 41244
rect 30716 41188 30772 41198
rect 30716 41094 30772 41132
rect 30604 40740 30660 40750
rect 30604 40402 30660 40684
rect 30604 40350 30606 40402
rect 30658 40350 30660 40402
rect 29820 36978 29876 36988
rect 30268 39452 30436 39508
rect 30492 39732 30548 39742
rect 29596 36542 29598 36594
rect 29650 36542 29652 36594
rect 29596 36530 29652 36542
rect 30268 36484 30324 39452
rect 30492 37828 30548 39676
rect 30492 37762 30548 37772
rect 30604 37492 30660 40350
rect 30828 38668 30884 41356
rect 31052 40516 31108 41580
rect 31276 41076 31332 42476
rect 31388 41860 31444 42700
rect 31724 42532 31780 43374
rect 31948 43314 32004 43326
rect 31948 43262 31950 43314
rect 32002 43262 32004 43314
rect 31948 42868 32004 43262
rect 31724 42466 31780 42476
rect 31836 42812 32004 42868
rect 31836 42420 31892 42812
rect 31836 42364 32004 42420
rect 31724 41860 31780 41870
rect 31388 41858 31780 41860
rect 31388 41806 31726 41858
rect 31778 41806 31780 41858
rect 31388 41804 31780 41806
rect 31612 41410 31668 41804
rect 31724 41794 31780 41804
rect 31612 41358 31614 41410
rect 31666 41358 31668 41410
rect 31612 41346 31668 41358
rect 31724 41636 31780 41646
rect 31948 41636 32004 42364
rect 32060 42082 32116 48188
rect 32172 48018 32228 48030
rect 32172 47966 32174 48018
rect 32226 47966 32228 48018
rect 32172 47460 32228 47966
rect 32172 47394 32228 47404
rect 32172 47236 32228 47246
rect 32172 47142 32228 47180
rect 32172 46900 32228 46910
rect 32172 46806 32228 46844
rect 32284 46674 32340 48860
rect 32508 48466 32564 48478
rect 32508 48414 32510 48466
rect 32562 48414 32564 48466
rect 32508 48244 32564 48414
rect 32508 48178 32564 48188
rect 32396 48018 32452 48030
rect 32396 47966 32398 48018
rect 32450 47966 32452 48018
rect 32396 46788 32452 47966
rect 32396 46722 32452 46732
rect 32620 47458 32676 51324
rect 32620 47406 32622 47458
rect 32674 47406 32676 47458
rect 32284 46622 32286 46674
rect 32338 46622 32340 46674
rect 32284 46340 32340 46622
rect 32620 46676 32676 47406
rect 32732 47012 32788 56590
rect 33628 56420 33684 57820
rect 33740 57810 33796 57820
rect 34076 57652 34132 57662
rect 34188 57652 34244 57820
rect 34356 57820 34804 57876
rect 34300 57782 34356 57820
rect 34636 57652 34692 57662
rect 34188 57650 34692 57652
rect 34188 57598 34638 57650
rect 34690 57598 34692 57650
rect 34188 57596 34692 57598
rect 34076 57558 34132 57596
rect 34636 57586 34692 57596
rect 34412 57428 34468 57438
rect 34412 57426 34692 57428
rect 34412 57374 34414 57426
rect 34466 57374 34692 57426
rect 34412 57372 34692 57374
rect 34412 57362 34468 57372
rect 33292 56364 33684 56420
rect 33740 56812 34468 56868
rect 33292 56084 33348 56364
rect 33292 55990 33348 56028
rect 33628 56084 33684 56094
rect 33628 54402 33684 56028
rect 33740 56082 33796 56812
rect 33852 56644 33908 56654
rect 33852 56550 33908 56588
rect 34300 56644 34356 56682
rect 34412 56644 34468 56812
rect 34636 56866 34692 57372
rect 34748 56980 34804 57820
rect 35196 57820 35364 57876
rect 34860 57316 34916 57326
rect 34860 57090 34916 57260
rect 34860 57038 34862 57090
rect 34914 57038 34916 57090
rect 34860 57026 34916 57038
rect 35196 56980 35252 57820
rect 35308 57650 35364 57662
rect 35308 57598 35310 57650
rect 35362 57598 35364 57650
rect 35308 57092 35364 57598
rect 35532 57316 35588 58268
rect 36876 58324 36932 58382
rect 35532 57250 35588 57260
rect 36428 58212 36484 58222
rect 35868 57092 35924 57102
rect 35308 57090 35924 57092
rect 35308 57038 35870 57090
rect 35922 57038 35924 57090
rect 35308 57036 35924 57038
rect 35868 57026 35924 57036
rect 36204 57092 36260 57102
rect 36204 56998 36260 57036
rect 35196 56924 35364 56980
rect 34748 56914 34804 56924
rect 34636 56814 34638 56866
rect 34690 56814 34692 56866
rect 34636 56802 34692 56814
rect 35084 56866 35140 56878
rect 35084 56814 35086 56866
rect 35138 56814 35140 56866
rect 34748 56644 34804 56654
rect 34412 56642 34804 56644
rect 34412 56590 34750 56642
rect 34802 56590 34804 56642
rect 34412 56588 34804 56590
rect 34300 56578 34356 56588
rect 34748 56578 34804 56588
rect 35084 56644 35140 56814
rect 35084 56578 35140 56588
rect 34008 56476 35208 56486
rect 34064 56474 34112 56476
rect 34168 56474 34216 56476
rect 34076 56422 34112 56474
rect 34200 56422 34216 56474
rect 34064 56420 34112 56422
rect 34168 56420 34216 56422
rect 34272 56474 34320 56476
rect 34376 56474 34424 56476
rect 34480 56474 34528 56476
rect 34376 56422 34396 56474
rect 34480 56422 34520 56474
rect 34272 56420 34320 56422
rect 34376 56420 34424 56422
rect 34480 56420 34528 56422
rect 34584 56420 34632 56476
rect 34688 56474 34736 56476
rect 34792 56474 34840 56476
rect 34896 56474 34944 56476
rect 34696 56422 34736 56474
rect 34820 56422 34840 56474
rect 34688 56420 34736 56422
rect 34792 56420 34840 56422
rect 34896 56420 34944 56422
rect 35000 56474 35048 56476
rect 35104 56474 35152 56476
rect 35000 56422 35016 56474
rect 35104 56422 35140 56474
rect 35000 56420 35048 56422
rect 35104 56420 35152 56422
rect 34008 56410 35208 56420
rect 35308 56308 35364 56924
rect 35980 56866 36036 56878
rect 35980 56814 35982 56866
rect 36034 56814 36036 56866
rect 35980 56644 36036 56814
rect 36428 56866 36484 58156
rect 36428 56814 36430 56866
rect 36482 56814 36484 56866
rect 36428 56802 36484 56814
rect 36764 56980 36820 56990
rect 35980 56578 36036 56588
rect 36428 56644 36484 56654
rect 35308 56242 35364 56252
rect 36204 56308 36260 56318
rect 36204 56214 36260 56252
rect 33740 56030 33742 56082
rect 33794 56030 33796 56082
rect 33740 56018 33796 56030
rect 33852 55972 33908 55982
rect 33852 54740 33908 55916
rect 35756 55972 35812 55982
rect 35756 55410 35812 55916
rect 35756 55358 35758 55410
rect 35810 55358 35812 55410
rect 35756 55346 35812 55358
rect 36428 55410 36484 56588
rect 36764 56306 36820 56924
rect 36876 56868 36932 58268
rect 37100 58212 37156 58222
rect 37100 58118 37156 58156
rect 36988 57092 37044 57102
rect 37212 57092 37268 59948
rect 37324 59910 37380 59948
rect 37324 58324 37380 58334
rect 37548 58324 37604 58334
rect 37324 58322 37492 58324
rect 37324 58270 37326 58322
rect 37378 58270 37492 58322
rect 37324 58268 37492 58270
rect 37324 58258 37380 58268
rect 37044 57036 37268 57092
rect 36988 56998 37044 57036
rect 37436 56980 37492 58268
rect 37548 58322 38388 58324
rect 37548 58270 37550 58322
rect 37602 58270 38388 58322
rect 37548 58268 38388 58270
rect 37548 58258 37604 58268
rect 37660 57874 37716 57886
rect 37660 57822 37662 57874
rect 37714 57822 37716 57874
rect 37212 56924 37604 56980
rect 36876 56812 37044 56868
rect 36764 56254 36766 56306
rect 36818 56254 36820 56306
rect 36764 56242 36820 56254
rect 36988 56756 37044 56812
rect 36988 56306 37044 56700
rect 36988 56254 36990 56306
rect 37042 56254 37044 56306
rect 36988 56242 37044 56254
rect 37212 56306 37268 56924
rect 37548 56866 37604 56924
rect 37548 56814 37550 56866
rect 37602 56814 37604 56866
rect 37548 56802 37604 56814
rect 37436 56756 37492 56766
rect 37436 56644 37492 56700
rect 37436 56588 37604 56644
rect 37212 56254 37214 56306
rect 37266 56254 37268 56306
rect 37100 55972 37156 55982
rect 37100 55878 37156 55916
rect 36428 55358 36430 55410
rect 36482 55358 36484 55410
rect 36428 55300 36484 55358
rect 36428 55234 36484 55244
rect 37100 55300 37156 55310
rect 37100 55206 37156 55244
rect 37212 55300 37268 56254
rect 37436 56194 37492 56206
rect 37436 56142 37438 56194
rect 37490 56142 37492 56194
rect 37436 55410 37492 56142
rect 37436 55358 37438 55410
rect 37490 55358 37492 55410
rect 37436 55346 37492 55358
rect 37212 55298 37380 55300
rect 37212 55246 37214 55298
rect 37266 55246 37380 55298
rect 37212 55244 37380 55246
rect 37212 55234 37268 55244
rect 37324 55188 37380 55244
rect 37548 55298 37604 56588
rect 37548 55246 37550 55298
rect 37602 55246 37604 55298
rect 37548 55234 37604 55246
rect 37660 56308 37716 57822
rect 37772 56866 37828 58268
rect 38332 57874 38388 58268
rect 38332 57822 38334 57874
rect 38386 57822 38388 57874
rect 38332 57810 38388 57822
rect 37772 56814 37774 56866
rect 37826 56814 37828 56866
rect 37772 56802 37828 56814
rect 37324 55132 37492 55188
rect 35644 55076 35700 55086
rect 35308 55074 35700 55076
rect 35308 55022 35646 55074
rect 35698 55022 35700 55074
rect 35308 55020 35700 55022
rect 34008 54908 35208 54918
rect 34064 54906 34112 54908
rect 34168 54906 34216 54908
rect 34076 54854 34112 54906
rect 34200 54854 34216 54906
rect 34064 54852 34112 54854
rect 34168 54852 34216 54854
rect 34272 54906 34320 54908
rect 34376 54906 34424 54908
rect 34480 54906 34528 54908
rect 34376 54854 34396 54906
rect 34480 54854 34520 54906
rect 34272 54852 34320 54854
rect 34376 54852 34424 54854
rect 34480 54852 34528 54854
rect 34584 54852 34632 54908
rect 34688 54906 34736 54908
rect 34792 54906 34840 54908
rect 34896 54906 34944 54908
rect 34696 54854 34736 54906
rect 34820 54854 34840 54906
rect 34688 54852 34736 54854
rect 34792 54852 34840 54854
rect 34896 54852 34944 54854
rect 35000 54906 35048 54908
rect 35104 54906 35152 54908
rect 35000 54854 35016 54906
rect 35104 54854 35140 54906
rect 35000 54852 35048 54854
rect 35104 54852 35152 54854
rect 34008 54842 35208 54852
rect 34076 54740 34132 54750
rect 33852 54738 34580 54740
rect 33852 54686 34078 54738
rect 34130 54686 34580 54738
rect 33852 54684 34580 54686
rect 34076 54674 34132 54684
rect 34524 54514 34580 54684
rect 34524 54462 34526 54514
rect 34578 54462 34580 54514
rect 34524 54450 34580 54462
rect 35196 54516 35252 54526
rect 35308 54516 35364 55020
rect 35644 55010 35700 55020
rect 35196 54514 35364 54516
rect 35196 54462 35198 54514
rect 35250 54462 35364 54514
rect 35196 54460 35364 54462
rect 37436 54516 37492 55132
rect 37660 55076 37716 56252
rect 37548 55020 37716 55076
rect 37548 54738 37604 55020
rect 37548 54686 37550 54738
rect 37602 54686 37604 54738
rect 37548 54674 37604 54686
rect 38220 54516 38276 54526
rect 37436 54514 38276 54516
rect 37436 54462 38222 54514
rect 38274 54462 38276 54514
rect 37436 54460 38276 54462
rect 35196 54450 35252 54460
rect 38220 54450 38276 54460
rect 33628 54350 33630 54402
rect 33682 54350 33684 54402
rect 33180 51940 33236 51950
rect 33628 51940 33684 54350
rect 34008 53340 35208 53350
rect 34064 53338 34112 53340
rect 34168 53338 34216 53340
rect 34076 53286 34112 53338
rect 34200 53286 34216 53338
rect 34064 53284 34112 53286
rect 34168 53284 34216 53286
rect 34272 53338 34320 53340
rect 34376 53338 34424 53340
rect 34480 53338 34528 53340
rect 34376 53286 34396 53338
rect 34480 53286 34520 53338
rect 34272 53284 34320 53286
rect 34376 53284 34424 53286
rect 34480 53284 34528 53286
rect 34584 53284 34632 53340
rect 34688 53338 34736 53340
rect 34792 53338 34840 53340
rect 34896 53338 34944 53340
rect 34696 53286 34736 53338
rect 34820 53286 34840 53338
rect 34688 53284 34736 53286
rect 34792 53284 34840 53286
rect 34896 53284 34944 53286
rect 35000 53338 35048 53340
rect 35104 53338 35152 53340
rect 35000 53286 35016 53338
rect 35104 53286 35140 53338
rect 35000 53284 35048 53286
rect 35104 53284 35152 53286
rect 34008 53274 35208 53284
rect 34076 51940 34132 51950
rect 33628 51938 34132 51940
rect 33628 51886 34078 51938
rect 34130 51886 34132 51938
rect 33628 51884 34132 51886
rect 33180 51380 33236 51884
rect 33180 51286 33236 51324
rect 33852 51604 33908 51884
rect 34076 51874 34132 51884
rect 34860 51940 34916 51978
rect 34860 51874 34916 51884
rect 34008 51772 35208 51782
rect 34064 51770 34112 51772
rect 34168 51770 34216 51772
rect 34076 51718 34112 51770
rect 34200 51718 34216 51770
rect 34064 51716 34112 51718
rect 34168 51716 34216 51718
rect 34272 51770 34320 51772
rect 34376 51770 34424 51772
rect 34480 51770 34528 51772
rect 34376 51718 34396 51770
rect 34480 51718 34520 51770
rect 34272 51716 34320 51718
rect 34376 51716 34424 51718
rect 34480 51716 34528 51718
rect 34584 51716 34632 51772
rect 34688 51770 34736 51772
rect 34792 51770 34840 51772
rect 34896 51770 34944 51772
rect 34696 51718 34736 51770
rect 34820 51718 34840 51770
rect 34688 51716 34736 51718
rect 34792 51716 34840 51718
rect 34896 51716 34944 51718
rect 35000 51770 35048 51772
rect 35104 51770 35152 51772
rect 35000 51718 35016 51770
rect 35104 51718 35140 51770
rect 35000 51716 35048 51718
rect 35104 51716 35152 51718
rect 34008 51706 35208 51716
rect 33852 50484 33908 51548
rect 33852 50418 33908 50428
rect 34524 50484 34580 50494
rect 34524 50390 34580 50428
rect 35308 50370 35364 50382
rect 35308 50318 35310 50370
rect 35362 50318 35364 50370
rect 34008 50204 35208 50214
rect 34064 50202 34112 50204
rect 34168 50202 34216 50204
rect 34076 50150 34112 50202
rect 34200 50150 34216 50202
rect 34064 50148 34112 50150
rect 34168 50148 34216 50150
rect 34272 50202 34320 50204
rect 34376 50202 34424 50204
rect 34480 50202 34528 50204
rect 34376 50150 34396 50202
rect 34480 50150 34520 50202
rect 34272 50148 34320 50150
rect 34376 50148 34424 50150
rect 34480 50148 34528 50150
rect 34584 50148 34632 50204
rect 34688 50202 34736 50204
rect 34792 50202 34840 50204
rect 34896 50202 34944 50204
rect 34696 50150 34736 50202
rect 34820 50150 34840 50202
rect 34688 50148 34736 50150
rect 34792 50148 34840 50150
rect 34896 50148 34944 50150
rect 35000 50202 35048 50204
rect 35104 50202 35152 50204
rect 35000 50150 35016 50202
rect 35104 50150 35140 50202
rect 35000 50148 35048 50150
rect 35104 50148 35152 50150
rect 34008 50138 35208 50148
rect 33180 49700 33236 49710
rect 33180 49606 33236 49644
rect 33740 49700 33796 49710
rect 33796 49644 33908 49700
rect 33740 49634 33796 49644
rect 33516 49252 33572 49262
rect 33516 49158 33572 49196
rect 32844 49026 32900 49038
rect 32844 48974 32846 49026
rect 32898 48974 32900 49026
rect 32844 48020 32900 48974
rect 33068 49028 33124 49038
rect 33068 48934 33124 48972
rect 33628 49028 33684 49038
rect 33628 48934 33684 48972
rect 33740 48804 33796 48814
rect 33628 48802 33796 48804
rect 33628 48750 33742 48802
rect 33794 48750 33796 48802
rect 33628 48748 33796 48750
rect 33068 48244 33124 48254
rect 33068 48242 33348 48244
rect 33068 48190 33070 48242
rect 33122 48190 33348 48242
rect 33068 48188 33348 48190
rect 33068 48178 33124 48188
rect 33180 48020 33236 48030
rect 32844 48018 33236 48020
rect 32844 47966 33182 48018
rect 33234 47966 33236 48018
rect 32844 47964 33236 47966
rect 33180 47346 33236 47964
rect 33180 47294 33182 47346
rect 33234 47294 33236 47346
rect 33180 47282 33236 47294
rect 32732 46946 32788 46956
rect 32620 46610 32676 46620
rect 33180 46564 33236 46574
rect 33292 46564 33348 48188
rect 33628 47460 33684 48748
rect 33740 48738 33796 48748
rect 33740 48244 33796 48254
rect 33852 48244 33908 49644
rect 34300 48804 34356 48842
rect 34300 48738 34356 48748
rect 34008 48636 35208 48646
rect 34064 48634 34112 48636
rect 34168 48634 34216 48636
rect 34076 48582 34112 48634
rect 34200 48582 34216 48634
rect 34064 48580 34112 48582
rect 34168 48580 34216 48582
rect 34272 48634 34320 48636
rect 34376 48634 34424 48636
rect 34480 48634 34528 48636
rect 34376 48582 34396 48634
rect 34480 48582 34520 48634
rect 34272 48580 34320 48582
rect 34376 48580 34424 48582
rect 34480 48580 34528 48582
rect 34584 48580 34632 48636
rect 34688 48634 34736 48636
rect 34792 48634 34840 48636
rect 34896 48634 34944 48636
rect 34696 48582 34736 48634
rect 34820 48582 34840 48634
rect 34688 48580 34736 48582
rect 34792 48580 34840 48582
rect 34896 48580 34944 48582
rect 35000 48634 35048 48636
rect 35104 48634 35152 48636
rect 35000 48582 35016 48634
rect 35104 48582 35140 48634
rect 35000 48580 35048 48582
rect 35104 48580 35152 48582
rect 34008 48570 35208 48580
rect 33740 48242 33908 48244
rect 33740 48190 33742 48242
rect 33794 48190 33908 48242
rect 33740 48188 33908 48190
rect 34076 48244 34132 48254
rect 33740 48178 33796 48188
rect 34076 48150 34132 48188
rect 33628 47404 33908 47460
rect 33628 47236 33684 47246
rect 33628 47234 33796 47236
rect 33628 47182 33630 47234
rect 33682 47182 33796 47234
rect 33628 47180 33796 47182
rect 33628 47170 33684 47180
rect 33628 46564 33684 46574
rect 33292 46562 33684 46564
rect 33292 46510 33630 46562
rect 33682 46510 33684 46562
rect 33292 46508 33684 46510
rect 33180 46470 33236 46508
rect 32284 44996 32340 46284
rect 33628 46452 33684 46508
rect 33180 45890 33236 45902
rect 33180 45838 33182 45890
rect 33234 45838 33236 45890
rect 33180 45668 33236 45838
rect 33180 45602 33236 45612
rect 33628 45444 33684 46396
rect 33628 45378 33684 45388
rect 32508 44996 32564 45006
rect 32284 44940 32508 44996
rect 32508 43428 32564 44940
rect 33740 44324 33796 47180
rect 33852 46900 33908 47404
rect 34008 47068 35208 47078
rect 34064 47066 34112 47068
rect 34168 47066 34216 47068
rect 34076 47014 34112 47066
rect 34200 47014 34216 47066
rect 34064 47012 34112 47014
rect 34168 47012 34216 47014
rect 34272 47066 34320 47068
rect 34376 47066 34424 47068
rect 34480 47066 34528 47068
rect 34376 47014 34396 47066
rect 34480 47014 34520 47066
rect 34272 47012 34320 47014
rect 34376 47012 34424 47014
rect 34480 47012 34528 47014
rect 34584 47012 34632 47068
rect 34688 47066 34736 47068
rect 34792 47066 34840 47068
rect 34896 47066 34944 47068
rect 34696 47014 34736 47066
rect 34820 47014 34840 47066
rect 34688 47012 34736 47014
rect 34792 47012 34840 47014
rect 34896 47012 34944 47014
rect 35000 47066 35048 47068
rect 35104 47066 35152 47068
rect 35000 47014 35016 47066
rect 35104 47014 35140 47066
rect 35000 47012 35048 47014
rect 35104 47012 35152 47014
rect 34008 47002 35208 47012
rect 34076 46900 34132 46910
rect 33852 46898 34132 46900
rect 33852 46846 34078 46898
rect 34130 46846 34132 46898
rect 33852 46844 34132 46846
rect 33852 45332 33908 46844
rect 34076 46834 34132 46844
rect 34524 46788 34580 46798
rect 34524 46694 34580 46732
rect 34188 46676 34244 46686
rect 34188 46582 34244 46620
rect 34636 46674 34692 46686
rect 34636 46622 34638 46674
rect 34690 46622 34692 46674
rect 34636 46340 34692 46622
rect 35196 46674 35252 46686
rect 35196 46622 35198 46674
rect 35250 46622 35252 46674
rect 34692 46284 34804 46340
rect 34636 46274 34692 46284
rect 34748 46114 34804 46284
rect 34748 46062 34750 46114
rect 34802 46062 34804 46114
rect 34748 46050 34804 46062
rect 35196 45780 35252 46622
rect 35308 46452 35364 50318
rect 36428 48692 36484 48702
rect 36428 48466 36484 48636
rect 36428 48414 36430 48466
rect 36482 48414 36484 48466
rect 36428 48402 36484 48414
rect 37212 48018 37268 48030
rect 37212 47966 37214 48018
rect 37266 47966 37268 48018
rect 36316 47458 36372 47470
rect 36316 47406 36318 47458
rect 36370 47406 36372 47458
rect 35756 47346 35812 47358
rect 35756 47294 35758 47346
rect 35810 47294 35812 47346
rect 35756 46564 35812 47294
rect 36316 46900 36372 47406
rect 37212 47460 37268 47966
rect 37548 47460 37604 47470
rect 37212 47458 37604 47460
rect 37212 47406 37550 47458
rect 37602 47406 37604 47458
rect 37212 47404 37604 47406
rect 37100 47234 37156 47246
rect 37100 47182 37102 47234
rect 37154 47182 37156 47234
rect 36316 46834 36372 46844
rect 36540 46900 36596 46910
rect 36540 46898 36932 46900
rect 36540 46846 36542 46898
rect 36594 46846 36932 46898
rect 36540 46844 36932 46846
rect 36540 46834 36596 46844
rect 35308 46386 35364 46396
rect 35644 46452 35700 46462
rect 35532 46340 35588 46350
rect 35532 46002 35588 46284
rect 35532 45950 35534 46002
rect 35586 45950 35588 46002
rect 35532 45938 35588 45950
rect 35420 45780 35476 45790
rect 35196 45724 35420 45780
rect 34008 45500 35208 45510
rect 34064 45498 34112 45500
rect 34168 45498 34216 45500
rect 34076 45446 34112 45498
rect 34200 45446 34216 45498
rect 34064 45444 34112 45446
rect 34168 45444 34216 45446
rect 34272 45498 34320 45500
rect 34376 45498 34424 45500
rect 34480 45498 34528 45500
rect 34376 45446 34396 45498
rect 34480 45446 34520 45498
rect 34272 45444 34320 45446
rect 34376 45444 34424 45446
rect 34480 45444 34528 45446
rect 34584 45444 34632 45500
rect 34688 45498 34736 45500
rect 34792 45498 34840 45500
rect 34896 45498 34944 45500
rect 34696 45446 34736 45498
rect 34820 45446 34840 45498
rect 34688 45444 34736 45446
rect 34792 45444 34840 45446
rect 34896 45444 34944 45446
rect 35000 45498 35048 45500
rect 35104 45498 35152 45500
rect 35000 45446 35016 45498
rect 35104 45446 35140 45498
rect 35000 45444 35048 45446
rect 35104 45444 35152 45446
rect 34008 45434 35208 45444
rect 34300 45332 34356 45342
rect 33852 45276 34244 45332
rect 34188 45218 34244 45276
rect 34356 45276 34468 45332
rect 34300 45266 34356 45276
rect 34188 45166 34190 45218
rect 34242 45166 34244 45218
rect 34188 45154 34244 45166
rect 34412 45218 34468 45276
rect 34412 45166 34414 45218
rect 34466 45166 34468 45218
rect 34412 45154 34468 45166
rect 34860 45220 34916 45230
rect 34860 45126 34916 45164
rect 34636 45106 34692 45118
rect 34636 45054 34638 45106
rect 34690 45054 34692 45106
rect 33852 44996 33908 45006
rect 33908 44940 34244 44996
rect 33852 44902 33908 44940
rect 34188 44434 34244 44940
rect 34188 44382 34190 44434
rect 34242 44382 34244 44434
rect 34188 44370 34244 44382
rect 33740 44258 33796 44268
rect 34524 44324 34580 44334
rect 34524 44230 34580 44268
rect 34636 44212 34692 45054
rect 35420 45106 35476 45724
rect 35644 45444 35700 46396
rect 35756 45892 35812 46508
rect 35980 46674 36036 46686
rect 35980 46622 35982 46674
rect 36034 46622 36036 46674
rect 35980 46452 36036 46622
rect 36204 46676 36260 46686
rect 36204 46582 36260 46620
rect 35980 46386 36036 46396
rect 35756 45798 35812 45836
rect 36316 46340 36372 46350
rect 35420 45054 35422 45106
rect 35474 45054 35476 45106
rect 35420 45042 35476 45054
rect 35532 45388 35700 45444
rect 35980 45666 36036 45678
rect 35980 45614 35982 45666
rect 36034 45614 36036 45666
rect 34748 44884 34804 44894
rect 34748 44790 34804 44828
rect 35308 44322 35364 44334
rect 35308 44270 35310 44322
rect 35362 44270 35364 44322
rect 34636 44118 34692 44156
rect 34860 44212 34916 44222
rect 35196 44212 35252 44222
rect 34860 44210 35252 44212
rect 34860 44158 34862 44210
rect 34914 44158 35198 44210
rect 35250 44158 35252 44210
rect 34860 44156 35252 44158
rect 34860 44146 34916 44156
rect 35196 44146 35252 44156
rect 33852 44100 33908 44110
rect 32508 43362 32564 43372
rect 33740 43426 33796 43438
rect 33740 43374 33742 43426
rect 33794 43374 33796 43426
rect 32284 43314 32340 43326
rect 32284 43262 32286 43314
rect 32338 43262 32340 43314
rect 32060 42030 32062 42082
rect 32114 42030 32116 42082
rect 32060 42018 32116 42030
rect 32172 42196 32228 42206
rect 32172 41970 32228 42140
rect 32172 41918 32174 41970
rect 32226 41918 32228 41970
rect 32172 41906 32228 41918
rect 31780 41580 32004 41636
rect 31724 41186 31780 41580
rect 32172 41412 32228 41422
rect 32172 41318 32228 41356
rect 31724 41134 31726 41186
rect 31778 41134 31780 41186
rect 31724 41122 31780 41134
rect 32060 41188 32116 41198
rect 32060 41094 32116 41132
rect 32284 41188 32340 43262
rect 33180 42754 33236 42766
rect 33180 42702 33182 42754
rect 33234 42702 33236 42754
rect 32396 42642 32452 42654
rect 32396 42590 32398 42642
rect 32450 42590 32452 42642
rect 32396 41300 32452 42590
rect 32396 41234 32452 41244
rect 32844 42530 32900 42542
rect 32844 42478 32846 42530
rect 32898 42478 32900 42530
rect 32284 41122 32340 41132
rect 31388 41076 31444 41086
rect 31276 41074 31444 41076
rect 31276 41022 31390 41074
rect 31442 41022 31444 41074
rect 31276 41020 31444 41022
rect 31388 41010 31444 41020
rect 32732 41074 32788 41086
rect 32732 41022 32734 41074
rect 32786 41022 32788 41074
rect 31612 40628 31668 40638
rect 31052 40514 31556 40516
rect 31052 40462 31054 40514
rect 31106 40462 31556 40514
rect 31052 40460 31556 40462
rect 31052 40450 31108 40460
rect 30940 40404 30996 40414
rect 30940 39956 30996 40348
rect 31500 40292 31556 40460
rect 30940 39900 31108 39956
rect 31052 39730 31108 39900
rect 31052 39678 31054 39730
rect 31106 39678 31108 39730
rect 31052 39666 31108 39678
rect 31500 39730 31556 40236
rect 31500 39678 31502 39730
rect 31554 39678 31556 39730
rect 31500 39666 31556 39678
rect 31612 38668 31668 40572
rect 32172 40404 32228 40414
rect 32172 40310 32228 40348
rect 32396 40180 32452 40190
rect 32396 40086 32452 40124
rect 31948 39732 32004 39742
rect 31948 39730 32564 39732
rect 31948 39678 31950 39730
rect 32002 39678 32564 39730
rect 31948 39676 32564 39678
rect 31948 39666 32004 39676
rect 30604 37426 30660 37436
rect 30716 38612 30884 38668
rect 31500 38612 31668 38668
rect 31836 38724 31892 38734
rect 30492 37268 30548 37278
rect 29484 36430 29486 36482
rect 29538 36430 29540 36482
rect 29484 36418 29540 36430
rect 30156 36428 30324 36484
rect 30380 37212 30492 37268
rect 30380 36482 30436 37212
rect 30492 37202 30548 37212
rect 30380 36430 30382 36482
rect 30434 36430 30436 36482
rect 28028 36318 28030 36370
rect 28082 36318 28084 36370
rect 27356 36260 27412 36270
rect 27356 36258 27636 36260
rect 27356 36206 27358 36258
rect 27410 36206 27636 36258
rect 27356 36204 27636 36206
rect 27356 36194 27412 36204
rect 27356 35812 27412 35822
rect 27244 35476 27300 35486
rect 27244 35382 27300 35420
rect 27356 35026 27412 35756
rect 27580 35698 27636 36204
rect 27804 35812 27860 35822
rect 27804 35718 27860 35756
rect 27580 35646 27582 35698
rect 27634 35646 27636 35698
rect 27580 35634 27636 35646
rect 27356 34974 27358 35026
rect 27410 34974 27412 35026
rect 27356 34962 27412 34974
rect 27804 34804 27860 34814
rect 27804 34710 27860 34748
rect 27132 34626 27188 34636
rect 26684 34078 26686 34130
rect 26738 34078 26740 34130
rect 26684 34066 26740 34078
rect 26236 33460 26292 33470
rect 26236 33366 26292 33404
rect 27020 33460 27076 33470
rect 25788 32788 25844 32798
rect 25788 32694 25844 32732
rect 26236 32676 26292 32686
rect 26236 32582 26292 32620
rect 27020 32562 27076 33404
rect 27244 32676 27300 32686
rect 27244 32582 27300 32620
rect 27804 32674 27860 32686
rect 27804 32622 27806 32674
rect 27858 32622 27860 32674
rect 27020 32510 27022 32562
rect 27074 32510 27076 32562
rect 27020 32498 27076 32510
rect 26236 32340 26292 32350
rect 26236 31778 26292 32284
rect 26684 32338 26740 32350
rect 26684 32286 26686 32338
rect 26738 32286 26740 32338
rect 26236 31726 26238 31778
rect 26290 31726 26292 31778
rect 26236 31714 26292 31726
rect 26348 31892 26404 31902
rect 25564 30994 25732 30996
rect 25564 30942 25566 30994
rect 25618 30942 25732 30994
rect 25564 30940 25732 30942
rect 25900 31556 25956 31566
rect 26348 31556 26404 31836
rect 25900 31554 26404 31556
rect 25900 31502 25902 31554
rect 25954 31502 26350 31554
rect 26402 31502 26404 31554
rect 25900 31500 26404 31502
rect 25564 30930 25620 30940
rect 25900 30324 25956 31500
rect 26348 31490 26404 31500
rect 26572 31556 26628 31566
rect 26572 31462 26628 31500
rect 26012 30996 26068 31006
rect 26012 30994 26628 30996
rect 26012 30942 26014 30994
rect 26066 30942 26628 30994
rect 26012 30940 26628 30942
rect 26012 30930 26068 30940
rect 26572 30434 26628 30940
rect 26572 30382 26574 30434
rect 26626 30382 26628 30434
rect 26572 30370 26628 30382
rect 26684 30436 26740 32286
rect 27692 31780 27748 31790
rect 27692 31686 27748 31724
rect 26908 31668 26964 31678
rect 27132 31668 27188 31678
rect 26908 31666 27132 31668
rect 26908 31614 26910 31666
rect 26962 31614 27132 31666
rect 26908 31612 27132 31614
rect 26908 31602 26964 31612
rect 27132 31602 27188 31612
rect 27356 31556 27412 31566
rect 27356 31462 27412 31500
rect 27804 31444 27860 32622
rect 28028 31668 28084 36318
rect 28476 36370 28532 36382
rect 28476 36318 28478 36370
rect 28530 36318 28532 36370
rect 28364 35810 28420 35822
rect 28364 35758 28366 35810
rect 28418 35758 28420 35810
rect 28252 34916 28308 34926
rect 28252 34690 28308 34860
rect 28252 34638 28254 34690
rect 28306 34638 28308 34690
rect 28252 33684 28308 34638
rect 28364 34356 28420 35758
rect 28476 35812 28532 36318
rect 29708 36260 29764 36270
rect 30044 36260 30100 36270
rect 29708 36258 30100 36260
rect 29708 36206 29710 36258
rect 29762 36206 30046 36258
rect 30098 36206 30100 36258
rect 29708 36204 30100 36206
rect 29708 36194 29764 36204
rect 30044 36194 30100 36204
rect 30156 36036 30212 36428
rect 30380 36418 30436 36430
rect 30268 36260 30324 36270
rect 30716 36260 30772 38612
rect 31388 37938 31444 37950
rect 31388 37886 31390 37938
rect 31442 37886 31444 37938
rect 31052 37828 31108 37838
rect 31388 37828 31444 37886
rect 31108 37772 31444 37828
rect 31052 37734 31108 37772
rect 31164 37492 31220 37502
rect 31164 37398 31220 37436
rect 31164 37156 31220 37166
rect 31164 36482 31220 37100
rect 31164 36430 31166 36482
rect 31218 36430 31220 36482
rect 31164 36418 31220 36430
rect 30828 36260 30884 36270
rect 30268 36258 30884 36260
rect 30268 36206 30270 36258
rect 30322 36206 30830 36258
rect 30882 36206 30884 36258
rect 30268 36204 30884 36206
rect 30268 36194 30324 36204
rect 30156 35980 30436 36036
rect 28476 35746 28532 35756
rect 29820 34692 29876 34702
rect 29596 34690 29876 34692
rect 29596 34638 29822 34690
rect 29874 34638 29876 34690
rect 29596 34636 29876 34638
rect 28364 34290 28420 34300
rect 29148 34356 29204 34366
rect 29596 34356 29652 34636
rect 29820 34626 29876 34636
rect 29148 34354 29652 34356
rect 29148 34302 29150 34354
rect 29202 34302 29652 34354
rect 29148 34300 29652 34302
rect 29708 34356 29764 34366
rect 29148 34290 29204 34300
rect 28252 33618 28308 33628
rect 28028 31574 28084 31612
rect 28476 31780 28532 31790
rect 28476 31666 28532 31724
rect 28476 31614 28478 31666
rect 28530 31614 28532 31666
rect 28476 31602 28532 31614
rect 27804 31378 27860 31388
rect 28364 31218 28420 31230
rect 28364 31166 28366 31218
rect 28418 31166 28420 31218
rect 27468 31108 27524 31118
rect 26908 30436 26964 30446
rect 26684 30434 26964 30436
rect 26684 30382 26910 30434
rect 26962 30382 26964 30434
rect 26684 30380 26964 30382
rect 26908 30370 26964 30380
rect 26012 30324 26068 30334
rect 25900 30268 26012 30324
rect 25452 29922 25508 29932
rect 24444 27748 24500 27758
rect 24444 27654 24500 27692
rect 24008 27468 25208 27478
rect 24064 27466 24112 27468
rect 24168 27466 24216 27468
rect 24076 27414 24112 27466
rect 24200 27414 24216 27466
rect 24064 27412 24112 27414
rect 24168 27412 24216 27414
rect 24272 27466 24320 27468
rect 24376 27466 24424 27468
rect 24480 27466 24528 27468
rect 24376 27414 24396 27466
rect 24480 27414 24520 27466
rect 24272 27412 24320 27414
rect 24376 27412 24424 27414
rect 24480 27412 24528 27414
rect 24584 27412 24632 27468
rect 24688 27466 24736 27468
rect 24792 27466 24840 27468
rect 24896 27466 24944 27468
rect 24696 27414 24736 27466
rect 24820 27414 24840 27466
rect 24688 27412 24736 27414
rect 24792 27412 24840 27414
rect 24896 27412 24944 27414
rect 25000 27466 25048 27468
rect 25104 27466 25152 27468
rect 25000 27414 25016 27466
rect 25104 27414 25140 27466
rect 25000 27412 25048 27414
rect 25104 27412 25152 27414
rect 24008 27402 25208 27412
rect 25340 27300 25396 28028
rect 24892 27244 25396 27300
rect 25452 29428 25508 29438
rect 25452 28644 25508 29372
rect 24892 26962 24948 27244
rect 24892 26910 24894 26962
rect 24946 26910 24948 26962
rect 23772 26852 23940 26908
rect 24892 26898 24948 26910
rect 25452 26908 25508 28588
rect 26012 28308 26068 30268
rect 26684 30212 26740 30222
rect 26124 29988 26180 29998
rect 26124 29894 26180 29932
rect 26684 29650 26740 30156
rect 27468 30098 27524 31052
rect 28364 30884 28420 31166
rect 29036 31108 29092 31118
rect 29036 31014 29092 31052
rect 28364 30324 28420 30828
rect 28364 30258 28420 30268
rect 29372 30884 29428 34300
rect 29708 34262 29764 34300
rect 30156 34356 30212 34366
rect 30156 34242 30212 34300
rect 30156 34190 30158 34242
rect 30210 34190 30212 34242
rect 30156 34178 30212 34190
rect 30268 34242 30324 34254
rect 30268 34190 30270 34242
rect 30322 34190 30324 34242
rect 30268 33908 30324 34190
rect 30156 33852 30324 33908
rect 29820 33124 29876 33134
rect 30156 33124 30212 33852
rect 29820 33122 30212 33124
rect 29820 33070 29822 33122
rect 29874 33070 30212 33122
rect 29820 33068 30212 33070
rect 30268 33684 30324 33694
rect 30268 33122 30324 33628
rect 30268 33070 30270 33122
rect 30322 33070 30324 33122
rect 29820 31892 29876 33068
rect 30156 32788 30212 32798
rect 29820 31826 29876 31836
rect 29932 32676 29988 32686
rect 29932 31778 29988 32620
rect 29932 31726 29934 31778
rect 29986 31726 29988 31778
rect 29932 31714 29988 31726
rect 30156 31778 30212 32732
rect 30156 31726 30158 31778
rect 30210 31726 30212 31778
rect 30156 31714 30212 31726
rect 27468 30046 27470 30098
rect 27522 30046 27524 30098
rect 27468 30034 27524 30046
rect 27692 30210 27748 30222
rect 27692 30158 27694 30210
rect 27746 30158 27748 30210
rect 27692 30100 27748 30158
rect 27692 30034 27748 30044
rect 28588 30100 28644 30110
rect 28588 30006 28644 30044
rect 26684 29598 26686 29650
rect 26738 29598 26740 29650
rect 26684 28754 26740 29598
rect 27580 29988 27636 29998
rect 27132 29428 27188 29438
rect 27132 29334 27188 29372
rect 27580 29426 27636 29932
rect 29260 29988 29316 29998
rect 29260 29894 29316 29932
rect 29372 29540 29428 30828
rect 29596 31556 29652 31566
rect 29596 30434 29652 31500
rect 29820 31554 29876 31566
rect 29820 31502 29822 31554
rect 29874 31502 29876 31554
rect 29820 31108 29876 31502
rect 29820 31052 29988 31108
rect 29596 30382 29598 30434
rect 29650 30382 29652 30434
rect 29596 30370 29652 30382
rect 29820 30882 29876 30894
rect 29820 30830 29822 30882
rect 29874 30830 29876 30882
rect 29820 30324 29876 30830
rect 29820 30258 29876 30268
rect 29820 30100 29876 30110
rect 29820 30006 29876 30044
rect 29820 29540 29876 29550
rect 29372 29538 29876 29540
rect 29372 29486 29822 29538
rect 29874 29486 29876 29538
rect 29372 29484 29876 29486
rect 27580 29374 27582 29426
rect 27634 29374 27636 29426
rect 27580 29362 27636 29374
rect 26684 28702 26686 28754
rect 26738 28702 26740 28754
rect 26684 28690 26740 28702
rect 28140 28644 28196 28654
rect 28140 28550 28196 28588
rect 29708 28644 29764 29484
rect 29820 29474 29876 29484
rect 26012 28252 26180 28308
rect 26012 28084 26068 28094
rect 25676 27860 25732 27870
rect 25676 27298 25732 27804
rect 25676 27246 25678 27298
rect 25730 27246 25732 27298
rect 25676 27188 25732 27246
rect 25788 27746 25844 27758
rect 25788 27694 25790 27746
rect 25842 27694 25844 27746
rect 25788 27300 25844 27694
rect 25900 27300 25956 27310
rect 25844 27298 25956 27300
rect 25844 27246 25902 27298
rect 25954 27246 25956 27298
rect 25844 27244 25956 27246
rect 25788 27206 25844 27244
rect 25900 27234 25956 27244
rect 25676 27122 25732 27132
rect 26012 27186 26068 28028
rect 26012 27134 26014 27186
rect 26066 27134 26068 27186
rect 26012 27122 26068 27134
rect 26124 26908 26180 28252
rect 29708 28082 29764 28588
rect 29708 28030 29710 28082
rect 29762 28030 29764 28082
rect 29708 28018 29764 28030
rect 26460 27298 26516 27310
rect 26460 27246 26462 27298
rect 26514 27246 26516 27298
rect 25452 26852 25620 26908
rect 23660 26674 23716 26684
rect 23772 26180 23828 26190
rect 23772 26086 23828 26124
rect 23772 25732 23828 25742
rect 23772 25638 23828 25676
rect 23772 23716 23828 23726
rect 23884 23716 23940 26852
rect 24008 25900 25208 25910
rect 24064 25898 24112 25900
rect 24168 25898 24216 25900
rect 24076 25846 24112 25898
rect 24200 25846 24216 25898
rect 24064 25844 24112 25846
rect 24168 25844 24216 25846
rect 24272 25898 24320 25900
rect 24376 25898 24424 25900
rect 24480 25898 24528 25900
rect 24376 25846 24396 25898
rect 24480 25846 24520 25898
rect 24272 25844 24320 25846
rect 24376 25844 24424 25846
rect 24480 25844 24528 25846
rect 24584 25844 24632 25900
rect 24688 25898 24736 25900
rect 24792 25898 24840 25900
rect 24896 25898 24944 25900
rect 24696 25846 24736 25898
rect 24820 25846 24840 25898
rect 24688 25844 24736 25846
rect 24792 25844 24840 25846
rect 24896 25844 24944 25846
rect 25000 25898 25048 25900
rect 25104 25898 25152 25900
rect 25000 25846 25016 25898
rect 25104 25846 25140 25898
rect 25000 25844 25048 25846
rect 25104 25844 25152 25846
rect 24008 25834 25208 25844
rect 24556 25284 24612 25294
rect 24556 25190 24612 25228
rect 24668 24836 24724 24846
rect 24668 24742 24724 24780
rect 25452 24836 25508 24846
rect 25452 24742 25508 24780
rect 25228 24500 25284 24538
rect 25228 24434 25284 24444
rect 24008 24332 25208 24342
rect 24064 24330 24112 24332
rect 24168 24330 24216 24332
rect 24076 24278 24112 24330
rect 24200 24278 24216 24330
rect 24064 24276 24112 24278
rect 24168 24276 24216 24278
rect 24272 24330 24320 24332
rect 24376 24330 24424 24332
rect 24480 24330 24528 24332
rect 24376 24278 24396 24330
rect 24480 24278 24520 24330
rect 24272 24276 24320 24278
rect 24376 24276 24424 24278
rect 24480 24276 24528 24278
rect 24584 24276 24632 24332
rect 24688 24330 24736 24332
rect 24792 24330 24840 24332
rect 24896 24330 24944 24332
rect 24696 24278 24736 24330
rect 24820 24278 24840 24330
rect 24688 24276 24736 24278
rect 24792 24276 24840 24278
rect 24896 24276 24944 24278
rect 25000 24330 25048 24332
rect 25104 24330 25152 24332
rect 25000 24278 25016 24330
rect 25104 24278 25140 24330
rect 25000 24276 25048 24278
rect 25104 24276 25152 24278
rect 24008 24266 25208 24276
rect 24556 24052 24612 24062
rect 24556 23958 24612 23996
rect 24444 23938 24500 23950
rect 24444 23886 24446 23938
rect 24498 23886 24500 23938
rect 24108 23716 24164 23726
rect 23884 23714 24164 23716
rect 23884 23662 24110 23714
rect 24162 23662 24164 23714
rect 23884 23660 24164 23662
rect 23660 23044 23716 23054
rect 23660 22950 23716 22988
rect 23772 22260 23828 23660
rect 24108 23268 24164 23660
rect 24444 23716 24500 23886
rect 24892 23940 24948 23950
rect 24892 23846 24948 23884
rect 25004 23938 25060 23950
rect 25004 23886 25006 23938
rect 25058 23886 25060 23938
rect 24444 23650 24500 23660
rect 24668 23716 24724 23726
rect 24668 23622 24724 23660
rect 24108 23202 24164 23212
rect 25004 22932 25060 23886
rect 25452 23938 25508 23950
rect 25452 23886 25454 23938
rect 25506 23886 25508 23938
rect 25340 23268 25396 23278
rect 25452 23268 25508 23886
rect 25396 23212 25508 23268
rect 25340 23174 25396 23212
rect 25004 22876 25396 22932
rect 24008 22764 25208 22774
rect 24064 22762 24112 22764
rect 24168 22762 24216 22764
rect 24076 22710 24112 22762
rect 24200 22710 24216 22762
rect 24064 22708 24112 22710
rect 24168 22708 24216 22710
rect 24272 22762 24320 22764
rect 24376 22762 24424 22764
rect 24480 22762 24528 22764
rect 24376 22710 24396 22762
rect 24480 22710 24520 22762
rect 24272 22708 24320 22710
rect 24376 22708 24424 22710
rect 24480 22708 24528 22710
rect 24584 22708 24632 22764
rect 24688 22762 24736 22764
rect 24792 22762 24840 22764
rect 24896 22762 24944 22764
rect 24696 22710 24736 22762
rect 24820 22710 24840 22762
rect 24688 22708 24736 22710
rect 24792 22708 24840 22710
rect 24896 22708 24944 22710
rect 25000 22762 25048 22764
rect 25104 22762 25152 22764
rect 25000 22710 25016 22762
rect 25104 22710 25140 22762
rect 25000 22708 25048 22710
rect 25104 22708 25152 22710
rect 24008 22698 25208 22708
rect 23996 22596 24052 22606
rect 23884 22484 23940 22494
rect 23884 22390 23940 22428
rect 23996 22370 24052 22540
rect 23996 22318 23998 22370
rect 24050 22318 24052 22370
rect 23996 22306 24052 22318
rect 24668 22370 24724 22382
rect 24668 22318 24670 22370
rect 24722 22318 24724 22370
rect 23772 22204 23940 22260
rect 23548 21746 23604 21756
rect 23324 21532 23604 21588
rect 23212 20738 23268 20748
rect 22988 20638 22990 20690
rect 23042 20638 23044 20690
rect 22988 20626 23044 20638
rect 23548 20356 23604 21532
rect 23884 20804 23940 22204
rect 23996 22148 24052 22158
rect 23996 21810 24052 22092
rect 23996 21758 23998 21810
rect 24050 21758 24052 21810
rect 23996 21746 24052 21758
rect 24668 21812 24724 22318
rect 24892 22260 24948 22270
rect 24892 22166 24948 22204
rect 25228 22260 25284 22270
rect 25340 22260 25396 22876
rect 25284 22204 25396 22260
rect 25452 22484 25508 22494
rect 25452 22370 25508 22428
rect 25452 22318 25454 22370
rect 25506 22318 25508 22370
rect 25228 22194 25284 22204
rect 25452 22148 25508 22318
rect 25452 22082 25508 22092
rect 24668 21588 24724 21756
rect 25340 21810 25396 21822
rect 25340 21758 25342 21810
rect 25394 21758 25396 21810
rect 25228 21588 25284 21598
rect 24668 21586 25284 21588
rect 24668 21534 25230 21586
rect 25282 21534 25284 21586
rect 24668 21532 25284 21534
rect 25228 21522 25284 21532
rect 24780 21364 24836 21402
rect 24780 21298 24836 21308
rect 24008 21196 25208 21206
rect 24064 21194 24112 21196
rect 24168 21194 24216 21196
rect 24076 21142 24112 21194
rect 24200 21142 24216 21194
rect 24064 21140 24112 21142
rect 24168 21140 24216 21142
rect 24272 21194 24320 21196
rect 24376 21194 24424 21196
rect 24480 21194 24528 21196
rect 24376 21142 24396 21194
rect 24480 21142 24520 21194
rect 24272 21140 24320 21142
rect 24376 21140 24424 21142
rect 24480 21140 24528 21142
rect 24584 21140 24632 21196
rect 24688 21194 24736 21196
rect 24792 21194 24840 21196
rect 24896 21194 24944 21196
rect 24696 21142 24736 21194
rect 24820 21142 24840 21194
rect 24688 21140 24736 21142
rect 24792 21140 24840 21142
rect 24896 21140 24944 21142
rect 25000 21194 25048 21196
rect 25104 21194 25152 21196
rect 25000 21142 25016 21194
rect 25104 21142 25140 21194
rect 25000 21140 25048 21142
rect 25104 21140 25152 21142
rect 24008 21130 25208 21140
rect 24220 21028 24276 21038
rect 24108 20916 24164 20926
rect 23996 20804 24052 20814
rect 23884 20802 24052 20804
rect 23884 20750 23998 20802
rect 24050 20750 24052 20802
rect 23884 20748 24052 20750
rect 23996 20738 24052 20748
rect 23660 20580 23716 20590
rect 23660 20486 23716 20524
rect 23884 20580 23940 20590
rect 24108 20580 24164 20860
rect 23884 20578 24164 20580
rect 23884 20526 23886 20578
rect 23938 20526 24164 20578
rect 23884 20524 24164 20526
rect 23884 20514 23940 20524
rect 23548 20300 23940 20356
rect 22540 19954 22596 19964
rect 23212 20020 23268 20030
rect 21420 19730 21476 19740
rect 21420 19460 21476 19470
rect 20524 18674 21364 18676
rect 20524 18622 20526 18674
rect 20578 18622 21364 18674
rect 20524 18620 21364 18622
rect 20524 18610 20580 18620
rect 21196 18452 21252 18462
rect 21196 18358 21252 18396
rect 21084 18228 21140 18238
rect 21084 18134 21140 18172
rect 20412 17668 20468 17678
rect 20412 17574 20468 17612
rect 20636 17668 20692 17678
rect 20636 17666 21028 17668
rect 20636 17614 20638 17666
rect 20690 17614 21028 17666
rect 20636 17612 21028 17614
rect 20636 17602 20692 17612
rect 19404 16718 19406 16770
rect 19458 16718 19460 16770
rect 19404 16706 19460 16718
rect 19740 16994 19796 17006
rect 19740 16942 19742 16994
rect 19794 16942 19796 16994
rect 19516 16660 19572 16670
rect 19516 16566 19572 16604
rect 19180 15262 19182 15314
rect 19234 15262 19236 15314
rect 19180 15250 19236 15262
rect 19740 15148 19796 16942
rect 20076 16994 20132 17052
rect 20860 17108 20916 17118
rect 20860 17014 20916 17052
rect 20076 16942 20078 16994
rect 20130 16942 20132 16994
rect 20076 16930 20132 16942
rect 20188 16882 20244 16894
rect 20188 16830 20190 16882
rect 20242 16830 20244 16882
rect 20188 16772 20244 16830
rect 20412 16884 20468 16894
rect 20972 16884 21028 17612
rect 21308 17444 21364 18620
rect 21420 18450 21476 19404
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18386 21476 18398
rect 21532 18562 21588 18574
rect 21532 18510 21534 18562
rect 21586 18510 21588 18562
rect 21532 17668 21588 18510
rect 21868 18450 21924 18462
rect 22540 18452 22596 18462
rect 21868 18398 21870 18450
rect 21922 18398 21924 18450
rect 21532 17602 21588 17612
rect 21644 17668 21700 17678
rect 21868 17668 21924 18398
rect 21644 17666 21924 17668
rect 21644 17614 21646 17666
rect 21698 17614 21924 17666
rect 21644 17612 21924 17614
rect 21420 17444 21476 17454
rect 21308 17442 21476 17444
rect 21308 17390 21422 17442
rect 21474 17390 21476 17442
rect 21308 17388 21476 17390
rect 21084 16884 21140 16894
rect 20972 16882 21140 16884
rect 20972 16830 21086 16882
rect 21138 16830 21140 16882
rect 20972 16828 21140 16830
rect 20412 16790 20468 16828
rect 20188 16706 20244 16716
rect 21084 16772 21140 16828
rect 21084 16706 21140 16716
rect 20748 16660 20804 16670
rect 20748 16566 20804 16604
rect 18060 14700 18172 14756
rect 18060 14642 18116 14700
rect 18172 14690 18228 14700
rect 19180 15092 19796 15148
rect 20524 15204 20580 15214
rect 18060 14590 18062 14642
rect 18114 14590 18116 14642
rect 18060 14578 18116 14590
rect 18620 14644 18676 14654
rect 18620 14550 18676 14588
rect 19180 14530 19236 15092
rect 19852 14644 19908 14654
rect 19852 14550 19908 14588
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 19180 14466 19236 14478
rect 18844 14418 18900 14430
rect 18844 14366 18846 14418
rect 18898 14366 18900 14418
rect 18060 13860 18116 13870
rect 18060 13766 18116 13804
rect 18620 13858 18676 13870
rect 18620 13806 18622 13858
rect 18674 13806 18676 13858
rect 17836 13694 17838 13746
rect 17890 13694 17892 13746
rect 17836 13682 17892 13694
rect 17500 13524 17556 13534
rect 16044 13458 16100 13468
rect 16940 13522 17556 13524
rect 16940 13470 17502 13522
rect 17554 13470 17556 13522
rect 16940 13468 17556 13470
rect 15484 12908 15596 12964
rect 15260 12674 15316 12684
rect 15372 12738 15428 12750
rect 15372 12686 15374 12738
rect 15426 12686 15428 12738
rect 14008 12572 15208 12582
rect 14064 12570 14112 12572
rect 14168 12570 14216 12572
rect 14076 12518 14112 12570
rect 14200 12518 14216 12570
rect 14064 12516 14112 12518
rect 14168 12516 14216 12518
rect 14272 12570 14320 12572
rect 14376 12570 14424 12572
rect 14480 12570 14528 12572
rect 14376 12518 14396 12570
rect 14480 12518 14520 12570
rect 14272 12516 14320 12518
rect 14376 12516 14424 12518
rect 14480 12516 14528 12518
rect 14584 12516 14632 12572
rect 14688 12570 14736 12572
rect 14792 12570 14840 12572
rect 14896 12570 14944 12572
rect 14696 12518 14736 12570
rect 14820 12518 14840 12570
rect 14688 12516 14736 12518
rect 14792 12516 14840 12518
rect 14896 12516 14944 12518
rect 15000 12570 15048 12572
rect 15104 12570 15152 12572
rect 15000 12518 15016 12570
rect 15104 12518 15140 12570
rect 15000 12516 15048 12518
rect 15104 12516 15152 12518
rect 14008 12506 15208 12516
rect 13916 12402 13972 12414
rect 13916 12350 13918 12402
rect 13970 12350 13972 12402
rect 13916 11620 13972 12350
rect 13916 11554 13972 11564
rect 14588 12404 14644 12414
rect 13916 11396 13972 11406
rect 13804 11394 13972 11396
rect 13804 11342 13918 11394
rect 13970 11342 13972 11394
rect 13804 11340 13972 11342
rect 13916 11330 13972 11340
rect 14588 11172 14644 12348
rect 14588 11106 14644 11116
rect 14008 11004 15208 11014
rect 14064 11002 14112 11004
rect 14168 11002 14216 11004
rect 14076 10950 14112 11002
rect 14200 10950 14216 11002
rect 14064 10948 14112 10950
rect 14168 10948 14216 10950
rect 14272 11002 14320 11004
rect 14376 11002 14424 11004
rect 14480 11002 14528 11004
rect 14376 10950 14396 11002
rect 14480 10950 14520 11002
rect 14272 10948 14320 10950
rect 14376 10948 14424 10950
rect 14480 10948 14528 10950
rect 14584 10948 14632 11004
rect 14688 11002 14736 11004
rect 14792 11002 14840 11004
rect 14896 11002 14944 11004
rect 14696 10950 14736 11002
rect 14820 10950 14840 11002
rect 14688 10948 14736 10950
rect 14792 10948 14840 10950
rect 14896 10948 14944 10950
rect 15000 11002 15048 11004
rect 15104 11002 15152 11004
rect 15000 10950 15016 11002
rect 15104 10950 15140 11002
rect 15000 10948 15048 10950
rect 15104 10948 15152 10950
rect 14008 10938 15208 10948
rect 14028 10836 14084 10846
rect 13692 10834 14084 10836
rect 13692 10782 14030 10834
rect 14082 10782 14084 10834
rect 13692 10780 14084 10782
rect 14028 10770 14084 10780
rect 14588 10836 14644 10846
rect 14588 10742 14644 10780
rect 15148 10836 15204 10846
rect 15372 10836 15428 12686
rect 15484 11844 15540 12908
rect 15596 12898 15652 12908
rect 15820 13188 15876 13198
rect 15820 12962 15876 13132
rect 15820 12910 15822 12962
rect 15874 12910 15876 12962
rect 15820 12898 15876 12910
rect 16380 12964 16436 12974
rect 16436 12908 16772 12964
rect 16380 12870 16436 12908
rect 15484 11778 15540 11788
rect 15596 12740 15652 12750
rect 15484 10836 15540 10846
rect 15372 10834 15540 10836
rect 15372 10782 15486 10834
rect 15538 10782 15540 10834
rect 15372 10780 15540 10782
rect 15148 10722 15204 10780
rect 15484 10770 15540 10780
rect 15596 10836 15652 12684
rect 15708 12738 15764 12750
rect 15708 12686 15710 12738
rect 15762 12686 15764 12738
rect 15708 12180 15764 12686
rect 16716 12404 16772 12908
rect 16940 12962 16996 13468
rect 17500 13458 17556 13468
rect 18620 13188 18676 13806
rect 18844 13188 18900 14366
rect 18956 14420 19012 14430
rect 18956 14326 19012 14364
rect 20524 14418 20580 15148
rect 20636 14644 20692 14654
rect 20636 14530 20692 14588
rect 20636 14478 20638 14530
rect 20690 14478 20692 14530
rect 20636 14466 20692 14478
rect 20524 14366 20526 14418
rect 20578 14366 20580 14418
rect 20524 14354 20580 14366
rect 19516 14308 19572 14318
rect 19516 14214 19572 14252
rect 20972 14308 21028 14318
rect 20188 13860 20244 13870
rect 20188 13766 20244 13804
rect 20972 13746 21028 14252
rect 21196 13860 21252 13870
rect 21196 13766 21252 13804
rect 20972 13694 20974 13746
rect 21026 13694 21028 13746
rect 20972 13682 21028 13694
rect 20636 13524 20692 13534
rect 20524 13522 20692 13524
rect 20524 13470 20638 13522
rect 20690 13470 20692 13522
rect 20524 13468 20692 13470
rect 19964 13188 20020 13198
rect 18620 13186 20020 13188
rect 18620 13134 19966 13186
rect 20018 13134 20020 13186
rect 18620 13132 20020 13134
rect 19964 13122 20020 13132
rect 16940 12910 16942 12962
rect 16994 12910 16996 12962
rect 16940 12898 16996 12910
rect 19180 12740 19236 12750
rect 17500 12404 17556 12414
rect 16268 12180 16324 12190
rect 15708 12178 16324 12180
rect 15708 12126 16270 12178
rect 16322 12126 16324 12178
rect 15708 12124 16324 12126
rect 16268 12114 16324 12124
rect 16716 12178 16772 12348
rect 16716 12126 16718 12178
rect 16770 12126 16772 12178
rect 16716 12114 16772 12126
rect 17388 12348 17500 12404
rect 17388 11506 17444 12348
rect 17500 12310 17556 12348
rect 17388 11454 17390 11506
rect 17442 11454 17444 11506
rect 17388 11442 17444 11454
rect 17948 12068 18004 12078
rect 16380 11284 16436 11294
rect 16380 11170 16436 11228
rect 17836 11284 17892 11294
rect 17948 11284 18004 12012
rect 19180 12068 19236 12684
rect 20300 12740 20356 12750
rect 20356 12684 20468 12740
rect 20300 12646 20356 12684
rect 20412 12402 20468 12684
rect 20412 12350 20414 12402
rect 20466 12350 20468 12402
rect 20412 12338 20468 12350
rect 19852 12180 19908 12190
rect 19852 12086 19908 12124
rect 19180 12002 19236 12012
rect 17892 11228 18004 11284
rect 17836 11190 17892 11228
rect 16380 11118 16382 11170
rect 16434 11118 16436 11170
rect 15932 10836 15988 10846
rect 15596 10834 15988 10836
rect 15596 10782 15934 10834
rect 15986 10782 15988 10834
rect 15596 10780 15988 10782
rect 15148 10670 15150 10722
rect 15202 10670 15204 10722
rect 15148 10658 15204 10670
rect 15260 10722 15316 10734
rect 15260 10670 15262 10722
rect 15314 10670 15316 10722
rect 15260 10612 15316 10670
rect 15596 10612 15652 10780
rect 15932 10770 15988 10780
rect 15260 10556 15652 10612
rect 15596 10388 15652 10398
rect 14008 9436 15208 9446
rect 14064 9434 14112 9436
rect 14168 9434 14216 9436
rect 14076 9382 14112 9434
rect 14200 9382 14216 9434
rect 14064 9380 14112 9382
rect 14168 9380 14216 9382
rect 14272 9434 14320 9436
rect 14376 9434 14424 9436
rect 14480 9434 14528 9436
rect 14376 9382 14396 9434
rect 14480 9382 14520 9434
rect 14272 9380 14320 9382
rect 14376 9380 14424 9382
rect 14480 9380 14528 9382
rect 14584 9380 14632 9436
rect 14688 9434 14736 9436
rect 14792 9434 14840 9436
rect 14896 9434 14944 9436
rect 14696 9382 14736 9434
rect 14820 9382 14840 9434
rect 14688 9380 14736 9382
rect 14792 9380 14840 9382
rect 14896 9380 14944 9382
rect 15000 9434 15048 9436
rect 15104 9434 15152 9436
rect 15000 9382 15016 9434
rect 15104 9382 15140 9434
rect 15000 9380 15048 9382
rect 15104 9380 15152 9382
rect 14008 9370 15208 9380
rect 14008 7868 15208 7878
rect 14064 7866 14112 7868
rect 14168 7866 14216 7868
rect 14076 7814 14112 7866
rect 14200 7814 14216 7866
rect 14064 7812 14112 7814
rect 14168 7812 14216 7814
rect 14272 7866 14320 7868
rect 14376 7866 14424 7868
rect 14480 7866 14528 7868
rect 14376 7814 14396 7866
rect 14480 7814 14520 7866
rect 14272 7812 14320 7814
rect 14376 7812 14424 7814
rect 14480 7812 14528 7814
rect 14584 7812 14632 7868
rect 14688 7866 14736 7868
rect 14792 7866 14840 7868
rect 14896 7866 14944 7868
rect 14696 7814 14736 7866
rect 14820 7814 14840 7866
rect 14688 7812 14736 7814
rect 14792 7812 14840 7814
rect 14896 7812 14944 7814
rect 15000 7866 15048 7868
rect 15104 7866 15152 7868
rect 15000 7814 15016 7866
rect 15104 7814 15140 7866
rect 15000 7812 15048 7814
rect 15104 7812 15152 7814
rect 14008 7802 15208 7812
rect 15596 7698 15652 10332
rect 16380 10388 16436 11118
rect 17052 11172 17108 11182
rect 17052 11078 17108 11116
rect 19740 10724 19796 10734
rect 19740 10610 19796 10668
rect 19740 10558 19742 10610
rect 19794 10558 19796 10610
rect 19740 10546 19796 10558
rect 20188 10612 20244 10622
rect 20524 10612 20580 13468
rect 20636 13458 20692 13468
rect 21308 12740 21364 17388
rect 21420 17378 21476 17388
rect 21420 17108 21476 17118
rect 21420 16882 21476 17052
rect 21420 16830 21422 16882
rect 21474 16830 21476 16882
rect 21420 16818 21476 16830
rect 21644 16884 21700 17612
rect 21868 17556 21924 17612
rect 22092 18450 22596 18452
rect 22092 18398 22542 18450
rect 22594 18398 22596 18450
rect 22092 18396 22596 18398
rect 22092 17666 22148 18396
rect 22428 18116 22484 18126
rect 22092 17614 22094 17666
rect 22146 17614 22148 17666
rect 22092 17602 22148 17614
rect 22316 17668 22372 17678
rect 22316 17574 22372 17612
rect 21868 17490 21924 17500
rect 22204 17442 22260 17454
rect 22204 17390 22206 17442
rect 22258 17390 22260 17442
rect 22204 17108 22260 17390
rect 22204 17042 22260 17052
rect 22428 17332 22484 18060
rect 22428 17106 22484 17276
rect 22428 17054 22430 17106
rect 22482 17054 22484 17106
rect 22428 17042 22484 17054
rect 22540 16996 22596 18396
rect 23212 18450 23268 19964
rect 23660 20020 23716 20030
rect 23660 19926 23716 19964
rect 23548 19908 23604 19918
rect 23548 19814 23604 19852
rect 23772 19796 23828 19806
rect 23772 18900 23828 19740
rect 23884 19458 23940 20300
rect 24220 19794 24276 20972
rect 24668 20916 24724 20926
rect 24556 20804 24612 20814
rect 24556 20710 24612 20748
rect 24668 20802 24724 20860
rect 24668 20750 24670 20802
rect 24722 20750 24724 20802
rect 24668 20738 24724 20750
rect 25228 20916 25284 20926
rect 25228 20802 25284 20860
rect 25228 20750 25230 20802
rect 25282 20750 25284 20802
rect 25228 20738 25284 20750
rect 24780 20692 24836 20702
rect 24780 20018 24836 20636
rect 24780 19966 24782 20018
rect 24834 19966 24836 20018
rect 24780 19954 24836 19966
rect 25340 20244 25396 21758
rect 25340 20018 25396 20188
rect 25452 20914 25508 20926
rect 25452 20862 25454 20914
rect 25506 20862 25508 20914
rect 25452 20132 25508 20862
rect 25564 20692 25620 26852
rect 25788 26852 26180 26908
rect 26348 27188 26404 27198
rect 25676 26180 25732 26190
rect 25788 26180 25844 26852
rect 26348 26402 26404 27132
rect 26460 27186 26516 27246
rect 26460 27134 26462 27186
rect 26514 27134 26516 27186
rect 26460 27122 26516 27134
rect 29708 27076 29764 27086
rect 29708 26982 29764 27020
rect 29932 27074 29988 31052
rect 30268 30324 30324 33070
rect 30380 31780 30436 35980
rect 30828 35364 30884 36204
rect 31388 36258 31444 36270
rect 31388 36206 31390 36258
rect 31442 36206 31444 36258
rect 31388 35700 31444 36206
rect 31388 35634 31444 35644
rect 30828 35298 30884 35308
rect 31164 35476 31220 35486
rect 30492 34132 30548 34142
rect 30492 34130 30772 34132
rect 30492 34078 30494 34130
rect 30546 34078 30772 34130
rect 30492 34076 30772 34078
rect 30492 34066 30548 34076
rect 30716 33460 30772 34076
rect 31164 34130 31220 35420
rect 31500 34132 31556 38612
rect 31724 38052 31780 38090
rect 31724 37986 31780 37996
rect 31724 37826 31780 37838
rect 31724 37774 31726 37826
rect 31778 37774 31780 37826
rect 31724 37268 31780 37774
rect 31724 37202 31780 37212
rect 31836 36932 31892 38668
rect 32060 38276 32116 39676
rect 32508 39618 32564 39676
rect 32508 39566 32510 39618
rect 32562 39566 32564 39618
rect 32508 39554 32564 39566
rect 32172 39506 32228 39518
rect 32172 39454 32174 39506
rect 32226 39454 32228 39506
rect 32172 39060 32228 39454
rect 32620 39506 32676 39518
rect 32620 39454 32622 39506
rect 32674 39454 32676 39506
rect 32284 39060 32340 39070
rect 32620 39060 32676 39454
rect 32172 39004 32284 39060
rect 32284 38946 32340 39004
rect 32508 39004 32676 39060
rect 32284 38894 32286 38946
rect 32338 38894 32340 38946
rect 32284 38882 32340 38894
rect 32396 38948 32452 38958
rect 32060 38210 32116 38220
rect 31612 36876 31892 36932
rect 31948 38164 32004 38174
rect 31948 37604 32004 38108
rect 32060 38050 32116 38062
rect 32060 37998 32062 38050
rect 32114 37998 32116 38050
rect 32060 37828 32116 37998
rect 32172 37828 32228 37838
rect 32060 37826 32228 37828
rect 32060 37774 32174 37826
rect 32226 37774 32228 37826
rect 32060 37772 32228 37774
rect 31948 37490 32004 37548
rect 31948 37438 31950 37490
rect 32002 37438 32004 37490
rect 31612 36370 31668 36876
rect 31948 36482 32004 37438
rect 32172 36596 32228 37772
rect 32172 36530 32228 36540
rect 32396 37826 32452 38892
rect 32508 38668 32564 39004
rect 32620 38836 32676 38846
rect 32620 38742 32676 38780
rect 32508 38612 32676 38668
rect 32620 38052 32676 38612
rect 32396 37774 32398 37826
rect 32450 37774 32452 37826
rect 32396 36932 32452 37774
rect 32508 37938 32564 37950
rect 32508 37886 32510 37938
rect 32562 37886 32564 37938
rect 32508 37268 32564 37886
rect 32508 37202 32564 37212
rect 31948 36430 31950 36482
rect 32002 36430 32004 36482
rect 31612 36318 31614 36370
rect 31666 36318 31668 36370
rect 31612 36306 31668 36318
rect 31724 36372 31780 36382
rect 31724 36278 31780 36316
rect 31724 36148 31780 36158
rect 31724 35476 31780 36092
rect 31724 35410 31780 35420
rect 31836 35812 31892 35822
rect 31948 35812 32004 36430
rect 32172 36370 32228 36382
rect 32172 36318 32174 36370
rect 32226 36318 32228 36370
rect 32172 36148 32228 36318
rect 32172 36082 32228 36092
rect 32396 35924 32452 36876
rect 32396 35858 32452 35868
rect 32620 36370 32676 37996
rect 32620 36318 32622 36370
rect 32674 36318 32676 36370
rect 31948 35756 32340 35812
rect 31836 35698 31892 35756
rect 31836 35646 31838 35698
rect 31890 35646 31892 35698
rect 31164 34078 31166 34130
rect 31218 34078 31220 34130
rect 31164 34066 31220 34078
rect 31276 34130 31556 34132
rect 31276 34078 31502 34130
rect 31554 34078 31556 34130
rect 31276 34076 31556 34078
rect 30716 33404 31220 33460
rect 31164 33346 31220 33404
rect 31164 33294 31166 33346
rect 31218 33294 31220 33346
rect 31164 33282 31220 33294
rect 30940 33122 30996 33134
rect 31276 33124 31332 34076
rect 31500 34066 31556 34076
rect 31612 35364 31668 35374
rect 31612 33908 31668 35308
rect 31836 35252 31892 35646
rect 31948 35586 32004 35598
rect 31948 35534 31950 35586
rect 32002 35534 32004 35586
rect 31948 35476 32004 35534
rect 32172 35476 32228 35486
rect 31948 35410 32004 35420
rect 32060 35420 32172 35476
rect 31836 35196 32004 35252
rect 31724 34020 31780 34030
rect 31724 34018 31892 34020
rect 31724 33966 31726 34018
rect 31778 33966 31892 34018
rect 31724 33964 31892 33966
rect 31724 33954 31780 33964
rect 31500 33852 31668 33908
rect 30940 33070 30942 33122
rect 30994 33070 30996 33122
rect 30940 33012 30996 33070
rect 30940 32946 30996 32956
rect 31052 33068 31332 33124
rect 31388 33572 31444 33582
rect 30940 32676 30996 32686
rect 31052 32676 31108 33068
rect 31164 32788 31220 32798
rect 31164 32694 31220 32732
rect 31388 32786 31444 33516
rect 31388 32734 31390 32786
rect 31442 32734 31444 32786
rect 30604 32674 31108 32676
rect 30604 32622 30942 32674
rect 30994 32622 31108 32674
rect 30604 32620 31108 32622
rect 31388 32676 31444 32734
rect 30380 31724 30548 31780
rect 30380 31554 30436 31566
rect 30380 31502 30382 31554
rect 30434 31502 30436 31554
rect 30380 31444 30436 31502
rect 30492 31556 30548 31724
rect 30604 31778 30660 32620
rect 30940 32610 30996 32620
rect 31388 32610 31444 32620
rect 30604 31726 30606 31778
rect 30658 31726 30660 31778
rect 30604 31714 30660 31726
rect 31052 32338 31108 32350
rect 31052 32286 31054 32338
rect 31106 32286 31108 32338
rect 31052 31778 31108 32286
rect 31052 31726 31054 31778
rect 31106 31726 31108 31778
rect 31052 31714 31108 31726
rect 30940 31666 30996 31678
rect 30940 31614 30942 31666
rect 30994 31614 30996 31666
rect 30492 31500 30660 31556
rect 30380 31378 30436 31388
rect 30492 31108 30548 31118
rect 30492 31014 30548 31052
rect 30604 30996 30660 31500
rect 30940 30996 30996 31614
rect 31500 31332 31556 33852
rect 31836 33346 31892 33964
rect 31948 33572 32004 35196
rect 31948 33506 32004 33516
rect 31836 33294 31838 33346
rect 31890 33294 31892 33346
rect 31836 33282 31892 33294
rect 31612 33122 31668 33134
rect 31612 33070 31614 33122
rect 31666 33070 31668 33122
rect 31612 33012 31668 33070
rect 31612 32946 31668 32956
rect 31724 33122 31780 33134
rect 31724 33070 31726 33122
rect 31778 33070 31780 33122
rect 31612 31778 31668 31790
rect 31612 31726 31614 31778
rect 31666 31726 31668 31778
rect 31612 31556 31668 31726
rect 31612 31490 31668 31500
rect 31500 31276 31668 31332
rect 31164 30996 31220 31006
rect 30604 30994 30884 30996
rect 30604 30942 30606 30994
rect 30658 30942 30884 30994
rect 30604 30940 30884 30942
rect 30940 30994 31220 30996
rect 30940 30942 31166 30994
rect 31218 30942 31220 30994
rect 30940 30940 31220 30942
rect 30604 30930 30660 30940
rect 30268 30258 30324 30268
rect 30716 30434 30772 30446
rect 30716 30382 30718 30434
rect 30770 30382 30772 30434
rect 30380 30098 30436 30110
rect 30380 30046 30382 30098
rect 30434 30046 30436 30098
rect 30268 29428 30324 29438
rect 30044 27972 30100 27982
rect 30044 27878 30100 27916
rect 29932 27022 29934 27074
rect 29986 27022 29988 27074
rect 29932 27010 29988 27022
rect 30156 27636 30212 27646
rect 30156 27076 30212 27580
rect 30156 27010 30212 27020
rect 30268 27074 30324 29372
rect 30380 29204 30436 30046
rect 30604 29204 30660 29214
rect 30380 29202 30660 29204
rect 30380 29150 30606 29202
rect 30658 29150 30660 29202
rect 30380 29148 30660 29150
rect 30268 27022 30270 27074
rect 30322 27022 30324 27074
rect 29372 26962 29428 26974
rect 29372 26910 29374 26962
rect 29426 26910 29428 26962
rect 26348 26350 26350 26402
rect 26402 26350 26404 26402
rect 26348 26338 26404 26350
rect 26460 26402 26516 26414
rect 26460 26350 26462 26402
rect 26514 26350 26516 26402
rect 26012 26180 26068 26190
rect 26460 26180 26516 26350
rect 25788 26178 26516 26180
rect 25788 26126 26014 26178
rect 26066 26126 26516 26178
rect 25788 26124 26516 26126
rect 26684 26290 26740 26302
rect 26684 26238 26686 26290
rect 26738 26238 26740 26290
rect 25676 20916 25732 26124
rect 26012 24836 26068 26124
rect 26684 25956 26740 26238
rect 29260 26180 29316 26190
rect 29260 26086 29316 26124
rect 29372 26066 29428 26910
rect 29820 26852 29876 26862
rect 29820 26758 29876 26796
rect 29372 26014 29374 26066
rect 29426 26014 29428 26066
rect 29372 26002 29428 26014
rect 29596 26292 29652 26302
rect 26684 25900 27076 25956
rect 26796 25508 26852 25518
rect 26124 25506 26852 25508
rect 26124 25454 26798 25506
rect 26850 25454 26852 25506
rect 26124 25452 26852 25454
rect 26124 24946 26180 25452
rect 26796 25442 26852 25452
rect 26796 25172 26852 25182
rect 26124 24894 26126 24946
rect 26178 24894 26180 24946
rect 26124 24882 26180 24894
rect 26684 25060 26740 25070
rect 26684 24946 26740 25004
rect 26684 24894 26686 24946
rect 26738 24894 26740 24946
rect 26684 24882 26740 24894
rect 26012 24770 26068 24780
rect 26460 24722 26516 24734
rect 26460 24670 26462 24722
rect 26514 24670 26516 24722
rect 25788 24612 25844 24622
rect 25788 24518 25844 24556
rect 26012 24498 26068 24510
rect 26012 24446 26014 24498
rect 26066 24446 26068 24498
rect 26012 24164 26068 24446
rect 26012 24098 26068 24108
rect 26348 23154 26404 23166
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 25788 22258 25844 22270
rect 25788 22206 25790 22258
rect 25842 22206 25844 22258
rect 25788 21028 25844 22206
rect 26348 22148 26404 23102
rect 26348 22082 26404 22092
rect 26460 22036 26516 24670
rect 26684 24500 26740 24510
rect 26684 23716 26740 24444
rect 26684 23042 26740 23660
rect 26684 22990 26686 23042
rect 26738 22990 26740 23042
rect 26684 22978 26740 22990
rect 26236 21700 26292 21710
rect 26460 21700 26516 21980
rect 26796 21812 26852 25116
rect 27020 25172 27076 25900
rect 27020 25106 27076 25116
rect 27356 25732 27412 25742
rect 27132 24948 27188 24958
rect 27132 24834 27188 24892
rect 27132 24782 27134 24834
rect 27186 24782 27188 24834
rect 27132 24770 27188 24782
rect 27244 24836 27300 24846
rect 27356 24836 27412 25676
rect 29372 25620 29428 25630
rect 29596 25620 29652 26236
rect 27468 25506 27524 25518
rect 29372 25508 29428 25564
rect 27468 25454 27470 25506
rect 27522 25454 27524 25506
rect 27468 25284 27524 25454
rect 29148 25506 29428 25508
rect 29148 25454 29374 25506
rect 29426 25454 29428 25506
rect 29148 25452 29428 25454
rect 27468 25218 27524 25228
rect 27580 25396 27636 25406
rect 27468 24836 27524 24846
rect 27356 24834 27524 24836
rect 27356 24782 27470 24834
rect 27522 24782 27524 24834
rect 27356 24780 27524 24782
rect 26908 24722 26964 24734
rect 26908 24670 26910 24722
rect 26962 24670 26964 24722
rect 26908 22596 26964 24670
rect 27020 24498 27076 24510
rect 27020 24446 27022 24498
rect 27074 24446 27076 24498
rect 27020 23940 27076 24446
rect 27244 24052 27300 24780
rect 27468 24770 27524 24780
rect 27244 23986 27300 23996
rect 27020 23874 27076 23884
rect 27020 23716 27076 23726
rect 27020 23266 27076 23660
rect 27580 23380 27636 25340
rect 27916 25396 27972 25406
rect 27916 25302 27972 25340
rect 28252 25284 28308 25294
rect 27804 24724 27860 24734
rect 27804 24630 27860 24668
rect 28140 24722 28196 24734
rect 28140 24670 28142 24722
rect 28194 24670 28196 24722
rect 27916 24612 27972 24622
rect 27916 24518 27972 24556
rect 27804 24220 28084 24276
rect 27804 24050 27860 24220
rect 27804 23998 27806 24050
rect 27858 23998 27860 24050
rect 27804 23986 27860 23998
rect 27916 24052 27972 24062
rect 27580 23314 27636 23324
rect 27804 23604 27860 23614
rect 27020 23214 27022 23266
rect 27074 23214 27076 23266
rect 27020 23202 27076 23214
rect 26908 22530 26964 22540
rect 27580 22930 27636 22942
rect 27580 22878 27582 22930
rect 27634 22878 27636 22930
rect 27580 22596 27636 22878
rect 27244 22482 27300 22494
rect 27244 22430 27246 22482
rect 27298 22430 27300 22482
rect 26796 21746 26852 21756
rect 27020 22148 27076 22158
rect 26236 21698 26516 21700
rect 26236 21646 26238 21698
rect 26290 21646 26516 21698
rect 26236 21644 26516 21646
rect 26236 21634 26292 21644
rect 27020 21586 27076 22092
rect 27020 21534 27022 21586
rect 27074 21534 27076 21586
rect 27020 21522 27076 21534
rect 25788 20962 25844 20972
rect 25676 20850 25732 20860
rect 25564 20636 26292 20692
rect 25452 20066 25508 20076
rect 25788 20130 25844 20142
rect 25788 20078 25790 20130
rect 25842 20078 25844 20130
rect 25340 19966 25342 20018
rect 25394 19966 25396 20018
rect 25340 19954 25396 19966
rect 25564 20020 25620 20030
rect 25620 19964 25732 20020
rect 25564 19954 25620 19964
rect 24220 19742 24222 19794
rect 24274 19742 24276 19794
rect 24220 19730 24276 19742
rect 25676 19684 25732 19964
rect 24008 19628 25208 19638
rect 24064 19626 24112 19628
rect 24168 19626 24216 19628
rect 24076 19574 24112 19626
rect 24200 19574 24216 19626
rect 24064 19572 24112 19574
rect 24168 19572 24216 19574
rect 24272 19626 24320 19628
rect 24376 19626 24424 19628
rect 24480 19626 24528 19628
rect 24376 19574 24396 19626
rect 24480 19574 24520 19626
rect 24272 19572 24320 19574
rect 24376 19572 24424 19574
rect 24480 19572 24528 19574
rect 24584 19572 24632 19628
rect 24688 19626 24736 19628
rect 24792 19626 24840 19628
rect 24896 19626 24944 19628
rect 24696 19574 24736 19626
rect 24820 19574 24840 19626
rect 24688 19572 24736 19574
rect 24792 19572 24840 19574
rect 24896 19572 24944 19574
rect 25000 19626 25048 19628
rect 25104 19626 25152 19628
rect 25000 19574 25016 19626
rect 25104 19574 25140 19626
rect 25000 19572 25048 19574
rect 25104 19572 25152 19574
rect 24008 19562 25208 19572
rect 23884 19406 23886 19458
rect 23938 19406 23940 19458
rect 23884 19394 23940 19406
rect 24668 19458 24724 19470
rect 24668 19406 24670 19458
rect 24722 19406 24724 19458
rect 24668 19346 24724 19406
rect 24668 19294 24670 19346
rect 24722 19294 24724 19346
rect 24668 19282 24724 19294
rect 25116 19236 25172 19246
rect 25116 19142 25172 19180
rect 25676 19234 25732 19628
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25676 19170 25732 19182
rect 24220 19010 24276 19022
rect 24220 18958 24222 19010
rect 24274 18958 24276 19010
rect 24220 18900 24276 18958
rect 23772 18844 24276 18900
rect 23772 18676 23828 18686
rect 23212 18398 23214 18450
rect 23266 18398 23268 18450
rect 22652 18228 22708 18238
rect 22652 17666 22708 18172
rect 22652 17614 22654 17666
rect 22706 17614 22708 17666
rect 22652 17602 22708 17614
rect 23100 18226 23156 18238
rect 23100 18174 23102 18226
rect 23154 18174 23156 18226
rect 23100 17892 23156 18174
rect 23212 18116 23268 18398
rect 23212 18050 23268 18060
rect 23660 18620 23772 18676
rect 23100 17836 23492 17892
rect 23100 17668 23156 17836
rect 23100 17602 23156 17612
rect 23324 17666 23380 17678
rect 23324 17614 23326 17666
rect 23378 17614 23380 17666
rect 22764 17556 22820 17566
rect 22764 17462 22820 17500
rect 22988 17444 23044 17454
rect 22988 17442 23156 17444
rect 22988 17390 22990 17442
rect 23042 17390 23156 17442
rect 22988 17388 23156 17390
rect 22988 17378 23044 17388
rect 23100 17220 23156 17388
rect 23324 17220 23380 17614
rect 23436 17668 23492 17836
rect 23548 17668 23604 17678
rect 23436 17666 23604 17668
rect 23436 17614 23550 17666
rect 23602 17614 23604 17666
rect 23436 17612 23604 17614
rect 23548 17602 23604 17612
rect 23100 17164 23324 17220
rect 23324 17126 23380 17164
rect 23548 17444 23604 17454
rect 22540 16930 22596 16940
rect 22652 16994 22708 17006
rect 22652 16942 22654 16994
rect 22706 16942 22708 16994
rect 21644 16322 21700 16828
rect 21644 16270 21646 16322
rect 21698 16270 21700 16322
rect 21644 16258 21700 16270
rect 22092 16882 22148 16894
rect 22092 16830 22094 16882
rect 22146 16830 22148 16882
rect 21644 15988 21700 15998
rect 21644 15538 21700 15932
rect 21644 15486 21646 15538
rect 21698 15486 21700 15538
rect 21644 14754 21700 15486
rect 21756 15988 21812 15998
rect 22092 15988 22148 16830
rect 22652 16884 22708 16942
rect 23212 16996 23268 17006
rect 23212 16902 23268 16940
rect 22652 16818 22708 16828
rect 23324 16884 23380 16894
rect 23380 16828 23492 16884
rect 23324 16790 23380 16828
rect 22316 16772 22372 16782
rect 22316 16678 22372 16716
rect 23436 16100 23492 16828
rect 23548 16212 23604 17388
rect 23660 17442 23716 18620
rect 23772 18610 23828 18620
rect 23884 17892 23940 18844
rect 25788 18676 25844 20078
rect 25788 18610 25844 18620
rect 26124 19458 26180 19470
rect 26124 19406 26126 19458
rect 26178 19406 26180 19458
rect 24008 18060 25208 18070
rect 24064 18058 24112 18060
rect 24168 18058 24216 18060
rect 24076 18006 24112 18058
rect 24200 18006 24216 18058
rect 24064 18004 24112 18006
rect 24168 18004 24216 18006
rect 24272 18058 24320 18060
rect 24376 18058 24424 18060
rect 24480 18058 24528 18060
rect 24376 18006 24396 18058
rect 24480 18006 24520 18058
rect 24272 18004 24320 18006
rect 24376 18004 24424 18006
rect 24480 18004 24528 18006
rect 24584 18004 24632 18060
rect 24688 18058 24736 18060
rect 24792 18058 24840 18060
rect 24896 18058 24944 18060
rect 24696 18006 24736 18058
rect 24820 18006 24840 18058
rect 24688 18004 24736 18006
rect 24792 18004 24840 18006
rect 24896 18004 24944 18006
rect 25000 18058 25048 18060
rect 25104 18058 25152 18060
rect 25000 18006 25016 18058
rect 25104 18006 25140 18058
rect 25000 18004 25048 18006
rect 25104 18004 25152 18006
rect 24008 17994 25208 18004
rect 23884 17836 24052 17892
rect 23660 17390 23662 17442
rect 23714 17390 23716 17442
rect 23660 17378 23716 17390
rect 23772 17666 23828 17678
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 23660 16996 23716 17006
rect 23660 16902 23716 16940
rect 23772 16884 23828 17614
rect 23884 17332 23940 17342
rect 23884 17106 23940 17276
rect 23884 17054 23886 17106
rect 23938 17054 23940 17106
rect 23884 17042 23940 17054
rect 23996 16884 24052 17836
rect 24892 17444 24948 17454
rect 24948 17388 25284 17444
rect 24892 17350 24948 17388
rect 24220 17220 24276 17230
rect 24108 17108 24164 17118
rect 24108 17014 24164 17052
rect 23772 16818 23828 16828
rect 23884 16828 24052 16884
rect 24220 16882 24276 17164
rect 25228 17220 25284 17388
rect 25228 16994 25284 17164
rect 25564 17108 25620 17118
rect 25228 16942 25230 16994
rect 25282 16942 25284 16994
rect 25228 16930 25284 16942
rect 25340 17106 25620 17108
rect 25340 17054 25566 17106
rect 25618 17054 25620 17106
rect 25340 17052 25620 17054
rect 24220 16830 24222 16882
rect 24274 16830 24276 16882
rect 23772 16660 23828 16670
rect 23772 16566 23828 16604
rect 23772 16212 23828 16222
rect 23548 16210 23828 16212
rect 23548 16158 23774 16210
rect 23826 16158 23828 16210
rect 23548 16156 23828 16158
rect 23436 16044 23604 16100
rect 21756 15986 22148 15988
rect 21756 15934 21758 15986
rect 21810 15934 22148 15986
rect 21756 15932 22148 15934
rect 21756 15204 21812 15932
rect 22204 15874 22260 15886
rect 22204 15822 22206 15874
rect 22258 15822 22260 15874
rect 22204 15540 22260 15822
rect 22204 15474 22260 15484
rect 22652 15876 22708 15886
rect 22316 15316 22372 15326
rect 22652 15316 22708 15820
rect 22372 15260 22708 15316
rect 22988 15540 23044 15550
rect 22988 15314 23044 15484
rect 22988 15262 22990 15314
rect 23042 15262 23044 15314
rect 21756 15138 21812 15148
rect 22204 15204 22260 15242
rect 22204 15138 22260 15148
rect 21644 14702 21646 14754
rect 21698 14702 21700 14754
rect 21644 14690 21700 14702
rect 21980 14644 22036 14654
rect 21980 14550 22036 14588
rect 21756 13858 21812 13870
rect 21756 13806 21758 13858
rect 21810 13806 21812 13858
rect 21756 12964 21812 13806
rect 21756 12898 21812 12908
rect 21308 12674 21364 12684
rect 20188 10610 20580 10612
rect 20188 10558 20190 10610
rect 20242 10558 20580 10610
rect 20188 10556 20580 10558
rect 22316 11394 22372 15260
rect 22988 15250 23044 15262
rect 23212 15426 23268 15438
rect 23212 15374 23214 15426
rect 23266 15374 23268 15426
rect 22652 15090 22708 15102
rect 22652 15038 22654 15090
rect 22706 15038 22708 15090
rect 22428 14754 22484 14766
rect 22428 14702 22430 14754
rect 22482 14702 22484 14754
rect 22428 14308 22484 14702
rect 22428 14306 22596 14308
rect 22428 14254 22430 14306
rect 22482 14254 22596 14306
rect 22428 14252 22596 14254
rect 22428 14242 22484 14252
rect 22428 13860 22484 13870
rect 22428 13076 22484 13804
rect 22428 12982 22484 13020
rect 22540 12180 22596 14252
rect 22652 13188 22708 15038
rect 23212 14644 23268 15374
rect 23548 15426 23604 16044
rect 23772 15652 23828 16156
rect 23884 15876 23940 16828
rect 24220 16818 24276 16830
rect 24008 16492 25208 16502
rect 24064 16490 24112 16492
rect 24168 16490 24216 16492
rect 24076 16438 24112 16490
rect 24200 16438 24216 16490
rect 24064 16436 24112 16438
rect 24168 16436 24216 16438
rect 24272 16490 24320 16492
rect 24376 16490 24424 16492
rect 24480 16490 24528 16492
rect 24376 16438 24396 16490
rect 24480 16438 24520 16490
rect 24272 16436 24320 16438
rect 24376 16436 24424 16438
rect 24480 16436 24528 16438
rect 24584 16436 24632 16492
rect 24688 16490 24736 16492
rect 24792 16490 24840 16492
rect 24896 16490 24944 16492
rect 24696 16438 24736 16490
rect 24820 16438 24840 16490
rect 24688 16436 24736 16438
rect 24792 16436 24840 16438
rect 24896 16436 24944 16438
rect 25000 16490 25048 16492
rect 25104 16490 25152 16492
rect 25000 16438 25016 16490
rect 25104 16438 25140 16490
rect 25000 16436 25048 16438
rect 25104 16436 25152 16438
rect 24008 16426 25208 16436
rect 25340 16324 25396 17052
rect 25564 17042 25620 17052
rect 26124 16996 26180 19406
rect 26236 18340 26292 20636
rect 26796 20132 26852 20142
rect 26348 20130 26852 20132
rect 26348 20078 26798 20130
rect 26850 20078 26852 20130
rect 26348 20076 26852 20078
rect 26348 19234 26404 20076
rect 26796 20066 26852 20076
rect 27020 19906 27076 19918
rect 27020 19854 27022 19906
rect 27074 19854 27076 19906
rect 26908 19460 26964 19470
rect 26908 19366 26964 19404
rect 26348 19182 26350 19234
rect 26402 19182 26404 19234
rect 26348 18564 26404 19182
rect 26460 19124 26516 19134
rect 26796 19124 26852 19134
rect 26460 19030 26516 19068
rect 26684 19122 26852 19124
rect 26684 19070 26798 19122
rect 26850 19070 26852 19122
rect 26684 19068 26852 19070
rect 26348 18498 26404 18508
rect 26236 18284 26404 18340
rect 26236 17556 26292 17566
rect 26236 17106 26292 17500
rect 26236 17054 26238 17106
rect 26290 17054 26292 17106
rect 26236 17042 26292 17054
rect 25900 16994 26180 16996
rect 25900 16942 26126 16994
rect 26178 16942 26180 16994
rect 25900 16940 26180 16942
rect 25452 16884 25508 16894
rect 25452 16790 25508 16828
rect 25900 16882 25956 16940
rect 26124 16930 26180 16940
rect 25900 16830 25902 16882
rect 25954 16830 25956 16882
rect 25900 16818 25956 16830
rect 26236 16660 26292 16670
rect 25900 16658 26292 16660
rect 25900 16606 26238 16658
rect 26290 16606 26292 16658
rect 25900 16604 26292 16606
rect 24780 16268 25396 16324
rect 25788 16324 25844 16334
rect 24556 16212 24612 16222
rect 24332 16100 24388 16110
rect 23884 15810 23940 15820
rect 24108 16098 24388 16100
rect 24108 16046 24334 16098
rect 24386 16046 24388 16098
rect 24108 16044 24388 16046
rect 24108 15652 24164 16044
rect 24332 16034 24388 16044
rect 24556 16098 24612 16156
rect 24556 16046 24558 16098
rect 24610 16046 24612 16098
rect 24556 16034 24612 16046
rect 24780 16098 24836 16268
rect 24780 16046 24782 16098
rect 24834 16046 24836 16098
rect 24780 16034 24836 16046
rect 25788 16098 25844 16268
rect 25788 16046 25790 16098
rect 25842 16046 25844 16098
rect 25788 16034 25844 16046
rect 25116 15988 25172 15998
rect 25116 15894 25172 15932
rect 23772 15596 24164 15652
rect 24220 15874 24276 15886
rect 24220 15822 24222 15874
rect 24274 15822 24276 15874
rect 23548 15374 23550 15426
rect 23602 15374 23604 15426
rect 23548 15148 23604 15374
rect 23548 15092 23940 15148
rect 23212 14578 23268 14588
rect 23772 14980 23828 14990
rect 23212 13188 23268 13198
rect 22652 13186 23268 13188
rect 22652 13134 23214 13186
rect 23266 13134 23268 13186
rect 22652 13132 23268 13134
rect 23212 13122 23268 13132
rect 23772 13188 23828 14924
rect 23884 14754 23940 15092
rect 24220 15092 24276 15822
rect 24220 15026 24276 15036
rect 24444 15874 24500 15886
rect 24444 15822 24446 15874
rect 24498 15822 24500 15874
rect 24444 15092 24500 15822
rect 25228 15874 25284 15886
rect 25228 15822 25230 15874
rect 25282 15822 25284 15874
rect 25228 15148 25284 15822
rect 25340 15876 25396 15886
rect 25900 15876 25956 16604
rect 26236 16594 26292 16604
rect 25340 15782 25396 15820
rect 25788 15820 25956 15876
rect 25564 15316 25620 15326
rect 25564 15222 25620 15260
rect 25228 15092 25508 15148
rect 24444 15026 24500 15036
rect 24008 14924 25208 14934
rect 24064 14922 24112 14924
rect 24168 14922 24216 14924
rect 24076 14870 24112 14922
rect 24200 14870 24216 14922
rect 24064 14868 24112 14870
rect 24168 14868 24216 14870
rect 24272 14922 24320 14924
rect 24376 14922 24424 14924
rect 24480 14922 24528 14924
rect 24376 14870 24396 14922
rect 24480 14870 24520 14922
rect 24272 14868 24320 14870
rect 24376 14868 24424 14870
rect 24480 14868 24528 14870
rect 24584 14868 24632 14924
rect 24688 14922 24736 14924
rect 24792 14922 24840 14924
rect 24896 14922 24944 14924
rect 24696 14870 24736 14922
rect 24820 14870 24840 14922
rect 24688 14868 24736 14870
rect 24792 14868 24840 14870
rect 24896 14868 24944 14870
rect 25000 14922 25048 14924
rect 25104 14922 25152 14924
rect 25000 14870 25016 14922
rect 25104 14870 25140 14922
rect 25000 14868 25048 14870
rect 25104 14868 25152 14870
rect 24008 14858 25208 14868
rect 23884 14702 23886 14754
rect 23938 14702 23940 14754
rect 23884 14690 23940 14702
rect 24668 14306 24724 14318
rect 24668 14254 24670 14306
rect 24722 14254 24724 14306
rect 24668 13748 24724 14254
rect 25452 13748 25508 15092
rect 25788 13970 25844 15820
rect 25788 13918 25790 13970
rect 25842 13918 25844 13970
rect 25788 13906 25844 13918
rect 25900 15314 25956 15326
rect 25900 15262 25902 15314
rect 25954 15262 25956 15314
rect 25900 13970 25956 15262
rect 25900 13918 25902 13970
rect 25954 13918 25956 13970
rect 25900 13906 25956 13918
rect 26012 13748 26068 13758
rect 25452 13746 26068 13748
rect 25452 13694 26014 13746
rect 26066 13694 26068 13746
rect 25452 13692 26068 13694
rect 24668 13682 24724 13692
rect 26012 13682 26068 13692
rect 26124 13636 26180 13646
rect 24008 13356 25208 13366
rect 24064 13354 24112 13356
rect 24168 13354 24216 13356
rect 24076 13302 24112 13354
rect 24200 13302 24216 13354
rect 24064 13300 24112 13302
rect 24168 13300 24216 13302
rect 24272 13354 24320 13356
rect 24376 13354 24424 13356
rect 24480 13354 24528 13356
rect 24376 13302 24396 13354
rect 24480 13302 24520 13354
rect 24272 13300 24320 13302
rect 24376 13300 24424 13302
rect 24480 13300 24528 13302
rect 24584 13300 24632 13356
rect 24688 13354 24736 13356
rect 24792 13354 24840 13356
rect 24896 13354 24944 13356
rect 24696 13302 24736 13354
rect 24820 13302 24840 13354
rect 24688 13300 24736 13302
rect 24792 13300 24840 13302
rect 24896 13300 24944 13302
rect 25000 13354 25048 13356
rect 25104 13354 25152 13356
rect 25000 13302 25016 13354
rect 25104 13302 25140 13354
rect 25000 13300 25048 13302
rect 25104 13300 25152 13302
rect 24008 13290 25208 13300
rect 23772 13122 23828 13132
rect 24556 13188 24612 13198
rect 26124 13188 26180 13580
rect 24556 13094 24612 13132
rect 25788 13132 26180 13188
rect 23436 13076 23492 13086
rect 23212 12964 23268 12974
rect 22428 12068 22484 12078
rect 22540 12068 22596 12124
rect 22428 12066 22596 12068
rect 22428 12014 22430 12066
rect 22482 12014 22596 12066
rect 22428 12012 22596 12014
rect 22428 12002 22484 12012
rect 22316 11342 22318 11394
rect 22370 11342 22372 11394
rect 22316 10724 22372 11342
rect 22540 10836 22596 12012
rect 22876 12738 22932 12750
rect 22876 12686 22878 12738
rect 22930 12686 22932 12738
rect 22764 11396 22820 11406
rect 22876 11396 22932 12686
rect 22764 11394 22932 11396
rect 22764 11342 22766 11394
rect 22818 11342 22932 11394
rect 22764 11340 22932 11342
rect 22764 11330 22820 11340
rect 22540 10742 22596 10780
rect 23212 10834 23268 12908
rect 23436 12850 23492 13020
rect 24444 12964 24500 12974
rect 24444 12870 24500 12908
rect 23436 12798 23438 12850
rect 23490 12798 23492 12850
rect 23436 12786 23492 12798
rect 23996 12852 24052 12862
rect 23996 12758 24052 12796
rect 25788 12852 25844 13132
rect 26348 13076 26404 18284
rect 26572 17220 26628 17230
rect 26572 15148 26628 17164
rect 26684 17108 26740 19068
rect 26796 19058 26852 19068
rect 26796 18564 26852 18574
rect 26796 18470 26852 18508
rect 26684 15988 26740 17052
rect 26796 17556 26852 17566
rect 26796 17106 26852 17500
rect 26796 17054 26798 17106
rect 26850 17054 26852 17106
rect 26796 16322 26852 17054
rect 27020 16996 27076 19854
rect 27244 19684 27300 22430
rect 27356 22484 27412 22494
rect 27356 22370 27412 22428
rect 27356 22318 27358 22370
rect 27410 22318 27412 22370
rect 27356 22260 27412 22318
rect 27356 22194 27412 22204
rect 27580 22036 27636 22540
rect 27580 21970 27636 21980
rect 27692 21364 27748 21374
rect 27468 20914 27524 20926
rect 27468 20862 27470 20914
rect 27522 20862 27524 20914
rect 27244 19618 27300 19628
rect 27356 20804 27412 20814
rect 27132 19236 27188 19246
rect 27132 18676 27188 19180
rect 27356 19234 27412 20748
rect 27356 19182 27358 19234
rect 27410 19182 27412 19234
rect 27356 19170 27412 19182
rect 27468 19684 27524 20862
rect 27468 19236 27524 19628
rect 27468 19170 27524 19180
rect 27692 19234 27748 21308
rect 27804 20802 27860 23548
rect 27804 20750 27806 20802
rect 27858 20750 27860 20802
rect 27804 19460 27860 20750
rect 27804 19394 27860 19404
rect 27916 19236 27972 23996
rect 28028 23716 28084 24220
rect 28140 23940 28196 24670
rect 28140 23874 28196 23884
rect 28252 23716 28308 25228
rect 28812 25172 28868 25182
rect 28868 25116 28980 25172
rect 28812 25106 28868 25116
rect 28476 24948 28532 24958
rect 28476 24854 28532 24892
rect 28812 24724 28868 24734
rect 28812 24630 28868 24668
rect 28924 23940 28980 25116
rect 29148 24948 29204 25452
rect 29372 25442 29428 25452
rect 29484 25618 29652 25620
rect 29484 25566 29598 25618
rect 29650 25566 29652 25618
rect 29484 25564 29652 25566
rect 29148 24882 29204 24892
rect 29372 24724 29428 24734
rect 29484 24724 29540 25564
rect 29596 25554 29652 25564
rect 29708 26178 29764 26190
rect 29708 26126 29710 26178
rect 29762 26126 29764 26178
rect 29708 25508 29764 26126
rect 29820 26068 29876 26078
rect 29820 26066 29988 26068
rect 29820 26014 29822 26066
rect 29874 26014 29988 26066
rect 29820 26012 29988 26014
rect 29820 26002 29876 26012
rect 29708 25442 29764 25452
rect 29932 25060 29988 26012
rect 30156 25620 30212 25630
rect 29932 24946 29988 25004
rect 29932 24894 29934 24946
rect 29986 24894 29988 24946
rect 29372 24722 29484 24724
rect 29372 24670 29374 24722
rect 29426 24670 29484 24722
rect 29372 24668 29484 24670
rect 29036 23940 29092 23950
rect 28924 23938 29092 23940
rect 28924 23886 29038 23938
rect 29090 23886 29092 23938
rect 28924 23884 29092 23886
rect 29036 23874 29092 23884
rect 29148 23940 29204 23950
rect 28476 23716 28532 23726
rect 28028 23714 28532 23716
rect 28028 23662 28478 23714
rect 28530 23662 28532 23714
rect 28028 23660 28532 23662
rect 28476 23604 28532 23660
rect 28476 23548 28644 23604
rect 28140 23380 28196 23390
rect 28140 23286 28196 23324
rect 28140 22596 28196 22606
rect 28140 22502 28196 22540
rect 28588 21924 28644 23548
rect 29148 22594 29204 23884
rect 29372 23604 29428 24668
rect 29484 24630 29540 24668
rect 29596 24722 29652 24734
rect 29596 24670 29598 24722
rect 29650 24670 29652 24722
rect 29596 24612 29652 24670
rect 29596 24546 29652 24556
rect 29484 24052 29540 24062
rect 29484 23938 29540 23996
rect 29484 23886 29486 23938
rect 29538 23886 29540 23938
rect 29484 23874 29540 23886
rect 29372 23538 29428 23548
rect 29596 23714 29652 23726
rect 29596 23662 29598 23714
rect 29650 23662 29652 23714
rect 29596 23380 29652 23662
rect 29708 23716 29764 23726
rect 29708 23622 29764 23660
rect 29596 23314 29652 23324
rect 29148 22542 29150 22594
rect 29202 22542 29204 22594
rect 29148 22530 29204 22542
rect 29484 22484 29540 22494
rect 29540 22428 29876 22484
rect 29484 22390 29540 22428
rect 28588 21858 28644 21868
rect 28924 22372 28980 22382
rect 28924 21700 28980 22316
rect 29708 22260 29764 22270
rect 29596 22204 29708 22260
rect 29260 22148 29316 22158
rect 29260 22054 29316 22092
rect 29148 21812 29204 21822
rect 28924 21698 29092 21700
rect 28924 21646 28926 21698
rect 28978 21646 29092 21698
rect 28924 21644 29092 21646
rect 28924 21634 28980 21644
rect 28588 21586 28644 21598
rect 28588 21534 28590 21586
rect 28642 21534 28644 21586
rect 28252 21362 28308 21374
rect 28252 21310 28254 21362
rect 28306 21310 28308 21362
rect 28252 20804 28308 21310
rect 28588 20916 28644 21534
rect 28588 20850 28644 20860
rect 28252 20710 28308 20748
rect 28028 20020 28084 20030
rect 28028 19346 28084 19964
rect 28028 19294 28030 19346
rect 28082 19294 28084 19346
rect 28028 19282 28084 19294
rect 28476 20018 28532 20030
rect 28476 19966 28478 20018
rect 28530 19966 28532 20018
rect 28476 19796 28532 19966
rect 29036 20020 29092 21644
rect 29148 20802 29204 21756
rect 29596 21364 29652 22204
rect 29708 22194 29764 22204
rect 29708 22036 29764 22046
rect 29708 21698 29764 21980
rect 29708 21646 29710 21698
rect 29762 21646 29764 21698
rect 29708 21634 29764 21646
rect 29820 21586 29876 22428
rect 29820 21534 29822 21586
rect 29874 21534 29876 21586
rect 29820 21522 29876 21534
rect 29932 22370 29988 24894
rect 30044 25564 30156 25620
rect 30044 22708 30100 25564
rect 30156 25526 30212 25564
rect 30268 25508 30324 27022
rect 30380 26404 30436 26414
rect 30492 26404 30548 29148
rect 30604 29138 30660 29148
rect 30604 27858 30660 27870
rect 30604 27806 30606 27858
rect 30658 27806 30660 27858
rect 30604 26628 30660 27806
rect 30716 27074 30772 30382
rect 30828 30324 30884 30940
rect 31164 30930 31220 30940
rect 31500 30772 31556 30782
rect 31388 30770 31556 30772
rect 31388 30718 31502 30770
rect 31554 30718 31556 30770
rect 31388 30716 31556 30718
rect 31388 30434 31444 30716
rect 31500 30706 31556 30716
rect 31388 30382 31390 30434
rect 31442 30382 31444 30434
rect 31388 30370 31444 30382
rect 30940 30324 30996 30334
rect 30828 30322 30996 30324
rect 30828 30270 30942 30322
rect 30994 30270 30996 30322
rect 30828 30268 30996 30270
rect 30828 28196 30884 30268
rect 30940 30258 30996 30268
rect 31500 30212 31556 30222
rect 31500 30118 31556 30156
rect 31612 29988 31668 31276
rect 31724 30884 31780 33070
rect 31836 33124 31892 33134
rect 31836 32786 31892 33068
rect 31836 32734 31838 32786
rect 31890 32734 31892 32786
rect 31836 32722 31892 32734
rect 31724 30818 31780 30828
rect 31836 30212 31892 30222
rect 31836 30118 31892 30156
rect 31612 29932 31892 29988
rect 31612 29764 31668 29774
rect 30940 29428 30996 29438
rect 30940 29334 30996 29372
rect 31612 29314 31668 29708
rect 31612 29262 31614 29314
rect 31666 29262 31668 29314
rect 31612 28644 31668 29262
rect 31612 28578 31668 28588
rect 31388 28532 31444 28542
rect 30828 28140 30996 28196
rect 30828 27970 30884 27982
rect 30828 27918 30830 27970
rect 30882 27918 30884 27970
rect 30828 27636 30884 27918
rect 30940 27748 30996 28140
rect 31388 27970 31444 28476
rect 31388 27918 31390 27970
rect 31442 27918 31444 27970
rect 31388 27906 31444 27918
rect 31724 28420 31780 28430
rect 31724 27970 31780 28364
rect 31724 27918 31726 27970
rect 31778 27918 31780 27970
rect 31724 27906 31780 27918
rect 30940 27692 31108 27748
rect 30828 27570 30884 27580
rect 30716 27022 30718 27074
rect 30770 27022 30772 27074
rect 30716 27010 30772 27022
rect 30940 26852 30996 26862
rect 30604 26572 30772 26628
rect 30380 26402 30548 26404
rect 30380 26350 30382 26402
rect 30434 26350 30548 26402
rect 30380 26348 30548 26350
rect 30604 26402 30660 26414
rect 30604 26350 30606 26402
rect 30658 26350 30660 26402
rect 30380 26338 30436 26348
rect 30268 25442 30324 25452
rect 30604 26180 30660 26350
rect 30716 26292 30772 26572
rect 30716 26226 30772 26236
rect 30940 26290 30996 26796
rect 30940 26238 30942 26290
rect 30994 26238 30996 26290
rect 30940 26226 30996 26238
rect 30604 26068 30660 26124
rect 31052 26068 31108 27692
rect 31276 26068 31332 26078
rect 30604 26012 31108 26068
rect 31164 26066 31332 26068
rect 31164 26014 31278 26066
rect 31330 26014 31332 26066
rect 31164 26012 31332 26014
rect 30268 24722 30324 24734
rect 30268 24670 30270 24722
rect 30322 24670 30324 24722
rect 30268 24612 30324 24670
rect 30044 22642 30100 22652
rect 30156 23938 30212 23950
rect 30156 23886 30158 23938
rect 30210 23886 30212 23938
rect 29932 22318 29934 22370
rect 29986 22318 29988 22370
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 29148 20738 29204 20750
rect 29260 21308 29652 21364
rect 29708 21476 29764 21486
rect 29260 20690 29316 21308
rect 29484 20804 29540 20814
rect 29484 20710 29540 20748
rect 29260 20638 29262 20690
rect 29314 20638 29316 20690
rect 29260 20626 29316 20638
rect 29596 20692 29652 20702
rect 29148 20020 29204 20030
rect 29036 20018 29204 20020
rect 29036 19966 29150 20018
rect 29202 19966 29204 20018
rect 29036 19964 29204 19966
rect 27692 19182 27694 19234
rect 27746 19182 27748 19234
rect 27692 19170 27748 19182
rect 27804 19234 27972 19236
rect 27804 19182 27918 19234
rect 27970 19182 27972 19234
rect 27804 19180 27972 19182
rect 27804 19012 27860 19180
rect 27916 19170 27972 19180
rect 28364 19236 28420 19246
rect 28364 19142 28420 19180
rect 28476 19124 28532 19740
rect 29148 19236 29204 19964
rect 29148 19142 29204 19180
rect 28532 19068 28644 19124
rect 28476 19058 28532 19068
rect 27132 18610 27188 18620
rect 27356 18956 27860 19012
rect 28140 19010 28196 19022
rect 28140 18958 28142 19010
rect 28194 18958 28196 19010
rect 27356 18674 27412 18956
rect 27356 18622 27358 18674
rect 27410 18622 27412 18674
rect 27356 18610 27412 18622
rect 27916 18676 27972 18686
rect 27916 18582 27972 18620
rect 28140 18676 28196 18958
rect 28140 18610 28196 18620
rect 28588 18450 28644 19068
rect 29596 19012 29652 20636
rect 29708 20580 29764 21420
rect 29708 20018 29764 20524
rect 29708 19966 29710 20018
rect 29762 19966 29764 20018
rect 29708 19954 29764 19966
rect 29820 19908 29876 19918
rect 29820 19814 29876 19852
rect 29932 19796 29988 22318
rect 30156 22372 30212 23886
rect 30268 23938 30324 24556
rect 30492 24724 30548 24734
rect 30492 24162 30548 24668
rect 30604 24500 30660 26012
rect 30716 25508 30772 25518
rect 30716 24612 30772 25452
rect 31164 25506 31220 26012
rect 31276 26002 31332 26012
rect 31164 25454 31166 25506
rect 31218 25454 31220 25506
rect 31164 25442 31220 25454
rect 31388 25284 31444 25294
rect 30940 24612 30996 24622
rect 30716 24610 30996 24612
rect 30716 24558 30942 24610
rect 30994 24558 30996 24610
rect 30716 24556 30996 24558
rect 30604 24444 30884 24500
rect 30492 24110 30494 24162
rect 30546 24110 30548 24162
rect 30492 24098 30548 24110
rect 30604 24164 30660 24174
rect 30604 24070 30660 24108
rect 30268 23886 30270 23938
rect 30322 23886 30324 23938
rect 30268 23716 30324 23886
rect 30268 23650 30324 23660
rect 30604 23380 30660 23390
rect 30604 23154 30660 23324
rect 30604 23102 30606 23154
rect 30658 23102 30660 23154
rect 30604 23090 30660 23102
rect 30492 22708 30548 22718
rect 30156 22316 30324 22372
rect 30044 22260 30100 22270
rect 30044 22166 30100 22204
rect 30156 22148 30212 22158
rect 30156 22054 30212 22092
rect 29932 19730 29988 19740
rect 30044 21924 30100 21934
rect 30268 21924 30324 22316
rect 30492 22148 30548 22652
rect 30828 22484 30884 24444
rect 30940 23156 30996 24556
rect 31388 24610 31444 25228
rect 31388 24558 31390 24610
rect 31442 24558 31444 24610
rect 31052 24052 31108 24062
rect 31052 23958 31108 23996
rect 31388 23492 31444 24558
rect 31836 24610 31892 29932
rect 32060 28420 32116 35420
rect 32172 35410 32228 35420
rect 32284 34132 32340 35756
rect 32508 35364 32564 35374
rect 32508 35138 32564 35308
rect 32508 35086 32510 35138
rect 32562 35086 32564 35138
rect 32508 35074 32564 35086
rect 32396 34804 32452 34814
rect 32396 34710 32452 34748
rect 32620 34580 32676 36318
rect 32732 34804 32788 41022
rect 32844 40628 32900 42478
rect 33180 42196 33236 42702
rect 33740 42756 33796 43374
rect 33852 43092 33908 44044
rect 35308 44100 35364 44270
rect 35308 44034 35364 44044
rect 34008 43932 35208 43942
rect 34064 43930 34112 43932
rect 34168 43930 34216 43932
rect 34076 43878 34112 43930
rect 34200 43878 34216 43930
rect 34064 43876 34112 43878
rect 34168 43876 34216 43878
rect 34272 43930 34320 43932
rect 34376 43930 34424 43932
rect 34480 43930 34528 43932
rect 34376 43878 34396 43930
rect 34480 43878 34520 43930
rect 34272 43876 34320 43878
rect 34376 43876 34424 43878
rect 34480 43876 34528 43878
rect 34584 43876 34632 43932
rect 34688 43930 34736 43932
rect 34792 43930 34840 43932
rect 34896 43930 34944 43932
rect 34696 43878 34736 43930
rect 34820 43878 34840 43930
rect 34688 43876 34736 43878
rect 34792 43876 34840 43878
rect 34896 43876 34944 43878
rect 35000 43930 35048 43932
rect 35104 43930 35152 43932
rect 35000 43878 35016 43930
rect 35104 43878 35140 43930
rect 35000 43876 35048 43878
rect 35104 43876 35152 43878
rect 35532 43876 35588 45388
rect 35980 45220 36036 45614
rect 34008 43866 35208 43876
rect 35308 43820 35588 43876
rect 35868 45164 35980 45220
rect 35868 44324 35924 45164
rect 35980 45154 36036 45164
rect 36316 45106 36372 46284
rect 36876 45220 36932 46844
rect 37100 46676 37156 47182
rect 37100 46582 37156 46620
rect 37212 46004 37268 47404
rect 37548 47394 37604 47404
rect 37996 47236 38052 47246
rect 37884 47234 38052 47236
rect 37884 47182 37998 47234
rect 38050 47182 38052 47234
rect 37884 47180 38052 47182
rect 37884 46676 37940 47180
rect 37996 47170 38052 47180
rect 37884 46610 37940 46620
rect 37548 46562 37604 46574
rect 37548 46510 37550 46562
rect 37602 46510 37604 46562
rect 37548 46452 37604 46510
rect 37548 46386 37604 46396
rect 37996 46562 38052 46574
rect 37996 46510 37998 46562
rect 38050 46510 38052 46562
rect 37996 46340 38052 46510
rect 37996 46274 38052 46284
rect 37548 46004 37604 46014
rect 37996 46004 38052 46014
rect 37212 46002 38052 46004
rect 37212 45950 37550 46002
rect 37602 45950 37998 46002
rect 38050 45950 38052 46002
rect 37212 45948 38052 45950
rect 37100 45892 37156 45902
rect 37212 45892 37268 45948
rect 37548 45938 37604 45948
rect 37996 45938 38052 45948
rect 37156 45836 37268 45892
rect 37100 45798 37156 45836
rect 36988 45780 37044 45790
rect 36988 45686 37044 45724
rect 36988 45220 37044 45230
rect 36316 45054 36318 45106
rect 36370 45054 36372 45106
rect 36316 45042 36372 45054
rect 36764 45218 37492 45220
rect 36764 45166 36990 45218
rect 37042 45166 37492 45218
rect 36764 45164 37492 45166
rect 35980 44884 36036 44894
rect 35980 44546 36036 44828
rect 35980 44494 35982 44546
rect 36034 44494 36036 44546
rect 35980 44482 36036 44494
rect 35196 43764 35252 43774
rect 35308 43764 35364 43820
rect 35196 43762 35364 43764
rect 35196 43710 35198 43762
rect 35250 43710 35364 43762
rect 35196 43708 35364 43710
rect 35196 43698 35252 43708
rect 35868 43650 35924 44268
rect 35868 43598 35870 43650
rect 35922 43598 35924 43650
rect 35868 43586 35924 43598
rect 36316 44098 36372 44110
rect 36316 44046 36318 44098
rect 36370 44046 36372 44098
rect 34636 43428 34692 43438
rect 34636 43334 34692 43372
rect 33852 43026 33908 43036
rect 34300 42868 34356 42878
rect 33964 42756 34020 42766
rect 33740 42690 33796 42700
rect 33852 42700 33964 42756
rect 33628 42644 33684 42654
rect 33180 42130 33236 42140
rect 33516 42532 33572 42542
rect 33516 42082 33572 42476
rect 33516 42030 33518 42082
rect 33570 42030 33572 42082
rect 33516 42018 33572 42030
rect 33292 41970 33348 41982
rect 33292 41918 33294 41970
rect 33346 41918 33348 41970
rect 33180 41746 33236 41758
rect 33180 41694 33182 41746
rect 33234 41694 33236 41746
rect 33180 41636 33236 41694
rect 33180 41570 33236 41580
rect 33292 41412 33348 41918
rect 32844 40562 32900 40572
rect 33180 40964 33236 40974
rect 33068 40404 33124 40414
rect 33068 40310 33124 40348
rect 33180 38274 33236 40908
rect 33292 40740 33348 41356
rect 33628 41074 33684 42588
rect 33852 42196 33908 42700
rect 33964 42690 34020 42700
rect 34300 42754 34356 42812
rect 34972 42868 35028 42878
rect 34300 42702 34302 42754
rect 34354 42702 34356 42754
rect 34300 42690 34356 42702
rect 34412 42756 34468 42766
rect 34412 42662 34468 42700
rect 34972 42754 35028 42812
rect 34972 42702 34974 42754
rect 35026 42702 35028 42754
rect 34972 42690 35028 42702
rect 35196 42866 35252 42878
rect 35196 42814 35198 42866
rect 35250 42814 35252 42866
rect 35084 42644 35140 42654
rect 35084 42550 35140 42588
rect 35196 42532 35252 42814
rect 36204 42756 36260 42766
rect 36316 42756 36372 44046
rect 36540 43762 36596 43774
rect 36540 43710 36542 43762
rect 36594 43710 36596 43762
rect 36428 43652 36484 43662
rect 36428 43558 36484 43596
rect 36204 42754 36316 42756
rect 36204 42702 36206 42754
rect 36258 42702 36316 42754
rect 36204 42700 36316 42702
rect 36204 42690 36260 42700
rect 36316 42662 36372 42700
rect 36428 42644 36484 42654
rect 36428 42550 36484 42588
rect 36092 42532 36148 42542
rect 35196 42476 35364 42532
rect 34008 42364 35208 42374
rect 34064 42362 34112 42364
rect 34168 42362 34216 42364
rect 34076 42310 34112 42362
rect 34200 42310 34216 42362
rect 34064 42308 34112 42310
rect 34168 42308 34216 42310
rect 34272 42362 34320 42364
rect 34376 42362 34424 42364
rect 34480 42362 34528 42364
rect 34376 42310 34396 42362
rect 34480 42310 34520 42362
rect 34272 42308 34320 42310
rect 34376 42308 34424 42310
rect 34480 42308 34528 42310
rect 34584 42308 34632 42364
rect 34688 42362 34736 42364
rect 34792 42362 34840 42364
rect 34896 42362 34944 42364
rect 34696 42310 34736 42362
rect 34820 42310 34840 42362
rect 34688 42308 34736 42310
rect 34792 42308 34840 42310
rect 34896 42308 34944 42310
rect 35000 42362 35048 42364
rect 35104 42362 35152 42364
rect 35000 42310 35016 42362
rect 35104 42310 35140 42362
rect 35000 42308 35048 42310
rect 35104 42308 35152 42310
rect 34008 42298 35208 42308
rect 33852 42140 34020 42196
rect 33852 41970 33908 41982
rect 33852 41918 33854 41970
rect 33906 41918 33908 41970
rect 33852 41636 33908 41918
rect 33964 41972 34020 42140
rect 35196 42084 35252 42094
rect 33964 41906 34020 41916
rect 34748 41970 34804 41982
rect 34748 41918 34750 41970
rect 34802 41918 34804 41970
rect 33852 41570 33908 41580
rect 33628 41022 33630 41074
rect 33682 41022 33684 41074
rect 33628 41010 33684 41022
rect 34748 41076 34804 41918
rect 35084 41972 35140 41982
rect 35084 41878 35140 41916
rect 34748 41010 34804 41020
rect 35196 40964 35252 42028
rect 35308 41972 35364 42476
rect 35532 42196 35588 42206
rect 35308 41906 35364 41916
rect 35420 42082 35476 42094
rect 35420 42030 35422 42082
rect 35474 42030 35476 42082
rect 35420 41300 35476 42030
rect 35532 41858 35588 42140
rect 35532 41806 35534 41858
rect 35586 41806 35588 41858
rect 35532 41794 35588 41806
rect 35756 41860 35812 41870
rect 35420 41244 35588 41300
rect 35308 41188 35364 41198
rect 35308 41094 35364 41132
rect 35196 40908 35364 40964
rect 34008 40796 35208 40806
rect 34064 40794 34112 40796
rect 34168 40794 34216 40796
rect 34076 40742 34112 40794
rect 34200 40742 34216 40794
rect 34064 40740 34112 40742
rect 34168 40740 34216 40742
rect 34272 40794 34320 40796
rect 34376 40794 34424 40796
rect 34480 40794 34528 40796
rect 34376 40742 34396 40794
rect 34480 40742 34520 40794
rect 34272 40740 34320 40742
rect 34376 40740 34424 40742
rect 34480 40740 34528 40742
rect 34584 40740 34632 40796
rect 34688 40794 34736 40796
rect 34792 40794 34840 40796
rect 34896 40794 34944 40796
rect 34696 40742 34736 40794
rect 34820 40742 34840 40794
rect 34688 40740 34736 40742
rect 34792 40740 34840 40742
rect 34896 40740 34944 40742
rect 35000 40794 35048 40796
rect 35104 40794 35152 40796
rect 35000 40742 35016 40794
rect 35104 40742 35140 40794
rect 35000 40740 35048 40742
rect 35104 40740 35152 40742
rect 33292 40684 33572 40740
rect 34008 40730 35208 40740
rect 33292 40516 33348 40526
rect 33292 40292 33348 40460
rect 33292 39058 33348 40236
rect 33292 39006 33294 39058
rect 33346 39006 33348 39058
rect 33292 38994 33348 39006
rect 33404 40180 33460 40190
rect 33180 38222 33182 38274
rect 33234 38222 33236 38274
rect 33180 38210 33236 38222
rect 32844 37938 32900 37950
rect 32844 37886 32846 37938
rect 32898 37886 32900 37938
rect 32844 35476 32900 37886
rect 33068 37826 33124 37838
rect 33068 37774 33070 37826
rect 33122 37774 33124 37826
rect 33068 36932 33124 37774
rect 33404 37604 33460 40124
rect 33516 40068 33572 40684
rect 33628 40628 33684 40638
rect 33628 40534 33684 40572
rect 33964 40628 34020 40638
rect 35308 40628 35364 40908
rect 33516 40012 33684 40068
rect 33516 39844 33572 39854
rect 33516 38834 33572 39788
rect 33516 38782 33518 38834
rect 33570 38782 33572 38834
rect 33516 38724 33572 38782
rect 33516 38658 33572 38668
rect 33628 38274 33684 40012
rect 33964 39844 34020 40572
rect 35084 40572 35364 40628
rect 34076 40516 34132 40526
rect 34076 40422 34132 40460
rect 33964 39778 34020 39788
rect 34188 40402 34244 40414
rect 34188 40350 34190 40402
rect 34242 40350 34244 40402
rect 34188 39620 34244 40350
rect 35084 40402 35140 40572
rect 35084 40350 35086 40402
rect 35138 40350 35140 40402
rect 35084 40338 35140 40350
rect 34636 39732 34692 39742
rect 34636 39638 34692 39676
rect 34524 39620 34580 39630
rect 34188 39618 34580 39620
rect 34188 39566 34526 39618
rect 34578 39566 34580 39618
rect 34188 39564 34580 39566
rect 34524 39554 34580 39564
rect 34008 39228 35208 39238
rect 34064 39226 34112 39228
rect 34168 39226 34216 39228
rect 34076 39174 34112 39226
rect 34200 39174 34216 39226
rect 34064 39172 34112 39174
rect 34168 39172 34216 39174
rect 34272 39226 34320 39228
rect 34376 39226 34424 39228
rect 34480 39226 34528 39228
rect 34376 39174 34396 39226
rect 34480 39174 34520 39226
rect 34272 39172 34320 39174
rect 34376 39172 34424 39174
rect 34480 39172 34528 39174
rect 34584 39172 34632 39228
rect 34688 39226 34736 39228
rect 34792 39226 34840 39228
rect 34896 39226 34944 39228
rect 34696 39174 34736 39226
rect 34820 39174 34840 39226
rect 34688 39172 34736 39174
rect 34792 39172 34840 39174
rect 34896 39172 34944 39174
rect 35000 39226 35048 39228
rect 35104 39226 35152 39228
rect 35000 39174 35016 39226
rect 35104 39174 35140 39226
rect 35000 39172 35048 39174
rect 35104 39172 35152 39174
rect 34008 39162 35208 39172
rect 33740 39060 33796 39070
rect 33740 38966 33796 39004
rect 34300 39060 34356 39070
rect 34300 38966 34356 39004
rect 34188 38948 34244 38958
rect 34188 38854 34244 38892
rect 34972 38948 35028 38958
rect 33964 38834 34020 38846
rect 33964 38782 33966 38834
rect 34018 38782 34020 38834
rect 33964 38668 34020 38782
rect 34748 38836 34804 38846
rect 34748 38742 34804 38780
rect 33964 38612 34132 38668
rect 33628 38222 33630 38274
rect 33682 38222 33684 38274
rect 33404 37548 33572 37604
rect 33068 36866 33124 36876
rect 33516 37380 33572 37548
rect 33516 36820 33572 37324
rect 33628 37156 33684 38222
rect 33740 38164 33796 38174
rect 33740 38070 33796 38108
rect 34076 38164 34132 38612
rect 34076 38098 34132 38108
rect 33852 38050 33908 38062
rect 33852 37998 33854 38050
rect 33906 37998 33908 38050
rect 33852 37940 33908 37998
rect 34972 38052 35028 38892
rect 35084 38948 35140 38958
rect 35084 38946 35364 38948
rect 35084 38894 35086 38946
rect 35138 38894 35364 38946
rect 35084 38892 35364 38894
rect 35084 38882 35140 38892
rect 35196 38724 35252 38734
rect 35196 38276 35252 38668
rect 35308 38668 35364 38892
rect 35532 38668 35588 41244
rect 35756 41186 35812 41804
rect 35756 41134 35758 41186
rect 35810 41134 35812 41186
rect 35756 41122 35812 41134
rect 36092 41186 36148 42476
rect 36092 41134 36094 41186
rect 36146 41134 36148 41186
rect 36092 41122 36148 41134
rect 36316 41076 36372 41086
rect 36316 41074 36484 41076
rect 36316 41022 36318 41074
rect 36370 41022 36484 41074
rect 36316 41020 36484 41022
rect 36316 41010 36372 41020
rect 35868 40964 35924 40974
rect 35868 40870 35924 40908
rect 35980 40962 36036 40974
rect 35980 40910 35982 40962
rect 36034 40910 36036 40962
rect 35980 40516 36036 40910
rect 35868 40460 36036 40516
rect 35644 40404 35700 40414
rect 35644 39506 35700 40348
rect 35644 39454 35646 39506
rect 35698 39454 35700 39506
rect 35644 39442 35700 39454
rect 35868 38724 35924 40460
rect 36316 40404 36372 40414
rect 35308 38612 35476 38668
rect 35532 38612 35812 38668
rect 35868 38658 35924 38668
rect 35980 40402 36372 40404
rect 35980 40350 36318 40402
rect 36370 40350 36372 40402
rect 35980 40348 36372 40350
rect 35980 38722 36036 40348
rect 36316 40338 36372 40348
rect 35980 38670 35982 38722
rect 36034 38670 36036 38722
rect 35980 38658 36036 38670
rect 36316 39844 36372 39854
rect 35196 38220 35364 38276
rect 35308 38162 35364 38220
rect 35308 38110 35310 38162
rect 35362 38110 35364 38162
rect 35308 38098 35364 38110
rect 35196 38052 35252 38062
rect 34972 38050 35252 38052
rect 34972 37998 35198 38050
rect 35250 37998 35252 38050
rect 34972 37996 35252 37998
rect 33628 37090 33684 37100
rect 33740 37884 33908 37940
rect 33740 36932 33796 37884
rect 35196 37828 35252 37996
rect 35196 37772 35364 37828
rect 33740 36866 33796 36876
rect 33852 37716 33908 37726
rect 33516 36764 33684 36820
rect 33628 36708 33684 36764
rect 33628 36652 33796 36708
rect 33292 36596 33348 36606
rect 33292 36502 33348 36540
rect 33628 36482 33684 36494
rect 33628 36430 33630 36482
rect 33682 36430 33684 36482
rect 33068 36148 33124 36158
rect 33068 35812 33124 36092
rect 33628 35924 33684 36430
rect 33740 36482 33796 36652
rect 33740 36430 33742 36482
rect 33794 36430 33796 36482
rect 33740 36418 33796 36430
rect 33740 35924 33796 35934
rect 33628 35868 33740 35924
rect 33740 35858 33796 35868
rect 33068 35718 33124 35756
rect 32844 35410 32900 35420
rect 33628 35700 33684 35710
rect 33292 35026 33348 35038
rect 33516 35028 33572 35038
rect 33292 34974 33294 35026
rect 33346 34974 33348 35026
rect 33180 34916 33236 34926
rect 32956 34914 33236 34916
rect 32956 34862 33182 34914
rect 33234 34862 33236 34914
rect 32956 34860 33236 34862
rect 32844 34804 32900 34814
rect 32732 34802 32900 34804
rect 32732 34750 32846 34802
rect 32898 34750 32900 34802
rect 32732 34748 32900 34750
rect 32844 34738 32900 34748
rect 32956 34580 33012 34860
rect 33180 34850 33236 34860
rect 32620 34524 33012 34580
rect 33068 34692 33124 34702
rect 32508 34244 32564 34254
rect 32508 34150 32564 34188
rect 33068 34242 33124 34636
rect 33292 34356 33348 34974
rect 33068 34190 33070 34242
rect 33122 34190 33124 34242
rect 32284 34130 32452 34132
rect 32284 34078 32286 34130
rect 32338 34078 32452 34130
rect 32284 34076 32452 34078
rect 32284 34066 32340 34076
rect 32172 33124 32228 33134
rect 32284 33124 32340 33134
rect 32228 33122 32340 33124
rect 32228 33070 32286 33122
rect 32338 33070 32340 33122
rect 32228 33068 32340 33070
rect 32172 32674 32228 33068
rect 32284 33058 32340 33068
rect 32172 32622 32174 32674
rect 32226 32622 32228 32674
rect 32172 32610 32228 32622
rect 32396 32788 32452 34076
rect 32956 33572 33012 33582
rect 32844 33348 32900 33358
rect 32732 33124 32788 33134
rect 32732 33030 32788 33068
rect 32396 32340 32452 32732
rect 32396 32274 32452 32284
rect 32508 32338 32564 32350
rect 32508 32286 32510 32338
rect 32562 32286 32564 32338
rect 32396 31556 32452 31566
rect 32284 31444 32340 31454
rect 32284 30994 32340 31388
rect 32284 30942 32286 30994
rect 32338 30942 32340 30994
rect 32284 30930 32340 30942
rect 32396 30996 32452 31500
rect 32508 31108 32564 32286
rect 32732 32004 32788 32014
rect 32844 32004 32900 33292
rect 32956 32564 33012 33516
rect 33068 33348 33124 34190
rect 33180 34300 33348 34356
rect 33404 34972 33516 35028
rect 33180 33572 33236 34300
rect 33292 34130 33348 34142
rect 33292 34078 33294 34130
rect 33346 34078 33348 34130
rect 33292 33684 33348 34078
rect 33404 34018 33460 34972
rect 33516 34962 33572 34972
rect 33404 33966 33406 34018
rect 33458 33966 33460 34018
rect 33404 33954 33460 33966
rect 33516 34242 33572 34254
rect 33516 34190 33518 34242
rect 33570 34190 33572 34242
rect 33516 33796 33572 34190
rect 33516 33730 33572 33740
rect 33292 33618 33348 33628
rect 33628 33572 33684 35644
rect 33740 35588 33796 35598
rect 33740 35494 33796 35532
rect 33852 35140 33908 37660
rect 34008 37660 35208 37670
rect 34064 37658 34112 37660
rect 34168 37658 34216 37660
rect 34076 37606 34112 37658
rect 34200 37606 34216 37658
rect 34064 37604 34112 37606
rect 34168 37604 34216 37606
rect 34272 37658 34320 37660
rect 34376 37658 34424 37660
rect 34480 37658 34528 37660
rect 34376 37606 34396 37658
rect 34480 37606 34520 37658
rect 34272 37604 34320 37606
rect 34376 37604 34424 37606
rect 34480 37604 34528 37606
rect 34584 37604 34632 37660
rect 34688 37658 34736 37660
rect 34792 37658 34840 37660
rect 34896 37658 34944 37660
rect 34696 37606 34736 37658
rect 34820 37606 34840 37658
rect 34688 37604 34736 37606
rect 34792 37604 34840 37606
rect 34896 37604 34944 37606
rect 35000 37658 35048 37660
rect 35104 37658 35152 37660
rect 35000 37606 35016 37658
rect 35104 37606 35140 37658
rect 35000 37604 35048 37606
rect 35104 37604 35152 37606
rect 34008 37594 35208 37604
rect 34524 37492 34580 37502
rect 34188 37378 34244 37390
rect 34188 37326 34190 37378
rect 34242 37326 34244 37378
rect 34188 36932 34244 37326
rect 34188 36260 34244 36876
rect 34524 36482 34580 37436
rect 35308 37490 35364 37772
rect 35308 37438 35310 37490
rect 35362 37438 35364 37490
rect 35308 37426 35364 37438
rect 34524 36430 34526 36482
rect 34578 36430 34580 36482
rect 34524 36418 34580 36430
rect 35196 37268 35252 37278
rect 35196 36260 35252 37212
rect 35420 36706 35476 38612
rect 35644 38276 35700 38286
rect 35644 37266 35700 38220
rect 35756 38274 35812 38612
rect 35756 38222 35758 38274
rect 35810 38222 35812 38274
rect 35756 38210 35812 38222
rect 36092 38164 36148 38174
rect 36092 38070 36148 38108
rect 36204 38052 36260 38062
rect 36316 38052 36372 39788
rect 36428 39172 36484 41020
rect 36428 39106 36484 39116
rect 36540 38668 36596 43710
rect 36764 43538 36820 45164
rect 36988 45154 37044 45164
rect 37436 44322 37492 45164
rect 37660 44884 37716 44894
rect 37660 44882 37828 44884
rect 37660 44830 37662 44882
rect 37714 44830 37828 44882
rect 37660 44828 37828 44830
rect 37660 44818 37716 44828
rect 37436 44270 37438 44322
rect 37490 44270 37492 44322
rect 37436 44258 37492 44270
rect 37548 44324 37604 44334
rect 37548 44230 37604 44268
rect 37660 44210 37716 44222
rect 37660 44158 37662 44210
rect 37714 44158 37716 44210
rect 36988 44100 37044 44110
rect 36988 44098 37268 44100
rect 36988 44046 36990 44098
rect 37042 44046 37268 44098
rect 36988 44044 37268 44046
rect 36988 44034 37044 44044
rect 36764 43486 36766 43538
rect 36818 43486 36820 43538
rect 36764 43474 36820 43486
rect 36988 42756 37044 42766
rect 36988 42662 37044 42700
rect 37100 42644 37156 42654
rect 37100 42530 37156 42588
rect 37100 42478 37102 42530
rect 37154 42478 37156 42530
rect 36988 41972 37044 41982
rect 36988 39732 37044 41916
rect 37100 41748 37156 42478
rect 37212 41972 37268 44044
rect 37660 43652 37716 44158
rect 37660 43586 37716 43596
rect 37660 43426 37716 43438
rect 37660 43374 37662 43426
rect 37714 43374 37716 43426
rect 37548 43314 37604 43326
rect 37548 43262 37550 43314
rect 37602 43262 37604 43314
rect 37212 41906 37268 41916
rect 37324 42530 37380 42542
rect 37324 42478 37326 42530
rect 37378 42478 37380 42530
rect 37324 41970 37380 42478
rect 37548 42084 37604 43262
rect 37660 42756 37716 43374
rect 37660 42690 37716 42700
rect 37660 42532 37716 42542
rect 37660 42438 37716 42476
rect 37548 42018 37604 42028
rect 37772 42420 37828 44828
rect 37884 43652 37940 43662
rect 37884 42532 37940 43596
rect 37884 42438 37940 42476
rect 37996 42642 38052 42654
rect 37996 42590 37998 42642
rect 38050 42590 38052 42642
rect 37772 41972 37828 42364
rect 37324 41918 37326 41970
rect 37378 41918 37380 41970
rect 37324 41906 37380 41918
rect 37660 41970 37828 41972
rect 37660 41918 37774 41970
rect 37826 41918 37828 41970
rect 37660 41916 37828 41918
rect 37660 41860 37716 41916
rect 37772 41906 37828 41916
rect 37436 41804 37716 41860
rect 37884 41860 37940 41870
rect 37100 41692 37380 41748
rect 37100 41412 37156 41422
rect 37100 41186 37156 41356
rect 37100 41134 37102 41186
rect 37154 41134 37156 41186
rect 37100 41122 37156 41134
rect 37212 41076 37268 41086
rect 37212 40982 37268 41020
rect 37324 40962 37380 41692
rect 37324 40910 37326 40962
rect 37378 40910 37380 40962
rect 37324 40898 37380 40910
rect 37100 39732 37156 39742
rect 36988 39730 37156 39732
rect 36988 39678 37102 39730
rect 37154 39678 37156 39730
rect 36988 39676 37156 39678
rect 37100 39666 37156 39676
rect 37212 39618 37268 39630
rect 37212 39566 37214 39618
rect 37266 39566 37268 39618
rect 36204 38050 36372 38052
rect 36204 37998 36206 38050
rect 36258 37998 36372 38050
rect 36204 37996 36372 37998
rect 36428 38612 36596 38668
rect 36988 39506 37044 39518
rect 36988 39454 36990 39506
rect 37042 39454 37044 39506
rect 36204 37986 36260 37996
rect 36428 37604 36484 38612
rect 35644 37214 35646 37266
rect 35698 37214 35700 37266
rect 35644 37202 35700 37214
rect 35980 37548 36484 37604
rect 35420 36654 35422 36706
rect 35474 36654 35476 36706
rect 35420 36642 35476 36654
rect 35644 36594 35700 36606
rect 35644 36542 35646 36594
rect 35698 36542 35700 36594
rect 35420 36482 35476 36494
rect 35420 36430 35422 36482
rect 35474 36430 35476 36482
rect 35196 36204 35364 36260
rect 34188 36194 34244 36204
rect 34008 36092 35208 36102
rect 34064 36090 34112 36092
rect 34168 36090 34216 36092
rect 34076 36038 34112 36090
rect 34200 36038 34216 36090
rect 34064 36036 34112 36038
rect 34168 36036 34216 36038
rect 34272 36090 34320 36092
rect 34376 36090 34424 36092
rect 34480 36090 34528 36092
rect 34376 36038 34396 36090
rect 34480 36038 34520 36090
rect 34272 36036 34320 36038
rect 34376 36036 34424 36038
rect 34480 36036 34528 36038
rect 34584 36036 34632 36092
rect 34688 36090 34736 36092
rect 34792 36090 34840 36092
rect 34896 36090 34944 36092
rect 34696 36038 34736 36090
rect 34820 36038 34840 36090
rect 34688 36036 34736 36038
rect 34792 36036 34840 36038
rect 34896 36036 34944 36038
rect 35000 36090 35048 36092
rect 35104 36090 35152 36092
rect 35000 36038 35016 36090
rect 35104 36038 35140 36090
rect 35000 36036 35048 36038
rect 35104 36036 35152 36038
rect 34008 36026 35208 36036
rect 34300 35924 34356 35934
rect 34300 35586 34356 35868
rect 34972 35922 35028 35934
rect 35196 35924 35252 35934
rect 34972 35870 34974 35922
rect 35026 35870 35028 35922
rect 34636 35812 34692 35822
rect 34636 35698 34692 35756
rect 34636 35646 34638 35698
rect 34690 35646 34692 35698
rect 34636 35634 34692 35646
rect 34860 35698 34916 35710
rect 34860 35646 34862 35698
rect 34914 35646 34916 35698
rect 34300 35534 34302 35586
rect 34354 35534 34356 35586
rect 34300 35476 34356 35534
rect 34860 35476 34916 35646
rect 34300 35410 34356 35420
rect 34524 35474 34916 35476
rect 34524 35422 34862 35474
rect 34914 35422 34916 35474
rect 34524 35420 34916 35422
rect 33180 33506 33236 33516
rect 33516 33516 33684 33572
rect 33740 35084 33908 35140
rect 33292 33348 33348 33358
rect 33068 33346 33348 33348
rect 33068 33294 33294 33346
rect 33346 33294 33348 33346
rect 33068 33292 33348 33294
rect 33292 33282 33348 33292
rect 33404 33124 33460 33134
rect 33180 32564 33236 32574
rect 33404 32564 33460 33068
rect 33516 32788 33572 33516
rect 33740 33460 33796 35084
rect 33852 34914 33908 34926
rect 33852 34862 33854 34914
rect 33906 34862 33908 34914
rect 33852 34356 33908 34862
rect 34524 34916 34580 35420
rect 34860 35410 34916 35420
rect 34524 34850 34580 34860
rect 34972 34804 35028 35870
rect 35084 35868 35196 35924
rect 35084 35028 35140 35868
rect 35196 35858 35252 35868
rect 35308 35700 35364 36204
rect 35196 35644 35364 35700
rect 35420 35700 35476 36430
rect 35196 35474 35252 35644
rect 35420 35634 35476 35644
rect 35196 35422 35198 35474
rect 35250 35422 35252 35474
rect 35196 35410 35252 35422
rect 35196 35028 35252 35038
rect 35084 35026 35252 35028
rect 35084 34974 35198 35026
rect 35250 34974 35252 35026
rect 35084 34972 35252 34974
rect 35196 34962 35252 34972
rect 35644 34914 35700 36542
rect 35980 35922 36036 37548
rect 36204 37380 36260 37390
rect 36204 37286 36260 37324
rect 36316 37156 36372 37166
rect 36204 37100 36316 37156
rect 35980 35870 35982 35922
rect 36034 35870 36036 35922
rect 35868 35028 35924 35038
rect 35868 34934 35924 34972
rect 35644 34862 35646 34914
rect 35698 34862 35700 34914
rect 35084 34804 35140 34814
rect 34972 34748 35084 34804
rect 35644 34804 35700 34862
rect 35980 34916 36036 35870
rect 36092 35924 36148 35934
rect 36204 35924 36260 37100
rect 36316 37090 36372 37100
rect 36988 37156 37044 39454
rect 37100 39172 37156 39182
rect 37100 38164 37156 39116
rect 37212 39060 37268 39566
rect 37436 39396 37492 41804
rect 37772 41748 37828 41758
rect 37548 41746 37828 41748
rect 37548 41694 37774 41746
rect 37826 41694 37828 41746
rect 37548 41692 37828 41694
rect 37548 39618 37604 41692
rect 37772 41682 37828 41692
rect 37660 41300 37716 41310
rect 37660 40626 37716 41244
rect 37660 40574 37662 40626
rect 37714 40574 37716 40626
rect 37660 40562 37716 40574
rect 37772 41074 37828 41086
rect 37772 41022 37774 41074
rect 37826 41022 37828 41074
rect 37772 40628 37828 41022
rect 37772 40562 37828 40572
rect 37884 40514 37940 41804
rect 37996 40964 38052 42590
rect 38220 42532 38276 42542
rect 37996 40898 38052 40908
rect 38108 41746 38164 41758
rect 38108 41694 38110 41746
rect 38162 41694 38164 41746
rect 37884 40462 37886 40514
rect 37938 40462 37940 40514
rect 37884 40450 37940 40462
rect 37548 39566 37550 39618
rect 37602 39566 37604 39618
rect 37548 39554 37604 39566
rect 37996 40402 38052 40414
rect 37996 40350 37998 40402
rect 38050 40350 38052 40402
rect 37996 39620 38052 40350
rect 38108 39844 38164 41694
rect 38220 40628 38276 42476
rect 38220 40562 38276 40572
rect 38220 39844 38276 39854
rect 38164 39842 38276 39844
rect 38164 39790 38222 39842
rect 38274 39790 38276 39842
rect 38164 39788 38276 39790
rect 38108 39750 38164 39788
rect 38220 39778 38276 39788
rect 37996 39564 38388 39620
rect 37884 39506 37940 39518
rect 37884 39454 37886 39506
rect 37938 39454 37940 39506
rect 37436 39340 37716 39396
rect 37212 38994 37268 39004
rect 37660 38834 37716 39340
rect 37660 38782 37662 38834
rect 37714 38782 37716 38834
rect 37324 38388 37380 38398
rect 37212 38164 37268 38174
rect 37100 38162 37268 38164
rect 37100 38110 37214 38162
rect 37266 38110 37268 38162
rect 37100 38108 37268 38110
rect 37212 38098 37268 38108
rect 37100 37828 37156 37838
rect 37100 37826 37268 37828
rect 37100 37774 37102 37826
rect 37154 37774 37268 37826
rect 37100 37772 37268 37774
rect 37100 37762 37156 37772
rect 36988 37090 37044 37100
rect 36540 36482 36596 36494
rect 36540 36430 36542 36482
rect 36594 36430 36596 36482
rect 36092 35922 36260 35924
rect 36092 35870 36094 35922
rect 36146 35870 36260 35922
rect 36092 35868 36260 35870
rect 36428 36260 36484 36270
rect 36092 35858 36148 35868
rect 36204 35698 36260 35710
rect 36204 35646 36206 35698
rect 36258 35646 36260 35698
rect 36204 35588 36260 35646
rect 36204 35522 36260 35532
rect 36316 35700 36372 35710
rect 36204 35028 36260 35038
rect 36316 35028 36372 35644
rect 36428 35698 36484 36204
rect 36428 35646 36430 35698
rect 36482 35646 36484 35698
rect 36428 35634 36484 35646
rect 36540 35588 36596 36430
rect 36988 36370 37044 36382
rect 36988 36318 36990 36370
rect 37042 36318 37044 36370
rect 36988 36148 37044 36318
rect 36988 36082 37044 36092
rect 37100 36258 37156 36270
rect 37100 36206 37102 36258
rect 37154 36206 37156 36258
rect 37100 35924 37156 36206
rect 36652 35868 37156 35924
rect 37212 35924 37268 37772
rect 37324 37826 37380 38332
rect 37660 38164 37716 38782
rect 37884 38388 37940 39454
rect 38108 39394 38164 39406
rect 38108 39342 38110 39394
rect 38162 39342 38164 39394
rect 38108 38948 38164 39342
rect 38108 38882 38164 38892
rect 38220 38834 38276 38846
rect 38220 38782 38222 38834
rect 38274 38782 38276 38834
rect 38220 38668 38276 38782
rect 37884 38322 37940 38332
rect 38108 38612 38276 38668
rect 37324 37774 37326 37826
rect 37378 37774 37380 37826
rect 37324 37492 37380 37774
rect 37324 37426 37380 37436
rect 37436 38050 37492 38062
rect 37436 37998 37438 38050
rect 37490 37998 37492 38050
rect 37436 37380 37492 37998
rect 37324 36372 37380 36382
rect 37324 36278 37380 36316
rect 37324 35924 37380 35934
rect 37212 35922 37380 35924
rect 37212 35870 37326 35922
rect 37378 35870 37380 35922
rect 37212 35868 37380 35870
rect 36652 35698 36708 35868
rect 37324 35858 37380 35868
rect 37436 35922 37492 37324
rect 37660 37266 37716 38108
rect 37996 38164 38052 38174
rect 37996 38070 38052 38108
rect 37772 38052 37828 38062
rect 37772 38050 37940 38052
rect 37772 37998 37774 38050
rect 37826 37998 37940 38050
rect 37772 37996 37940 37998
rect 37772 37986 37828 37996
rect 37660 37214 37662 37266
rect 37714 37214 37716 37266
rect 37660 37202 37716 37214
rect 37772 37490 37828 37502
rect 37772 37438 37774 37490
rect 37826 37438 37828 37490
rect 37548 36484 37604 36494
rect 37772 36484 37828 37438
rect 37548 36482 37828 36484
rect 37548 36430 37550 36482
rect 37602 36430 37828 36482
rect 37548 36428 37828 36430
rect 37884 37042 37940 37996
rect 37884 36990 37886 37042
rect 37938 36990 37940 37042
rect 37548 36418 37604 36428
rect 37436 35870 37438 35922
rect 37490 35870 37492 35922
rect 36652 35646 36654 35698
rect 36706 35646 36708 35698
rect 36652 35634 36708 35646
rect 36988 35698 37044 35710
rect 36988 35646 36990 35698
rect 37042 35646 37044 35698
rect 36540 35522 36596 35532
rect 36988 35364 37044 35646
rect 37212 35700 37268 35710
rect 37212 35606 37268 35644
rect 36988 35298 37044 35308
rect 37324 35140 37380 35150
rect 37436 35140 37492 35870
rect 37660 35700 37716 35710
rect 37660 35698 37828 35700
rect 37660 35646 37662 35698
rect 37714 35646 37828 35698
rect 37660 35644 37828 35646
rect 37660 35634 37716 35644
rect 37772 35252 37828 35644
rect 37772 35186 37828 35196
rect 37884 35140 37940 36990
rect 37996 37380 38052 37390
rect 37996 37044 38052 37324
rect 38108 37044 38164 38612
rect 37996 37042 38164 37044
rect 37996 36990 38110 37042
rect 38162 36990 38164 37042
rect 37996 36988 38164 36990
rect 37996 36370 38052 36988
rect 38108 36978 38164 36988
rect 37996 36318 37998 36370
rect 38050 36318 38052 36370
rect 37996 36306 38052 36318
rect 38220 36370 38276 36382
rect 38220 36318 38222 36370
rect 38274 36318 38276 36370
rect 38108 36260 38164 36270
rect 38108 36166 38164 36204
rect 38108 35812 38164 35822
rect 38220 35812 38276 36318
rect 38332 35922 38388 39564
rect 38332 35870 38334 35922
rect 38386 35870 38388 35922
rect 38332 35858 38388 35870
rect 38108 35810 38276 35812
rect 38108 35758 38110 35810
rect 38162 35758 38276 35810
rect 38108 35756 38276 35758
rect 37436 35084 37716 35140
rect 37324 35046 37380 35084
rect 36204 35026 36372 35028
rect 36204 34974 36206 35026
rect 36258 34974 36372 35026
rect 36204 34972 36372 34974
rect 37660 35028 37716 35084
rect 37884 35074 37940 35084
rect 37996 35698 38052 35710
rect 37996 35646 37998 35698
rect 38050 35646 38052 35698
rect 37660 34972 37828 35028
rect 36204 34962 36260 34972
rect 36092 34916 36148 34926
rect 35980 34914 36148 34916
rect 35980 34862 36094 34914
rect 36146 34862 36148 34914
rect 35980 34860 36148 34862
rect 35644 34748 35924 34804
rect 34860 34692 34916 34730
rect 35084 34710 35140 34748
rect 34860 34626 34916 34636
rect 35308 34692 35364 34702
rect 35308 34690 35812 34692
rect 35308 34638 35310 34690
rect 35362 34638 35812 34690
rect 35308 34636 35812 34638
rect 35308 34626 35364 34636
rect 34008 34524 35208 34534
rect 34064 34522 34112 34524
rect 34168 34522 34216 34524
rect 34076 34470 34112 34522
rect 34200 34470 34216 34522
rect 34064 34468 34112 34470
rect 34168 34468 34216 34470
rect 34272 34522 34320 34524
rect 34376 34522 34424 34524
rect 34480 34522 34528 34524
rect 34376 34470 34396 34522
rect 34480 34470 34520 34522
rect 34272 34468 34320 34470
rect 34376 34468 34424 34470
rect 34480 34468 34528 34470
rect 34584 34468 34632 34524
rect 34688 34522 34736 34524
rect 34792 34522 34840 34524
rect 34896 34522 34944 34524
rect 34696 34470 34736 34522
rect 34820 34470 34840 34522
rect 34688 34468 34736 34470
rect 34792 34468 34840 34470
rect 34896 34468 34944 34470
rect 35000 34522 35048 34524
rect 35104 34522 35152 34524
rect 35000 34470 35016 34522
rect 35104 34470 35140 34522
rect 35000 34468 35048 34470
rect 35104 34468 35152 34470
rect 34008 34458 35208 34468
rect 33852 34300 34020 34356
rect 33516 32722 33572 32732
rect 33628 33404 33796 33460
rect 33852 34130 33908 34142
rect 33852 34078 33854 34130
rect 33906 34078 33908 34130
rect 33516 32564 33572 32574
rect 32956 32562 33236 32564
rect 32956 32510 33182 32562
rect 33234 32510 33236 32562
rect 32956 32508 33236 32510
rect 33180 32498 33236 32508
rect 33292 32508 33516 32564
rect 33068 32340 33124 32350
rect 32732 32002 32900 32004
rect 32732 31950 32734 32002
rect 32786 31950 32900 32002
rect 32732 31948 32900 31950
rect 32956 32338 33124 32340
rect 32956 32286 33070 32338
rect 33122 32286 33124 32338
rect 32956 32284 33124 32286
rect 32732 31938 32788 31948
rect 32620 31780 32676 31790
rect 32620 31686 32676 31724
rect 32956 31778 33012 32284
rect 33068 32274 33124 32284
rect 33292 32116 33348 32508
rect 33516 32470 33572 32508
rect 33404 32340 33460 32350
rect 33404 32246 33460 32284
rect 32956 31726 32958 31778
rect 33010 31726 33012 31778
rect 32956 31714 33012 31726
rect 33180 32060 33348 32116
rect 32508 31042 32564 31052
rect 33180 31218 33236 32060
rect 33516 31780 33572 31790
rect 33180 31166 33182 31218
rect 33234 31166 33236 31218
rect 32396 30882 32452 30940
rect 32396 30830 32398 30882
rect 32450 30830 32452 30882
rect 32396 30818 32452 30830
rect 32508 30884 32564 30894
rect 32508 30210 32564 30828
rect 32508 30158 32510 30210
rect 32562 30158 32564 30210
rect 32508 30146 32564 30158
rect 33068 29428 33124 29438
rect 32060 28354 32116 28364
rect 32956 29372 33068 29428
rect 32956 27972 33012 29372
rect 33068 29334 33124 29372
rect 32956 25732 33012 27916
rect 33068 28644 33124 28654
rect 33068 26962 33124 28588
rect 33180 28308 33236 31166
rect 33292 31444 33348 31454
rect 33292 29426 33348 31388
rect 33292 29374 33294 29426
rect 33346 29374 33348 29426
rect 33292 28532 33348 29374
rect 33516 30994 33572 31724
rect 33516 30942 33518 30994
rect 33570 30942 33572 30994
rect 33516 29428 33572 30942
rect 33628 30996 33684 33404
rect 33852 33346 33908 34078
rect 33964 33796 34020 34300
rect 35756 34354 35812 34636
rect 35756 34302 35758 34354
rect 35810 34302 35812 34354
rect 35756 34290 35812 34302
rect 35868 34580 35924 34748
rect 34076 34244 34132 34254
rect 34412 34244 34468 34254
rect 34076 34242 34244 34244
rect 34076 34190 34078 34242
rect 34130 34190 34244 34242
rect 34076 34188 34244 34190
rect 34076 34178 34132 34188
rect 34188 34020 34244 34188
rect 34468 34188 34580 34244
rect 34412 34178 34468 34188
rect 34524 34130 34580 34188
rect 34524 34078 34526 34130
rect 34578 34078 34580 34130
rect 34524 34066 34580 34078
rect 35196 34130 35252 34142
rect 35196 34078 35198 34130
rect 35250 34078 35252 34130
rect 33964 33740 34132 33796
rect 34076 33684 34132 33740
rect 34076 33618 34132 33628
rect 33964 33572 34020 33582
rect 33964 33458 34020 33516
rect 33964 33406 33966 33458
rect 34018 33406 34020 33458
rect 33964 33394 34020 33406
rect 33852 33294 33854 33346
rect 33906 33294 33908 33346
rect 33740 33236 33796 33274
rect 33740 33170 33796 33180
rect 33740 33012 33796 33022
rect 33740 31554 33796 32956
rect 33740 31502 33742 31554
rect 33794 31502 33796 31554
rect 33740 31490 33796 31502
rect 33628 30940 33796 30996
rect 33516 29362 33572 29372
rect 33740 29316 33796 30940
rect 33852 29538 33908 33294
rect 34076 33236 34132 33246
rect 34188 33236 34244 33964
rect 34972 33906 35028 33918
rect 34972 33854 34974 33906
rect 35026 33854 35028 33906
rect 34972 33796 35028 33854
rect 35084 33796 35140 33806
rect 34972 33740 35084 33796
rect 35084 33730 35140 33740
rect 35084 33460 35140 33470
rect 35196 33460 35252 34078
rect 35420 33572 35476 33582
rect 35140 33404 35364 33460
rect 35084 33394 35140 33404
rect 34748 33348 34804 33358
rect 34748 33254 34804 33292
rect 34132 33180 34244 33236
rect 34076 33170 34132 33180
rect 34008 32956 35208 32966
rect 34064 32954 34112 32956
rect 34168 32954 34216 32956
rect 34076 32902 34112 32954
rect 34200 32902 34216 32954
rect 34064 32900 34112 32902
rect 34168 32900 34216 32902
rect 34272 32954 34320 32956
rect 34376 32954 34424 32956
rect 34480 32954 34528 32956
rect 34376 32902 34396 32954
rect 34480 32902 34520 32954
rect 34272 32900 34320 32902
rect 34376 32900 34424 32902
rect 34480 32900 34528 32902
rect 34584 32900 34632 32956
rect 34688 32954 34736 32956
rect 34792 32954 34840 32956
rect 34896 32954 34944 32956
rect 34696 32902 34736 32954
rect 34820 32902 34840 32954
rect 34688 32900 34736 32902
rect 34792 32900 34840 32902
rect 34896 32900 34944 32902
rect 35000 32954 35048 32956
rect 35104 32954 35152 32956
rect 35000 32902 35016 32954
rect 35104 32902 35140 32954
rect 35000 32900 35048 32902
rect 35104 32900 35152 32902
rect 34008 32890 35208 32900
rect 34076 32788 34132 32798
rect 34076 32694 34132 32732
rect 34524 32674 34580 32686
rect 34524 32622 34526 32674
rect 34578 32622 34580 32674
rect 34076 32562 34132 32574
rect 34076 32510 34078 32562
rect 34130 32510 34132 32562
rect 33964 31778 34020 31790
rect 33964 31726 33966 31778
rect 34018 31726 34020 31778
rect 33964 31556 34020 31726
rect 34076 31780 34132 32510
rect 34524 32564 34580 32622
rect 34580 32508 34804 32564
rect 34524 32498 34580 32508
rect 34748 31892 34804 32508
rect 34188 31780 34244 31790
rect 34076 31724 34188 31780
rect 34188 31686 34244 31724
rect 34748 31666 34804 31836
rect 34748 31614 34750 31666
rect 34802 31614 34804 31666
rect 34748 31602 34804 31614
rect 35308 32004 35364 33404
rect 35420 33458 35476 33516
rect 35868 33570 35924 34524
rect 36092 34468 36148 34860
rect 36428 34916 36484 34926
rect 36316 34804 36372 34814
rect 36428 34804 36484 34860
rect 36316 34802 36484 34804
rect 36316 34750 36318 34802
rect 36370 34750 36484 34802
rect 36316 34748 36484 34750
rect 36876 34916 36932 34926
rect 36316 34738 36372 34748
rect 36092 34412 36708 34468
rect 36652 34242 36708 34412
rect 36652 34190 36654 34242
rect 36706 34190 36708 34242
rect 36652 34178 36708 34190
rect 36876 34130 36932 34860
rect 37548 34916 37604 34926
rect 37604 34860 37716 34916
rect 37548 34850 37604 34860
rect 36988 34802 37044 34814
rect 36988 34750 36990 34802
rect 37042 34750 37044 34802
rect 36988 34580 37044 34750
rect 37212 34804 37268 34814
rect 37212 34710 37268 34748
rect 37548 34692 37604 34702
rect 37548 34598 37604 34636
rect 36988 34514 37044 34524
rect 36876 34078 36878 34130
rect 36930 34078 36932 34130
rect 36876 34066 36932 34078
rect 37436 34356 37492 34366
rect 35868 33518 35870 33570
rect 35922 33518 35924 33570
rect 35868 33506 35924 33518
rect 36092 33906 36148 33918
rect 36092 33854 36094 33906
rect 36146 33854 36148 33906
rect 35420 33406 35422 33458
rect 35474 33406 35476 33458
rect 35420 33394 35476 33406
rect 35532 33460 35588 33470
rect 35532 33346 35588 33404
rect 35532 33294 35534 33346
rect 35586 33294 35588 33346
rect 35532 33282 35588 33294
rect 36092 32788 36148 33854
rect 36988 33796 37044 33806
rect 36092 32722 36148 32732
rect 36876 33572 36932 33582
rect 36876 32786 36932 33516
rect 36988 33458 37044 33740
rect 37212 33572 37268 33582
rect 36988 33406 36990 33458
rect 37042 33406 37044 33458
rect 36988 33394 37044 33406
rect 37100 33460 37156 33470
rect 36876 32734 36878 32786
rect 36930 32734 36932 32786
rect 36876 32722 36932 32734
rect 36988 32788 37044 32798
rect 36988 32694 37044 32732
rect 37100 32786 37156 33404
rect 37100 32734 37102 32786
rect 37154 32734 37156 32786
rect 37100 32722 37156 32734
rect 37212 33346 37268 33516
rect 37212 33294 37214 33346
rect 37266 33294 37268 33346
rect 33964 31490 34020 31500
rect 34008 31388 35208 31398
rect 34064 31386 34112 31388
rect 34168 31386 34216 31388
rect 34076 31334 34112 31386
rect 34200 31334 34216 31386
rect 34064 31332 34112 31334
rect 34168 31332 34216 31334
rect 34272 31386 34320 31388
rect 34376 31386 34424 31388
rect 34480 31386 34528 31388
rect 34376 31334 34396 31386
rect 34480 31334 34520 31386
rect 34272 31332 34320 31334
rect 34376 31332 34424 31334
rect 34480 31332 34528 31334
rect 34584 31332 34632 31388
rect 34688 31386 34736 31388
rect 34792 31386 34840 31388
rect 34896 31386 34944 31388
rect 34696 31334 34736 31386
rect 34820 31334 34840 31386
rect 34688 31332 34736 31334
rect 34792 31332 34840 31334
rect 34896 31332 34944 31334
rect 35000 31386 35048 31388
rect 35104 31386 35152 31388
rect 35000 31334 35016 31386
rect 35104 31334 35140 31386
rect 35000 31332 35048 31334
rect 35104 31332 35152 31334
rect 34008 31322 35208 31332
rect 35308 31220 35364 31948
rect 35084 31164 35364 31220
rect 35756 32450 35812 32462
rect 37212 32452 37268 33294
rect 37324 33348 37380 33358
rect 37324 32562 37380 33292
rect 37324 32510 37326 32562
rect 37378 32510 37380 32562
rect 37324 32498 37380 32510
rect 37436 32674 37492 34300
rect 37548 33572 37604 33582
rect 37660 33572 37716 34860
rect 37772 34802 37828 34972
rect 37996 34916 38052 35646
rect 38108 35588 38164 35756
rect 38108 35522 38164 35532
rect 37996 34850 38052 34860
rect 38108 35252 38164 35262
rect 37772 34750 37774 34802
rect 37826 34750 37828 34802
rect 37772 34738 37828 34750
rect 37884 34802 37940 34814
rect 37884 34750 37886 34802
rect 37938 34750 37940 34802
rect 37884 34692 37940 34750
rect 38108 34692 38164 35196
rect 37884 34636 38164 34692
rect 37772 34356 37828 34366
rect 37884 34356 37940 34636
rect 37828 34300 37940 34356
rect 37772 34290 37828 34300
rect 37884 34020 37940 34030
rect 37884 33926 37940 33964
rect 37548 33570 37716 33572
rect 37548 33518 37550 33570
rect 37602 33518 37716 33570
rect 37548 33516 37716 33518
rect 37548 33506 37604 33516
rect 37996 33458 38052 34636
rect 37996 33406 37998 33458
rect 38050 33406 38052 33458
rect 37996 33394 38052 33406
rect 37436 32622 37438 32674
rect 37490 32622 37492 32674
rect 35756 32398 35758 32450
rect 35810 32398 35812 32450
rect 34076 31108 34132 31118
rect 34076 31014 34132 31052
rect 35084 31106 35140 31164
rect 35084 31054 35086 31106
rect 35138 31054 35140 31106
rect 35084 31042 35140 31054
rect 35196 30996 35252 31006
rect 35756 30996 35812 32398
rect 36876 32396 37268 32452
rect 35252 30940 35812 30996
rect 36092 32004 36148 32014
rect 35196 30902 35252 30940
rect 36092 30436 36148 31948
rect 36204 31892 36260 31902
rect 36204 31798 36260 31836
rect 36876 31106 36932 32396
rect 37212 31892 37268 31902
rect 37436 31892 37492 32622
rect 37212 31890 37492 31892
rect 37212 31838 37214 31890
rect 37266 31838 37492 31890
rect 37212 31836 37492 31838
rect 37212 31826 37268 31836
rect 36876 31054 36878 31106
rect 36930 31054 36932 31106
rect 36876 31042 36932 31054
rect 36204 30436 36260 30446
rect 36092 30434 36260 30436
rect 36092 30382 36206 30434
rect 36258 30382 36260 30434
rect 36092 30380 36260 30382
rect 36204 30370 36260 30380
rect 34636 30210 34692 30222
rect 34636 30158 34638 30210
rect 34690 30158 34692 30210
rect 34636 29988 34692 30158
rect 34636 29922 34692 29932
rect 34008 29820 35208 29830
rect 34064 29818 34112 29820
rect 34168 29818 34216 29820
rect 34076 29766 34112 29818
rect 34200 29766 34216 29818
rect 34064 29764 34112 29766
rect 34168 29764 34216 29766
rect 34272 29818 34320 29820
rect 34376 29818 34424 29820
rect 34480 29818 34528 29820
rect 34376 29766 34396 29818
rect 34480 29766 34520 29818
rect 34272 29764 34320 29766
rect 34376 29764 34424 29766
rect 34480 29764 34528 29766
rect 34584 29764 34632 29820
rect 34688 29818 34736 29820
rect 34792 29818 34840 29820
rect 34896 29818 34944 29820
rect 34696 29766 34736 29818
rect 34820 29766 34840 29818
rect 34688 29764 34736 29766
rect 34792 29764 34840 29766
rect 34896 29764 34944 29766
rect 35000 29818 35048 29820
rect 35104 29818 35152 29820
rect 35000 29766 35016 29818
rect 35104 29766 35140 29818
rect 35000 29764 35048 29766
rect 35104 29764 35152 29766
rect 34008 29754 35208 29764
rect 33852 29486 33854 29538
rect 33906 29486 33908 29538
rect 33852 29474 33908 29486
rect 33740 29260 33908 29316
rect 33292 28466 33348 28476
rect 33180 28252 33572 28308
rect 33516 27860 33572 28252
rect 33516 27804 33684 27860
rect 33068 26910 33070 26962
rect 33122 26910 33124 26962
rect 33068 26898 33124 26910
rect 33628 26908 33684 27804
rect 33628 26852 33796 26908
rect 32956 25666 33012 25676
rect 33740 25620 33796 26852
rect 33740 25554 33796 25564
rect 33404 25284 33460 25294
rect 33404 25190 33460 25228
rect 31836 24558 31838 24610
rect 31890 24558 31892 24610
rect 31388 23426 31444 23436
rect 31500 23716 31556 23726
rect 31836 23716 31892 24558
rect 31948 23716 32004 23726
rect 31836 23660 31948 23716
rect 31052 23156 31108 23166
rect 30940 23154 31108 23156
rect 30940 23102 31054 23154
rect 31106 23102 31108 23154
rect 30940 23100 31108 23102
rect 30940 22484 30996 22494
rect 30828 22482 30996 22484
rect 30828 22430 30942 22482
rect 30994 22430 30996 22482
rect 30828 22428 30996 22430
rect 30940 22418 30996 22428
rect 30492 22082 30548 22092
rect 30604 22370 30660 22382
rect 30604 22318 30606 22370
rect 30658 22318 30660 22370
rect 30044 20802 30100 21868
rect 30156 21868 30324 21924
rect 30156 21476 30212 21868
rect 30156 21410 30212 21420
rect 30044 20750 30046 20802
rect 30098 20750 30100 20802
rect 30044 19236 30100 20750
rect 30380 20804 30436 20814
rect 30380 20710 30436 20748
rect 30268 20132 30324 20142
rect 30156 20020 30212 20030
rect 30156 19926 30212 19964
rect 30268 20018 30324 20076
rect 30268 19966 30270 20018
rect 30322 19966 30324 20018
rect 30268 19954 30324 19966
rect 30604 20020 30660 22318
rect 31052 21924 31108 23100
rect 31388 22708 31444 22718
rect 31388 22482 31444 22652
rect 31388 22430 31390 22482
rect 31442 22430 31444 22482
rect 31388 22418 31444 22430
rect 31052 21858 31108 21868
rect 30828 20132 30884 20142
rect 30716 20020 30772 20030
rect 30604 20018 30772 20020
rect 30604 19966 30718 20018
rect 30770 19966 30772 20018
rect 30604 19964 30772 19966
rect 30268 19796 30324 19806
rect 30268 19702 30324 19740
rect 29820 19012 29876 19022
rect 29260 19010 29876 19012
rect 29260 18958 29822 19010
rect 29874 18958 29876 19010
rect 29260 18956 29876 18958
rect 29036 18564 29092 18574
rect 29036 18470 29092 18508
rect 28588 18398 28590 18450
rect 28642 18398 28644 18450
rect 28588 18386 28644 18398
rect 28252 18340 28308 18350
rect 28364 18340 28420 18350
rect 28252 18338 28364 18340
rect 28252 18286 28254 18338
rect 28306 18286 28364 18338
rect 28252 18284 28364 18286
rect 28252 18274 28308 18284
rect 28252 17444 28308 17454
rect 28252 17350 28308 17388
rect 27020 16930 27076 16940
rect 26796 16270 26798 16322
rect 26850 16270 26852 16322
rect 26796 16100 26852 16270
rect 26796 16034 26852 16044
rect 26684 15922 26740 15932
rect 27580 15316 27636 15326
rect 26572 15092 26852 15148
rect 26796 13972 26852 15092
rect 26908 15092 26964 15102
rect 26908 14530 26964 15036
rect 26908 14478 26910 14530
rect 26962 14478 26964 14530
rect 26908 14466 26964 14478
rect 27580 14532 27636 15260
rect 28252 15316 28308 15326
rect 28364 15316 28420 18284
rect 29260 17778 29316 18956
rect 29820 18946 29876 18956
rect 29596 18676 29652 18686
rect 29596 18582 29652 18620
rect 29260 17726 29262 17778
rect 29314 17726 29316 17778
rect 29036 15876 29092 15886
rect 28308 15260 28420 15316
rect 28476 15540 28532 15550
rect 28252 15250 28308 15260
rect 27580 14530 28084 14532
rect 27580 14478 27582 14530
rect 27634 14478 28084 14530
rect 27580 14476 28084 14478
rect 27580 14466 27636 14476
rect 27916 14308 27972 14318
rect 28028 14308 28084 14476
rect 28364 14308 28420 14318
rect 28028 14306 28420 14308
rect 28028 14254 28366 14306
rect 28418 14254 28420 14306
rect 28028 14252 28420 14254
rect 27356 13972 27412 13982
rect 26796 13970 27412 13972
rect 26796 13918 26798 13970
rect 26850 13918 27358 13970
rect 27410 13918 27412 13970
rect 26796 13916 27412 13918
rect 26796 13878 26852 13916
rect 27356 13906 27412 13916
rect 26460 13746 26516 13758
rect 26460 13694 26462 13746
rect 26514 13694 26516 13746
rect 26460 13524 26516 13694
rect 26684 13746 26740 13758
rect 26684 13694 26686 13746
rect 26738 13694 26740 13746
rect 26684 13636 26740 13694
rect 26684 13570 26740 13580
rect 26908 13748 26964 13758
rect 26460 13458 26516 13468
rect 26796 13524 26852 13534
rect 26796 13430 26852 13468
rect 26908 13300 26964 13692
rect 27916 13748 27972 14252
rect 27916 13682 27972 13692
rect 26796 13244 26964 13300
rect 26796 13188 26852 13244
rect 26684 13132 26852 13188
rect 27356 13188 27412 13198
rect 26572 13076 26628 13086
rect 26348 13020 26572 13076
rect 26572 12982 26628 13020
rect 25452 11954 25508 11966
rect 25452 11902 25454 11954
rect 25506 11902 25508 11954
rect 24008 11788 25208 11798
rect 24064 11786 24112 11788
rect 24168 11786 24216 11788
rect 24076 11734 24112 11786
rect 24200 11734 24216 11786
rect 24064 11732 24112 11734
rect 24168 11732 24216 11734
rect 24272 11786 24320 11788
rect 24376 11786 24424 11788
rect 24480 11786 24528 11788
rect 24376 11734 24396 11786
rect 24480 11734 24520 11786
rect 24272 11732 24320 11734
rect 24376 11732 24424 11734
rect 24480 11732 24528 11734
rect 24584 11732 24632 11788
rect 24688 11786 24736 11788
rect 24792 11786 24840 11788
rect 24896 11786 24944 11788
rect 24696 11734 24736 11786
rect 24820 11734 24840 11786
rect 24688 11732 24736 11734
rect 24792 11732 24840 11734
rect 24896 11732 24944 11734
rect 25000 11786 25048 11788
rect 25104 11786 25152 11788
rect 25000 11734 25016 11786
rect 25104 11734 25140 11786
rect 25000 11732 25048 11734
rect 25104 11732 25152 11734
rect 24008 11722 25208 11732
rect 25452 11508 25508 11902
rect 25788 11618 25844 12796
rect 25788 11566 25790 11618
rect 25842 11566 25844 11618
rect 25788 11554 25844 11566
rect 25004 11172 25060 11182
rect 25452 11172 25508 11452
rect 26124 11508 26180 11518
rect 26124 11414 26180 11452
rect 26684 11508 26740 13132
rect 27356 12404 27412 13132
rect 27804 12964 27860 12974
rect 27356 12178 27412 12348
rect 27356 12126 27358 12178
rect 27410 12126 27412 12178
rect 27356 12114 27412 12126
rect 27468 12962 27860 12964
rect 27468 12910 27806 12962
rect 27858 12910 27860 12962
rect 27468 12908 27860 12910
rect 26684 11442 26740 11452
rect 25004 11170 25508 11172
rect 25004 11118 25006 11170
rect 25058 11118 25508 11170
rect 25004 11116 25508 11118
rect 26572 11170 26628 11182
rect 26572 11118 26574 11170
rect 26626 11118 26628 11170
rect 23212 10782 23214 10834
rect 23266 10782 23268 10834
rect 23212 10770 23268 10782
rect 23660 10836 23716 10846
rect 23660 10742 23716 10780
rect 25004 10836 25060 11116
rect 25004 10770 25060 10780
rect 20188 10546 20244 10556
rect 16380 10322 16436 10332
rect 18956 9154 19012 9166
rect 18956 9102 18958 9154
rect 19010 9102 19012 9154
rect 18732 9044 18788 9054
rect 18396 9042 18788 9044
rect 18396 8990 18734 9042
rect 18786 8990 18788 9042
rect 18396 8988 18788 8990
rect 17612 8484 17668 8494
rect 17612 8146 17668 8428
rect 17948 8260 18004 8270
rect 17612 8094 17614 8146
rect 17666 8094 17668 8146
rect 15596 7646 15598 7698
rect 15650 7646 15652 7698
rect 15596 7634 15652 7646
rect 16828 7700 16884 7710
rect 16828 7606 16884 7644
rect 13580 7410 13636 7420
rect 14252 7474 14308 7486
rect 14252 7422 14254 7474
rect 14306 7422 14308 7474
rect 14252 6804 14308 7422
rect 14588 7476 14644 7486
rect 14588 7382 14644 7420
rect 15148 7476 15204 7486
rect 15148 7382 15204 7420
rect 17500 7474 17556 7486
rect 17500 7422 17502 7474
rect 17554 7422 17556 7474
rect 14252 6738 14308 6748
rect 15036 6804 15092 6814
rect 15036 6710 15092 6748
rect 13244 6692 13300 6702
rect 12236 6580 12292 6590
rect 13020 6580 13076 6590
rect 11900 6578 12404 6580
rect 11900 6526 12238 6578
rect 12290 6526 12404 6578
rect 11900 6524 12404 6526
rect 10108 5684 10164 5694
rect 9884 5124 9940 5134
rect 9772 5122 9940 5124
rect 9772 5070 9886 5122
rect 9938 5070 9940 5122
rect 9772 5068 9940 5070
rect 8764 4452 8820 4462
rect 8652 4450 8820 4452
rect 8652 4398 8766 4450
rect 8818 4398 8820 4450
rect 8652 4396 8820 4398
rect 8764 4386 8820 4396
rect 6972 4286 6974 4338
rect 7026 4286 7028 4338
rect 6412 3666 6468 4284
rect 6972 4274 7028 4286
rect 7532 4338 8148 4340
rect 7532 4286 8094 4338
rect 8146 4286 8148 4338
rect 7532 4284 8148 4286
rect 7308 4228 7364 4238
rect 7532 4228 7588 4284
rect 8092 4274 8148 4284
rect 7308 4226 7588 4228
rect 7308 4174 7310 4226
rect 7362 4174 7588 4226
rect 7308 4172 7588 4174
rect 7308 4162 7364 4172
rect 6412 3614 6414 3666
rect 6466 3614 6468 3666
rect 6412 3602 6468 3614
rect 8316 3668 8372 3678
rect 8316 3574 8372 3612
rect 9324 3668 9380 5068
rect 9884 5058 9940 5068
rect 9660 4340 9716 4350
rect 9660 4246 9716 4284
rect 10108 4338 10164 5628
rect 11340 5236 11396 5246
rect 11340 5142 11396 5180
rect 11900 5236 11956 6524
rect 12236 6514 12292 6524
rect 12348 6130 12404 6524
rect 13020 6486 13076 6524
rect 12348 6078 12350 6130
rect 12402 6078 12404 6130
rect 12348 6066 12404 6078
rect 13244 6130 13300 6636
rect 16716 6692 16772 6702
rect 13916 6580 13972 6590
rect 13916 6486 13972 6524
rect 16716 6578 16772 6636
rect 17052 6692 17108 6702
rect 17500 6692 17556 7422
rect 17052 6690 17556 6692
rect 17052 6638 17054 6690
rect 17106 6638 17556 6690
rect 17052 6636 17556 6638
rect 16716 6526 16718 6578
rect 16770 6526 16772 6578
rect 16716 6514 16772 6526
rect 16828 6580 16884 6590
rect 16828 6486 16884 6524
rect 16492 6468 16548 6478
rect 16492 6374 16548 6412
rect 14008 6300 15208 6310
rect 14064 6298 14112 6300
rect 14168 6298 14216 6300
rect 14076 6246 14112 6298
rect 14200 6246 14216 6298
rect 14064 6244 14112 6246
rect 14168 6244 14216 6246
rect 14272 6298 14320 6300
rect 14376 6298 14424 6300
rect 14480 6298 14528 6300
rect 14376 6246 14396 6298
rect 14480 6246 14520 6298
rect 14272 6244 14320 6246
rect 14376 6244 14424 6246
rect 14480 6244 14528 6246
rect 14584 6244 14632 6300
rect 14688 6298 14736 6300
rect 14792 6298 14840 6300
rect 14896 6298 14944 6300
rect 14696 6246 14736 6298
rect 14820 6246 14840 6298
rect 14688 6244 14736 6246
rect 14792 6244 14840 6246
rect 14896 6244 14944 6246
rect 15000 6298 15048 6300
rect 15104 6298 15152 6300
rect 15000 6246 15016 6298
rect 15104 6246 15140 6298
rect 15000 6244 15048 6246
rect 15104 6244 15152 6246
rect 14008 6234 15208 6244
rect 13244 6078 13246 6130
rect 13298 6078 13300 6130
rect 13244 6066 13300 6078
rect 13804 6130 13860 6142
rect 13804 6078 13806 6130
rect 13858 6078 13860 6130
rect 13132 5684 13188 5694
rect 13132 5590 13188 5628
rect 11900 5170 11956 5180
rect 13580 5236 13636 5246
rect 13580 5142 13636 5180
rect 10332 5124 10388 5134
rect 10332 5030 10388 5068
rect 10892 5124 10948 5134
rect 10892 5030 10948 5068
rect 13244 5012 13300 5022
rect 12572 4564 12628 4574
rect 12572 4470 12628 4508
rect 10108 4286 10110 4338
rect 10162 4286 10164 4338
rect 10108 4274 10164 4286
rect 13244 4340 13300 4956
rect 13804 4900 13860 6078
rect 16380 5908 16436 5918
rect 16380 5814 16436 5852
rect 16828 5908 16884 5918
rect 17052 5908 17108 6636
rect 17500 6468 17556 6478
rect 17500 6130 17556 6412
rect 17500 6078 17502 6130
rect 17554 6078 17556 6130
rect 17500 6066 17556 6078
rect 17612 6018 17668 8094
rect 17724 8258 18004 8260
rect 17724 8206 17950 8258
rect 18002 8206 18004 8258
rect 17724 8204 18004 8206
rect 17724 6690 17780 8204
rect 17948 8194 18004 8204
rect 18396 8258 18452 8988
rect 18732 8978 18788 8988
rect 18956 8372 19012 9102
rect 19068 9044 19124 9054
rect 19068 9042 19572 9044
rect 19068 8990 19070 9042
rect 19122 8990 19572 9042
rect 19068 8988 19572 8990
rect 19068 8978 19124 8988
rect 19404 8484 19460 8494
rect 19404 8390 19460 8428
rect 18956 8306 19012 8316
rect 18396 8206 18398 8258
rect 18450 8206 18452 8258
rect 18396 8194 18452 8206
rect 18620 8260 18676 8270
rect 18060 8148 18116 8158
rect 18060 8054 18116 8092
rect 17724 6638 17726 6690
rect 17778 6638 17780 6690
rect 17724 6626 17780 6638
rect 17836 8034 17892 8046
rect 17836 7982 17838 8034
rect 17890 7982 17892 8034
rect 17612 5966 17614 6018
rect 17666 5966 17668 6018
rect 17612 5954 17668 5966
rect 16828 5906 17108 5908
rect 16828 5854 16830 5906
rect 16882 5854 17108 5906
rect 16828 5852 17108 5854
rect 17276 5908 17332 5918
rect 17836 5908 17892 7982
rect 18508 8034 18564 8046
rect 18508 7982 18510 8034
rect 18562 7982 18564 8034
rect 18172 7476 18228 7486
rect 18508 7476 18564 7982
rect 18172 7474 18564 7476
rect 18172 7422 18174 7474
rect 18226 7422 18564 7474
rect 18172 7420 18564 7422
rect 18172 7410 18228 7420
rect 18620 6804 18676 8204
rect 19292 8258 19348 8270
rect 19292 8206 19294 8258
rect 19346 8206 19348 8258
rect 18732 8148 18788 8158
rect 18732 8054 18788 8092
rect 18956 8148 19012 8158
rect 18956 8146 19236 8148
rect 18956 8094 18958 8146
rect 19010 8094 19236 8146
rect 18956 8092 19236 8094
rect 18956 8082 19012 8092
rect 18508 6748 18676 6804
rect 18508 6692 18564 6748
rect 18396 6636 18564 6692
rect 18060 6580 18116 6590
rect 18116 6524 18340 6580
rect 18060 6514 18116 6524
rect 18284 6130 18340 6524
rect 18284 6078 18286 6130
rect 18338 6078 18340 6130
rect 18284 6066 18340 6078
rect 18396 6130 18452 6636
rect 18396 6078 18398 6130
rect 18450 6078 18452 6130
rect 18396 6066 18452 6078
rect 18620 6132 18676 6142
rect 18620 6038 18676 6076
rect 18172 5908 18228 5918
rect 17836 5906 18228 5908
rect 17836 5854 18174 5906
rect 18226 5854 18228 5906
rect 17836 5852 18228 5854
rect 14028 5236 14084 5246
rect 14028 5142 14084 5180
rect 15372 5012 15428 5022
rect 15372 4918 15428 4956
rect 16828 5012 16884 5852
rect 17276 5814 17332 5852
rect 16828 4946 16884 4956
rect 13804 4564 13860 4844
rect 14008 4732 15208 4742
rect 14064 4730 14112 4732
rect 14168 4730 14216 4732
rect 14076 4678 14112 4730
rect 14200 4678 14216 4730
rect 14064 4676 14112 4678
rect 14168 4676 14216 4678
rect 14272 4730 14320 4732
rect 14376 4730 14424 4732
rect 14480 4730 14528 4732
rect 14376 4678 14396 4730
rect 14480 4678 14520 4730
rect 14272 4676 14320 4678
rect 14376 4676 14424 4678
rect 14480 4676 14528 4678
rect 14584 4676 14632 4732
rect 14688 4730 14736 4732
rect 14792 4730 14840 4732
rect 14896 4730 14944 4732
rect 14696 4678 14736 4730
rect 14820 4678 14840 4730
rect 14688 4676 14736 4678
rect 14792 4676 14840 4678
rect 14896 4676 14944 4678
rect 15000 4730 15048 4732
rect 15104 4730 15152 4732
rect 15000 4678 15016 4730
rect 15104 4678 15140 4730
rect 15000 4676 15048 4678
rect 15104 4676 15152 4678
rect 14008 4666 15208 4676
rect 13804 4498 13860 4508
rect 16380 4564 16436 4574
rect 16380 4470 16436 4508
rect 18060 4452 18116 4462
rect 18060 4358 18116 4396
rect 13244 4246 13300 4284
rect 13916 4338 13972 4350
rect 13916 4286 13918 4338
rect 13970 4286 13972 4338
rect 13132 4116 13188 4126
rect 13132 4022 13188 4060
rect 9324 3602 9380 3612
rect 13916 3668 13972 4286
rect 16940 4114 16996 4126
rect 16940 4062 16942 4114
rect 16994 4062 16996 4114
rect 16940 4004 16996 4062
rect 16940 3938 16996 3948
rect 17276 4114 17332 4126
rect 17276 4062 17278 4114
rect 17330 4062 17332 4114
rect 17276 3780 17332 4062
rect 17276 3714 17332 3724
rect 17948 4116 18004 4126
rect 13916 3602 13972 3612
rect 16940 3668 16996 3678
rect 16940 3574 16996 3612
rect 9884 3444 9940 3454
rect 9884 800 9940 3388
rect 13244 3444 13300 3482
rect 13244 3378 13300 3388
rect 13692 3444 13748 3482
rect 13692 3378 13748 3388
rect 16156 3444 16212 3482
rect 16156 3378 16212 3388
rect 17948 3442 18004 4060
rect 18172 4004 18228 5852
rect 19180 5796 19236 8092
rect 19292 7700 19348 8206
rect 19516 8260 19572 8988
rect 19516 8194 19572 8204
rect 19740 8372 19796 8382
rect 19516 8036 19572 8046
rect 19516 7942 19572 7980
rect 19740 8034 19796 8316
rect 21196 8260 21252 8270
rect 19964 8148 20020 8158
rect 19964 8054 20020 8092
rect 20300 8146 20356 8158
rect 20300 8094 20302 8146
rect 20354 8094 20356 8146
rect 19740 7982 19742 8034
rect 19794 7982 19796 8034
rect 19292 7634 19348 7644
rect 19740 7700 19796 7982
rect 19740 7634 19796 7644
rect 20188 8034 20244 8046
rect 20188 7982 20190 8034
rect 20242 7982 20244 8034
rect 20076 7588 20132 7598
rect 20076 6466 20132 7532
rect 20076 6414 20078 6466
rect 20130 6414 20132 6466
rect 19180 5740 19796 5796
rect 18172 3938 18228 3948
rect 19068 4452 19124 4462
rect 17948 3390 17950 3442
rect 18002 3390 18004 3442
rect 17948 3378 18004 3390
rect 18732 3444 18788 3482
rect 18732 3378 18788 3388
rect 19068 3442 19124 4396
rect 19740 3778 19796 5740
rect 20076 4564 20132 6414
rect 20188 6132 20244 7982
rect 20300 8036 20356 8094
rect 20300 6916 20356 7980
rect 20636 7698 20692 7710
rect 20636 7646 20638 7698
rect 20690 7646 20692 7698
rect 20636 7588 20692 7646
rect 21196 7700 21252 8204
rect 22316 8258 22372 10668
rect 23996 10724 24052 10734
rect 23996 10630 24052 10668
rect 26572 10724 26628 11118
rect 24008 10220 25208 10230
rect 24064 10218 24112 10220
rect 24168 10218 24216 10220
rect 24076 10166 24112 10218
rect 24200 10166 24216 10218
rect 24064 10164 24112 10166
rect 24168 10164 24216 10166
rect 24272 10218 24320 10220
rect 24376 10218 24424 10220
rect 24480 10218 24528 10220
rect 24376 10166 24396 10218
rect 24480 10166 24520 10218
rect 24272 10164 24320 10166
rect 24376 10164 24424 10166
rect 24480 10164 24528 10166
rect 24584 10164 24632 10220
rect 24688 10218 24736 10220
rect 24792 10218 24840 10220
rect 24896 10218 24944 10220
rect 24696 10166 24736 10218
rect 24820 10166 24840 10218
rect 24688 10164 24736 10166
rect 24792 10164 24840 10166
rect 24896 10164 24944 10166
rect 25000 10218 25048 10220
rect 25104 10218 25152 10220
rect 25000 10166 25016 10218
rect 25104 10166 25140 10218
rect 25000 10164 25048 10166
rect 25104 10164 25152 10166
rect 24008 10154 25208 10164
rect 25788 9940 25844 9950
rect 25340 9044 25396 9054
rect 25340 8950 25396 8988
rect 25788 9042 25844 9884
rect 25788 8990 25790 9042
rect 25842 8990 25844 9042
rect 25788 8978 25844 8990
rect 25900 9716 25956 9726
rect 22988 8820 23044 8830
rect 22316 8206 22318 8258
rect 22370 8206 22372 8258
rect 22316 8194 22372 8206
rect 22876 8818 23044 8820
rect 22876 8766 22990 8818
rect 23042 8766 23044 8818
rect 22876 8764 23044 8766
rect 22876 8258 22932 8764
rect 22988 8754 23044 8764
rect 24008 8652 25208 8662
rect 24064 8650 24112 8652
rect 24168 8650 24216 8652
rect 24076 8598 24112 8650
rect 24200 8598 24216 8650
rect 24064 8596 24112 8598
rect 24168 8596 24216 8598
rect 24272 8650 24320 8652
rect 24376 8650 24424 8652
rect 24480 8650 24528 8652
rect 24376 8598 24396 8650
rect 24480 8598 24520 8650
rect 24272 8596 24320 8598
rect 24376 8596 24424 8598
rect 24480 8596 24528 8598
rect 24584 8596 24632 8652
rect 24688 8650 24736 8652
rect 24792 8650 24840 8652
rect 24896 8650 24944 8652
rect 24696 8598 24736 8650
rect 24820 8598 24840 8650
rect 24688 8596 24736 8598
rect 24792 8596 24840 8598
rect 24896 8596 24944 8598
rect 25000 8650 25048 8652
rect 25104 8650 25152 8652
rect 25000 8598 25016 8650
rect 25104 8598 25140 8650
rect 25000 8596 25048 8598
rect 25104 8596 25152 8598
rect 24008 8586 25208 8596
rect 25900 8370 25956 9660
rect 25900 8318 25902 8370
rect 25954 8318 25956 8370
rect 25900 8306 25956 8318
rect 26348 8372 26404 8382
rect 26572 8372 26628 10668
rect 27020 9940 27076 9950
rect 27020 9846 27076 9884
rect 27468 8428 27524 12908
rect 27804 12898 27860 12908
rect 28252 12404 28308 12414
rect 28252 12310 28308 12348
rect 28028 9716 28084 9726
rect 28028 9622 28084 9660
rect 28028 9156 28084 9166
rect 26348 8370 26628 8372
rect 26348 8318 26350 8370
rect 26402 8318 26628 8370
rect 26348 8316 26628 8318
rect 27244 8372 27524 8428
rect 27580 9154 28084 9156
rect 27580 9102 28030 9154
rect 28082 9102 28084 9154
rect 27580 9100 28084 9102
rect 27580 8482 27636 9100
rect 28028 9090 28084 9100
rect 28252 9156 28308 9166
rect 27580 8430 27582 8482
rect 27634 8430 27636 8482
rect 27244 8370 27300 8372
rect 27244 8318 27246 8370
rect 27298 8318 27300 8370
rect 26348 8306 26404 8316
rect 27244 8306 27300 8318
rect 22876 8206 22878 8258
rect 22930 8206 22932 8258
rect 22876 8194 22932 8206
rect 25340 8034 25396 8046
rect 25340 7982 25342 8034
rect 25394 7982 25396 8034
rect 25340 7812 25396 7982
rect 21420 7700 21476 7710
rect 21196 7698 21364 7700
rect 21196 7646 21198 7698
rect 21250 7646 21364 7698
rect 21196 7644 21364 7646
rect 21196 7634 21252 7644
rect 20636 7522 20692 7532
rect 21308 7140 21364 7644
rect 21420 7606 21476 7644
rect 24668 7586 24724 7598
rect 24668 7534 24670 7586
rect 24722 7534 24724 7586
rect 21532 7362 21588 7374
rect 21532 7310 21534 7362
rect 21586 7310 21588 7362
rect 21308 7084 21476 7140
rect 20300 6850 20356 6860
rect 21308 6916 21364 6926
rect 21308 6822 21364 6860
rect 21420 6802 21476 7084
rect 21420 6750 21422 6802
rect 21474 6750 21476 6802
rect 21420 6738 21476 6750
rect 21084 6692 21140 6702
rect 20188 6066 20244 6076
rect 20748 6466 20804 6478
rect 20748 6414 20750 6466
rect 20802 6414 20804 6466
rect 20748 6132 20804 6414
rect 20748 6066 20804 6076
rect 20412 5124 20468 5134
rect 20412 5030 20468 5068
rect 20076 4498 20132 4508
rect 20412 4338 20468 4350
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4116 20468 4286
rect 20972 4340 21028 4350
rect 21084 4340 21140 6636
rect 21532 6132 21588 7310
rect 24668 7252 24724 7534
rect 24668 7186 24724 7196
rect 24008 7084 25208 7094
rect 24064 7082 24112 7084
rect 24168 7082 24216 7084
rect 24076 7030 24112 7082
rect 24200 7030 24216 7082
rect 24064 7028 24112 7030
rect 24168 7028 24216 7030
rect 24272 7082 24320 7084
rect 24376 7082 24424 7084
rect 24480 7082 24528 7084
rect 24376 7030 24396 7082
rect 24480 7030 24520 7082
rect 24272 7028 24320 7030
rect 24376 7028 24424 7030
rect 24480 7028 24528 7030
rect 24584 7028 24632 7084
rect 24688 7082 24736 7084
rect 24792 7082 24840 7084
rect 24896 7082 24944 7084
rect 24696 7030 24736 7082
rect 24820 7030 24840 7082
rect 24688 7028 24736 7030
rect 24792 7028 24840 7030
rect 24896 7028 24944 7030
rect 25000 7082 25048 7084
rect 25104 7082 25152 7084
rect 25000 7030 25016 7082
rect 25104 7030 25140 7082
rect 25000 7028 25048 7030
rect 25104 7028 25152 7030
rect 24008 7018 25208 7028
rect 25340 6916 25396 7756
rect 26348 7812 26404 7822
rect 26012 7588 26068 7598
rect 26012 7494 26068 7532
rect 26348 7474 26404 7756
rect 26348 7422 26350 7474
rect 26402 7422 26404 7474
rect 26348 7410 26404 7422
rect 26908 7812 26964 7822
rect 25004 6860 25396 6916
rect 25676 7252 25732 7262
rect 22092 6692 22148 6702
rect 22428 6692 22484 6702
rect 22092 6598 22148 6636
rect 22204 6690 22484 6692
rect 22204 6638 22430 6690
rect 22482 6638 22484 6690
rect 22204 6636 22484 6638
rect 21532 6066 21588 6076
rect 22204 5346 22260 6636
rect 22428 6626 22484 6636
rect 25004 6466 25060 6860
rect 25004 6414 25006 6466
rect 25058 6414 25060 6466
rect 25004 6402 25060 6414
rect 25340 6692 25396 6702
rect 24332 5908 24388 5918
rect 24332 5814 24388 5852
rect 25340 5906 25396 6636
rect 25564 6580 25620 6590
rect 25564 6486 25620 6524
rect 25340 5854 25342 5906
rect 25394 5854 25396 5906
rect 22204 5294 22206 5346
rect 22258 5294 22260 5346
rect 22204 5282 22260 5294
rect 22316 5794 22372 5806
rect 22316 5742 22318 5794
rect 22370 5742 22372 5794
rect 21308 5236 21364 5246
rect 20972 4338 21140 4340
rect 20972 4286 20974 4338
rect 21026 4286 21086 4338
rect 21138 4286 21140 4338
rect 20972 4284 21140 4286
rect 20972 4274 21028 4284
rect 21084 4274 21140 4284
rect 21196 5234 21364 5236
rect 21196 5182 21310 5234
rect 21362 5182 21364 5234
rect 21196 5180 21364 5182
rect 21196 4116 21252 5180
rect 21308 5170 21364 5180
rect 22316 5124 22372 5742
rect 24008 5516 25208 5526
rect 24064 5514 24112 5516
rect 24168 5514 24216 5516
rect 24076 5462 24112 5514
rect 24200 5462 24216 5514
rect 24064 5460 24112 5462
rect 24168 5460 24216 5462
rect 24272 5514 24320 5516
rect 24376 5514 24424 5516
rect 24480 5514 24528 5516
rect 24376 5462 24396 5514
rect 24480 5462 24520 5514
rect 24272 5460 24320 5462
rect 24376 5460 24424 5462
rect 24480 5460 24528 5462
rect 24584 5460 24632 5516
rect 24688 5514 24736 5516
rect 24792 5514 24840 5516
rect 24896 5514 24944 5516
rect 24696 5462 24736 5514
rect 24820 5462 24840 5514
rect 24688 5460 24736 5462
rect 24792 5460 24840 5462
rect 24896 5460 24944 5462
rect 25000 5514 25048 5516
rect 25104 5514 25152 5516
rect 25000 5462 25016 5514
rect 25104 5462 25140 5514
rect 25000 5460 25048 5462
rect 25104 5460 25152 5462
rect 24008 5450 25208 5460
rect 25340 5234 25396 5854
rect 25340 5182 25342 5234
rect 25394 5182 25396 5234
rect 25340 5170 25396 5182
rect 22540 5124 22596 5134
rect 22372 5122 22596 5124
rect 22372 5070 22542 5122
rect 22594 5070 22596 5122
rect 22372 5068 22596 5070
rect 22316 5030 22372 5068
rect 22540 5058 22596 5068
rect 23996 4452 24052 4462
rect 23996 4358 24052 4396
rect 24780 4452 24836 4462
rect 24780 4358 24836 4396
rect 20412 4060 21252 4116
rect 21756 4338 21812 4350
rect 21756 4286 21758 4338
rect 21810 4286 21812 4338
rect 19740 3726 19742 3778
rect 19794 3726 19796 3778
rect 19740 3714 19796 3726
rect 19852 4004 19908 4014
rect 19852 3666 19908 3948
rect 19852 3614 19854 3666
rect 19906 3614 19908 3666
rect 19852 3602 19908 3614
rect 20860 3780 20916 3790
rect 19068 3390 19070 3442
rect 19122 3390 19124 3442
rect 19068 3378 19124 3390
rect 20860 3442 20916 3724
rect 21756 3668 21812 4286
rect 25676 4340 25732 7196
rect 26796 6804 26852 6814
rect 25788 6802 26852 6804
rect 25788 6750 26798 6802
rect 26850 6750 26852 6802
rect 25788 6748 26852 6750
rect 25788 5906 25844 6748
rect 26796 6738 26852 6748
rect 25788 5854 25790 5906
rect 25842 5854 25844 5906
rect 25788 5842 25844 5854
rect 26012 6468 26068 6478
rect 26012 5908 26068 6412
rect 26012 5842 26068 5852
rect 26908 4562 26964 7756
rect 27580 7812 27636 8430
rect 28252 8258 28308 9100
rect 28364 9044 28420 14252
rect 28476 14308 28532 15484
rect 29036 15538 29092 15820
rect 29036 15486 29038 15538
rect 29090 15486 29092 15538
rect 29036 15474 29092 15486
rect 29260 15540 29316 17726
rect 29708 18450 29764 18462
rect 29708 18398 29710 18450
rect 29762 18398 29764 18450
rect 29708 17444 29764 18398
rect 30044 18340 30100 19180
rect 30604 18676 30660 19964
rect 30716 19954 30772 19964
rect 30604 18610 30660 18620
rect 30828 18564 30884 20076
rect 30940 19908 30996 19918
rect 30940 19814 30996 19852
rect 31500 19906 31556 23660
rect 31948 23622 32004 23660
rect 31612 23492 31668 23502
rect 31612 23380 31668 23436
rect 31612 23378 31892 23380
rect 31612 23326 31614 23378
rect 31666 23326 31892 23378
rect 31612 23324 31892 23326
rect 31612 23314 31668 23324
rect 31836 21810 31892 23324
rect 31836 21758 31838 21810
rect 31890 21758 31892 21810
rect 31836 20692 31892 21758
rect 33628 22708 33684 22718
rect 33516 21028 33572 21038
rect 33628 21028 33684 22652
rect 33852 22596 33908 29260
rect 34008 28252 35208 28262
rect 34064 28250 34112 28252
rect 34168 28250 34216 28252
rect 34076 28198 34112 28250
rect 34200 28198 34216 28250
rect 34064 28196 34112 28198
rect 34168 28196 34216 28198
rect 34272 28250 34320 28252
rect 34376 28250 34424 28252
rect 34480 28250 34528 28252
rect 34376 28198 34396 28250
rect 34480 28198 34520 28250
rect 34272 28196 34320 28198
rect 34376 28196 34424 28198
rect 34480 28196 34528 28198
rect 34584 28196 34632 28252
rect 34688 28250 34736 28252
rect 34792 28250 34840 28252
rect 34896 28250 34944 28252
rect 34696 28198 34736 28250
rect 34820 28198 34840 28250
rect 34688 28196 34736 28198
rect 34792 28196 34840 28198
rect 34896 28196 34944 28198
rect 35000 28250 35048 28252
rect 35104 28250 35152 28252
rect 35000 28198 35016 28250
rect 35104 28198 35140 28250
rect 35000 28196 35048 28198
rect 35104 28196 35152 28198
rect 34008 28186 35208 28196
rect 33964 28084 34020 28094
rect 33964 27074 34020 28028
rect 33964 27022 33966 27074
rect 34018 27022 34020 27074
rect 33964 27010 34020 27022
rect 34008 26684 35208 26694
rect 34064 26682 34112 26684
rect 34168 26682 34216 26684
rect 34076 26630 34112 26682
rect 34200 26630 34216 26682
rect 34064 26628 34112 26630
rect 34168 26628 34216 26630
rect 34272 26682 34320 26684
rect 34376 26682 34424 26684
rect 34480 26682 34528 26684
rect 34376 26630 34396 26682
rect 34480 26630 34520 26682
rect 34272 26628 34320 26630
rect 34376 26628 34424 26630
rect 34480 26628 34528 26630
rect 34584 26628 34632 26684
rect 34688 26682 34736 26684
rect 34792 26682 34840 26684
rect 34896 26682 34944 26684
rect 34696 26630 34736 26682
rect 34820 26630 34840 26682
rect 34688 26628 34736 26630
rect 34792 26628 34840 26630
rect 34896 26628 34944 26630
rect 35000 26682 35048 26684
rect 35104 26682 35152 26684
rect 35000 26630 35016 26682
rect 35104 26630 35140 26682
rect 35000 26628 35048 26630
rect 35104 26628 35152 26630
rect 34008 26618 35208 26628
rect 34188 25732 34244 25742
rect 34188 25638 34244 25676
rect 34008 25116 35208 25126
rect 34064 25114 34112 25116
rect 34168 25114 34216 25116
rect 34076 25062 34112 25114
rect 34200 25062 34216 25114
rect 34064 25060 34112 25062
rect 34168 25060 34216 25062
rect 34272 25114 34320 25116
rect 34376 25114 34424 25116
rect 34480 25114 34528 25116
rect 34376 25062 34396 25114
rect 34480 25062 34520 25114
rect 34272 25060 34320 25062
rect 34376 25060 34424 25062
rect 34480 25060 34528 25062
rect 34584 25060 34632 25116
rect 34688 25114 34736 25116
rect 34792 25114 34840 25116
rect 34896 25114 34944 25116
rect 34696 25062 34736 25114
rect 34820 25062 34840 25114
rect 34688 25060 34736 25062
rect 34792 25060 34840 25062
rect 34896 25060 34944 25062
rect 35000 25114 35048 25116
rect 35104 25114 35152 25116
rect 35000 25062 35016 25114
rect 35104 25062 35140 25114
rect 35000 25060 35048 25062
rect 35104 25060 35152 25062
rect 34008 25050 35208 25060
rect 34008 23548 35208 23558
rect 34064 23546 34112 23548
rect 34168 23546 34216 23548
rect 34076 23494 34112 23546
rect 34200 23494 34216 23546
rect 34064 23492 34112 23494
rect 34168 23492 34216 23494
rect 34272 23546 34320 23548
rect 34376 23546 34424 23548
rect 34480 23546 34528 23548
rect 34376 23494 34396 23546
rect 34480 23494 34520 23546
rect 34272 23492 34320 23494
rect 34376 23492 34424 23494
rect 34480 23492 34528 23494
rect 34584 23492 34632 23548
rect 34688 23546 34736 23548
rect 34792 23546 34840 23548
rect 34896 23546 34944 23548
rect 34696 23494 34736 23546
rect 34820 23494 34840 23546
rect 34688 23492 34736 23494
rect 34792 23492 34840 23494
rect 34896 23492 34944 23494
rect 35000 23546 35048 23548
rect 35104 23546 35152 23548
rect 35000 23494 35016 23546
rect 35104 23494 35140 23546
rect 35000 23492 35048 23494
rect 35104 23492 35152 23494
rect 34008 23482 35208 23492
rect 33852 22530 33908 22540
rect 34008 21980 35208 21990
rect 34064 21978 34112 21980
rect 34168 21978 34216 21980
rect 34076 21926 34112 21978
rect 34200 21926 34216 21978
rect 34064 21924 34112 21926
rect 34168 21924 34216 21926
rect 34272 21978 34320 21980
rect 34376 21978 34424 21980
rect 34480 21978 34528 21980
rect 34376 21926 34396 21978
rect 34480 21926 34520 21978
rect 34272 21924 34320 21926
rect 34376 21924 34424 21926
rect 34480 21924 34528 21926
rect 34584 21924 34632 21980
rect 34688 21978 34736 21980
rect 34792 21978 34840 21980
rect 34896 21978 34944 21980
rect 34696 21926 34736 21978
rect 34820 21926 34840 21978
rect 34688 21924 34736 21926
rect 34792 21924 34840 21926
rect 34896 21924 34944 21926
rect 35000 21978 35048 21980
rect 35104 21978 35152 21980
rect 35000 21926 35016 21978
rect 35104 21926 35140 21978
rect 35000 21924 35048 21926
rect 35104 21924 35152 21926
rect 34008 21914 35208 21924
rect 33516 21026 33684 21028
rect 33516 20974 33518 21026
rect 33570 20974 33684 21026
rect 33516 20972 33684 20974
rect 33516 20962 33572 20972
rect 31836 20626 31892 20636
rect 32732 20692 32788 20702
rect 32732 20598 32788 20636
rect 31948 20132 32004 20142
rect 31948 20038 32004 20076
rect 33628 20132 33684 20972
rect 34008 20412 35208 20422
rect 34064 20410 34112 20412
rect 34168 20410 34216 20412
rect 34076 20358 34112 20410
rect 34200 20358 34216 20410
rect 34064 20356 34112 20358
rect 34168 20356 34216 20358
rect 34272 20410 34320 20412
rect 34376 20410 34424 20412
rect 34480 20410 34528 20412
rect 34376 20358 34396 20410
rect 34480 20358 34520 20410
rect 34272 20356 34320 20358
rect 34376 20356 34424 20358
rect 34480 20356 34528 20358
rect 34584 20356 34632 20412
rect 34688 20410 34736 20412
rect 34792 20410 34840 20412
rect 34896 20410 34944 20412
rect 34696 20358 34736 20410
rect 34820 20358 34840 20410
rect 34688 20356 34736 20358
rect 34792 20356 34840 20358
rect 34896 20356 34944 20358
rect 35000 20410 35048 20412
rect 35104 20410 35152 20412
rect 35000 20358 35016 20410
rect 35104 20358 35140 20410
rect 35000 20356 35048 20358
rect 35104 20356 35152 20358
rect 34008 20346 35208 20356
rect 33628 20066 33684 20076
rect 31500 19854 31502 19906
rect 31554 19854 31556 19906
rect 31500 19684 31556 19854
rect 31500 19618 31556 19628
rect 32284 19796 32340 19806
rect 32284 19234 32340 19740
rect 32284 19182 32286 19234
rect 32338 19182 32340 19234
rect 32284 19170 32340 19182
rect 32732 19236 32788 19246
rect 32732 19142 32788 19180
rect 34008 18844 35208 18854
rect 34064 18842 34112 18844
rect 34168 18842 34216 18844
rect 34076 18790 34112 18842
rect 34200 18790 34216 18842
rect 34064 18788 34112 18790
rect 34168 18788 34216 18790
rect 34272 18842 34320 18844
rect 34376 18842 34424 18844
rect 34480 18842 34528 18844
rect 34376 18790 34396 18842
rect 34480 18790 34520 18842
rect 34272 18788 34320 18790
rect 34376 18788 34424 18790
rect 34480 18788 34528 18790
rect 34584 18788 34632 18844
rect 34688 18842 34736 18844
rect 34792 18842 34840 18844
rect 34896 18842 34944 18844
rect 34696 18790 34736 18842
rect 34820 18790 34840 18842
rect 34688 18788 34736 18790
rect 34792 18788 34840 18790
rect 34896 18788 34944 18790
rect 35000 18842 35048 18844
rect 35104 18842 35152 18844
rect 35000 18790 35016 18842
rect 35104 18790 35140 18842
rect 35000 18788 35048 18790
rect 35104 18788 35152 18790
rect 34008 18778 35208 18788
rect 30716 18452 30772 18462
rect 30828 18452 30884 18508
rect 30716 18450 30884 18452
rect 30716 18398 30718 18450
rect 30770 18398 30884 18450
rect 30716 18396 30884 18398
rect 30716 18386 30772 18396
rect 30156 18340 30212 18350
rect 30044 18284 30156 18340
rect 30156 18246 30212 18284
rect 29372 16324 29428 16334
rect 29372 16210 29428 16268
rect 29372 16158 29374 16210
rect 29426 16158 29428 16210
rect 29372 16146 29428 16158
rect 29708 16100 29764 17388
rect 34008 17276 35208 17286
rect 34064 17274 34112 17276
rect 34168 17274 34216 17276
rect 34076 17222 34112 17274
rect 34200 17222 34216 17274
rect 34064 17220 34112 17222
rect 34168 17220 34216 17222
rect 34272 17274 34320 17276
rect 34376 17274 34424 17276
rect 34480 17274 34528 17276
rect 34376 17222 34396 17274
rect 34480 17222 34520 17274
rect 34272 17220 34320 17222
rect 34376 17220 34424 17222
rect 34480 17220 34528 17222
rect 34584 17220 34632 17276
rect 34688 17274 34736 17276
rect 34792 17274 34840 17276
rect 34896 17274 34944 17276
rect 34696 17222 34736 17274
rect 34820 17222 34840 17274
rect 34688 17220 34736 17222
rect 34792 17220 34840 17222
rect 34896 17220 34944 17222
rect 35000 17274 35048 17276
rect 35104 17274 35152 17276
rect 35000 17222 35016 17274
rect 35104 17222 35140 17274
rect 35000 17220 35048 17222
rect 35104 17220 35152 17222
rect 34008 17210 35208 17220
rect 30380 16324 30436 16334
rect 30380 16230 30436 16268
rect 29932 16100 29988 16110
rect 30268 16100 30324 16110
rect 29708 16098 30324 16100
rect 29708 16046 29934 16098
rect 29986 16046 30270 16098
rect 30322 16046 30324 16098
rect 29708 16044 30324 16046
rect 29932 16034 29988 16044
rect 30268 16034 30324 16044
rect 34008 15708 35208 15718
rect 34064 15706 34112 15708
rect 34168 15706 34216 15708
rect 34076 15654 34112 15706
rect 34200 15654 34216 15706
rect 34064 15652 34112 15654
rect 34168 15652 34216 15654
rect 34272 15706 34320 15708
rect 34376 15706 34424 15708
rect 34480 15706 34528 15708
rect 34376 15654 34396 15706
rect 34480 15654 34520 15706
rect 34272 15652 34320 15654
rect 34376 15652 34424 15654
rect 34480 15652 34528 15654
rect 34584 15652 34632 15708
rect 34688 15706 34736 15708
rect 34792 15706 34840 15708
rect 34896 15706 34944 15708
rect 34696 15654 34736 15706
rect 34820 15654 34840 15706
rect 34688 15652 34736 15654
rect 34792 15652 34840 15654
rect 34896 15652 34944 15654
rect 35000 15706 35048 15708
rect 35104 15706 35152 15708
rect 35000 15654 35016 15706
rect 35104 15654 35140 15706
rect 35000 15652 35048 15654
rect 35104 15652 35152 15654
rect 34008 15642 35208 15652
rect 29596 15540 29652 15550
rect 29316 15538 29652 15540
rect 29316 15486 29598 15538
rect 29650 15486 29652 15538
rect 29316 15484 29652 15486
rect 29260 15474 29316 15484
rect 29596 15474 29652 15484
rect 30044 15426 30100 15438
rect 30044 15374 30046 15426
rect 30098 15374 30100 15426
rect 29932 15316 29988 15326
rect 30044 15316 30100 15374
rect 29988 15260 30100 15316
rect 29932 15250 29988 15260
rect 28476 14242 28532 14252
rect 34008 14140 35208 14150
rect 34064 14138 34112 14140
rect 34168 14138 34216 14140
rect 34076 14086 34112 14138
rect 34200 14086 34216 14138
rect 34064 14084 34112 14086
rect 34168 14084 34216 14086
rect 34272 14138 34320 14140
rect 34376 14138 34424 14140
rect 34480 14138 34528 14140
rect 34376 14086 34396 14138
rect 34480 14086 34520 14138
rect 34272 14084 34320 14086
rect 34376 14084 34424 14086
rect 34480 14084 34528 14086
rect 34584 14084 34632 14140
rect 34688 14138 34736 14140
rect 34792 14138 34840 14140
rect 34896 14138 34944 14140
rect 34696 14086 34736 14138
rect 34820 14086 34840 14138
rect 34688 14084 34736 14086
rect 34792 14084 34840 14086
rect 34896 14084 34944 14086
rect 35000 14138 35048 14140
rect 35104 14138 35152 14140
rect 35000 14086 35016 14138
rect 35104 14086 35140 14138
rect 35000 14084 35048 14086
rect 35104 14084 35152 14086
rect 34008 14074 35208 14084
rect 34008 12572 35208 12582
rect 34064 12570 34112 12572
rect 34168 12570 34216 12572
rect 34076 12518 34112 12570
rect 34200 12518 34216 12570
rect 34064 12516 34112 12518
rect 34168 12516 34216 12518
rect 34272 12570 34320 12572
rect 34376 12570 34424 12572
rect 34480 12570 34528 12572
rect 34376 12518 34396 12570
rect 34480 12518 34520 12570
rect 34272 12516 34320 12518
rect 34376 12516 34424 12518
rect 34480 12516 34528 12518
rect 34584 12516 34632 12572
rect 34688 12570 34736 12572
rect 34792 12570 34840 12572
rect 34896 12570 34944 12572
rect 34696 12518 34736 12570
rect 34820 12518 34840 12570
rect 34688 12516 34736 12518
rect 34792 12516 34840 12518
rect 34896 12516 34944 12518
rect 35000 12570 35048 12572
rect 35104 12570 35152 12572
rect 35000 12518 35016 12570
rect 35104 12518 35140 12570
rect 35000 12516 35048 12518
rect 35104 12516 35152 12518
rect 34008 12506 35208 12516
rect 34008 11004 35208 11014
rect 34064 11002 34112 11004
rect 34168 11002 34216 11004
rect 34076 10950 34112 11002
rect 34200 10950 34216 11002
rect 34064 10948 34112 10950
rect 34168 10948 34216 10950
rect 34272 11002 34320 11004
rect 34376 11002 34424 11004
rect 34480 11002 34528 11004
rect 34376 10950 34396 11002
rect 34480 10950 34520 11002
rect 34272 10948 34320 10950
rect 34376 10948 34424 10950
rect 34480 10948 34528 10950
rect 34584 10948 34632 11004
rect 34688 11002 34736 11004
rect 34792 11002 34840 11004
rect 34896 11002 34944 11004
rect 34696 10950 34736 11002
rect 34820 10950 34840 11002
rect 34688 10948 34736 10950
rect 34792 10948 34840 10950
rect 34896 10948 34944 10950
rect 35000 11002 35048 11004
rect 35104 11002 35152 11004
rect 35000 10950 35016 11002
rect 35104 10950 35140 11002
rect 35000 10948 35048 10950
rect 35104 10948 35152 10950
rect 34008 10938 35208 10948
rect 34008 9436 35208 9446
rect 34064 9434 34112 9436
rect 34168 9434 34216 9436
rect 34076 9382 34112 9434
rect 34200 9382 34216 9434
rect 34064 9380 34112 9382
rect 34168 9380 34216 9382
rect 34272 9434 34320 9436
rect 34376 9434 34424 9436
rect 34480 9434 34528 9436
rect 34376 9382 34396 9434
rect 34480 9382 34520 9434
rect 34272 9380 34320 9382
rect 34376 9380 34424 9382
rect 34480 9380 34528 9382
rect 34584 9380 34632 9436
rect 34688 9434 34736 9436
rect 34792 9434 34840 9436
rect 34896 9434 34944 9436
rect 34696 9382 34736 9434
rect 34820 9382 34840 9434
rect 34688 9380 34736 9382
rect 34792 9380 34840 9382
rect 34896 9380 34944 9382
rect 35000 9434 35048 9436
rect 35104 9434 35152 9436
rect 35000 9382 35016 9434
rect 35104 9382 35140 9434
rect 35000 9380 35048 9382
rect 35104 9380 35152 9382
rect 34008 9370 35208 9380
rect 29036 9156 29092 9166
rect 29036 9062 29092 9100
rect 28364 8978 28420 8988
rect 29596 9044 29652 9054
rect 29596 8950 29652 8988
rect 28812 8818 28868 8830
rect 28812 8766 28814 8818
rect 28866 8766 28868 8818
rect 28812 8428 28868 8766
rect 28252 8206 28254 8258
rect 28306 8206 28308 8258
rect 28252 8194 28308 8206
rect 28364 8372 28868 8428
rect 28364 8146 28420 8372
rect 28364 8094 28366 8146
rect 28418 8094 28420 8146
rect 28364 8082 28420 8094
rect 34008 7868 35208 7878
rect 34064 7866 34112 7868
rect 34168 7866 34216 7868
rect 27580 7746 27636 7756
rect 28140 7812 28196 7822
rect 34076 7814 34112 7866
rect 34200 7814 34216 7866
rect 34064 7812 34112 7814
rect 34168 7812 34216 7814
rect 34272 7866 34320 7868
rect 34376 7866 34424 7868
rect 34480 7866 34528 7868
rect 34376 7814 34396 7866
rect 34480 7814 34520 7866
rect 34272 7812 34320 7814
rect 34376 7812 34424 7814
rect 34480 7812 34528 7814
rect 34584 7812 34632 7868
rect 34688 7866 34736 7868
rect 34792 7866 34840 7868
rect 34896 7866 34944 7868
rect 34696 7814 34736 7866
rect 34820 7814 34840 7866
rect 34688 7812 34736 7814
rect 34792 7812 34840 7814
rect 34896 7812 34944 7814
rect 35000 7866 35048 7868
rect 35104 7866 35152 7868
rect 35000 7814 35016 7866
rect 35104 7814 35140 7866
rect 35000 7812 35048 7814
rect 35104 7812 35152 7814
rect 34008 7802 35208 7812
rect 27020 7586 27076 7598
rect 27020 7534 27022 7586
rect 27074 7534 27076 7586
rect 27020 6132 27076 7534
rect 27580 7586 27636 7598
rect 27580 7534 27582 7586
rect 27634 7534 27636 7586
rect 27132 7476 27188 7486
rect 27580 7476 27636 7534
rect 27132 7474 27636 7476
rect 27132 7422 27134 7474
rect 27186 7422 27636 7474
rect 27132 7420 27636 7422
rect 27132 7410 27188 7420
rect 27804 6580 27860 6590
rect 27804 6486 27860 6524
rect 27020 6066 27076 6076
rect 28140 6130 28196 7756
rect 29820 6468 29876 6478
rect 28140 6078 28142 6130
rect 28194 6078 28196 6130
rect 28140 6066 28196 6078
rect 28812 6132 28868 6142
rect 28812 6038 28868 6076
rect 26908 4510 26910 4562
rect 26962 4510 26964 4562
rect 26908 4498 26964 4510
rect 25900 4452 25956 4462
rect 25900 4358 25956 4396
rect 25788 4340 25844 4350
rect 25676 4338 25844 4340
rect 25676 4286 25790 4338
rect 25842 4286 25844 4338
rect 25676 4284 25844 4286
rect 25788 4274 25844 4284
rect 25452 4226 25508 4238
rect 25452 4174 25454 4226
rect 25506 4174 25508 4226
rect 25452 4116 25508 4174
rect 24008 3948 25208 3958
rect 24064 3946 24112 3948
rect 24168 3946 24216 3948
rect 24076 3894 24112 3946
rect 24200 3894 24216 3946
rect 24064 3892 24112 3894
rect 24168 3892 24216 3894
rect 24272 3946 24320 3948
rect 24376 3946 24424 3948
rect 24480 3946 24528 3948
rect 24376 3894 24396 3946
rect 24480 3894 24520 3946
rect 24272 3892 24320 3894
rect 24376 3892 24424 3894
rect 24480 3892 24528 3894
rect 24584 3892 24632 3948
rect 24688 3946 24736 3948
rect 24792 3946 24840 3948
rect 24896 3946 24944 3948
rect 24696 3894 24736 3946
rect 24820 3894 24840 3946
rect 24688 3892 24736 3894
rect 24792 3892 24840 3894
rect 24896 3892 24944 3894
rect 25000 3946 25048 3948
rect 25104 3946 25152 3948
rect 25000 3894 25016 3946
rect 25104 3894 25140 3946
rect 25000 3892 25048 3894
rect 25104 3892 25152 3894
rect 24008 3882 25208 3892
rect 21980 3668 22036 3678
rect 21756 3666 22036 3668
rect 21756 3614 21982 3666
rect 22034 3614 22036 3666
rect 21756 3612 22036 3614
rect 21980 3602 22036 3612
rect 25452 3556 25508 4060
rect 26572 4116 26628 4126
rect 26572 4022 26628 4060
rect 25452 3490 25508 3500
rect 20860 3390 20862 3442
rect 20914 3390 20916 3442
rect 20860 3378 20916 3390
rect 14008 3164 15208 3174
rect 14064 3162 14112 3164
rect 14168 3162 14216 3164
rect 14076 3110 14112 3162
rect 14200 3110 14216 3162
rect 14064 3108 14112 3110
rect 14168 3108 14216 3110
rect 14272 3162 14320 3164
rect 14376 3162 14424 3164
rect 14480 3162 14528 3164
rect 14376 3110 14396 3162
rect 14480 3110 14520 3162
rect 14272 3108 14320 3110
rect 14376 3108 14424 3110
rect 14480 3108 14528 3110
rect 14584 3108 14632 3164
rect 14688 3162 14736 3164
rect 14792 3162 14840 3164
rect 14896 3162 14944 3164
rect 14696 3110 14736 3162
rect 14820 3110 14840 3162
rect 14688 3108 14736 3110
rect 14792 3108 14840 3110
rect 14896 3108 14944 3110
rect 15000 3162 15048 3164
rect 15104 3162 15152 3164
rect 15000 3110 15016 3162
rect 15104 3110 15140 3162
rect 15000 3108 15048 3110
rect 15104 3108 15152 3110
rect 14008 3098 15208 3108
rect 29820 800 29876 6412
rect 34008 6300 35208 6310
rect 34064 6298 34112 6300
rect 34168 6298 34216 6300
rect 34076 6246 34112 6298
rect 34200 6246 34216 6298
rect 34064 6244 34112 6246
rect 34168 6244 34216 6246
rect 34272 6298 34320 6300
rect 34376 6298 34424 6300
rect 34480 6298 34528 6300
rect 34376 6246 34396 6298
rect 34480 6246 34520 6298
rect 34272 6244 34320 6246
rect 34376 6244 34424 6246
rect 34480 6244 34528 6246
rect 34584 6244 34632 6300
rect 34688 6298 34736 6300
rect 34792 6298 34840 6300
rect 34896 6298 34944 6300
rect 34696 6246 34736 6298
rect 34820 6246 34840 6298
rect 34688 6244 34736 6246
rect 34792 6244 34840 6246
rect 34896 6244 34944 6246
rect 35000 6298 35048 6300
rect 35104 6298 35152 6300
rect 35000 6246 35016 6298
rect 35104 6246 35140 6298
rect 35000 6244 35048 6246
rect 35104 6244 35152 6246
rect 34008 6234 35208 6244
rect 34008 4732 35208 4742
rect 34064 4730 34112 4732
rect 34168 4730 34216 4732
rect 34076 4678 34112 4730
rect 34200 4678 34216 4730
rect 34064 4676 34112 4678
rect 34168 4676 34216 4678
rect 34272 4730 34320 4732
rect 34376 4730 34424 4732
rect 34480 4730 34528 4732
rect 34376 4678 34396 4730
rect 34480 4678 34520 4730
rect 34272 4676 34320 4678
rect 34376 4676 34424 4678
rect 34480 4676 34528 4678
rect 34584 4676 34632 4732
rect 34688 4730 34736 4732
rect 34792 4730 34840 4732
rect 34896 4730 34944 4732
rect 34696 4678 34736 4730
rect 34820 4678 34840 4730
rect 34688 4676 34736 4678
rect 34792 4676 34840 4678
rect 34896 4676 34944 4678
rect 35000 4730 35048 4732
rect 35104 4730 35152 4732
rect 35000 4678 35016 4730
rect 35104 4678 35140 4730
rect 35000 4676 35048 4678
rect 35104 4676 35152 4678
rect 34008 4666 35208 4676
rect 34008 3164 35208 3174
rect 34064 3162 34112 3164
rect 34168 3162 34216 3164
rect 34076 3110 34112 3162
rect 34200 3110 34216 3162
rect 34064 3108 34112 3110
rect 34168 3108 34216 3110
rect 34272 3162 34320 3164
rect 34376 3162 34424 3164
rect 34480 3162 34528 3164
rect 34376 3110 34396 3162
rect 34480 3110 34520 3162
rect 34272 3108 34320 3110
rect 34376 3108 34424 3110
rect 34480 3108 34528 3110
rect 34584 3108 34632 3164
rect 34688 3162 34736 3164
rect 34792 3162 34840 3164
rect 34896 3162 34944 3164
rect 34696 3110 34736 3162
rect 34820 3110 34840 3162
rect 34688 3108 34736 3110
rect 34792 3108 34840 3110
rect 34896 3108 34944 3110
rect 35000 3162 35048 3164
rect 35104 3162 35152 3164
rect 35000 3110 35016 3162
rect 35104 3110 35140 3162
rect 35000 3108 35048 3110
rect 35104 3108 35152 3110
rect 34008 3098 35208 3108
rect 9856 0 9968 800
rect 29792 0 29904 800
<< via2 >>
rect 4008 96458 4064 96460
rect 4112 96458 4168 96460
rect 4008 96406 4024 96458
rect 4024 96406 4064 96458
rect 4112 96406 4148 96458
rect 4148 96406 4168 96458
rect 4008 96404 4064 96406
rect 4112 96404 4168 96406
rect 4216 96404 4272 96460
rect 4320 96458 4376 96460
rect 4424 96458 4480 96460
rect 4528 96458 4584 96460
rect 4320 96406 4324 96458
rect 4324 96406 4376 96458
rect 4424 96406 4448 96458
rect 4448 96406 4480 96458
rect 4528 96406 4572 96458
rect 4572 96406 4584 96458
rect 4320 96404 4376 96406
rect 4424 96404 4480 96406
rect 4528 96404 4584 96406
rect 4632 96458 4688 96460
rect 4736 96458 4792 96460
rect 4840 96458 4896 96460
rect 4632 96406 4644 96458
rect 4644 96406 4688 96458
rect 4736 96406 4768 96458
rect 4768 96406 4792 96458
rect 4840 96406 4892 96458
rect 4892 96406 4896 96458
rect 4632 96404 4688 96406
rect 4736 96404 4792 96406
rect 4840 96404 4896 96406
rect 4944 96404 5000 96460
rect 5048 96458 5104 96460
rect 5152 96458 5208 96460
rect 5048 96406 5068 96458
rect 5068 96406 5104 96458
rect 5152 96406 5192 96458
rect 5192 96406 5208 96458
rect 5048 96404 5104 96406
rect 5152 96404 5208 96406
rect 1708 95228 1764 95284
rect 4008 94890 4064 94892
rect 4112 94890 4168 94892
rect 4008 94838 4024 94890
rect 4024 94838 4064 94890
rect 4112 94838 4148 94890
rect 4148 94838 4168 94890
rect 4008 94836 4064 94838
rect 4112 94836 4168 94838
rect 4216 94836 4272 94892
rect 4320 94890 4376 94892
rect 4424 94890 4480 94892
rect 4528 94890 4584 94892
rect 4320 94838 4324 94890
rect 4324 94838 4376 94890
rect 4424 94838 4448 94890
rect 4448 94838 4480 94890
rect 4528 94838 4572 94890
rect 4572 94838 4584 94890
rect 4320 94836 4376 94838
rect 4424 94836 4480 94838
rect 4528 94836 4584 94838
rect 4632 94890 4688 94892
rect 4736 94890 4792 94892
rect 4840 94890 4896 94892
rect 4632 94838 4644 94890
rect 4644 94838 4688 94890
rect 4736 94838 4768 94890
rect 4768 94838 4792 94890
rect 4840 94838 4892 94890
rect 4892 94838 4896 94890
rect 4632 94836 4688 94838
rect 4736 94836 4792 94838
rect 4840 94836 4896 94838
rect 4944 94836 5000 94892
rect 5048 94890 5104 94892
rect 5152 94890 5208 94892
rect 5048 94838 5068 94890
rect 5068 94838 5104 94890
rect 5152 94838 5192 94890
rect 5192 94838 5208 94890
rect 5048 94836 5104 94838
rect 5152 94836 5208 94838
rect 1708 94274 1764 94276
rect 1708 94222 1710 94274
rect 1710 94222 1762 94274
rect 1762 94222 1764 94274
rect 1708 94220 1764 94222
rect 24008 96458 24064 96460
rect 24112 96458 24168 96460
rect 24008 96406 24024 96458
rect 24024 96406 24064 96458
rect 24112 96406 24148 96458
rect 24148 96406 24168 96458
rect 24008 96404 24064 96406
rect 24112 96404 24168 96406
rect 24216 96404 24272 96460
rect 24320 96458 24376 96460
rect 24424 96458 24480 96460
rect 24528 96458 24584 96460
rect 24320 96406 24324 96458
rect 24324 96406 24376 96458
rect 24424 96406 24448 96458
rect 24448 96406 24480 96458
rect 24528 96406 24572 96458
rect 24572 96406 24584 96458
rect 24320 96404 24376 96406
rect 24424 96404 24480 96406
rect 24528 96404 24584 96406
rect 24632 96458 24688 96460
rect 24736 96458 24792 96460
rect 24840 96458 24896 96460
rect 24632 96406 24644 96458
rect 24644 96406 24688 96458
rect 24736 96406 24768 96458
rect 24768 96406 24792 96458
rect 24840 96406 24892 96458
rect 24892 96406 24896 96458
rect 24632 96404 24688 96406
rect 24736 96404 24792 96406
rect 24840 96404 24896 96406
rect 24944 96404 25000 96460
rect 25048 96458 25104 96460
rect 25152 96458 25208 96460
rect 25048 96406 25068 96458
rect 25068 96406 25104 96458
rect 25152 96406 25192 96458
rect 25192 96406 25208 96458
rect 25048 96404 25104 96406
rect 25152 96404 25208 96406
rect 14008 95674 14064 95676
rect 14112 95674 14168 95676
rect 14008 95622 14024 95674
rect 14024 95622 14064 95674
rect 14112 95622 14148 95674
rect 14148 95622 14168 95674
rect 14008 95620 14064 95622
rect 14112 95620 14168 95622
rect 14216 95620 14272 95676
rect 14320 95674 14376 95676
rect 14424 95674 14480 95676
rect 14528 95674 14584 95676
rect 14320 95622 14324 95674
rect 14324 95622 14376 95674
rect 14424 95622 14448 95674
rect 14448 95622 14480 95674
rect 14528 95622 14572 95674
rect 14572 95622 14584 95674
rect 14320 95620 14376 95622
rect 14424 95620 14480 95622
rect 14528 95620 14584 95622
rect 14632 95674 14688 95676
rect 14736 95674 14792 95676
rect 14840 95674 14896 95676
rect 14632 95622 14644 95674
rect 14644 95622 14688 95674
rect 14736 95622 14768 95674
rect 14768 95622 14792 95674
rect 14840 95622 14892 95674
rect 14892 95622 14896 95674
rect 14632 95620 14688 95622
rect 14736 95620 14792 95622
rect 14840 95620 14896 95622
rect 14944 95620 15000 95676
rect 15048 95674 15104 95676
rect 15152 95674 15208 95676
rect 15048 95622 15068 95674
rect 15068 95622 15104 95674
rect 15152 95622 15192 95674
rect 15192 95622 15208 95674
rect 15048 95620 15104 95622
rect 15152 95620 15208 95622
rect 24008 94890 24064 94892
rect 24112 94890 24168 94892
rect 24008 94838 24024 94890
rect 24024 94838 24064 94890
rect 24112 94838 24148 94890
rect 24148 94838 24168 94890
rect 24008 94836 24064 94838
rect 24112 94836 24168 94838
rect 24216 94836 24272 94892
rect 24320 94890 24376 94892
rect 24424 94890 24480 94892
rect 24528 94890 24584 94892
rect 24320 94838 24324 94890
rect 24324 94838 24376 94890
rect 24424 94838 24448 94890
rect 24448 94838 24480 94890
rect 24528 94838 24572 94890
rect 24572 94838 24584 94890
rect 24320 94836 24376 94838
rect 24424 94836 24480 94838
rect 24528 94836 24584 94838
rect 24632 94890 24688 94892
rect 24736 94890 24792 94892
rect 24840 94890 24896 94892
rect 24632 94838 24644 94890
rect 24644 94838 24688 94890
rect 24736 94838 24768 94890
rect 24768 94838 24792 94890
rect 24840 94838 24892 94890
rect 24892 94838 24896 94890
rect 24632 94836 24688 94838
rect 24736 94836 24792 94838
rect 24840 94836 24896 94838
rect 24944 94836 25000 94892
rect 25048 94890 25104 94892
rect 25152 94890 25208 94892
rect 25048 94838 25068 94890
rect 25068 94838 25104 94890
rect 25152 94838 25192 94890
rect 25192 94838 25208 94890
rect 25048 94836 25104 94838
rect 25152 94836 25208 94838
rect 9884 94108 9940 94164
rect 12908 94108 12964 94164
rect 4008 93322 4064 93324
rect 4112 93322 4168 93324
rect 4008 93270 4024 93322
rect 4024 93270 4064 93322
rect 4112 93270 4148 93322
rect 4148 93270 4168 93322
rect 4008 93268 4064 93270
rect 4112 93268 4168 93270
rect 4216 93268 4272 93324
rect 4320 93322 4376 93324
rect 4424 93322 4480 93324
rect 4528 93322 4584 93324
rect 4320 93270 4324 93322
rect 4324 93270 4376 93322
rect 4424 93270 4448 93322
rect 4448 93270 4480 93322
rect 4528 93270 4572 93322
rect 4572 93270 4584 93322
rect 4320 93268 4376 93270
rect 4424 93268 4480 93270
rect 4528 93268 4584 93270
rect 4632 93322 4688 93324
rect 4736 93322 4792 93324
rect 4840 93322 4896 93324
rect 4632 93270 4644 93322
rect 4644 93270 4688 93322
rect 4736 93270 4768 93322
rect 4768 93270 4792 93322
rect 4840 93270 4892 93322
rect 4892 93270 4896 93322
rect 4632 93268 4688 93270
rect 4736 93268 4792 93270
rect 4840 93268 4896 93270
rect 4944 93268 5000 93324
rect 5048 93322 5104 93324
rect 5152 93322 5208 93324
rect 5048 93270 5068 93322
rect 5068 93270 5104 93322
rect 5152 93270 5192 93322
rect 5192 93270 5208 93322
rect 5048 93268 5104 93270
rect 5152 93268 5208 93270
rect 1708 92988 1764 93044
rect 1708 91868 1764 91924
rect 4008 91754 4064 91756
rect 4112 91754 4168 91756
rect 4008 91702 4024 91754
rect 4024 91702 4064 91754
rect 4112 91702 4148 91754
rect 4148 91702 4168 91754
rect 4008 91700 4064 91702
rect 4112 91700 4168 91702
rect 4216 91700 4272 91756
rect 4320 91754 4376 91756
rect 4424 91754 4480 91756
rect 4528 91754 4584 91756
rect 4320 91702 4324 91754
rect 4324 91702 4376 91754
rect 4424 91702 4448 91754
rect 4448 91702 4480 91754
rect 4528 91702 4572 91754
rect 4572 91702 4584 91754
rect 4320 91700 4376 91702
rect 4424 91700 4480 91702
rect 4528 91700 4584 91702
rect 4632 91754 4688 91756
rect 4736 91754 4792 91756
rect 4840 91754 4896 91756
rect 4632 91702 4644 91754
rect 4644 91702 4688 91754
rect 4736 91702 4768 91754
rect 4768 91702 4792 91754
rect 4840 91702 4892 91754
rect 4892 91702 4896 91754
rect 4632 91700 4688 91702
rect 4736 91700 4792 91702
rect 4840 91700 4896 91702
rect 4944 91700 5000 91756
rect 5048 91754 5104 91756
rect 5152 91754 5208 91756
rect 5048 91702 5068 91754
rect 5068 91702 5104 91754
rect 5152 91702 5192 91754
rect 5192 91702 5208 91754
rect 5048 91700 5104 91702
rect 5152 91700 5208 91702
rect 1708 90748 1764 90804
rect 4008 90186 4064 90188
rect 4112 90186 4168 90188
rect 4008 90134 4024 90186
rect 4024 90134 4064 90186
rect 4112 90134 4148 90186
rect 4148 90134 4168 90186
rect 4008 90132 4064 90134
rect 4112 90132 4168 90134
rect 4216 90132 4272 90188
rect 4320 90186 4376 90188
rect 4424 90186 4480 90188
rect 4528 90186 4584 90188
rect 4320 90134 4324 90186
rect 4324 90134 4376 90186
rect 4424 90134 4448 90186
rect 4448 90134 4480 90186
rect 4528 90134 4572 90186
rect 4572 90134 4584 90186
rect 4320 90132 4376 90134
rect 4424 90132 4480 90134
rect 4528 90132 4584 90134
rect 4632 90186 4688 90188
rect 4736 90186 4792 90188
rect 4840 90186 4896 90188
rect 4632 90134 4644 90186
rect 4644 90134 4688 90186
rect 4736 90134 4768 90186
rect 4768 90134 4792 90186
rect 4840 90134 4892 90186
rect 4892 90134 4896 90186
rect 4632 90132 4688 90134
rect 4736 90132 4792 90134
rect 4840 90132 4896 90134
rect 4944 90132 5000 90188
rect 5048 90186 5104 90188
rect 5152 90186 5208 90188
rect 5048 90134 5068 90186
rect 5068 90134 5104 90186
rect 5152 90134 5192 90186
rect 5192 90134 5208 90186
rect 5048 90132 5104 90134
rect 5152 90132 5208 90134
rect 1708 89682 1764 89684
rect 1708 89630 1710 89682
rect 1710 89630 1762 89682
rect 1762 89630 1764 89682
rect 1708 89628 1764 89630
rect 1708 88508 1764 88564
rect 4008 88618 4064 88620
rect 4112 88618 4168 88620
rect 4008 88566 4024 88618
rect 4024 88566 4064 88618
rect 4112 88566 4148 88618
rect 4148 88566 4168 88618
rect 4008 88564 4064 88566
rect 4112 88564 4168 88566
rect 4216 88564 4272 88620
rect 4320 88618 4376 88620
rect 4424 88618 4480 88620
rect 4528 88618 4584 88620
rect 4320 88566 4324 88618
rect 4324 88566 4376 88618
rect 4424 88566 4448 88618
rect 4448 88566 4480 88618
rect 4528 88566 4572 88618
rect 4572 88566 4584 88618
rect 4320 88564 4376 88566
rect 4424 88564 4480 88566
rect 4528 88564 4584 88566
rect 4632 88618 4688 88620
rect 4736 88618 4792 88620
rect 4840 88618 4896 88620
rect 4632 88566 4644 88618
rect 4644 88566 4688 88618
rect 4736 88566 4768 88618
rect 4768 88566 4792 88618
rect 4840 88566 4892 88618
rect 4892 88566 4896 88618
rect 4632 88564 4688 88566
rect 4736 88564 4792 88566
rect 4840 88564 4896 88566
rect 4944 88564 5000 88620
rect 5048 88618 5104 88620
rect 5152 88618 5208 88620
rect 5048 88566 5068 88618
rect 5068 88566 5104 88618
rect 5152 88566 5192 88618
rect 5192 88566 5208 88618
rect 5048 88564 5104 88566
rect 5152 88564 5208 88566
rect 8428 88002 8484 88004
rect 8428 87950 8430 88002
rect 8430 87950 8482 88002
rect 8482 87950 8484 88002
rect 8428 87948 8484 87950
rect 9772 88226 9828 88228
rect 9772 88174 9774 88226
rect 9774 88174 9826 88226
rect 9826 88174 9828 88226
rect 9772 88172 9828 88174
rect 1708 87388 1764 87444
rect 5628 87442 5684 87444
rect 5628 87390 5630 87442
rect 5630 87390 5682 87442
rect 5682 87390 5684 87442
rect 5628 87388 5684 87390
rect 4008 87050 4064 87052
rect 4112 87050 4168 87052
rect 4008 86998 4024 87050
rect 4024 86998 4064 87050
rect 4112 86998 4148 87050
rect 4148 86998 4168 87050
rect 4008 86996 4064 86998
rect 4112 86996 4168 86998
rect 4216 86996 4272 87052
rect 4320 87050 4376 87052
rect 4424 87050 4480 87052
rect 4528 87050 4584 87052
rect 4320 86998 4324 87050
rect 4324 86998 4376 87050
rect 4424 86998 4448 87050
rect 4448 86998 4480 87050
rect 4528 86998 4572 87050
rect 4572 86998 4584 87050
rect 4320 86996 4376 86998
rect 4424 86996 4480 86998
rect 4528 86996 4584 86998
rect 4632 87050 4688 87052
rect 4736 87050 4792 87052
rect 4840 87050 4896 87052
rect 4632 86998 4644 87050
rect 4644 86998 4688 87050
rect 4736 86998 4768 87050
rect 4768 86998 4792 87050
rect 4840 86998 4892 87050
rect 4892 86998 4896 87050
rect 4632 86996 4688 86998
rect 4736 86996 4792 86998
rect 4840 86996 4896 86998
rect 4944 86996 5000 87052
rect 5048 87050 5104 87052
rect 5152 87050 5208 87052
rect 5048 86998 5068 87050
rect 5068 86998 5104 87050
rect 5152 86998 5192 87050
rect 5192 86998 5208 87050
rect 5048 86996 5104 86998
rect 5152 86996 5208 86998
rect 6076 86828 6132 86884
rect 6524 87388 6580 87444
rect 1708 86434 1764 86436
rect 1708 86382 1710 86434
rect 1710 86382 1762 86434
rect 1762 86382 1764 86434
rect 1708 86380 1764 86382
rect 4008 85482 4064 85484
rect 4112 85482 4168 85484
rect 4008 85430 4024 85482
rect 4024 85430 4064 85482
rect 4112 85430 4148 85482
rect 4148 85430 4168 85482
rect 4008 85428 4064 85430
rect 4112 85428 4168 85430
rect 4216 85428 4272 85484
rect 4320 85482 4376 85484
rect 4424 85482 4480 85484
rect 4528 85482 4584 85484
rect 4320 85430 4324 85482
rect 4324 85430 4376 85482
rect 4424 85430 4448 85482
rect 4448 85430 4480 85482
rect 4528 85430 4572 85482
rect 4572 85430 4584 85482
rect 4320 85428 4376 85430
rect 4424 85428 4480 85430
rect 4528 85428 4584 85430
rect 4632 85482 4688 85484
rect 4736 85482 4792 85484
rect 4840 85482 4896 85484
rect 4632 85430 4644 85482
rect 4644 85430 4688 85482
rect 4736 85430 4768 85482
rect 4768 85430 4792 85482
rect 4840 85430 4892 85482
rect 4892 85430 4896 85482
rect 4632 85428 4688 85430
rect 4736 85428 4792 85430
rect 4840 85428 4896 85430
rect 4944 85428 5000 85484
rect 5048 85482 5104 85484
rect 5152 85482 5208 85484
rect 5048 85430 5068 85482
rect 5068 85430 5104 85482
rect 5152 85430 5192 85482
rect 5192 85430 5208 85482
rect 5048 85428 5104 85430
rect 5152 85428 5208 85430
rect 1708 85148 1764 85204
rect 4844 85202 4900 85204
rect 4844 85150 4846 85202
rect 4846 85150 4898 85202
rect 4898 85150 4900 85202
rect 4844 85148 4900 85150
rect 5404 85148 5460 85204
rect 3836 85036 3892 85092
rect 1708 84028 1764 84084
rect 4008 83914 4064 83916
rect 4112 83914 4168 83916
rect 4008 83862 4024 83914
rect 4024 83862 4064 83914
rect 4112 83862 4148 83914
rect 4148 83862 4168 83914
rect 4008 83860 4064 83862
rect 4112 83860 4168 83862
rect 4216 83860 4272 83916
rect 4320 83914 4376 83916
rect 4424 83914 4480 83916
rect 4528 83914 4584 83916
rect 4320 83862 4324 83914
rect 4324 83862 4376 83914
rect 4424 83862 4448 83914
rect 4448 83862 4480 83914
rect 4528 83862 4572 83914
rect 4572 83862 4584 83914
rect 4320 83860 4376 83862
rect 4424 83860 4480 83862
rect 4528 83860 4584 83862
rect 4632 83914 4688 83916
rect 4736 83914 4792 83916
rect 4840 83914 4896 83916
rect 4632 83862 4644 83914
rect 4644 83862 4688 83914
rect 4736 83862 4768 83914
rect 4768 83862 4792 83914
rect 4840 83862 4892 83914
rect 4892 83862 4896 83914
rect 4632 83860 4688 83862
rect 4736 83860 4792 83862
rect 4840 83860 4896 83862
rect 4944 83860 5000 83916
rect 5048 83914 5104 83916
rect 5152 83914 5208 83916
rect 5048 83862 5068 83914
rect 5068 83862 5104 83914
rect 5152 83862 5192 83914
rect 5192 83862 5208 83914
rect 5048 83860 5104 83862
rect 5152 83860 5208 83862
rect 3836 83692 3892 83748
rect 1708 82908 1764 82964
rect 2268 83244 2324 83300
rect 1708 81842 1764 81844
rect 1708 81790 1710 81842
rect 1710 81790 1762 81842
rect 1762 81790 1764 81842
rect 1708 81788 1764 81790
rect 1708 80668 1764 80724
rect 3388 83298 3444 83300
rect 3388 83246 3390 83298
rect 3390 83246 3442 83298
rect 3442 83246 3444 83298
rect 3388 83244 3444 83246
rect 4284 83522 4340 83524
rect 4284 83470 4286 83522
rect 4286 83470 4338 83522
rect 4338 83470 4340 83522
rect 4284 83468 4340 83470
rect 3612 82012 3668 82068
rect 1820 80556 1876 80612
rect 1708 79548 1764 79604
rect 1708 78594 1764 78596
rect 1708 78542 1710 78594
rect 1710 78542 1762 78594
rect 1762 78542 1764 78594
rect 1708 78540 1764 78542
rect 3388 78930 3444 78932
rect 3388 78878 3390 78930
rect 3390 78878 3442 78930
rect 3442 78878 3444 78930
rect 3388 78876 3444 78878
rect 3612 77756 3668 77812
rect 1708 77308 1764 77364
rect 9884 87666 9940 87668
rect 9884 87614 9886 87666
rect 9886 87614 9938 87666
rect 9938 87614 9940 87666
rect 9884 87612 9940 87614
rect 8876 87388 8932 87444
rect 7644 86882 7700 86884
rect 7644 86830 7646 86882
rect 7646 86830 7698 86882
rect 7698 86830 7700 86882
rect 7644 86828 7700 86830
rect 7308 86546 7364 86548
rect 7308 86494 7310 86546
rect 7310 86494 7362 86546
rect 7362 86494 7364 86546
rect 7308 86492 7364 86494
rect 8764 86658 8820 86660
rect 8764 86606 8766 86658
rect 8766 86606 8818 86658
rect 8818 86606 8820 86658
rect 8764 86604 8820 86606
rect 7980 86380 8036 86436
rect 8540 86546 8596 86548
rect 8540 86494 8542 86546
rect 8542 86494 8594 86546
rect 8594 86494 8596 86546
rect 8540 86492 8596 86494
rect 8540 86156 8596 86212
rect 12348 88844 12404 88900
rect 10332 88172 10388 88228
rect 10444 87948 10500 88004
rect 9324 86658 9380 86660
rect 9324 86606 9326 86658
rect 9326 86606 9378 86658
rect 9378 86606 9380 86658
rect 9324 86604 9380 86606
rect 9884 86658 9940 86660
rect 9884 86606 9886 86658
rect 9886 86606 9938 86658
rect 9938 86606 9940 86658
rect 9884 86604 9940 86606
rect 9100 86380 9156 86436
rect 9660 86098 9716 86100
rect 9660 86046 9662 86098
rect 9662 86046 9714 86098
rect 9714 86046 9716 86098
rect 9660 86044 9716 86046
rect 10220 86546 10276 86548
rect 10220 86494 10222 86546
rect 10222 86494 10274 86546
rect 10274 86494 10276 86546
rect 10220 86492 10276 86494
rect 10220 86098 10276 86100
rect 10220 86046 10222 86098
rect 10222 86046 10274 86098
rect 10274 86046 10276 86098
rect 10220 86044 10276 86046
rect 6524 85090 6580 85092
rect 6524 85038 6526 85090
rect 6526 85038 6578 85090
rect 6578 85038 6580 85090
rect 6524 85036 6580 85038
rect 6748 84924 6804 84980
rect 6972 84476 7028 84532
rect 7196 85036 7252 85092
rect 5852 84028 5908 84084
rect 6860 84028 6916 84084
rect 5964 83746 6020 83748
rect 5964 83694 5966 83746
rect 5966 83694 6018 83746
rect 6018 83694 6020 83746
rect 5964 83692 6020 83694
rect 6300 83746 6356 83748
rect 6300 83694 6302 83746
rect 6302 83694 6354 83746
rect 6354 83694 6356 83746
rect 6300 83692 6356 83694
rect 5404 83468 5460 83524
rect 5628 83580 5684 83636
rect 4508 83410 4564 83412
rect 4508 83358 4510 83410
rect 4510 83358 4562 83410
rect 4562 83358 4564 83410
rect 4508 83356 4564 83358
rect 5292 83356 5348 83412
rect 4732 82796 4788 82852
rect 7084 83244 7140 83300
rect 5068 82796 5124 82852
rect 6300 82572 6356 82628
rect 4008 82346 4064 82348
rect 4112 82346 4168 82348
rect 4008 82294 4024 82346
rect 4024 82294 4064 82346
rect 4112 82294 4148 82346
rect 4148 82294 4168 82346
rect 4008 82292 4064 82294
rect 4112 82292 4168 82294
rect 4216 82292 4272 82348
rect 4320 82346 4376 82348
rect 4424 82346 4480 82348
rect 4528 82346 4584 82348
rect 4320 82294 4324 82346
rect 4324 82294 4376 82346
rect 4424 82294 4448 82346
rect 4448 82294 4480 82346
rect 4528 82294 4572 82346
rect 4572 82294 4584 82346
rect 4320 82292 4376 82294
rect 4424 82292 4480 82294
rect 4528 82292 4584 82294
rect 4632 82346 4688 82348
rect 4736 82346 4792 82348
rect 4840 82346 4896 82348
rect 4632 82294 4644 82346
rect 4644 82294 4688 82346
rect 4736 82294 4768 82346
rect 4768 82294 4792 82346
rect 4840 82294 4892 82346
rect 4892 82294 4896 82346
rect 4632 82292 4688 82294
rect 4736 82292 4792 82294
rect 4840 82292 4896 82294
rect 4944 82292 5000 82348
rect 5048 82346 5104 82348
rect 5152 82346 5208 82348
rect 5048 82294 5068 82346
rect 5068 82294 5104 82346
rect 5152 82294 5192 82346
rect 5192 82294 5208 82346
rect 5048 82292 5104 82294
rect 5152 82292 5208 82294
rect 4844 82124 4900 82180
rect 4508 82066 4564 82068
rect 4508 82014 4510 82066
rect 4510 82014 4562 82066
rect 4562 82014 4564 82066
rect 4508 82012 4564 82014
rect 4396 81730 4452 81732
rect 4396 81678 4398 81730
rect 4398 81678 4450 81730
rect 4450 81678 4452 81730
rect 4396 81676 4452 81678
rect 4620 81004 4676 81060
rect 5180 81676 5236 81732
rect 4008 80778 4064 80780
rect 4112 80778 4168 80780
rect 4008 80726 4024 80778
rect 4024 80726 4064 80778
rect 4112 80726 4148 80778
rect 4148 80726 4168 80778
rect 4008 80724 4064 80726
rect 4112 80724 4168 80726
rect 4216 80724 4272 80780
rect 4320 80778 4376 80780
rect 4424 80778 4480 80780
rect 4528 80778 4584 80780
rect 4320 80726 4324 80778
rect 4324 80726 4376 80778
rect 4424 80726 4448 80778
rect 4448 80726 4480 80778
rect 4528 80726 4572 80778
rect 4572 80726 4584 80778
rect 4320 80724 4376 80726
rect 4424 80724 4480 80726
rect 4528 80724 4584 80726
rect 4632 80778 4688 80780
rect 4736 80778 4792 80780
rect 4840 80778 4896 80780
rect 4632 80726 4644 80778
rect 4644 80726 4688 80778
rect 4736 80726 4768 80778
rect 4768 80726 4792 80778
rect 4840 80726 4892 80778
rect 4892 80726 4896 80778
rect 4632 80724 4688 80726
rect 4736 80724 4792 80726
rect 4840 80724 4896 80726
rect 4944 80724 5000 80780
rect 5048 80778 5104 80780
rect 5152 80778 5208 80780
rect 5048 80726 5068 80778
rect 5068 80726 5104 80778
rect 5152 80726 5192 80778
rect 5192 80726 5208 80778
rect 5048 80724 5104 80726
rect 5152 80724 5208 80726
rect 4732 79826 4788 79828
rect 4732 79774 4734 79826
rect 4734 79774 4786 79826
rect 4786 79774 4788 79826
rect 4732 79772 4788 79774
rect 4008 79210 4064 79212
rect 4112 79210 4168 79212
rect 4008 79158 4024 79210
rect 4024 79158 4064 79210
rect 4112 79158 4148 79210
rect 4148 79158 4168 79210
rect 4008 79156 4064 79158
rect 4112 79156 4168 79158
rect 4216 79156 4272 79212
rect 4320 79210 4376 79212
rect 4424 79210 4480 79212
rect 4528 79210 4584 79212
rect 4320 79158 4324 79210
rect 4324 79158 4376 79210
rect 4424 79158 4448 79210
rect 4448 79158 4480 79210
rect 4528 79158 4572 79210
rect 4572 79158 4584 79210
rect 4320 79156 4376 79158
rect 4424 79156 4480 79158
rect 4528 79156 4584 79158
rect 4632 79210 4688 79212
rect 4736 79210 4792 79212
rect 4840 79210 4896 79212
rect 4632 79158 4644 79210
rect 4644 79158 4688 79210
rect 4736 79158 4768 79210
rect 4768 79158 4792 79210
rect 4840 79158 4892 79210
rect 4892 79158 4896 79210
rect 4632 79156 4688 79158
rect 4736 79156 4792 79158
rect 4840 79156 4896 79158
rect 4944 79156 5000 79212
rect 5048 79210 5104 79212
rect 5152 79210 5208 79212
rect 5048 79158 5068 79210
rect 5068 79158 5104 79210
rect 5152 79158 5192 79210
rect 5192 79158 5208 79210
rect 5048 79156 5104 79158
rect 5152 79156 5208 79158
rect 4508 78930 4564 78932
rect 4508 78878 4510 78930
rect 4510 78878 4562 78930
rect 4562 78878 4564 78930
rect 4508 78876 4564 78878
rect 5516 80892 5572 80948
rect 5852 82236 5908 82292
rect 6188 82348 6244 82404
rect 6412 82460 6468 82516
rect 5628 80556 5684 80612
rect 6300 82236 6356 82292
rect 5964 80892 6020 80948
rect 6076 80386 6132 80388
rect 6076 80334 6078 80386
rect 6078 80334 6130 80386
rect 6130 80334 6132 80386
rect 6076 80332 6132 80334
rect 5404 79324 5460 79380
rect 5404 78876 5460 78932
rect 6636 82572 6692 82628
rect 8316 84530 8372 84532
rect 8316 84478 8318 84530
rect 8318 84478 8370 84530
rect 8370 84478 8372 84530
rect 8316 84476 8372 84478
rect 7308 83692 7364 83748
rect 8204 83410 8260 83412
rect 8204 83358 8206 83410
rect 8206 83358 8258 83410
rect 8258 83358 8260 83410
rect 8204 83356 8260 83358
rect 12012 88002 12068 88004
rect 12012 87950 12014 88002
rect 12014 87950 12066 88002
rect 12066 87950 12068 88002
rect 12012 87948 12068 87950
rect 12572 87948 12628 88004
rect 11452 87612 11508 87668
rect 10668 87218 10724 87220
rect 10668 87166 10670 87218
rect 10670 87166 10722 87218
rect 10722 87166 10724 87218
rect 10668 87164 10724 87166
rect 10892 86658 10948 86660
rect 10892 86606 10894 86658
rect 10894 86606 10946 86658
rect 10946 86606 10948 86658
rect 10892 86604 10948 86606
rect 11004 86492 11060 86548
rect 9212 84978 9268 84980
rect 9212 84926 9214 84978
rect 9214 84926 9266 84978
rect 9266 84926 9268 84978
rect 9212 84924 9268 84926
rect 10444 84924 10500 84980
rect 7644 83298 7700 83300
rect 7644 83246 7646 83298
rect 7646 83246 7698 83298
rect 7698 83246 7700 83298
rect 7644 83244 7700 83246
rect 8428 83244 8484 83300
rect 8764 83356 8820 83412
rect 8204 82796 8260 82852
rect 7644 82348 7700 82404
rect 6636 81676 6692 81732
rect 9212 83298 9268 83300
rect 9212 83246 9214 83298
rect 9214 83246 9266 83298
rect 9266 83246 9268 83298
rect 9212 83244 9268 83246
rect 8764 82460 8820 82516
rect 4620 78818 4676 78820
rect 4620 78766 4622 78818
rect 4622 78766 4674 78818
rect 4674 78766 4676 78818
rect 4620 78764 4676 78766
rect 5852 78764 5908 78820
rect 4172 78594 4228 78596
rect 4172 78542 4174 78594
rect 4174 78542 4226 78594
rect 4226 78542 4228 78594
rect 4172 78540 4228 78542
rect 4508 78316 4564 78372
rect 4732 78258 4788 78260
rect 4732 78206 4734 78258
rect 4734 78206 4786 78258
rect 4786 78206 4788 78258
rect 4732 78204 4788 78206
rect 4844 77868 4900 77924
rect 5292 78316 5348 78372
rect 4008 77642 4064 77644
rect 4112 77642 4168 77644
rect 4008 77590 4024 77642
rect 4024 77590 4064 77642
rect 4112 77590 4148 77642
rect 4148 77590 4168 77642
rect 4008 77588 4064 77590
rect 4112 77588 4168 77590
rect 4216 77588 4272 77644
rect 4320 77642 4376 77644
rect 4424 77642 4480 77644
rect 4528 77642 4584 77644
rect 4320 77590 4324 77642
rect 4324 77590 4376 77642
rect 4424 77590 4448 77642
rect 4448 77590 4480 77642
rect 4528 77590 4572 77642
rect 4572 77590 4584 77642
rect 4320 77588 4376 77590
rect 4424 77588 4480 77590
rect 4528 77588 4584 77590
rect 4632 77642 4688 77644
rect 4736 77642 4792 77644
rect 4840 77642 4896 77644
rect 4632 77590 4644 77642
rect 4644 77590 4688 77642
rect 4736 77590 4768 77642
rect 4768 77590 4792 77642
rect 4840 77590 4892 77642
rect 4892 77590 4896 77642
rect 4632 77588 4688 77590
rect 4736 77588 4792 77590
rect 4840 77588 4896 77590
rect 4944 77588 5000 77644
rect 5048 77642 5104 77644
rect 5152 77642 5208 77644
rect 5048 77590 5068 77642
rect 5068 77590 5104 77642
rect 5152 77590 5192 77642
rect 5192 77590 5208 77642
rect 5048 77588 5104 77590
rect 5152 77588 5208 77590
rect 4284 77420 4340 77476
rect 5292 77420 5348 77476
rect 5404 78204 5460 78260
rect 5068 77250 5124 77252
rect 5068 77198 5070 77250
rect 5070 77198 5122 77250
rect 5122 77198 5124 77250
rect 5068 77196 5124 77198
rect 3836 76636 3892 76692
rect 4732 76690 4788 76692
rect 4732 76638 4734 76690
rect 4734 76638 4786 76690
rect 4786 76638 4788 76690
rect 4732 76636 4788 76638
rect 5628 77810 5684 77812
rect 5628 77758 5630 77810
rect 5630 77758 5682 77810
rect 5682 77758 5684 77810
rect 5628 77756 5684 77758
rect 6076 79324 6132 79380
rect 6300 78988 6356 79044
rect 7308 80386 7364 80388
rect 7308 80334 7310 80386
rect 7310 80334 7362 80386
rect 7362 80334 7364 80386
rect 7308 80332 7364 80334
rect 6748 80220 6804 80276
rect 8204 80220 8260 80276
rect 6748 79826 6804 79828
rect 6748 79774 6750 79826
rect 6750 79774 6802 79826
rect 6802 79774 6804 79826
rect 6748 79772 6804 79774
rect 7420 80108 7476 80164
rect 8092 80162 8148 80164
rect 8092 80110 8094 80162
rect 8094 80110 8146 80162
rect 8146 80110 8148 80162
rect 8092 80108 8148 80110
rect 6524 79324 6580 79380
rect 5964 78540 6020 78596
rect 1708 76188 1764 76244
rect 5852 77980 5908 78036
rect 7980 79378 8036 79380
rect 7980 79326 7982 79378
rect 7982 79326 8034 79378
rect 8034 79326 8036 79378
rect 7980 79324 8036 79326
rect 6748 78988 6804 79044
rect 6076 77868 6132 77924
rect 6188 78540 6244 78596
rect 5964 77308 6020 77364
rect 6076 77644 6132 77700
rect 5740 76300 5796 76356
rect 4008 76074 4064 76076
rect 4112 76074 4168 76076
rect 4008 76022 4024 76074
rect 4024 76022 4064 76074
rect 4112 76022 4148 76074
rect 4148 76022 4168 76074
rect 4008 76020 4064 76022
rect 4112 76020 4168 76022
rect 4216 76020 4272 76076
rect 4320 76074 4376 76076
rect 4424 76074 4480 76076
rect 4528 76074 4584 76076
rect 4320 76022 4324 76074
rect 4324 76022 4376 76074
rect 4424 76022 4448 76074
rect 4448 76022 4480 76074
rect 4528 76022 4572 76074
rect 4572 76022 4584 76074
rect 4320 76020 4376 76022
rect 4424 76020 4480 76022
rect 4528 76020 4584 76022
rect 4632 76074 4688 76076
rect 4736 76074 4792 76076
rect 4840 76074 4896 76076
rect 4632 76022 4644 76074
rect 4644 76022 4688 76074
rect 4736 76022 4768 76074
rect 4768 76022 4792 76074
rect 4840 76022 4892 76074
rect 4892 76022 4896 76074
rect 4632 76020 4688 76022
rect 4736 76020 4792 76022
rect 4840 76020 4896 76022
rect 4944 76020 5000 76076
rect 5048 76074 5104 76076
rect 5152 76074 5208 76076
rect 5048 76022 5068 76074
rect 5068 76022 5104 76074
rect 5152 76022 5192 76074
rect 5192 76022 5208 76074
rect 5048 76020 5104 76022
rect 5152 76020 5208 76022
rect 4396 75794 4452 75796
rect 4396 75742 4398 75794
rect 4398 75742 4450 75794
rect 4450 75742 4452 75794
rect 4396 75740 4452 75742
rect 1708 75068 1764 75124
rect 1820 74172 1876 74228
rect 4008 74506 4064 74508
rect 4112 74506 4168 74508
rect 4008 74454 4024 74506
rect 4024 74454 4064 74506
rect 4112 74454 4148 74506
rect 4148 74454 4168 74506
rect 4008 74452 4064 74454
rect 4112 74452 4168 74454
rect 4216 74452 4272 74508
rect 4320 74506 4376 74508
rect 4424 74506 4480 74508
rect 4528 74506 4584 74508
rect 4320 74454 4324 74506
rect 4324 74454 4376 74506
rect 4424 74454 4448 74506
rect 4448 74454 4480 74506
rect 4528 74454 4572 74506
rect 4572 74454 4584 74506
rect 4320 74452 4376 74454
rect 4424 74452 4480 74454
rect 4528 74452 4584 74454
rect 4632 74506 4688 74508
rect 4736 74506 4792 74508
rect 4840 74506 4896 74508
rect 4632 74454 4644 74506
rect 4644 74454 4688 74506
rect 4736 74454 4768 74506
rect 4768 74454 4792 74506
rect 4840 74454 4892 74506
rect 4892 74454 4896 74506
rect 4632 74452 4688 74454
rect 4736 74452 4792 74454
rect 4840 74452 4896 74454
rect 4944 74452 5000 74508
rect 5048 74506 5104 74508
rect 5152 74506 5208 74508
rect 5048 74454 5068 74506
rect 5068 74454 5104 74506
rect 5152 74454 5192 74506
rect 5192 74454 5208 74506
rect 5048 74452 5104 74454
rect 5152 74452 5208 74454
rect 3164 74172 3220 74228
rect 4060 74284 4116 74340
rect 2156 73948 2212 74004
rect 2492 73948 2548 74004
rect 3500 74002 3556 74004
rect 3500 73950 3502 74002
rect 3502 73950 3554 74002
rect 3554 73950 3556 74002
rect 3500 73948 3556 73950
rect 1708 72828 1764 72884
rect 4060 74060 4116 74116
rect 4620 74002 4676 74004
rect 4620 73950 4622 74002
rect 4622 73950 4674 74002
rect 4674 73950 4676 74002
rect 4620 73948 4676 73950
rect 5852 75794 5908 75796
rect 5852 75742 5854 75794
rect 5854 75742 5906 75794
rect 5906 75742 5908 75794
rect 5852 75740 5908 75742
rect 5292 73948 5348 74004
rect 5740 74226 5796 74228
rect 5740 74174 5742 74226
rect 5742 74174 5794 74226
rect 5794 74174 5796 74226
rect 5740 74172 5796 74174
rect 4732 73836 4788 73892
rect 4008 72938 4064 72940
rect 4112 72938 4168 72940
rect 4008 72886 4024 72938
rect 4024 72886 4064 72938
rect 4112 72886 4148 72938
rect 4148 72886 4168 72938
rect 4008 72884 4064 72886
rect 4112 72884 4168 72886
rect 4216 72884 4272 72940
rect 4320 72938 4376 72940
rect 4424 72938 4480 72940
rect 4528 72938 4584 72940
rect 4320 72886 4324 72938
rect 4324 72886 4376 72938
rect 4424 72886 4448 72938
rect 4448 72886 4480 72938
rect 4528 72886 4572 72938
rect 4572 72886 4584 72938
rect 4320 72884 4376 72886
rect 4424 72884 4480 72886
rect 4528 72884 4584 72886
rect 4632 72938 4688 72940
rect 4736 72938 4792 72940
rect 4840 72938 4896 72940
rect 4632 72886 4644 72938
rect 4644 72886 4688 72938
rect 4736 72886 4768 72938
rect 4768 72886 4792 72938
rect 4840 72886 4892 72938
rect 4892 72886 4896 72938
rect 4632 72884 4688 72886
rect 4736 72884 4792 72886
rect 4840 72884 4896 72886
rect 4944 72884 5000 72940
rect 5048 72938 5104 72940
rect 5152 72938 5208 72940
rect 5048 72886 5068 72938
rect 5068 72886 5104 72938
rect 5152 72886 5192 72938
rect 5192 72886 5208 72938
rect 5048 72884 5104 72886
rect 5152 72884 5208 72886
rect 4956 72716 5012 72772
rect 3164 72492 3220 72548
rect 1708 71708 1764 71764
rect 1708 70754 1764 70756
rect 1708 70702 1710 70754
rect 1710 70702 1762 70754
rect 1762 70702 1764 70754
rect 1708 70700 1764 70702
rect 4172 72546 4228 72548
rect 4172 72494 4174 72546
rect 4174 72494 4226 72546
rect 4226 72494 4228 72546
rect 4172 72492 4228 72494
rect 4732 72380 4788 72436
rect 5292 72380 5348 72436
rect 4008 71370 4064 71372
rect 4112 71370 4168 71372
rect 4008 71318 4024 71370
rect 4024 71318 4064 71370
rect 4112 71318 4148 71370
rect 4148 71318 4168 71370
rect 4008 71316 4064 71318
rect 4112 71316 4168 71318
rect 4216 71316 4272 71372
rect 4320 71370 4376 71372
rect 4424 71370 4480 71372
rect 4528 71370 4584 71372
rect 4320 71318 4324 71370
rect 4324 71318 4376 71370
rect 4424 71318 4448 71370
rect 4448 71318 4480 71370
rect 4528 71318 4572 71370
rect 4572 71318 4584 71370
rect 4320 71316 4376 71318
rect 4424 71316 4480 71318
rect 4528 71316 4584 71318
rect 4632 71370 4688 71372
rect 4736 71370 4792 71372
rect 4840 71370 4896 71372
rect 4632 71318 4644 71370
rect 4644 71318 4688 71370
rect 4736 71318 4768 71370
rect 4768 71318 4792 71370
rect 4840 71318 4892 71370
rect 4892 71318 4896 71370
rect 4632 71316 4688 71318
rect 4736 71316 4792 71318
rect 4840 71316 4896 71318
rect 4944 71316 5000 71372
rect 5048 71370 5104 71372
rect 5152 71370 5208 71372
rect 5048 71318 5068 71370
rect 5068 71318 5104 71370
rect 5152 71318 5192 71370
rect 5192 71318 5208 71370
rect 5048 71316 5104 71318
rect 5152 71316 5208 71318
rect 1708 69468 1764 69524
rect 1708 68348 1764 68404
rect 1708 67228 1764 67284
rect 4008 69802 4064 69804
rect 4112 69802 4168 69804
rect 4008 69750 4024 69802
rect 4024 69750 4064 69802
rect 4112 69750 4148 69802
rect 4148 69750 4168 69802
rect 4008 69748 4064 69750
rect 4112 69748 4168 69750
rect 4216 69748 4272 69804
rect 4320 69802 4376 69804
rect 4424 69802 4480 69804
rect 4528 69802 4584 69804
rect 4320 69750 4324 69802
rect 4324 69750 4376 69802
rect 4424 69750 4448 69802
rect 4448 69750 4480 69802
rect 4528 69750 4572 69802
rect 4572 69750 4584 69802
rect 4320 69748 4376 69750
rect 4424 69748 4480 69750
rect 4528 69748 4584 69750
rect 4632 69802 4688 69804
rect 4736 69802 4792 69804
rect 4840 69802 4896 69804
rect 4632 69750 4644 69802
rect 4644 69750 4688 69802
rect 4736 69750 4768 69802
rect 4768 69750 4792 69802
rect 4840 69750 4892 69802
rect 4892 69750 4896 69802
rect 4632 69748 4688 69750
rect 4736 69748 4792 69750
rect 4840 69748 4896 69750
rect 4944 69748 5000 69804
rect 5048 69802 5104 69804
rect 5152 69802 5208 69804
rect 5048 69750 5068 69802
rect 5068 69750 5104 69802
rect 5152 69750 5192 69802
rect 5192 69750 5208 69802
rect 5048 69748 5104 69750
rect 5152 69748 5208 69750
rect 3052 67842 3108 67844
rect 3052 67790 3054 67842
rect 3054 67790 3106 67842
rect 3106 67790 3108 67842
rect 3052 67788 3108 67790
rect 1932 65212 1988 65268
rect 1708 64988 1764 65044
rect 1708 63868 1764 63924
rect 1708 62914 1764 62916
rect 1708 62862 1710 62914
rect 1710 62862 1762 62914
rect 1762 62862 1764 62914
rect 1708 62860 1764 62862
rect 1708 61628 1764 61684
rect 1708 60508 1764 60564
rect 1708 59388 1764 59444
rect 2268 66780 2324 66836
rect 2156 66162 2212 66164
rect 2156 66110 2158 66162
rect 2158 66110 2210 66162
rect 2210 66110 2212 66162
rect 2156 66108 2212 66110
rect 2380 63308 2436 63364
rect 1820 55356 1876 55412
rect 2044 52668 2100 52724
rect 1932 51548 1988 51604
rect 2268 61292 2324 61348
rect 2492 58322 2548 58324
rect 2492 58270 2494 58322
rect 2494 58270 2546 58322
rect 2546 58270 2548 58322
rect 2492 58268 2548 58270
rect 2940 58268 2996 58324
rect 2604 57148 2660 57204
rect 2268 56588 2324 56644
rect 2380 56082 2436 56084
rect 2380 56030 2382 56082
rect 2382 56030 2434 56082
rect 2434 56030 2436 56082
rect 2380 56028 2436 56030
rect 2828 56082 2884 56084
rect 2828 56030 2830 56082
rect 2830 56030 2882 56082
rect 2882 56030 2884 56082
rect 2828 56028 2884 56030
rect 3500 66892 3556 66948
rect 3388 66834 3444 66836
rect 3388 66782 3390 66834
rect 3390 66782 3442 66834
rect 3442 66782 3444 66834
rect 3388 66780 3444 66782
rect 4008 68234 4064 68236
rect 4112 68234 4168 68236
rect 4008 68182 4024 68234
rect 4024 68182 4064 68234
rect 4112 68182 4148 68234
rect 4148 68182 4168 68234
rect 4008 68180 4064 68182
rect 4112 68180 4168 68182
rect 4216 68180 4272 68236
rect 4320 68234 4376 68236
rect 4424 68234 4480 68236
rect 4528 68234 4584 68236
rect 4320 68182 4324 68234
rect 4324 68182 4376 68234
rect 4424 68182 4448 68234
rect 4448 68182 4480 68234
rect 4528 68182 4572 68234
rect 4572 68182 4584 68234
rect 4320 68180 4376 68182
rect 4424 68180 4480 68182
rect 4528 68180 4584 68182
rect 4632 68234 4688 68236
rect 4736 68234 4792 68236
rect 4840 68234 4896 68236
rect 4632 68182 4644 68234
rect 4644 68182 4688 68234
rect 4736 68182 4768 68234
rect 4768 68182 4792 68234
rect 4840 68182 4892 68234
rect 4892 68182 4896 68234
rect 4632 68180 4688 68182
rect 4736 68180 4792 68182
rect 4840 68180 4896 68182
rect 4944 68180 5000 68236
rect 5048 68234 5104 68236
rect 5152 68234 5208 68236
rect 5048 68182 5068 68234
rect 5068 68182 5104 68234
rect 5152 68182 5192 68234
rect 5192 68182 5208 68234
rect 5048 68180 5104 68182
rect 5152 68180 5208 68182
rect 4172 67842 4228 67844
rect 4172 67790 4174 67842
rect 4174 67790 4226 67842
rect 4226 67790 4228 67842
rect 4172 67788 4228 67790
rect 6524 77756 6580 77812
rect 6300 77138 6356 77140
rect 6300 77086 6302 77138
rect 6302 77086 6354 77138
rect 6354 77086 6356 77138
rect 6300 77084 6356 77086
rect 6524 77196 6580 77252
rect 6636 77084 6692 77140
rect 6748 77868 6804 77924
rect 7532 78988 7588 79044
rect 8204 78818 8260 78820
rect 8204 78766 8206 78818
rect 8206 78766 8258 78818
rect 8258 78766 8260 78818
rect 8204 78764 8260 78766
rect 9212 80274 9268 80276
rect 9212 80222 9214 80274
rect 9214 80222 9266 80274
rect 9266 80222 9268 80274
rect 9212 80220 9268 80222
rect 9100 80108 9156 80164
rect 8764 79436 8820 79492
rect 7084 78594 7140 78596
rect 7084 78542 7086 78594
rect 7086 78542 7138 78594
rect 7138 78542 7140 78594
rect 7084 78540 7140 78542
rect 6860 77196 6916 77252
rect 7308 77810 7364 77812
rect 7308 77758 7310 77810
rect 7310 77758 7362 77810
rect 7362 77758 7364 77810
rect 7308 77756 7364 77758
rect 7756 78034 7812 78036
rect 7756 77982 7758 78034
rect 7758 77982 7810 78034
rect 7810 77982 7812 78034
rect 7756 77980 7812 77982
rect 7420 77308 7476 77364
rect 8652 77980 8708 78036
rect 8316 77644 8372 77700
rect 6524 76354 6580 76356
rect 6524 76302 6526 76354
rect 6526 76302 6578 76354
rect 6578 76302 6580 76354
rect 6524 76300 6580 76302
rect 6748 76300 6804 76356
rect 6076 75292 6132 75348
rect 6188 74620 6244 74676
rect 6188 74060 6244 74116
rect 6636 75292 6692 75348
rect 6636 74284 6692 74340
rect 6076 73330 6132 73332
rect 6076 73278 6078 73330
rect 6078 73278 6130 73330
rect 6130 73278 6132 73330
rect 6076 73276 6132 73278
rect 5964 72546 6020 72548
rect 5964 72494 5966 72546
rect 5966 72494 6018 72546
rect 6018 72494 6020 72546
rect 5964 72492 6020 72494
rect 6300 72492 6356 72548
rect 6412 72380 6468 72436
rect 6188 70028 6244 70084
rect 3612 66108 3668 66164
rect 4508 67170 4564 67172
rect 4508 67118 4510 67170
rect 4510 67118 4562 67170
rect 4562 67118 4564 67170
rect 4508 67116 4564 67118
rect 4956 67228 5012 67284
rect 5292 67564 5348 67620
rect 4732 66892 4788 66948
rect 4008 66666 4064 66668
rect 4112 66666 4168 66668
rect 4008 66614 4024 66666
rect 4024 66614 4064 66666
rect 4112 66614 4148 66666
rect 4148 66614 4168 66666
rect 4008 66612 4064 66614
rect 4112 66612 4168 66614
rect 4216 66612 4272 66668
rect 4320 66666 4376 66668
rect 4424 66666 4480 66668
rect 4528 66666 4584 66668
rect 4320 66614 4324 66666
rect 4324 66614 4376 66666
rect 4424 66614 4448 66666
rect 4448 66614 4480 66666
rect 4528 66614 4572 66666
rect 4572 66614 4584 66666
rect 4320 66612 4376 66614
rect 4424 66612 4480 66614
rect 4528 66612 4584 66614
rect 4632 66666 4688 66668
rect 4736 66666 4792 66668
rect 4840 66666 4896 66668
rect 4632 66614 4644 66666
rect 4644 66614 4688 66666
rect 4736 66614 4768 66666
rect 4768 66614 4792 66666
rect 4840 66614 4892 66666
rect 4892 66614 4896 66666
rect 4632 66612 4688 66614
rect 4736 66612 4792 66614
rect 4840 66612 4896 66614
rect 4944 66612 5000 66668
rect 5048 66666 5104 66668
rect 5152 66666 5208 66668
rect 5048 66614 5068 66666
rect 5068 66614 5104 66666
rect 5152 66614 5192 66666
rect 5192 66614 5208 66666
rect 5048 66612 5104 66614
rect 5152 66612 5208 66614
rect 5852 68012 5908 68068
rect 5628 67618 5684 67620
rect 5628 67566 5630 67618
rect 5630 67566 5682 67618
rect 5682 67566 5684 67618
rect 5628 67564 5684 67566
rect 5404 67116 5460 67172
rect 5404 66946 5460 66948
rect 5404 66894 5406 66946
rect 5406 66894 5458 66946
rect 5458 66894 5460 66946
rect 5404 66892 5460 66894
rect 4508 66162 4564 66164
rect 4508 66110 4510 66162
rect 4510 66110 4562 66162
rect 4562 66110 4564 66162
rect 4508 66108 4564 66110
rect 4396 66050 4452 66052
rect 4396 65998 4398 66050
rect 4398 65998 4450 66050
rect 4450 65998 4452 66050
rect 4396 65996 4452 65998
rect 4060 65548 4116 65604
rect 4732 65714 4788 65716
rect 4732 65662 4734 65714
rect 4734 65662 4786 65714
rect 4786 65662 4788 65714
rect 4732 65660 4788 65662
rect 6076 67452 6132 67508
rect 6412 67618 6468 67620
rect 6412 67566 6414 67618
rect 6414 67566 6466 67618
rect 6466 67566 6468 67618
rect 6412 67564 6468 67566
rect 7980 74898 8036 74900
rect 7980 74846 7982 74898
rect 7982 74846 8034 74898
rect 8034 74846 8036 74898
rect 7980 74844 8036 74846
rect 7420 74674 7476 74676
rect 7420 74622 7422 74674
rect 7422 74622 7474 74674
rect 7474 74622 7476 74674
rect 7420 74620 7476 74622
rect 8092 74620 8148 74676
rect 6972 74172 7028 74228
rect 7868 73500 7924 73556
rect 6636 72716 6692 72772
rect 7756 73276 7812 73332
rect 7868 72546 7924 72548
rect 7868 72494 7870 72546
rect 7870 72494 7922 72546
rect 7922 72494 7924 72546
rect 7868 72492 7924 72494
rect 7644 72322 7700 72324
rect 7644 72270 7646 72322
rect 7646 72270 7698 72322
rect 7698 72270 7700 72322
rect 7644 72268 7700 72270
rect 6972 70700 7028 70756
rect 8316 72380 8372 72436
rect 8540 76636 8596 76692
rect 9436 82348 9492 82404
rect 10220 83692 10276 83748
rect 9772 81116 9828 81172
rect 9884 81058 9940 81060
rect 9884 81006 9886 81058
rect 9886 81006 9938 81058
rect 9938 81006 9940 81058
rect 9884 81004 9940 81006
rect 10892 83692 10948 83748
rect 10332 82348 10388 82404
rect 10668 82738 10724 82740
rect 10668 82686 10670 82738
rect 10670 82686 10722 82738
rect 10722 82686 10724 82738
rect 10668 82684 10724 82686
rect 10444 82066 10500 82068
rect 10444 82014 10446 82066
rect 10446 82014 10498 82066
rect 10498 82014 10500 82066
rect 10444 82012 10500 82014
rect 11900 86546 11956 86548
rect 11900 86494 11902 86546
rect 11902 86494 11954 86546
rect 11954 86494 11956 86546
rect 11900 86492 11956 86494
rect 11116 86380 11172 86436
rect 12796 87164 12852 87220
rect 12460 86658 12516 86660
rect 12460 86606 12462 86658
rect 12462 86606 12514 86658
rect 12514 86606 12516 86658
rect 12460 86604 12516 86606
rect 14008 94106 14064 94108
rect 14112 94106 14168 94108
rect 14008 94054 14024 94106
rect 14024 94054 14064 94106
rect 14112 94054 14148 94106
rect 14148 94054 14168 94106
rect 14008 94052 14064 94054
rect 14112 94052 14168 94054
rect 14216 94052 14272 94108
rect 14320 94106 14376 94108
rect 14424 94106 14480 94108
rect 14528 94106 14584 94108
rect 14320 94054 14324 94106
rect 14324 94054 14376 94106
rect 14424 94054 14448 94106
rect 14448 94054 14480 94106
rect 14528 94054 14572 94106
rect 14572 94054 14584 94106
rect 14320 94052 14376 94054
rect 14424 94052 14480 94054
rect 14528 94052 14584 94054
rect 14632 94106 14688 94108
rect 14736 94106 14792 94108
rect 14840 94106 14896 94108
rect 14632 94054 14644 94106
rect 14644 94054 14688 94106
rect 14736 94054 14768 94106
rect 14768 94054 14792 94106
rect 14840 94054 14892 94106
rect 14892 94054 14896 94106
rect 14632 94052 14688 94054
rect 14736 94052 14792 94054
rect 14840 94052 14896 94054
rect 14944 94052 15000 94108
rect 15048 94106 15104 94108
rect 15152 94106 15208 94108
rect 15048 94054 15068 94106
rect 15068 94054 15104 94106
rect 15152 94054 15192 94106
rect 15192 94054 15208 94106
rect 15048 94052 15104 94054
rect 15152 94052 15208 94054
rect 24008 93322 24064 93324
rect 24112 93322 24168 93324
rect 24008 93270 24024 93322
rect 24024 93270 24064 93322
rect 24112 93270 24148 93322
rect 24148 93270 24168 93322
rect 24008 93268 24064 93270
rect 24112 93268 24168 93270
rect 24216 93268 24272 93324
rect 24320 93322 24376 93324
rect 24424 93322 24480 93324
rect 24528 93322 24584 93324
rect 24320 93270 24324 93322
rect 24324 93270 24376 93322
rect 24424 93270 24448 93322
rect 24448 93270 24480 93322
rect 24528 93270 24572 93322
rect 24572 93270 24584 93322
rect 24320 93268 24376 93270
rect 24424 93268 24480 93270
rect 24528 93268 24584 93270
rect 24632 93322 24688 93324
rect 24736 93322 24792 93324
rect 24840 93322 24896 93324
rect 24632 93270 24644 93322
rect 24644 93270 24688 93322
rect 24736 93270 24768 93322
rect 24768 93270 24792 93322
rect 24840 93270 24892 93322
rect 24892 93270 24896 93322
rect 24632 93268 24688 93270
rect 24736 93268 24792 93270
rect 24840 93268 24896 93270
rect 24944 93268 25000 93324
rect 25048 93322 25104 93324
rect 25152 93322 25208 93324
rect 25048 93270 25068 93322
rect 25068 93270 25104 93322
rect 25152 93270 25192 93322
rect 25192 93270 25208 93322
rect 25048 93268 25104 93270
rect 25152 93268 25208 93270
rect 14008 92538 14064 92540
rect 14112 92538 14168 92540
rect 14008 92486 14024 92538
rect 14024 92486 14064 92538
rect 14112 92486 14148 92538
rect 14148 92486 14168 92538
rect 14008 92484 14064 92486
rect 14112 92484 14168 92486
rect 14216 92484 14272 92540
rect 14320 92538 14376 92540
rect 14424 92538 14480 92540
rect 14528 92538 14584 92540
rect 14320 92486 14324 92538
rect 14324 92486 14376 92538
rect 14424 92486 14448 92538
rect 14448 92486 14480 92538
rect 14528 92486 14572 92538
rect 14572 92486 14584 92538
rect 14320 92484 14376 92486
rect 14424 92484 14480 92486
rect 14528 92484 14584 92486
rect 14632 92538 14688 92540
rect 14736 92538 14792 92540
rect 14840 92538 14896 92540
rect 14632 92486 14644 92538
rect 14644 92486 14688 92538
rect 14736 92486 14768 92538
rect 14768 92486 14792 92538
rect 14840 92486 14892 92538
rect 14892 92486 14896 92538
rect 14632 92484 14688 92486
rect 14736 92484 14792 92486
rect 14840 92484 14896 92486
rect 14944 92484 15000 92540
rect 15048 92538 15104 92540
rect 15152 92538 15208 92540
rect 15048 92486 15068 92538
rect 15068 92486 15104 92538
rect 15152 92486 15192 92538
rect 15192 92486 15208 92538
rect 15048 92484 15104 92486
rect 15152 92484 15208 92486
rect 24008 91754 24064 91756
rect 24112 91754 24168 91756
rect 24008 91702 24024 91754
rect 24024 91702 24064 91754
rect 24112 91702 24148 91754
rect 24148 91702 24168 91754
rect 24008 91700 24064 91702
rect 24112 91700 24168 91702
rect 24216 91700 24272 91756
rect 24320 91754 24376 91756
rect 24424 91754 24480 91756
rect 24528 91754 24584 91756
rect 24320 91702 24324 91754
rect 24324 91702 24376 91754
rect 24424 91702 24448 91754
rect 24448 91702 24480 91754
rect 24528 91702 24572 91754
rect 24572 91702 24584 91754
rect 24320 91700 24376 91702
rect 24424 91700 24480 91702
rect 24528 91700 24584 91702
rect 24632 91754 24688 91756
rect 24736 91754 24792 91756
rect 24840 91754 24896 91756
rect 24632 91702 24644 91754
rect 24644 91702 24688 91754
rect 24736 91702 24768 91754
rect 24768 91702 24792 91754
rect 24840 91702 24892 91754
rect 24892 91702 24896 91754
rect 24632 91700 24688 91702
rect 24736 91700 24792 91702
rect 24840 91700 24896 91702
rect 24944 91700 25000 91756
rect 25048 91754 25104 91756
rect 25152 91754 25208 91756
rect 25048 91702 25068 91754
rect 25068 91702 25104 91754
rect 25152 91702 25192 91754
rect 25192 91702 25208 91754
rect 25048 91700 25104 91702
rect 25152 91700 25208 91702
rect 14008 90970 14064 90972
rect 14112 90970 14168 90972
rect 14008 90918 14024 90970
rect 14024 90918 14064 90970
rect 14112 90918 14148 90970
rect 14148 90918 14168 90970
rect 14008 90916 14064 90918
rect 14112 90916 14168 90918
rect 14216 90916 14272 90972
rect 14320 90970 14376 90972
rect 14424 90970 14480 90972
rect 14528 90970 14584 90972
rect 14320 90918 14324 90970
rect 14324 90918 14376 90970
rect 14424 90918 14448 90970
rect 14448 90918 14480 90970
rect 14528 90918 14572 90970
rect 14572 90918 14584 90970
rect 14320 90916 14376 90918
rect 14424 90916 14480 90918
rect 14528 90916 14584 90918
rect 14632 90970 14688 90972
rect 14736 90970 14792 90972
rect 14840 90970 14896 90972
rect 14632 90918 14644 90970
rect 14644 90918 14688 90970
rect 14736 90918 14768 90970
rect 14768 90918 14792 90970
rect 14840 90918 14892 90970
rect 14892 90918 14896 90970
rect 14632 90916 14688 90918
rect 14736 90916 14792 90918
rect 14840 90916 14896 90918
rect 14944 90916 15000 90972
rect 15048 90970 15104 90972
rect 15152 90970 15208 90972
rect 15048 90918 15068 90970
rect 15068 90918 15104 90970
rect 15152 90918 15192 90970
rect 15192 90918 15208 90970
rect 15048 90916 15104 90918
rect 15152 90916 15208 90918
rect 24008 90186 24064 90188
rect 24112 90186 24168 90188
rect 24008 90134 24024 90186
rect 24024 90134 24064 90186
rect 24112 90134 24148 90186
rect 24148 90134 24168 90186
rect 24008 90132 24064 90134
rect 24112 90132 24168 90134
rect 24216 90132 24272 90188
rect 24320 90186 24376 90188
rect 24424 90186 24480 90188
rect 24528 90186 24584 90188
rect 24320 90134 24324 90186
rect 24324 90134 24376 90186
rect 24424 90134 24448 90186
rect 24448 90134 24480 90186
rect 24528 90134 24572 90186
rect 24572 90134 24584 90186
rect 24320 90132 24376 90134
rect 24424 90132 24480 90134
rect 24528 90132 24584 90134
rect 24632 90186 24688 90188
rect 24736 90186 24792 90188
rect 24840 90186 24896 90188
rect 24632 90134 24644 90186
rect 24644 90134 24688 90186
rect 24736 90134 24768 90186
rect 24768 90134 24792 90186
rect 24840 90134 24892 90186
rect 24892 90134 24896 90186
rect 24632 90132 24688 90134
rect 24736 90132 24792 90134
rect 24840 90132 24896 90134
rect 24944 90132 25000 90188
rect 25048 90186 25104 90188
rect 25152 90186 25208 90188
rect 25048 90134 25068 90186
rect 25068 90134 25104 90186
rect 25152 90134 25192 90186
rect 25192 90134 25208 90186
rect 25048 90132 25104 90134
rect 25152 90132 25208 90134
rect 14008 89402 14064 89404
rect 14112 89402 14168 89404
rect 14008 89350 14024 89402
rect 14024 89350 14064 89402
rect 14112 89350 14148 89402
rect 14148 89350 14168 89402
rect 14008 89348 14064 89350
rect 14112 89348 14168 89350
rect 14216 89348 14272 89404
rect 14320 89402 14376 89404
rect 14424 89402 14480 89404
rect 14528 89402 14584 89404
rect 14320 89350 14324 89402
rect 14324 89350 14376 89402
rect 14424 89350 14448 89402
rect 14448 89350 14480 89402
rect 14528 89350 14572 89402
rect 14572 89350 14584 89402
rect 14320 89348 14376 89350
rect 14424 89348 14480 89350
rect 14528 89348 14584 89350
rect 14632 89402 14688 89404
rect 14736 89402 14792 89404
rect 14840 89402 14896 89404
rect 14632 89350 14644 89402
rect 14644 89350 14688 89402
rect 14736 89350 14768 89402
rect 14768 89350 14792 89402
rect 14840 89350 14892 89402
rect 14892 89350 14896 89402
rect 14632 89348 14688 89350
rect 14736 89348 14792 89350
rect 14840 89348 14896 89350
rect 14944 89348 15000 89404
rect 15048 89402 15104 89404
rect 15152 89402 15208 89404
rect 15048 89350 15068 89402
rect 15068 89350 15104 89402
rect 15152 89350 15192 89402
rect 15192 89350 15208 89402
rect 15048 89348 15104 89350
rect 15152 89348 15208 89350
rect 13916 88898 13972 88900
rect 13916 88846 13918 88898
rect 13918 88846 13970 88898
rect 13970 88846 13972 88898
rect 13916 88844 13972 88846
rect 14252 88844 14308 88900
rect 13244 88172 13300 88228
rect 12908 86604 12964 86660
rect 12348 85820 12404 85876
rect 11004 82124 11060 82180
rect 11788 84252 11844 84308
rect 11228 82292 11284 82348
rect 11788 82572 11844 82628
rect 11900 82124 11956 82180
rect 10220 81452 10276 81508
rect 10108 80498 10164 80500
rect 10108 80446 10110 80498
rect 10110 80446 10162 80498
rect 10162 80446 10164 80498
rect 10108 80444 10164 80446
rect 9660 80162 9716 80164
rect 9660 80110 9662 80162
rect 9662 80110 9714 80162
rect 9714 80110 9716 80162
rect 9660 80108 9716 80110
rect 9212 78092 9268 78148
rect 9660 79100 9716 79156
rect 9660 77868 9716 77924
rect 8876 77308 8932 77364
rect 9772 78876 9828 78932
rect 11452 81788 11508 81844
rect 10332 80668 10388 80724
rect 10668 81004 10724 81060
rect 11676 81170 11732 81172
rect 11676 81118 11678 81170
rect 11678 81118 11730 81170
rect 11730 81118 11732 81170
rect 11676 81116 11732 81118
rect 11004 80780 11060 80836
rect 10780 80668 10836 80724
rect 10556 80332 10612 80388
rect 10556 80108 10612 80164
rect 10556 79436 10612 79492
rect 9884 78764 9940 78820
rect 9996 78540 10052 78596
rect 10108 78034 10164 78036
rect 10108 77982 10110 78034
rect 10110 77982 10162 78034
rect 10162 77982 10164 78034
rect 10108 77980 10164 77982
rect 10108 77644 10164 77700
rect 9324 76636 9380 76692
rect 8876 75628 8932 75684
rect 8652 74844 8708 74900
rect 8540 73164 8596 73220
rect 8988 74898 9044 74900
rect 8988 74846 8990 74898
rect 8990 74846 9042 74898
rect 9042 74846 9044 74898
rect 8988 74844 9044 74846
rect 8876 74674 8932 74676
rect 8876 74622 8878 74674
rect 8878 74622 8930 74674
rect 8930 74622 8932 74674
rect 8876 74620 8932 74622
rect 8652 72322 8708 72324
rect 8652 72270 8654 72322
rect 8654 72270 8706 72322
rect 8706 72270 8708 72322
rect 8652 72268 8708 72270
rect 8428 70194 8484 70196
rect 8428 70142 8430 70194
rect 8430 70142 8482 70194
rect 8482 70142 8484 70194
rect 8428 70140 8484 70142
rect 7420 70082 7476 70084
rect 7420 70030 7422 70082
rect 7422 70030 7474 70082
rect 7474 70030 7476 70082
rect 7420 70028 7476 70030
rect 6860 68012 6916 68068
rect 6524 67340 6580 67396
rect 6300 67116 6356 67172
rect 6524 67116 6580 67172
rect 5740 66050 5796 66052
rect 5740 65998 5742 66050
rect 5742 65998 5794 66050
rect 5794 65998 5796 66050
rect 5740 65996 5796 65998
rect 3276 65212 3332 65268
rect 4008 65098 4064 65100
rect 4112 65098 4168 65100
rect 4008 65046 4024 65098
rect 4024 65046 4064 65098
rect 4112 65046 4148 65098
rect 4148 65046 4168 65098
rect 4008 65044 4064 65046
rect 4112 65044 4168 65046
rect 4216 65044 4272 65100
rect 4320 65098 4376 65100
rect 4424 65098 4480 65100
rect 4528 65098 4584 65100
rect 4320 65046 4324 65098
rect 4324 65046 4376 65098
rect 4424 65046 4448 65098
rect 4448 65046 4480 65098
rect 4528 65046 4572 65098
rect 4572 65046 4584 65098
rect 4320 65044 4376 65046
rect 4424 65044 4480 65046
rect 4528 65044 4584 65046
rect 4632 65098 4688 65100
rect 4736 65098 4792 65100
rect 4840 65098 4896 65100
rect 4632 65046 4644 65098
rect 4644 65046 4688 65098
rect 4736 65046 4768 65098
rect 4768 65046 4792 65098
rect 4840 65046 4892 65098
rect 4892 65046 4896 65098
rect 4632 65044 4688 65046
rect 4736 65044 4792 65046
rect 4840 65044 4896 65046
rect 4944 65044 5000 65100
rect 5048 65098 5104 65100
rect 5152 65098 5208 65100
rect 5048 65046 5068 65098
rect 5068 65046 5104 65098
rect 5152 65046 5192 65098
rect 5192 65046 5208 65098
rect 5048 65044 5104 65046
rect 5152 65044 5208 65046
rect 3164 64594 3220 64596
rect 3164 64542 3166 64594
rect 3166 64542 3218 64594
rect 3218 64542 3220 64594
rect 3164 64540 3220 64542
rect 3724 64594 3780 64596
rect 3724 64542 3726 64594
rect 3726 64542 3778 64594
rect 3778 64542 3780 64594
rect 3724 64540 3780 64542
rect 4844 63980 4900 64036
rect 5292 64092 5348 64148
rect 4008 63530 4064 63532
rect 4112 63530 4168 63532
rect 4008 63478 4024 63530
rect 4024 63478 4064 63530
rect 4112 63478 4148 63530
rect 4148 63478 4168 63530
rect 4008 63476 4064 63478
rect 4112 63476 4168 63478
rect 4216 63476 4272 63532
rect 4320 63530 4376 63532
rect 4424 63530 4480 63532
rect 4528 63530 4584 63532
rect 4320 63478 4324 63530
rect 4324 63478 4376 63530
rect 4424 63478 4448 63530
rect 4448 63478 4480 63530
rect 4528 63478 4572 63530
rect 4572 63478 4584 63530
rect 4320 63476 4376 63478
rect 4424 63476 4480 63478
rect 4528 63476 4584 63478
rect 4632 63530 4688 63532
rect 4736 63530 4792 63532
rect 4840 63530 4896 63532
rect 4632 63478 4644 63530
rect 4644 63478 4688 63530
rect 4736 63478 4768 63530
rect 4768 63478 4792 63530
rect 4840 63478 4892 63530
rect 4892 63478 4896 63530
rect 4632 63476 4688 63478
rect 4736 63476 4792 63478
rect 4840 63476 4896 63478
rect 4944 63476 5000 63532
rect 5048 63530 5104 63532
rect 5152 63530 5208 63532
rect 5048 63478 5068 63530
rect 5068 63478 5104 63530
rect 5152 63478 5192 63530
rect 5192 63478 5208 63530
rect 5048 63476 5104 63478
rect 5152 63476 5208 63478
rect 3836 63362 3892 63364
rect 3836 63310 3838 63362
rect 3838 63310 3890 63362
rect 3890 63310 3892 63362
rect 3836 63308 3892 63310
rect 4732 63308 4788 63364
rect 4172 63250 4228 63252
rect 4172 63198 4174 63250
rect 4174 63198 4226 63250
rect 4226 63198 4228 63250
rect 4172 63196 4228 63198
rect 3500 62972 3556 63028
rect 4956 63138 5012 63140
rect 4956 63086 4958 63138
rect 4958 63086 5010 63138
rect 5010 63086 5012 63138
rect 4956 63084 5012 63086
rect 4732 63026 4788 63028
rect 4732 62974 4734 63026
rect 4734 62974 4786 63026
rect 4786 62974 4788 63026
rect 4732 62972 4788 62974
rect 4396 62354 4452 62356
rect 4396 62302 4398 62354
rect 4398 62302 4450 62354
rect 4450 62302 4452 62354
rect 4396 62300 4452 62302
rect 4844 62466 4900 62468
rect 4844 62414 4846 62466
rect 4846 62414 4898 62466
rect 4898 62414 4900 62466
rect 4844 62412 4900 62414
rect 4844 62188 4900 62244
rect 5404 63922 5460 63924
rect 5404 63870 5406 63922
rect 5406 63870 5458 63922
rect 5458 63870 5460 63922
rect 5404 63868 5460 63870
rect 5404 63196 5460 63252
rect 5628 65490 5684 65492
rect 5628 65438 5630 65490
rect 5630 65438 5682 65490
rect 5682 65438 5684 65490
rect 5628 65436 5684 65438
rect 5740 65100 5796 65156
rect 6412 66274 6468 66276
rect 6412 66222 6414 66274
rect 6414 66222 6466 66274
rect 6466 66222 6468 66274
rect 6412 66220 6468 66222
rect 5852 63980 5908 64036
rect 6076 65996 6132 66052
rect 5628 63756 5684 63812
rect 6188 65660 6244 65716
rect 6300 65436 6356 65492
rect 6188 64146 6244 64148
rect 6188 64094 6190 64146
rect 6190 64094 6242 64146
rect 6242 64094 6244 64146
rect 6188 64092 6244 64094
rect 6188 63138 6244 63140
rect 6188 63086 6190 63138
rect 6190 63086 6242 63138
rect 6242 63086 6244 63138
rect 6188 63084 6244 63086
rect 5516 62412 5572 62468
rect 4956 62076 5012 62132
rect 5292 62076 5348 62132
rect 4008 61962 4064 61964
rect 4112 61962 4168 61964
rect 4008 61910 4024 61962
rect 4024 61910 4064 61962
rect 4112 61910 4148 61962
rect 4148 61910 4168 61962
rect 4008 61908 4064 61910
rect 4112 61908 4168 61910
rect 4216 61908 4272 61964
rect 4320 61962 4376 61964
rect 4424 61962 4480 61964
rect 4528 61962 4584 61964
rect 4320 61910 4324 61962
rect 4324 61910 4376 61962
rect 4424 61910 4448 61962
rect 4448 61910 4480 61962
rect 4528 61910 4572 61962
rect 4572 61910 4584 61962
rect 4320 61908 4376 61910
rect 4424 61908 4480 61910
rect 4528 61908 4584 61910
rect 4632 61962 4688 61964
rect 4736 61962 4792 61964
rect 4840 61962 4896 61964
rect 4632 61910 4644 61962
rect 4644 61910 4688 61962
rect 4736 61910 4768 61962
rect 4768 61910 4792 61962
rect 4840 61910 4892 61962
rect 4892 61910 4896 61962
rect 4632 61908 4688 61910
rect 4736 61908 4792 61910
rect 4840 61908 4896 61910
rect 4944 61908 5000 61964
rect 5048 61962 5104 61964
rect 5152 61962 5208 61964
rect 5048 61910 5068 61962
rect 5068 61910 5104 61962
rect 5152 61910 5192 61962
rect 5192 61910 5208 61962
rect 5048 61908 5104 61910
rect 5152 61908 5208 61910
rect 4060 61570 4116 61572
rect 4060 61518 4062 61570
rect 4062 61518 4114 61570
rect 4114 61518 4116 61570
rect 4060 61516 4116 61518
rect 3836 61404 3892 61460
rect 3724 61346 3780 61348
rect 3724 61294 3726 61346
rect 3726 61294 3778 61346
rect 3778 61294 3780 61346
rect 3724 61292 3780 61294
rect 3276 56642 3332 56644
rect 3276 56590 3278 56642
rect 3278 56590 3330 56642
rect 3330 56590 3332 56642
rect 3276 56588 3332 56590
rect 3276 55970 3332 55972
rect 3276 55918 3278 55970
rect 3278 55918 3330 55970
rect 3330 55918 3332 55970
rect 3276 55916 3332 55918
rect 2604 54908 2660 54964
rect 2492 53788 2548 53844
rect 2492 52946 2548 52948
rect 2492 52894 2494 52946
rect 2494 52894 2546 52946
rect 2546 52894 2548 52946
rect 2492 52892 2548 52894
rect 2828 52668 2884 52724
rect 3276 55244 3332 55300
rect 3276 53842 3332 53844
rect 3276 53790 3278 53842
rect 3278 53790 3330 53842
rect 3330 53790 3332 53842
rect 3276 53788 3332 53790
rect 3276 53228 3332 53284
rect 3164 52556 3220 52612
rect 2380 51324 2436 51380
rect 2156 50428 2212 50484
rect 3724 58492 3780 58548
rect 4620 61404 4676 61460
rect 4732 61292 4788 61348
rect 4008 60394 4064 60396
rect 4112 60394 4168 60396
rect 4008 60342 4024 60394
rect 4024 60342 4064 60394
rect 4112 60342 4148 60394
rect 4148 60342 4168 60394
rect 4008 60340 4064 60342
rect 4112 60340 4168 60342
rect 4216 60340 4272 60396
rect 4320 60394 4376 60396
rect 4424 60394 4480 60396
rect 4528 60394 4584 60396
rect 4320 60342 4324 60394
rect 4324 60342 4376 60394
rect 4424 60342 4448 60394
rect 4448 60342 4480 60394
rect 4528 60342 4572 60394
rect 4572 60342 4584 60394
rect 4320 60340 4376 60342
rect 4424 60340 4480 60342
rect 4528 60340 4584 60342
rect 4632 60394 4688 60396
rect 4736 60394 4792 60396
rect 4840 60394 4896 60396
rect 4632 60342 4644 60394
rect 4644 60342 4688 60394
rect 4736 60342 4768 60394
rect 4768 60342 4792 60394
rect 4840 60342 4892 60394
rect 4892 60342 4896 60394
rect 4632 60340 4688 60342
rect 4736 60340 4792 60342
rect 4840 60340 4896 60342
rect 4944 60340 5000 60396
rect 5048 60394 5104 60396
rect 5152 60394 5208 60396
rect 5048 60342 5068 60394
rect 5068 60342 5104 60394
rect 5152 60342 5192 60394
rect 5192 60342 5208 60394
rect 5048 60340 5104 60342
rect 5152 60340 5208 60342
rect 5628 61516 5684 61572
rect 5964 61628 6020 61684
rect 5740 61346 5796 61348
rect 5740 61294 5742 61346
rect 5742 61294 5794 61346
rect 5794 61294 5796 61346
rect 5740 61292 5796 61294
rect 5852 60844 5908 60900
rect 5740 60114 5796 60116
rect 5740 60062 5742 60114
rect 5742 60062 5794 60114
rect 5794 60062 5796 60114
rect 5740 60060 5796 60062
rect 4008 58826 4064 58828
rect 4112 58826 4168 58828
rect 4008 58774 4024 58826
rect 4024 58774 4064 58826
rect 4112 58774 4148 58826
rect 4148 58774 4168 58826
rect 4008 58772 4064 58774
rect 4112 58772 4168 58774
rect 4216 58772 4272 58828
rect 4320 58826 4376 58828
rect 4424 58826 4480 58828
rect 4528 58826 4584 58828
rect 4320 58774 4324 58826
rect 4324 58774 4376 58826
rect 4424 58774 4448 58826
rect 4448 58774 4480 58826
rect 4528 58774 4572 58826
rect 4572 58774 4584 58826
rect 4320 58772 4376 58774
rect 4424 58772 4480 58774
rect 4528 58772 4584 58774
rect 4632 58826 4688 58828
rect 4736 58826 4792 58828
rect 4840 58826 4896 58828
rect 4632 58774 4644 58826
rect 4644 58774 4688 58826
rect 4736 58774 4768 58826
rect 4768 58774 4792 58826
rect 4840 58774 4892 58826
rect 4892 58774 4896 58826
rect 4632 58772 4688 58774
rect 4736 58772 4792 58774
rect 4840 58772 4896 58774
rect 4944 58772 5000 58828
rect 5048 58826 5104 58828
rect 5152 58826 5208 58828
rect 5048 58774 5068 58826
rect 5068 58774 5104 58826
rect 5152 58774 5192 58826
rect 5192 58774 5208 58826
rect 5048 58772 5104 58774
rect 5152 58772 5208 58774
rect 3948 58546 4004 58548
rect 3948 58494 3950 58546
rect 3950 58494 4002 58546
rect 4002 58494 4004 58546
rect 3948 58492 4004 58494
rect 4008 57258 4064 57260
rect 4112 57258 4168 57260
rect 4008 57206 4024 57258
rect 4024 57206 4064 57258
rect 4112 57206 4148 57258
rect 4148 57206 4168 57258
rect 4008 57204 4064 57206
rect 4112 57204 4168 57206
rect 4216 57204 4272 57260
rect 4320 57258 4376 57260
rect 4424 57258 4480 57260
rect 4528 57258 4584 57260
rect 4320 57206 4324 57258
rect 4324 57206 4376 57258
rect 4424 57206 4448 57258
rect 4448 57206 4480 57258
rect 4528 57206 4572 57258
rect 4572 57206 4584 57258
rect 4320 57204 4376 57206
rect 4424 57204 4480 57206
rect 4528 57204 4584 57206
rect 4632 57258 4688 57260
rect 4736 57258 4792 57260
rect 4840 57258 4896 57260
rect 4632 57206 4644 57258
rect 4644 57206 4688 57258
rect 4736 57206 4768 57258
rect 4768 57206 4792 57258
rect 4840 57206 4892 57258
rect 4892 57206 4896 57258
rect 4632 57204 4688 57206
rect 4736 57204 4792 57206
rect 4840 57204 4896 57206
rect 4944 57204 5000 57260
rect 5048 57258 5104 57260
rect 5152 57258 5208 57260
rect 5048 57206 5068 57258
rect 5068 57206 5104 57258
rect 5152 57206 5192 57258
rect 5192 57206 5208 57258
rect 5048 57204 5104 57206
rect 5152 57204 5208 57206
rect 4396 56754 4452 56756
rect 4396 56702 4398 56754
rect 4398 56702 4450 56754
rect 4450 56702 4452 56754
rect 4396 56700 4452 56702
rect 5292 56700 5348 56756
rect 4284 56588 4340 56644
rect 4956 56642 5012 56644
rect 4956 56590 4958 56642
rect 4958 56590 5010 56642
rect 5010 56590 5012 56642
rect 4956 56588 5012 56590
rect 4172 56252 4228 56308
rect 4008 55690 4064 55692
rect 4112 55690 4168 55692
rect 4008 55638 4024 55690
rect 4024 55638 4064 55690
rect 4112 55638 4148 55690
rect 4148 55638 4168 55690
rect 4008 55636 4064 55638
rect 4112 55636 4168 55638
rect 4216 55636 4272 55692
rect 4320 55690 4376 55692
rect 4424 55690 4480 55692
rect 4528 55690 4584 55692
rect 4320 55638 4324 55690
rect 4324 55638 4376 55690
rect 4424 55638 4448 55690
rect 4448 55638 4480 55690
rect 4528 55638 4572 55690
rect 4572 55638 4584 55690
rect 4320 55636 4376 55638
rect 4424 55636 4480 55638
rect 4528 55636 4584 55638
rect 4632 55690 4688 55692
rect 4736 55690 4792 55692
rect 4840 55690 4896 55692
rect 4632 55638 4644 55690
rect 4644 55638 4688 55690
rect 4736 55638 4768 55690
rect 4768 55638 4792 55690
rect 4840 55638 4892 55690
rect 4892 55638 4896 55690
rect 4632 55636 4688 55638
rect 4736 55636 4792 55638
rect 4840 55636 4896 55638
rect 4944 55636 5000 55692
rect 5048 55690 5104 55692
rect 5152 55690 5208 55692
rect 5048 55638 5068 55690
rect 5068 55638 5104 55690
rect 5152 55638 5192 55690
rect 5192 55638 5208 55690
rect 5048 55636 5104 55638
rect 5152 55636 5208 55638
rect 3724 55356 3780 55412
rect 3500 53116 3556 53172
rect 3612 55244 3668 55300
rect 3724 54684 3780 54740
rect 4844 55298 4900 55300
rect 4844 55246 4846 55298
rect 4846 55246 4898 55298
rect 4898 55246 4900 55298
rect 4844 55244 4900 55246
rect 4956 55186 5012 55188
rect 4956 55134 4958 55186
rect 4958 55134 5010 55186
rect 5010 55134 5012 55186
rect 4956 55132 5012 55134
rect 5740 56252 5796 56308
rect 5740 55074 5796 55076
rect 5740 55022 5742 55074
rect 5742 55022 5794 55074
rect 5794 55022 5796 55074
rect 5740 55020 5796 55022
rect 5628 54738 5684 54740
rect 5628 54686 5630 54738
rect 5630 54686 5682 54738
rect 5682 54686 5684 54738
rect 5628 54684 5684 54686
rect 4732 54236 4788 54292
rect 4008 54122 4064 54124
rect 4112 54122 4168 54124
rect 4008 54070 4024 54122
rect 4024 54070 4064 54122
rect 4112 54070 4148 54122
rect 4148 54070 4168 54122
rect 4008 54068 4064 54070
rect 4112 54068 4168 54070
rect 4216 54068 4272 54124
rect 4320 54122 4376 54124
rect 4424 54122 4480 54124
rect 4528 54122 4584 54124
rect 4320 54070 4324 54122
rect 4324 54070 4376 54122
rect 4424 54070 4448 54122
rect 4448 54070 4480 54122
rect 4528 54070 4572 54122
rect 4572 54070 4584 54122
rect 4320 54068 4376 54070
rect 4424 54068 4480 54070
rect 4528 54068 4584 54070
rect 4632 54122 4688 54124
rect 4736 54122 4792 54124
rect 4840 54122 4896 54124
rect 4632 54070 4644 54122
rect 4644 54070 4688 54122
rect 4736 54070 4768 54122
rect 4768 54070 4792 54122
rect 4840 54070 4892 54122
rect 4892 54070 4896 54122
rect 4632 54068 4688 54070
rect 4736 54068 4792 54070
rect 4840 54068 4896 54070
rect 4944 54068 5000 54124
rect 5048 54122 5104 54124
rect 5152 54122 5208 54124
rect 5048 54070 5068 54122
rect 5068 54070 5104 54122
rect 5152 54070 5192 54122
rect 5192 54070 5208 54122
rect 5048 54068 5104 54070
rect 5152 54068 5208 54070
rect 4060 53676 4116 53732
rect 3388 51884 3444 51940
rect 3500 52892 3556 52948
rect 3276 51324 3332 51380
rect 3388 51660 3444 51716
rect 2492 49308 2548 49364
rect 3276 48524 3332 48580
rect 2492 48242 2548 48244
rect 2492 48190 2494 48242
rect 2494 48190 2546 48242
rect 2546 48190 2548 48242
rect 2492 48188 2548 48190
rect 2940 48242 2996 48244
rect 2940 48190 2942 48242
rect 2942 48190 2994 48242
rect 2994 48190 2996 48242
rect 2940 48188 2996 48190
rect 3388 47516 3444 47572
rect 3276 47404 3332 47460
rect 2604 47346 2660 47348
rect 2604 47294 2606 47346
rect 2606 47294 2658 47346
rect 2658 47294 2660 47346
rect 2604 47292 2660 47294
rect 3388 47292 3444 47348
rect 2156 47068 2212 47124
rect 2828 47068 2884 47124
rect 2492 46674 2548 46676
rect 2492 46622 2494 46674
rect 2494 46622 2546 46674
rect 2546 46622 2548 46674
rect 2492 46620 2548 46622
rect 2492 46002 2548 46004
rect 2492 45950 2494 46002
rect 2494 45950 2546 46002
rect 2546 45950 2548 46002
rect 2492 45948 2548 45950
rect 3276 46002 3332 46004
rect 3276 45950 3278 46002
rect 3278 45950 3330 46002
rect 3330 45950 3332 46002
rect 3276 45948 3332 45950
rect 3276 45164 3332 45220
rect 2492 44828 2548 44884
rect 1820 43708 1876 43764
rect 2268 44044 2324 44100
rect 3388 43820 3444 43876
rect 3388 43596 3444 43652
rect 3164 42700 3220 42756
rect 2604 41468 2660 41524
rect 2604 40348 2660 40404
rect 2268 39788 2324 39844
rect 3164 39452 3220 39508
rect 2492 39228 2548 39284
rect 3164 39058 3220 39060
rect 3164 39006 3166 39058
rect 3166 39006 3218 39058
rect 3218 39006 3220 39058
rect 3164 39004 3220 39006
rect 3276 38892 3332 38948
rect 3612 51772 3668 51828
rect 5180 53170 5236 53172
rect 5180 53118 5182 53170
rect 5182 53118 5234 53170
rect 5234 53118 5236 53170
rect 5180 53116 5236 53118
rect 4732 52834 4788 52836
rect 4732 52782 4734 52834
rect 4734 52782 4786 52834
rect 4786 52782 4788 52834
rect 4732 52780 4788 52782
rect 4008 52554 4064 52556
rect 4112 52554 4168 52556
rect 4008 52502 4024 52554
rect 4024 52502 4064 52554
rect 4112 52502 4148 52554
rect 4148 52502 4168 52554
rect 4008 52500 4064 52502
rect 4112 52500 4168 52502
rect 4216 52500 4272 52556
rect 4320 52554 4376 52556
rect 4424 52554 4480 52556
rect 4528 52554 4584 52556
rect 4320 52502 4324 52554
rect 4324 52502 4376 52554
rect 4424 52502 4448 52554
rect 4448 52502 4480 52554
rect 4528 52502 4572 52554
rect 4572 52502 4584 52554
rect 4320 52500 4376 52502
rect 4424 52500 4480 52502
rect 4528 52500 4584 52502
rect 4632 52554 4688 52556
rect 4736 52554 4792 52556
rect 4840 52554 4896 52556
rect 4632 52502 4644 52554
rect 4644 52502 4688 52554
rect 4736 52502 4768 52554
rect 4768 52502 4792 52554
rect 4840 52502 4892 52554
rect 4892 52502 4896 52554
rect 4632 52500 4688 52502
rect 4736 52500 4792 52502
rect 4840 52500 4896 52502
rect 4944 52500 5000 52556
rect 5048 52554 5104 52556
rect 5152 52554 5208 52556
rect 5048 52502 5068 52554
rect 5068 52502 5104 52554
rect 5152 52502 5192 52554
rect 5192 52502 5208 52554
rect 5048 52500 5104 52502
rect 5152 52500 5208 52502
rect 5740 54236 5796 54292
rect 5628 53730 5684 53732
rect 5628 53678 5630 53730
rect 5630 53678 5682 53730
rect 5682 53678 5684 53730
rect 5628 53676 5684 53678
rect 5740 53618 5796 53620
rect 5740 53566 5742 53618
rect 5742 53566 5794 53618
rect 5794 53566 5796 53618
rect 5740 53564 5796 53566
rect 6188 59724 6244 59780
rect 6076 57484 6132 57540
rect 6972 67618 7028 67620
rect 6972 67566 6974 67618
rect 6974 67566 7026 67618
rect 7026 67566 7028 67618
rect 6972 67564 7028 67566
rect 6860 66892 6916 66948
rect 6972 66668 7028 66724
rect 6972 66274 7028 66276
rect 6972 66222 6974 66274
rect 6974 66222 7026 66274
rect 7026 66222 7028 66274
rect 6972 66220 7028 66222
rect 7420 67452 7476 67508
rect 7308 66780 7364 66836
rect 8092 66892 8148 66948
rect 7644 66556 7700 66612
rect 8428 66556 8484 66612
rect 8204 66274 8260 66276
rect 8204 66222 8206 66274
rect 8206 66222 8258 66274
rect 8258 66222 8260 66274
rect 8204 66220 8260 66222
rect 7196 65436 7252 65492
rect 8540 65436 8596 65492
rect 7756 65324 7812 65380
rect 8428 64316 8484 64372
rect 8316 63756 8372 63812
rect 7532 63362 7588 63364
rect 7532 63310 7534 63362
rect 7534 63310 7586 63362
rect 7586 63310 7588 63362
rect 7532 63308 7588 63310
rect 6860 63250 6916 63252
rect 6860 63198 6862 63250
rect 6862 63198 6914 63250
rect 6914 63198 6916 63250
rect 6860 63196 6916 63198
rect 7084 62412 7140 62468
rect 6636 61180 6692 61236
rect 7420 62300 7476 62356
rect 7084 61180 7140 61236
rect 7196 62188 7252 62244
rect 6636 60060 6692 60116
rect 6524 58716 6580 58772
rect 7532 60898 7588 60900
rect 7532 60846 7534 60898
rect 7534 60846 7586 60898
rect 7586 60846 7588 60898
rect 7532 60844 7588 60846
rect 7420 60786 7476 60788
rect 7420 60734 7422 60786
rect 7422 60734 7474 60786
rect 7474 60734 7476 60786
rect 7420 60732 7476 60734
rect 8316 62188 8372 62244
rect 7084 60002 7140 60004
rect 7084 59950 7086 60002
rect 7086 59950 7138 60002
rect 7138 59950 7140 60002
rect 7084 59948 7140 59950
rect 8316 61292 8372 61348
rect 8204 60620 8260 60676
rect 7420 58604 7476 58660
rect 6972 57538 7028 57540
rect 6972 57486 6974 57538
rect 6974 57486 7026 57538
rect 7026 57486 7028 57538
rect 6972 57484 7028 57486
rect 6860 57260 6916 57316
rect 7532 58156 7588 58212
rect 7084 57148 7140 57204
rect 7868 57148 7924 57204
rect 6636 56754 6692 56756
rect 6636 56702 6638 56754
rect 6638 56702 6690 56754
rect 6690 56702 6692 56754
rect 6636 56700 6692 56702
rect 6524 56588 6580 56644
rect 6188 55298 6244 55300
rect 6188 55246 6190 55298
rect 6190 55246 6242 55298
rect 6242 55246 6244 55298
rect 6188 55244 6244 55246
rect 6300 54626 6356 54628
rect 6300 54574 6302 54626
rect 6302 54574 6354 54626
rect 6354 54574 6356 54626
rect 6300 54572 6356 54574
rect 6188 54514 6244 54516
rect 6188 54462 6190 54514
rect 6190 54462 6242 54514
rect 6242 54462 6244 54514
rect 6188 54460 6244 54462
rect 6300 54236 6356 54292
rect 4060 51660 4116 51716
rect 4732 51602 4788 51604
rect 4732 51550 4734 51602
rect 4734 51550 4786 51602
rect 4786 51550 4788 51602
rect 4732 51548 4788 51550
rect 4956 52050 5012 52052
rect 4956 51998 4958 52050
rect 4958 51998 5010 52050
rect 5010 51998 5012 52050
rect 4956 51996 5012 51998
rect 4008 50986 4064 50988
rect 4112 50986 4168 50988
rect 4008 50934 4024 50986
rect 4024 50934 4064 50986
rect 4112 50934 4148 50986
rect 4148 50934 4168 50986
rect 4008 50932 4064 50934
rect 4112 50932 4168 50934
rect 4216 50932 4272 50988
rect 4320 50986 4376 50988
rect 4424 50986 4480 50988
rect 4528 50986 4584 50988
rect 4320 50934 4324 50986
rect 4324 50934 4376 50986
rect 4424 50934 4448 50986
rect 4448 50934 4480 50986
rect 4528 50934 4572 50986
rect 4572 50934 4584 50986
rect 4320 50932 4376 50934
rect 4424 50932 4480 50934
rect 4528 50932 4584 50934
rect 4632 50986 4688 50988
rect 4736 50986 4792 50988
rect 4840 50986 4896 50988
rect 4632 50934 4644 50986
rect 4644 50934 4688 50986
rect 4736 50934 4768 50986
rect 4768 50934 4792 50986
rect 4840 50934 4892 50986
rect 4892 50934 4896 50986
rect 4632 50932 4688 50934
rect 4736 50932 4792 50934
rect 4840 50932 4896 50934
rect 4944 50932 5000 50988
rect 5048 50986 5104 50988
rect 5152 50986 5208 50988
rect 5048 50934 5068 50986
rect 5068 50934 5104 50986
rect 5152 50934 5192 50986
rect 5192 50934 5208 50986
rect 5048 50932 5104 50934
rect 5152 50932 5208 50934
rect 3612 49868 3668 49924
rect 6188 53564 6244 53620
rect 4956 50482 5012 50484
rect 4956 50430 4958 50482
rect 4958 50430 5010 50482
rect 5010 50430 5012 50482
rect 4956 50428 5012 50430
rect 5852 53170 5908 53172
rect 5852 53118 5854 53170
rect 5854 53118 5906 53170
rect 5906 53118 5908 53170
rect 5852 53116 5908 53118
rect 6076 53058 6132 53060
rect 6076 53006 6078 53058
rect 6078 53006 6130 53058
rect 6130 53006 6132 53058
rect 6076 53004 6132 53006
rect 6188 52556 6244 52612
rect 5852 51996 5908 52052
rect 6188 51884 6244 51940
rect 6188 51548 6244 51604
rect 6076 51378 6132 51380
rect 6076 51326 6078 51378
rect 6078 51326 6130 51378
rect 6130 51326 6132 51378
rect 6076 51324 6132 51326
rect 6300 51660 6356 51716
rect 4508 49980 4564 50036
rect 5516 50034 5572 50036
rect 5516 49982 5518 50034
rect 5518 49982 5570 50034
rect 5570 49982 5572 50034
rect 5516 49980 5572 49982
rect 4008 49418 4064 49420
rect 4112 49418 4168 49420
rect 4008 49366 4024 49418
rect 4024 49366 4064 49418
rect 4112 49366 4148 49418
rect 4148 49366 4168 49418
rect 4008 49364 4064 49366
rect 4112 49364 4168 49366
rect 4216 49364 4272 49420
rect 4320 49418 4376 49420
rect 4424 49418 4480 49420
rect 4528 49418 4584 49420
rect 4320 49366 4324 49418
rect 4324 49366 4376 49418
rect 4424 49366 4448 49418
rect 4448 49366 4480 49418
rect 4528 49366 4572 49418
rect 4572 49366 4584 49418
rect 4320 49364 4376 49366
rect 4424 49364 4480 49366
rect 4528 49364 4584 49366
rect 4632 49418 4688 49420
rect 4736 49418 4792 49420
rect 4840 49418 4896 49420
rect 4632 49366 4644 49418
rect 4644 49366 4688 49418
rect 4736 49366 4768 49418
rect 4768 49366 4792 49418
rect 4840 49366 4892 49418
rect 4892 49366 4896 49418
rect 4632 49364 4688 49366
rect 4736 49364 4792 49366
rect 4840 49364 4896 49366
rect 4944 49364 5000 49420
rect 5048 49418 5104 49420
rect 5152 49418 5208 49420
rect 5048 49366 5068 49418
rect 5068 49366 5104 49418
rect 5152 49366 5192 49418
rect 5192 49366 5208 49418
rect 5048 49364 5104 49366
rect 5152 49364 5208 49366
rect 3836 48860 3892 48916
rect 3724 47346 3780 47348
rect 3724 47294 3726 47346
rect 3726 47294 3778 47346
rect 3778 47294 3780 47346
rect 3724 47292 3780 47294
rect 5628 48914 5684 48916
rect 5628 48862 5630 48914
rect 5630 48862 5682 48914
rect 5682 48862 5684 48914
rect 5628 48860 5684 48862
rect 5740 48802 5796 48804
rect 5740 48750 5742 48802
rect 5742 48750 5794 48802
rect 5794 48750 5796 48802
rect 5740 48748 5796 48750
rect 4620 48130 4676 48132
rect 4620 48078 4622 48130
rect 4622 48078 4674 48130
rect 4674 48078 4676 48130
rect 4620 48076 4676 48078
rect 4008 47850 4064 47852
rect 4112 47850 4168 47852
rect 4008 47798 4024 47850
rect 4024 47798 4064 47850
rect 4112 47798 4148 47850
rect 4148 47798 4168 47850
rect 4008 47796 4064 47798
rect 4112 47796 4168 47798
rect 4216 47796 4272 47852
rect 4320 47850 4376 47852
rect 4424 47850 4480 47852
rect 4528 47850 4584 47852
rect 4320 47798 4324 47850
rect 4324 47798 4376 47850
rect 4424 47798 4448 47850
rect 4448 47798 4480 47850
rect 4528 47798 4572 47850
rect 4572 47798 4584 47850
rect 4320 47796 4376 47798
rect 4424 47796 4480 47798
rect 4528 47796 4584 47798
rect 4632 47850 4688 47852
rect 4736 47850 4792 47852
rect 4840 47850 4896 47852
rect 4632 47798 4644 47850
rect 4644 47798 4688 47850
rect 4736 47798 4768 47850
rect 4768 47798 4792 47850
rect 4840 47798 4892 47850
rect 4892 47798 4896 47850
rect 4632 47796 4688 47798
rect 4736 47796 4792 47798
rect 4840 47796 4896 47798
rect 4944 47796 5000 47852
rect 5048 47850 5104 47852
rect 5152 47850 5208 47852
rect 5048 47798 5068 47850
rect 5068 47798 5104 47850
rect 5152 47798 5192 47850
rect 5192 47798 5208 47850
rect 5048 47796 5104 47798
rect 5152 47796 5208 47798
rect 4956 47068 5012 47124
rect 4844 46956 4900 47012
rect 5628 46956 5684 47012
rect 5516 46898 5572 46900
rect 5516 46846 5518 46898
rect 5518 46846 5570 46898
rect 5570 46846 5572 46898
rect 5516 46844 5572 46846
rect 3836 46620 3892 46676
rect 3500 42588 3556 42644
rect 4008 46282 4064 46284
rect 4112 46282 4168 46284
rect 4008 46230 4024 46282
rect 4024 46230 4064 46282
rect 4112 46230 4148 46282
rect 4148 46230 4168 46282
rect 4008 46228 4064 46230
rect 4112 46228 4168 46230
rect 4216 46228 4272 46284
rect 4320 46282 4376 46284
rect 4424 46282 4480 46284
rect 4528 46282 4584 46284
rect 4320 46230 4324 46282
rect 4324 46230 4376 46282
rect 4424 46230 4448 46282
rect 4448 46230 4480 46282
rect 4528 46230 4572 46282
rect 4572 46230 4584 46282
rect 4320 46228 4376 46230
rect 4424 46228 4480 46230
rect 4528 46228 4584 46230
rect 4632 46282 4688 46284
rect 4736 46282 4792 46284
rect 4840 46282 4896 46284
rect 4632 46230 4644 46282
rect 4644 46230 4688 46282
rect 4736 46230 4768 46282
rect 4768 46230 4792 46282
rect 4840 46230 4892 46282
rect 4892 46230 4896 46282
rect 4632 46228 4688 46230
rect 4736 46228 4792 46230
rect 4840 46228 4896 46230
rect 4944 46228 5000 46284
rect 5048 46282 5104 46284
rect 5152 46282 5208 46284
rect 5048 46230 5068 46282
rect 5068 46230 5104 46282
rect 5152 46230 5192 46282
rect 5192 46230 5208 46282
rect 5048 46228 5104 46230
rect 5152 46228 5208 46230
rect 4172 45164 4228 45220
rect 4956 45778 5012 45780
rect 4956 45726 4958 45778
rect 4958 45726 5010 45778
rect 5010 45726 5012 45778
rect 4956 45724 5012 45726
rect 5740 46786 5796 46788
rect 5740 46734 5742 46786
rect 5742 46734 5794 46786
rect 5794 46734 5796 46786
rect 5740 46732 5796 46734
rect 5516 45724 5572 45780
rect 5628 45218 5684 45220
rect 5628 45166 5630 45218
rect 5630 45166 5682 45218
rect 5682 45166 5684 45218
rect 5628 45164 5684 45166
rect 4396 44828 4452 44884
rect 5292 44828 5348 44884
rect 5852 45388 5908 45444
rect 6076 44940 6132 44996
rect 4008 44714 4064 44716
rect 4112 44714 4168 44716
rect 4008 44662 4024 44714
rect 4024 44662 4064 44714
rect 4112 44662 4148 44714
rect 4148 44662 4168 44714
rect 4008 44660 4064 44662
rect 4112 44660 4168 44662
rect 4216 44660 4272 44716
rect 4320 44714 4376 44716
rect 4424 44714 4480 44716
rect 4528 44714 4584 44716
rect 4320 44662 4324 44714
rect 4324 44662 4376 44714
rect 4424 44662 4448 44714
rect 4448 44662 4480 44714
rect 4528 44662 4572 44714
rect 4572 44662 4584 44714
rect 4320 44660 4376 44662
rect 4424 44660 4480 44662
rect 4528 44660 4584 44662
rect 4632 44714 4688 44716
rect 4736 44714 4792 44716
rect 4840 44714 4896 44716
rect 4632 44662 4644 44714
rect 4644 44662 4688 44714
rect 4736 44662 4768 44714
rect 4768 44662 4792 44714
rect 4840 44662 4892 44714
rect 4892 44662 4896 44714
rect 4632 44660 4688 44662
rect 4736 44660 4792 44662
rect 4840 44660 4896 44662
rect 4944 44660 5000 44716
rect 5048 44714 5104 44716
rect 5152 44714 5208 44716
rect 5048 44662 5068 44714
rect 5068 44662 5104 44714
rect 5152 44662 5192 44714
rect 5192 44662 5208 44714
rect 5048 44660 5104 44662
rect 5152 44660 5208 44662
rect 5964 44882 6020 44884
rect 5964 44830 5966 44882
rect 5966 44830 6018 44882
rect 6018 44830 6020 44882
rect 5964 44828 6020 44830
rect 4396 44492 4452 44548
rect 3836 44098 3892 44100
rect 3836 44046 3838 44098
rect 3838 44046 3890 44098
rect 3890 44046 3892 44098
rect 3836 44044 3892 44046
rect 4956 44210 5012 44212
rect 4956 44158 4958 44210
rect 4958 44158 5010 44210
rect 5010 44158 5012 44210
rect 4956 44156 5012 44158
rect 5292 44156 5348 44212
rect 4732 43820 4788 43876
rect 6076 43820 6132 43876
rect 5628 43708 5684 43764
rect 4172 43372 4228 43428
rect 4008 43146 4064 43148
rect 4112 43146 4168 43148
rect 4008 43094 4024 43146
rect 4024 43094 4064 43146
rect 4112 43094 4148 43146
rect 4148 43094 4168 43146
rect 4008 43092 4064 43094
rect 4112 43092 4168 43094
rect 4216 43092 4272 43148
rect 4320 43146 4376 43148
rect 4424 43146 4480 43148
rect 4528 43146 4584 43148
rect 4320 43094 4324 43146
rect 4324 43094 4376 43146
rect 4424 43094 4448 43146
rect 4448 43094 4480 43146
rect 4528 43094 4572 43146
rect 4572 43094 4584 43146
rect 4320 43092 4376 43094
rect 4424 43092 4480 43094
rect 4528 43092 4584 43094
rect 4632 43146 4688 43148
rect 4736 43146 4792 43148
rect 4840 43146 4896 43148
rect 4632 43094 4644 43146
rect 4644 43094 4688 43146
rect 4736 43094 4768 43146
rect 4768 43094 4792 43146
rect 4840 43094 4892 43146
rect 4892 43094 4896 43146
rect 4632 43092 4688 43094
rect 4736 43092 4792 43094
rect 4840 43092 4896 43094
rect 4944 43092 5000 43148
rect 5048 43146 5104 43148
rect 5152 43146 5208 43148
rect 5048 43094 5068 43146
rect 5068 43094 5104 43146
rect 5152 43094 5192 43146
rect 5192 43094 5208 43146
rect 5048 43092 5104 43094
rect 5152 43092 5208 43094
rect 5068 42812 5124 42868
rect 4008 41578 4064 41580
rect 4112 41578 4168 41580
rect 4008 41526 4024 41578
rect 4024 41526 4064 41578
rect 4112 41526 4148 41578
rect 4148 41526 4168 41578
rect 4008 41524 4064 41526
rect 4112 41524 4168 41526
rect 4216 41524 4272 41580
rect 4320 41578 4376 41580
rect 4424 41578 4480 41580
rect 4528 41578 4584 41580
rect 4320 41526 4324 41578
rect 4324 41526 4376 41578
rect 4424 41526 4448 41578
rect 4448 41526 4480 41578
rect 4528 41526 4572 41578
rect 4572 41526 4584 41578
rect 4320 41524 4376 41526
rect 4424 41524 4480 41526
rect 4528 41524 4584 41526
rect 4632 41578 4688 41580
rect 4736 41578 4792 41580
rect 4840 41578 4896 41580
rect 4632 41526 4644 41578
rect 4644 41526 4688 41578
rect 4736 41526 4768 41578
rect 4768 41526 4792 41578
rect 4840 41526 4892 41578
rect 4892 41526 4896 41578
rect 4632 41524 4688 41526
rect 4736 41524 4792 41526
rect 4840 41524 4896 41526
rect 4944 41524 5000 41580
rect 5048 41578 5104 41580
rect 5152 41578 5208 41580
rect 5048 41526 5068 41578
rect 5068 41526 5104 41578
rect 5152 41526 5192 41578
rect 5192 41526 5208 41578
rect 5048 41524 5104 41526
rect 5152 41524 5208 41526
rect 5292 40908 5348 40964
rect 4732 40684 4788 40740
rect 3948 40460 4004 40516
rect 3724 39842 3780 39844
rect 3724 39790 3726 39842
rect 3726 39790 3778 39842
rect 3778 39790 3780 39842
rect 3724 39788 3780 39790
rect 4008 40010 4064 40012
rect 4112 40010 4168 40012
rect 4008 39958 4024 40010
rect 4024 39958 4064 40010
rect 4112 39958 4148 40010
rect 4148 39958 4168 40010
rect 4008 39956 4064 39958
rect 4112 39956 4168 39958
rect 4216 39956 4272 40012
rect 4320 40010 4376 40012
rect 4424 40010 4480 40012
rect 4528 40010 4584 40012
rect 4320 39958 4324 40010
rect 4324 39958 4376 40010
rect 4424 39958 4448 40010
rect 4448 39958 4480 40010
rect 4528 39958 4572 40010
rect 4572 39958 4584 40010
rect 4320 39956 4376 39958
rect 4424 39956 4480 39958
rect 4528 39956 4584 39958
rect 4632 40010 4688 40012
rect 4736 40010 4792 40012
rect 4840 40010 4896 40012
rect 4632 39958 4644 40010
rect 4644 39958 4688 40010
rect 4736 39958 4768 40010
rect 4768 39958 4792 40010
rect 4840 39958 4892 40010
rect 4892 39958 4896 40010
rect 4632 39956 4688 39958
rect 4736 39956 4792 39958
rect 4840 39956 4896 39958
rect 4944 39956 5000 40012
rect 5048 40010 5104 40012
rect 5152 40010 5208 40012
rect 5048 39958 5068 40010
rect 5068 39958 5104 40010
rect 5152 39958 5192 40010
rect 5192 39958 5208 40010
rect 5048 39956 5104 39958
rect 5152 39956 5208 39958
rect 4284 39564 4340 39620
rect 2492 38108 2548 38164
rect 3164 37378 3220 37380
rect 3164 37326 3166 37378
rect 3166 37326 3218 37378
rect 3218 37326 3220 37378
rect 3164 37324 3220 37326
rect 2492 36988 2548 37044
rect 2492 35868 2548 35924
rect 2268 34636 2324 34692
rect 3164 35420 3220 35476
rect 3052 35084 3108 35140
rect 2604 34748 2660 34804
rect 3276 34188 3332 34244
rect 2492 33404 2548 33460
rect 3164 33234 3220 33236
rect 3164 33182 3166 33234
rect 3166 33182 3218 33234
rect 3218 33182 3220 33234
rect 3164 33180 3220 33182
rect 1820 32732 1876 32788
rect 5740 43372 5796 43428
rect 6076 42866 6132 42868
rect 6076 42814 6078 42866
rect 6078 42814 6130 42866
rect 6130 42814 6132 42866
rect 6076 42812 6132 42814
rect 6636 55020 6692 55076
rect 7532 56588 7588 56644
rect 7196 55522 7252 55524
rect 7196 55470 7198 55522
rect 7198 55470 7250 55522
rect 7250 55470 7252 55522
rect 7196 55468 7252 55470
rect 7084 55132 7140 55188
rect 6860 55074 6916 55076
rect 6860 55022 6862 55074
rect 6862 55022 6914 55074
rect 6914 55022 6916 55074
rect 6860 55020 6916 55022
rect 6524 54348 6580 54404
rect 6524 53170 6580 53172
rect 6524 53118 6526 53170
rect 6526 53118 6578 53170
rect 6578 53118 6580 53170
rect 6524 53116 6580 53118
rect 6748 54684 6804 54740
rect 7196 54572 7252 54628
rect 7196 54348 7252 54404
rect 7420 54402 7476 54404
rect 7420 54350 7422 54402
rect 7422 54350 7474 54402
rect 7474 54350 7476 54402
rect 7420 54348 7476 54350
rect 6636 51324 6692 51380
rect 6748 50540 6804 50596
rect 6636 50482 6692 50484
rect 6636 50430 6638 50482
rect 6638 50430 6690 50482
rect 6690 50430 6692 50482
rect 6636 50428 6692 50430
rect 6412 46786 6468 46788
rect 6412 46734 6414 46786
rect 6414 46734 6466 46786
rect 6466 46734 6468 46786
rect 6412 46732 6468 46734
rect 6412 44210 6468 44212
rect 6412 44158 6414 44210
rect 6414 44158 6466 44210
rect 6466 44158 6468 44210
rect 6412 44156 6468 44158
rect 6972 50428 7028 50484
rect 7308 53116 7364 53172
rect 7308 50428 7364 50484
rect 7756 56082 7812 56084
rect 7756 56030 7758 56082
rect 7758 56030 7810 56082
rect 7810 56030 7812 56082
rect 7756 56028 7812 56030
rect 7868 55468 7924 55524
rect 7980 57036 8036 57092
rect 8204 58210 8260 58212
rect 8204 58158 8206 58210
rect 8206 58158 8258 58210
rect 8258 58158 8260 58210
rect 8204 58156 8260 58158
rect 8540 64092 8596 64148
rect 8540 60786 8596 60788
rect 8540 60734 8542 60786
rect 8542 60734 8594 60786
rect 8594 60734 8596 60786
rect 8540 60732 8596 60734
rect 8204 57148 8260 57204
rect 8204 55356 8260 55412
rect 7868 54684 7924 54740
rect 7644 54514 7700 54516
rect 7644 54462 7646 54514
rect 7646 54462 7698 54514
rect 7698 54462 7700 54514
rect 7644 54460 7700 54462
rect 7868 53730 7924 53732
rect 7868 53678 7870 53730
rect 7870 53678 7922 53730
rect 7922 53678 7924 53730
rect 7868 53676 7924 53678
rect 8428 56028 8484 56084
rect 8092 54572 8148 54628
rect 8540 54012 8596 54068
rect 8540 51938 8596 51940
rect 8540 51886 8542 51938
rect 8542 51886 8594 51938
rect 8594 51886 8596 51938
rect 8540 51884 8596 51886
rect 8540 51378 8596 51380
rect 8540 51326 8542 51378
rect 8542 51326 8594 51378
rect 8594 51326 8596 51378
rect 8540 51324 8596 51326
rect 7980 50540 8036 50596
rect 8316 50428 8372 50484
rect 6860 48412 6916 48468
rect 7644 49532 7700 49588
rect 8988 70082 9044 70084
rect 8988 70030 8990 70082
rect 8990 70030 9042 70082
rect 9042 70030 9044 70082
rect 8988 70028 9044 70030
rect 9100 67228 9156 67284
rect 8764 66780 8820 66836
rect 9772 76690 9828 76692
rect 9772 76638 9774 76690
rect 9774 76638 9826 76690
rect 9826 76638 9828 76690
rect 9772 76636 9828 76638
rect 10780 79212 10836 79268
rect 10556 78034 10612 78036
rect 10556 77982 10558 78034
rect 10558 77982 10610 78034
rect 10610 77982 10612 78034
rect 10556 77980 10612 77982
rect 10668 77868 10724 77924
rect 10668 76354 10724 76356
rect 10668 76302 10670 76354
rect 10670 76302 10722 76354
rect 10722 76302 10724 76354
rect 10668 76300 10724 76302
rect 9436 74172 9492 74228
rect 11004 79602 11060 79604
rect 11004 79550 11006 79602
rect 11006 79550 11058 79602
rect 11058 79550 11060 79602
rect 11004 79548 11060 79550
rect 10892 79100 10948 79156
rect 13580 88002 13636 88004
rect 13580 87950 13582 88002
rect 13582 87950 13634 88002
rect 13634 87950 13636 88002
rect 13580 87948 13636 87950
rect 13580 86658 13636 86660
rect 13580 86606 13582 86658
rect 13582 86606 13634 86658
rect 13634 86606 13636 86658
rect 13580 86604 13636 86606
rect 13580 86156 13636 86212
rect 13468 85820 13524 85876
rect 13020 84866 13076 84868
rect 13020 84814 13022 84866
rect 13022 84814 13074 84866
rect 13074 84814 13076 84866
rect 13020 84812 13076 84814
rect 12572 84306 12628 84308
rect 12572 84254 12574 84306
rect 12574 84254 12626 84306
rect 12626 84254 12628 84306
rect 12572 84252 12628 84254
rect 12572 82908 12628 82964
rect 13020 84252 13076 84308
rect 13580 85708 13636 85764
rect 13916 88226 13972 88228
rect 13916 88174 13918 88226
rect 13918 88174 13970 88226
rect 13970 88174 13972 88226
rect 13916 88172 13972 88174
rect 24008 88618 24064 88620
rect 24112 88618 24168 88620
rect 24008 88566 24024 88618
rect 24024 88566 24064 88618
rect 24112 88566 24148 88618
rect 24148 88566 24168 88618
rect 24008 88564 24064 88566
rect 24112 88564 24168 88566
rect 24216 88564 24272 88620
rect 24320 88618 24376 88620
rect 24424 88618 24480 88620
rect 24528 88618 24584 88620
rect 24320 88566 24324 88618
rect 24324 88566 24376 88618
rect 24424 88566 24448 88618
rect 24448 88566 24480 88618
rect 24528 88566 24572 88618
rect 24572 88566 24584 88618
rect 24320 88564 24376 88566
rect 24424 88564 24480 88566
rect 24528 88564 24584 88566
rect 24632 88618 24688 88620
rect 24736 88618 24792 88620
rect 24840 88618 24896 88620
rect 24632 88566 24644 88618
rect 24644 88566 24688 88618
rect 24736 88566 24768 88618
rect 24768 88566 24792 88618
rect 24840 88566 24892 88618
rect 24892 88566 24896 88618
rect 24632 88564 24688 88566
rect 24736 88564 24792 88566
rect 24840 88564 24896 88566
rect 24944 88564 25000 88620
rect 25048 88618 25104 88620
rect 25152 88618 25208 88620
rect 25048 88566 25068 88618
rect 25068 88566 25104 88618
rect 25152 88566 25192 88618
rect 25192 88566 25208 88618
rect 25048 88564 25104 88566
rect 25152 88564 25208 88566
rect 14700 88114 14756 88116
rect 14700 88062 14702 88114
rect 14702 88062 14754 88114
rect 14754 88062 14756 88114
rect 14700 88060 14756 88062
rect 15596 88060 15652 88116
rect 14252 87948 14308 88004
rect 14008 87834 14064 87836
rect 14112 87834 14168 87836
rect 14008 87782 14024 87834
rect 14024 87782 14064 87834
rect 14112 87782 14148 87834
rect 14148 87782 14168 87834
rect 14008 87780 14064 87782
rect 14112 87780 14168 87782
rect 14216 87780 14272 87836
rect 14320 87834 14376 87836
rect 14424 87834 14480 87836
rect 14528 87834 14584 87836
rect 14320 87782 14324 87834
rect 14324 87782 14376 87834
rect 14424 87782 14448 87834
rect 14448 87782 14480 87834
rect 14528 87782 14572 87834
rect 14572 87782 14584 87834
rect 14320 87780 14376 87782
rect 14424 87780 14480 87782
rect 14528 87780 14584 87782
rect 14632 87834 14688 87836
rect 14736 87834 14792 87836
rect 14840 87834 14896 87836
rect 14632 87782 14644 87834
rect 14644 87782 14688 87834
rect 14736 87782 14768 87834
rect 14768 87782 14792 87834
rect 14840 87782 14892 87834
rect 14892 87782 14896 87834
rect 14632 87780 14688 87782
rect 14736 87780 14792 87782
rect 14840 87780 14896 87782
rect 14944 87780 15000 87836
rect 15048 87834 15104 87836
rect 15152 87834 15208 87836
rect 15048 87782 15068 87834
rect 15068 87782 15104 87834
rect 15152 87782 15192 87834
rect 15192 87782 15208 87834
rect 15048 87780 15104 87782
rect 15152 87780 15208 87782
rect 15372 87724 15428 87780
rect 17276 87948 17332 88004
rect 16380 87666 16436 87668
rect 16380 87614 16382 87666
rect 16382 87614 16434 87666
rect 16434 87614 16436 87666
rect 16380 87612 16436 87614
rect 16716 87612 16772 87668
rect 14364 86658 14420 86660
rect 14364 86606 14366 86658
rect 14366 86606 14418 86658
rect 14418 86606 14420 86658
rect 14364 86604 14420 86606
rect 13692 85484 13748 85540
rect 13692 85148 13748 85204
rect 13692 84306 13748 84308
rect 13692 84254 13694 84306
rect 13694 84254 13746 84306
rect 13746 84254 13748 84306
rect 13692 84252 13748 84254
rect 13580 84028 13636 84084
rect 13468 83522 13524 83524
rect 13468 83470 13470 83522
rect 13470 83470 13522 83522
rect 13522 83470 13524 83522
rect 13468 83468 13524 83470
rect 13692 83132 13748 83188
rect 13020 82850 13076 82852
rect 13020 82798 13022 82850
rect 13022 82798 13074 82850
rect 13074 82798 13076 82850
rect 13020 82796 13076 82798
rect 12796 82684 12852 82740
rect 12572 82626 12628 82628
rect 12572 82574 12574 82626
rect 12574 82574 12626 82626
rect 12626 82574 12628 82626
rect 12572 82572 12628 82574
rect 13356 82626 13412 82628
rect 13356 82574 13358 82626
rect 13358 82574 13410 82626
rect 13410 82574 13412 82626
rect 13356 82572 13412 82574
rect 12348 82012 12404 82068
rect 14008 86266 14064 86268
rect 14112 86266 14168 86268
rect 14008 86214 14024 86266
rect 14024 86214 14064 86266
rect 14112 86214 14148 86266
rect 14148 86214 14168 86266
rect 14008 86212 14064 86214
rect 14112 86212 14168 86214
rect 14216 86212 14272 86268
rect 14320 86266 14376 86268
rect 14424 86266 14480 86268
rect 14528 86266 14584 86268
rect 14320 86214 14324 86266
rect 14324 86214 14376 86266
rect 14424 86214 14448 86266
rect 14448 86214 14480 86266
rect 14528 86214 14572 86266
rect 14572 86214 14584 86266
rect 14320 86212 14376 86214
rect 14424 86212 14480 86214
rect 14528 86212 14584 86214
rect 14632 86266 14688 86268
rect 14736 86266 14792 86268
rect 14840 86266 14896 86268
rect 14632 86214 14644 86266
rect 14644 86214 14688 86266
rect 14736 86214 14768 86266
rect 14768 86214 14792 86266
rect 14840 86214 14892 86266
rect 14892 86214 14896 86266
rect 14632 86212 14688 86214
rect 14736 86212 14792 86214
rect 14840 86212 14896 86214
rect 14944 86212 15000 86268
rect 15048 86266 15104 86268
rect 15152 86266 15208 86268
rect 15048 86214 15068 86266
rect 15068 86214 15104 86266
rect 15152 86214 15192 86266
rect 15192 86214 15208 86266
rect 15048 86212 15104 86214
rect 15152 86212 15208 86214
rect 14140 85874 14196 85876
rect 14140 85822 14142 85874
rect 14142 85822 14194 85874
rect 14194 85822 14196 85874
rect 14140 85820 14196 85822
rect 14476 85820 14532 85876
rect 14252 85708 14308 85764
rect 15036 85874 15092 85876
rect 15036 85822 15038 85874
rect 15038 85822 15090 85874
rect 15090 85822 15092 85874
rect 15036 85820 15092 85822
rect 14252 85148 14308 85204
rect 14812 85762 14868 85764
rect 14812 85710 14814 85762
rect 14814 85710 14866 85762
rect 14866 85710 14868 85762
rect 14812 85708 14868 85710
rect 15372 85708 15428 85764
rect 14812 85484 14868 85540
rect 13916 84978 13972 84980
rect 13916 84926 13918 84978
rect 13918 84926 13970 84978
rect 13970 84926 13972 84978
rect 13916 84924 13972 84926
rect 14476 84812 14532 84868
rect 14008 84698 14064 84700
rect 14112 84698 14168 84700
rect 14008 84646 14024 84698
rect 14024 84646 14064 84698
rect 14112 84646 14148 84698
rect 14148 84646 14168 84698
rect 14008 84644 14064 84646
rect 14112 84644 14168 84646
rect 14216 84644 14272 84700
rect 14320 84698 14376 84700
rect 14424 84698 14480 84700
rect 14528 84698 14584 84700
rect 14320 84646 14324 84698
rect 14324 84646 14376 84698
rect 14424 84646 14448 84698
rect 14448 84646 14480 84698
rect 14528 84646 14572 84698
rect 14572 84646 14584 84698
rect 14320 84644 14376 84646
rect 14424 84644 14480 84646
rect 14528 84644 14584 84646
rect 14632 84698 14688 84700
rect 14736 84698 14792 84700
rect 14840 84698 14896 84700
rect 14632 84646 14644 84698
rect 14644 84646 14688 84698
rect 14736 84646 14768 84698
rect 14768 84646 14792 84698
rect 14840 84646 14892 84698
rect 14892 84646 14896 84698
rect 14632 84644 14688 84646
rect 14736 84644 14792 84646
rect 14840 84644 14896 84646
rect 14944 84644 15000 84700
rect 15048 84698 15104 84700
rect 15152 84698 15208 84700
rect 15048 84646 15068 84698
rect 15068 84646 15104 84698
rect 15152 84646 15192 84698
rect 15192 84646 15208 84698
rect 15048 84644 15104 84646
rect 15152 84644 15208 84646
rect 14588 84476 14644 84532
rect 14476 84418 14532 84420
rect 14476 84366 14478 84418
rect 14478 84366 14530 84418
rect 14530 84366 14532 84418
rect 14476 84364 14532 84366
rect 16044 86604 16100 86660
rect 16156 85762 16212 85764
rect 16156 85710 16158 85762
rect 16158 85710 16210 85762
rect 16210 85710 16212 85762
rect 16156 85708 16212 85710
rect 16604 85986 16660 85988
rect 16604 85934 16606 85986
rect 16606 85934 16658 85986
rect 16658 85934 16660 85986
rect 16604 85932 16660 85934
rect 15596 84476 15652 84532
rect 15036 84418 15092 84420
rect 15036 84366 15038 84418
rect 15038 84366 15090 84418
rect 15090 84366 15092 84418
rect 15036 84364 15092 84366
rect 14476 83356 14532 83412
rect 15260 83356 15316 83412
rect 14028 83244 14084 83300
rect 14008 83130 14064 83132
rect 14112 83130 14168 83132
rect 14008 83078 14024 83130
rect 14024 83078 14064 83130
rect 14112 83078 14148 83130
rect 14148 83078 14168 83130
rect 14008 83076 14064 83078
rect 14112 83076 14168 83078
rect 14216 83076 14272 83132
rect 14320 83130 14376 83132
rect 14424 83130 14480 83132
rect 14528 83130 14584 83132
rect 14320 83078 14324 83130
rect 14324 83078 14376 83130
rect 14424 83078 14448 83130
rect 14448 83078 14480 83130
rect 14528 83078 14572 83130
rect 14572 83078 14584 83130
rect 14320 83076 14376 83078
rect 14424 83076 14480 83078
rect 14528 83076 14584 83078
rect 14632 83130 14688 83132
rect 14736 83130 14792 83132
rect 14840 83130 14896 83132
rect 14632 83078 14644 83130
rect 14644 83078 14688 83130
rect 14736 83078 14768 83130
rect 14768 83078 14792 83130
rect 14840 83078 14892 83130
rect 14892 83078 14896 83130
rect 14632 83076 14688 83078
rect 14736 83076 14792 83078
rect 14840 83076 14896 83078
rect 14944 83076 15000 83132
rect 15048 83130 15104 83132
rect 15152 83130 15208 83132
rect 15048 83078 15068 83130
rect 15068 83078 15104 83130
rect 15152 83078 15192 83130
rect 15192 83078 15208 83130
rect 15048 83076 15104 83078
rect 15152 83076 15208 83078
rect 15148 82908 15204 82964
rect 14140 82738 14196 82740
rect 14140 82686 14142 82738
rect 14142 82686 14194 82738
rect 14194 82686 14196 82738
rect 14140 82684 14196 82686
rect 13468 81788 13524 81844
rect 12124 81058 12180 81060
rect 12124 81006 12126 81058
rect 12126 81006 12178 81058
rect 12178 81006 12180 81058
rect 12124 81004 12180 81006
rect 12796 80946 12852 80948
rect 12796 80894 12798 80946
rect 12798 80894 12850 80946
rect 12850 80894 12852 80946
rect 12796 80892 12852 80894
rect 11900 80386 11956 80388
rect 11900 80334 11902 80386
rect 11902 80334 11954 80386
rect 11954 80334 11956 80386
rect 11900 80332 11956 80334
rect 11228 79212 11284 79268
rect 11676 80162 11732 80164
rect 11676 80110 11678 80162
rect 11678 80110 11730 80162
rect 11730 80110 11732 80162
rect 11676 80108 11732 80110
rect 11900 79772 11956 79828
rect 12908 80162 12964 80164
rect 12908 80110 12910 80162
rect 12910 80110 12962 80162
rect 12962 80110 12964 80162
rect 12908 80108 12964 80110
rect 13468 80108 13524 80164
rect 11452 78594 11508 78596
rect 11452 78542 11454 78594
rect 11454 78542 11506 78594
rect 11506 78542 11508 78594
rect 11452 78540 11508 78542
rect 11340 77922 11396 77924
rect 11340 77870 11342 77922
rect 11342 77870 11394 77922
rect 11394 77870 11396 77922
rect 11340 77868 11396 77870
rect 11116 76466 11172 76468
rect 11116 76414 11118 76466
rect 11118 76414 11170 76466
rect 11170 76414 11172 76466
rect 11116 76412 11172 76414
rect 10892 75682 10948 75684
rect 10892 75630 10894 75682
rect 10894 75630 10946 75682
rect 10946 75630 10948 75682
rect 10892 75628 10948 75630
rect 10780 75292 10836 75348
rect 9660 73554 9716 73556
rect 9660 73502 9662 73554
rect 9662 73502 9714 73554
rect 9714 73502 9716 73554
rect 9660 73500 9716 73502
rect 9548 73164 9604 73220
rect 9996 75010 10052 75012
rect 9996 74958 9998 75010
rect 9998 74958 10050 75010
rect 10050 74958 10052 75010
rect 9996 74956 10052 74958
rect 9884 73164 9940 73220
rect 10108 73276 10164 73332
rect 9772 72492 9828 72548
rect 10892 74956 10948 75012
rect 11004 73330 11060 73332
rect 11004 73278 11006 73330
rect 11006 73278 11058 73330
rect 11058 73278 11060 73330
rect 11004 73276 11060 73278
rect 10556 73218 10612 73220
rect 10556 73166 10558 73218
rect 10558 73166 10610 73218
rect 10610 73166 10612 73218
rect 10556 73164 10612 73166
rect 9884 72380 9940 72436
rect 9660 70306 9716 70308
rect 9660 70254 9662 70306
rect 9662 70254 9714 70306
rect 9714 70254 9716 70306
rect 9660 70252 9716 70254
rect 9436 70194 9492 70196
rect 9436 70142 9438 70194
rect 9438 70142 9490 70194
rect 9490 70142 9492 70194
rect 9436 70140 9492 70142
rect 9772 70028 9828 70084
rect 10556 70252 10612 70308
rect 10332 70082 10388 70084
rect 10332 70030 10334 70082
rect 10334 70030 10386 70082
rect 10386 70030 10388 70082
rect 10332 70028 10388 70030
rect 11228 74226 11284 74228
rect 11228 74174 11230 74226
rect 11230 74174 11282 74226
rect 11282 74174 11284 74226
rect 11228 74172 11284 74174
rect 11676 76972 11732 77028
rect 12012 78930 12068 78932
rect 12012 78878 12014 78930
rect 12014 78878 12066 78930
rect 12066 78878 12068 78930
rect 12012 78876 12068 78878
rect 12908 78204 12964 78260
rect 12460 77868 12516 77924
rect 12012 76972 12068 77028
rect 13020 77308 13076 77364
rect 12572 77196 12628 77252
rect 12460 76636 12516 76692
rect 12012 76524 12068 76580
rect 12460 76300 12516 76356
rect 12348 75740 12404 75796
rect 12236 74898 12292 74900
rect 12236 74846 12238 74898
rect 12238 74846 12290 74898
rect 12290 74846 12292 74898
rect 12236 74844 12292 74846
rect 13356 79100 13412 79156
rect 13244 78876 13300 78932
rect 12796 75740 12852 75796
rect 12684 75068 12740 75124
rect 12572 74844 12628 74900
rect 11340 73836 11396 73892
rect 11340 73276 11396 73332
rect 11676 73164 11732 73220
rect 11116 70754 11172 70756
rect 11116 70702 11118 70754
rect 11118 70702 11170 70754
rect 11170 70702 11172 70754
rect 11116 70700 11172 70702
rect 10444 69132 10500 69188
rect 9884 67452 9940 67508
rect 9660 67228 9716 67284
rect 9324 65436 9380 65492
rect 8988 65212 9044 65268
rect 8988 64146 9044 64148
rect 8988 64094 8990 64146
rect 8990 64094 9042 64146
rect 9042 64094 9044 64146
rect 8988 64092 9044 64094
rect 9212 64988 9268 65044
rect 9884 66108 9940 66164
rect 9212 63308 9268 63364
rect 8764 63196 8820 63252
rect 8876 62412 8932 62468
rect 8764 58210 8820 58212
rect 8764 58158 8766 58210
rect 8766 58158 8818 58210
rect 8818 58158 8820 58210
rect 8764 58156 8820 58158
rect 8764 56028 8820 56084
rect 8764 55468 8820 55524
rect 9548 63138 9604 63140
rect 9548 63086 9550 63138
rect 9550 63086 9602 63138
rect 9602 63086 9604 63138
rect 9548 63084 9604 63086
rect 9772 62300 9828 62356
rect 10892 68514 10948 68516
rect 10892 68462 10894 68514
rect 10894 68462 10946 68514
rect 10946 68462 10948 68514
rect 10892 68460 10948 68462
rect 10780 66780 10836 66836
rect 10220 66386 10276 66388
rect 10220 66334 10222 66386
rect 10222 66334 10274 66386
rect 10274 66334 10276 66386
rect 10220 66332 10276 66334
rect 9996 65660 10052 65716
rect 9996 65490 10052 65492
rect 9996 65438 9998 65490
rect 9998 65438 10050 65490
rect 10050 65438 10052 65490
rect 9996 65436 10052 65438
rect 10220 65436 10276 65492
rect 10108 64988 10164 65044
rect 9884 63084 9940 63140
rect 10108 63196 10164 63252
rect 8988 60674 9044 60676
rect 8988 60622 8990 60674
rect 8990 60622 9042 60674
rect 9042 60622 9044 60674
rect 8988 60620 9044 60622
rect 9100 60508 9156 60564
rect 9884 61346 9940 61348
rect 9884 61294 9886 61346
rect 9886 61294 9938 61346
rect 9938 61294 9940 61346
rect 9884 61292 9940 61294
rect 9660 60060 9716 60116
rect 9324 59276 9380 59332
rect 9100 57538 9156 57540
rect 9100 57486 9102 57538
rect 9102 57486 9154 57538
rect 9154 57486 9156 57538
rect 9100 57484 9156 57486
rect 8988 54626 9044 54628
rect 8988 54574 8990 54626
rect 8990 54574 9042 54626
rect 9042 54574 9044 54626
rect 8988 54572 9044 54574
rect 8876 54460 8932 54516
rect 9212 54572 9268 54628
rect 9436 58156 9492 58212
rect 9436 57708 9492 57764
rect 9660 57148 9716 57204
rect 9660 56924 9716 56980
rect 9436 52946 9492 52948
rect 9436 52894 9438 52946
rect 9438 52894 9490 52946
rect 9490 52894 9492 52946
rect 9436 52892 9492 52894
rect 9212 51660 9268 51716
rect 8652 50034 8708 50036
rect 8652 49982 8654 50034
rect 8654 49982 8706 50034
rect 8706 49982 8708 50034
rect 8652 49980 8708 49982
rect 8540 49586 8596 49588
rect 8540 49534 8542 49586
rect 8542 49534 8594 49586
rect 8594 49534 8596 49586
rect 8540 49532 8596 49534
rect 8540 48188 8596 48244
rect 7084 47180 7140 47236
rect 6860 46732 6916 46788
rect 7420 46844 7476 46900
rect 6748 44434 6804 44436
rect 6748 44382 6750 44434
rect 6750 44382 6802 44434
rect 6802 44382 6804 44434
rect 6748 44380 6804 44382
rect 6524 44044 6580 44100
rect 6300 42812 6356 42868
rect 6748 42642 6804 42644
rect 6748 42590 6750 42642
rect 6750 42590 6802 42642
rect 6802 42590 6804 42642
rect 6748 42588 6804 42590
rect 5740 40684 5796 40740
rect 5740 40514 5796 40516
rect 5740 40462 5742 40514
rect 5742 40462 5794 40514
rect 5794 40462 5796 40514
rect 5740 40460 5796 40462
rect 5404 38892 5460 38948
rect 4620 38834 4676 38836
rect 4620 38782 4622 38834
rect 4622 38782 4674 38834
rect 4674 38782 4676 38834
rect 4620 38780 4676 38782
rect 5740 38780 5796 38836
rect 6748 40572 6804 40628
rect 6636 40514 6692 40516
rect 6636 40462 6638 40514
rect 6638 40462 6690 40514
rect 6690 40462 6692 40514
rect 6636 40460 6692 40462
rect 6188 39564 6244 39620
rect 6076 39004 6132 39060
rect 6188 39340 6244 39396
rect 4008 38442 4064 38444
rect 4112 38442 4168 38444
rect 4008 38390 4024 38442
rect 4024 38390 4064 38442
rect 4112 38390 4148 38442
rect 4148 38390 4168 38442
rect 4008 38388 4064 38390
rect 4112 38388 4168 38390
rect 4216 38388 4272 38444
rect 4320 38442 4376 38444
rect 4424 38442 4480 38444
rect 4528 38442 4584 38444
rect 4320 38390 4324 38442
rect 4324 38390 4376 38442
rect 4424 38390 4448 38442
rect 4448 38390 4480 38442
rect 4528 38390 4572 38442
rect 4572 38390 4584 38442
rect 4320 38388 4376 38390
rect 4424 38388 4480 38390
rect 4528 38388 4584 38390
rect 4632 38442 4688 38444
rect 4736 38442 4792 38444
rect 4840 38442 4896 38444
rect 4632 38390 4644 38442
rect 4644 38390 4688 38442
rect 4736 38390 4768 38442
rect 4768 38390 4792 38442
rect 4840 38390 4892 38442
rect 4892 38390 4896 38442
rect 4632 38388 4688 38390
rect 4736 38388 4792 38390
rect 4840 38388 4896 38390
rect 4944 38388 5000 38444
rect 5048 38442 5104 38444
rect 5152 38442 5208 38444
rect 5048 38390 5068 38442
rect 5068 38390 5104 38442
rect 5152 38390 5192 38442
rect 5192 38390 5208 38442
rect 5048 38388 5104 38390
rect 5152 38388 5208 38390
rect 4008 36874 4064 36876
rect 4112 36874 4168 36876
rect 4008 36822 4024 36874
rect 4024 36822 4064 36874
rect 4112 36822 4148 36874
rect 4148 36822 4168 36874
rect 4008 36820 4064 36822
rect 4112 36820 4168 36822
rect 4216 36820 4272 36876
rect 4320 36874 4376 36876
rect 4424 36874 4480 36876
rect 4528 36874 4584 36876
rect 4320 36822 4324 36874
rect 4324 36822 4376 36874
rect 4424 36822 4448 36874
rect 4448 36822 4480 36874
rect 4528 36822 4572 36874
rect 4572 36822 4584 36874
rect 4320 36820 4376 36822
rect 4424 36820 4480 36822
rect 4528 36820 4584 36822
rect 4632 36874 4688 36876
rect 4736 36874 4792 36876
rect 4840 36874 4896 36876
rect 4632 36822 4644 36874
rect 4644 36822 4688 36874
rect 4736 36822 4768 36874
rect 4768 36822 4792 36874
rect 4840 36822 4892 36874
rect 4892 36822 4896 36874
rect 4632 36820 4688 36822
rect 4736 36820 4792 36822
rect 4840 36820 4896 36822
rect 4944 36820 5000 36876
rect 5048 36874 5104 36876
rect 5152 36874 5208 36876
rect 5048 36822 5068 36874
rect 5068 36822 5104 36874
rect 5152 36822 5192 36874
rect 5192 36822 5208 36874
rect 5048 36820 5104 36822
rect 5152 36820 5208 36822
rect 4060 36258 4116 36260
rect 4060 36206 4062 36258
rect 4062 36206 4114 36258
rect 4114 36206 4116 36258
rect 4060 36204 4116 36206
rect 5180 36370 5236 36372
rect 5180 36318 5182 36370
rect 5182 36318 5234 36370
rect 5234 36318 5236 36370
rect 5180 36316 5236 36318
rect 5852 36370 5908 36372
rect 5852 36318 5854 36370
rect 5854 36318 5906 36370
rect 5906 36318 5908 36370
rect 5852 36316 5908 36318
rect 4956 36258 5012 36260
rect 4956 36206 4958 36258
rect 4958 36206 5010 36258
rect 5010 36206 5012 36258
rect 4956 36204 5012 36206
rect 4844 35980 4900 36036
rect 4956 35922 5012 35924
rect 4956 35870 4958 35922
rect 4958 35870 5010 35922
rect 5010 35870 5012 35922
rect 4956 35868 5012 35870
rect 5292 35868 5348 35924
rect 3612 32060 3668 32116
rect 2156 31388 2212 31444
rect 2828 31388 2884 31444
rect 3164 31106 3220 31108
rect 3164 31054 3166 31106
rect 3166 31054 3218 31106
rect 3218 31054 3220 31106
rect 3164 31052 3220 31054
rect 3164 30716 3220 30772
rect 2828 30380 2884 30436
rect 2604 30156 2660 30212
rect 4008 35306 4064 35308
rect 4112 35306 4168 35308
rect 4008 35254 4024 35306
rect 4024 35254 4064 35306
rect 4112 35254 4148 35306
rect 4148 35254 4168 35306
rect 4008 35252 4064 35254
rect 4112 35252 4168 35254
rect 4216 35252 4272 35308
rect 4320 35306 4376 35308
rect 4424 35306 4480 35308
rect 4528 35306 4584 35308
rect 4320 35254 4324 35306
rect 4324 35254 4376 35306
rect 4424 35254 4448 35306
rect 4448 35254 4480 35306
rect 4528 35254 4572 35306
rect 4572 35254 4584 35306
rect 4320 35252 4376 35254
rect 4424 35252 4480 35254
rect 4528 35252 4584 35254
rect 4632 35306 4688 35308
rect 4736 35306 4792 35308
rect 4840 35306 4896 35308
rect 4632 35254 4644 35306
rect 4644 35254 4688 35306
rect 4736 35254 4768 35306
rect 4768 35254 4792 35306
rect 4840 35254 4892 35306
rect 4892 35254 4896 35306
rect 4632 35252 4688 35254
rect 4736 35252 4792 35254
rect 4840 35252 4896 35254
rect 4944 35252 5000 35308
rect 5048 35306 5104 35308
rect 5152 35306 5208 35308
rect 5048 35254 5068 35306
rect 5068 35254 5104 35306
rect 5152 35254 5192 35306
rect 5192 35254 5208 35306
rect 5048 35252 5104 35254
rect 5152 35252 5208 35254
rect 4732 35084 4788 35140
rect 4620 34972 4676 35028
rect 4172 34914 4228 34916
rect 4172 34862 4174 34914
rect 4174 34862 4226 34914
rect 4226 34862 4228 34914
rect 4172 34860 4228 34862
rect 3836 34690 3892 34692
rect 3836 34638 3838 34690
rect 3838 34638 3890 34690
rect 3890 34638 3892 34690
rect 3836 34636 3892 34638
rect 5292 34972 5348 35028
rect 4956 34802 5012 34804
rect 4956 34750 4958 34802
rect 4958 34750 5010 34802
rect 5010 34750 5012 34802
rect 4956 34748 5012 34750
rect 5404 35420 5460 35476
rect 5292 34748 5348 34804
rect 4008 33738 4064 33740
rect 4112 33738 4168 33740
rect 4008 33686 4024 33738
rect 4024 33686 4064 33738
rect 4112 33686 4148 33738
rect 4148 33686 4168 33738
rect 4008 33684 4064 33686
rect 4112 33684 4168 33686
rect 4216 33684 4272 33740
rect 4320 33738 4376 33740
rect 4424 33738 4480 33740
rect 4528 33738 4584 33740
rect 4320 33686 4324 33738
rect 4324 33686 4376 33738
rect 4424 33686 4448 33738
rect 4448 33686 4480 33738
rect 4528 33686 4572 33738
rect 4572 33686 4584 33738
rect 4320 33684 4376 33686
rect 4424 33684 4480 33686
rect 4528 33684 4584 33686
rect 4632 33738 4688 33740
rect 4736 33738 4792 33740
rect 4840 33738 4896 33740
rect 4632 33686 4644 33738
rect 4644 33686 4688 33738
rect 4736 33686 4768 33738
rect 4768 33686 4792 33738
rect 4840 33686 4892 33738
rect 4892 33686 4896 33738
rect 4632 33684 4688 33686
rect 4736 33684 4792 33686
rect 4840 33684 4896 33686
rect 4944 33684 5000 33740
rect 5048 33738 5104 33740
rect 5152 33738 5208 33740
rect 5048 33686 5068 33738
rect 5068 33686 5104 33738
rect 5152 33686 5192 33738
rect 5192 33686 5208 33738
rect 5048 33684 5104 33686
rect 5152 33684 5208 33686
rect 5292 33516 5348 33572
rect 5068 33458 5124 33460
rect 5068 33406 5070 33458
rect 5070 33406 5122 33458
rect 5122 33406 5124 33458
rect 5068 33404 5124 33406
rect 4172 33122 4228 33124
rect 4172 33070 4174 33122
rect 4174 33070 4226 33122
rect 4226 33070 4228 33122
rect 4172 33068 4228 33070
rect 5180 33292 5236 33348
rect 5180 32956 5236 33012
rect 4732 32786 4788 32788
rect 4732 32734 4734 32786
rect 4734 32734 4786 32786
rect 4786 32734 4788 32786
rect 4732 32732 4788 32734
rect 3836 32396 3892 32452
rect 6524 39618 6580 39620
rect 6524 39566 6526 39618
rect 6526 39566 6578 39618
rect 6578 39566 6580 39618
rect 6524 39564 6580 39566
rect 6188 36204 6244 36260
rect 6300 35922 6356 35924
rect 6300 35870 6302 35922
rect 6302 35870 6354 35922
rect 6354 35870 6356 35922
rect 6300 35868 6356 35870
rect 5628 34860 5684 34916
rect 5740 34690 5796 34692
rect 5740 34638 5742 34690
rect 5742 34638 5794 34690
rect 5794 34638 5796 34690
rect 5740 34636 5796 34638
rect 5516 33964 5572 34020
rect 6076 34802 6132 34804
rect 6076 34750 6078 34802
rect 6078 34750 6130 34802
rect 6130 34750 6132 34802
rect 6076 34748 6132 34750
rect 6188 34690 6244 34692
rect 6188 34638 6190 34690
rect 6190 34638 6242 34690
rect 6242 34638 6244 34690
rect 6188 34636 6244 34638
rect 6188 34300 6244 34356
rect 5516 32396 5572 32452
rect 4008 32170 4064 32172
rect 4112 32170 4168 32172
rect 4008 32118 4024 32170
rect 4024 32118 4064 32170
rect 4112 32118 4148 32170
rect 4148 32118 4168 32170
rect 4008 32116 4064 32118
rect 4112 32116 4168 32118
rect 4216 32116 4272 32172
rect 4320 32170 4376 32172
rect 4424 32170 4480 32172
rect 4528 32170 4584 32172
rect 4320 32118 4324 32170
rect 4324 32118 4376 32170
rect 4424 32118 4448 32170
rect 4448 32118 4480 32170
rect 4528 32118 4572 32170
rect 4572 32118 4584 32170
rect 4320 32116 4376 32118
rect 4424 32116 4480 32118
rect 4528 32116 4584 32118
rect 4632 32170 4688 32172
rect 4736 32170 4792 32172
rect 4840 32170 4896 32172
rect 4632 32118 4644 32170
rect 4644 32118 4688 32170
rect 4736 32118 4768 32170
rect 4768 32118 4792 32170
rect 4840 32118 4892 32170
rect 4892 32118 4896 32170
rect 4632 32116 4688 32118
rect 4736 32116 4792 32118
rect 4840 32116 4896 32118
rect 4944 32116 5000 32172
rect 5048 32170 5104 32172
rect 5152 32170 5208 32172
rect 5048 32118 5068 32170
rect 5068 32118 5104 32170
rect 5152 32118 5192 32170
rect 5192 32118 5208 32170
rect 5048 32116 5104 32118
rect 5152 32116 5208 32118
rect 5740 32956 5796 33012
rect 5404 31836 5460 31892
rect 5852 31836 5908 31892
rect 5964 33068 6020 33124
rect 5068 31778 5124 31780
rect 5068 31726 5070 31778
rect 5070 31726 5122 31778
rect 5122 31726 5124 31778
rect 5068 31724 5124 31726
rect 4508 30940 4564 30996
rect 4008 30602 4064 30604
rect 4112 30602 4168 30604
rect 4008 30550 4024 30602
rect 4024 30550 4064 30602
rect 4112 30550 4148 30602
rect 4148 30550 4168 30602
rect 4008 30548 4064 30550
rect 4112 30548 4168 30550
rect 4216 30548 4272 30604
rect 4320 30602 4376 30604
rect 4424 30602 4480 30604
rect 4528 30602 4584 30604
rect 4320 30550 4324 30602
rect 4324 30550 4376 30602
rect 4424 30550 4448 30602
rect 4448 30550 4480 30602
rect 4528 30550 4572 30602
rect 4572 30550 4584 30602
rect 4320 30548 4376 30550
rect 4424 30548 4480 30550
rect 4528 30548 4584 30550
rect 4632 30602 4688 30604
rect 4736 30602 4792 30604
rect 4840 30602 4896 30604
rect 4632 30550 4644 30602
rect 4644 30550 4688 30602
rect 4736 30550 4768 30602
rect 4768 30550 4792 30602
rect 4840 30550 4892 30602
rect 4892 30550 4896 30602
rect 4632 30548 4688 30550
rect 4736 30548 4792 30550
rect 4840 30548 4896 30550
rect 4944 30548 5000 30604
rect 5048 30602 5104 30604
rect 5152 30602 5208 30604
rect 5048 30550 5068 30602
rect 5068 30550 5104 30602
rect 5152 30550 5192 30602
rect 5192 30550 5208 30602
rect 5048 30548 5104 30550
rect 5152 30548 5208 30550
rect 3724 30156 3780 30212
rect 3948 30098 4004 30100
rect 3948 30046 3950 30098
rect 3950 30046 4002 30098
rect 4002 30046 4004 30098
rect 3948 30044 4004 30046
rect 2156 29820 2212 29876
rect 2044 29484 2100 29540
rect 2156 29148 2212 29204
rect 2492 28924 2548 28980
rect 1596 28476 1652 28532
rect 1820 27916 1876 27972
rect 1708 25788 1764 25844
rect 3276 29932 3332 29988
rect 3164 28866 3220 28868
rect 3164 28814 3166 28866
rect 3166 28814 3218 28866
rect 3218 28814 3220 28866
rect 3164 28812 3220 28814
rect 2828 28588 2884 28644
rect 3724 29986 3780 29988
rect 3724 29934 3726 29986
rect 3726 29934 3778 29986
rect 3778 29934 3780 29986
rect 3724 29932 3780 29934
rect 4732 30156 4788 30212
rect 4060 29820 4116 29876
rect 3948 29596 4004 29652
rect 3836 29372 3892 29428
rect 3500 29260 3556 29316
rect 2940 28364 2996 28420
rect 3388 27244 3444 27300
rect 4620 29484 4676 29540
rect 4508 29372 4564 29428
rect 4732 29260 4788 29316
rect 3948 29148 4004 29204
rect 4844 29148 4900 29204
rect 5180 30268 5236 30324
rect 5516 30994 5572 30996
rect 5516 30942 5518 30994
rect 5518 30942 5570 30994
rect 5570 30942 5572 30994
rect 5516 30940 5572 30942
rect 5852 30210 5908 30212
rect 5852 30158 5854 30210
rect 5854 30158 5906 30210
rect 5906 30158 5908 30210
rect 5852 30156 5908 30158
rect 4008 29034 4064 29036
rect 4112 29034 4168 29036
rect 4008 28982 4024 29034
rect 4024 28982 4064 29034
rect 4112 28982 4148 29034
rect 4148 28982 4168 29034
rect 4008 28980 4064 28982
rect 4112 28980 4168 28982
rect 4216 28980 4272 29036
rect 4320 29034 4376 29036
rect 4424 29034 4480 29036
rect 4528 29034 4584 29036
rect 4320 28982 4324 29034
rect 4324 28982 4376 29034
rect 4424 28982 4448 29034
rect 4448 28982 4480 29034
rect 4528 28982 4572 29034
rect 4572 28982 4584 29034
rect 4320 28980 4376 28982
rect 4424 28980 4480 28982
rect 4528 28980 4584 28982
rect 4632 29034 4688 29036
rect 4736 29034 4792 29036
rect 4840 29034 4896 29036
rect 4632 28982 4644 29034
rect 4644 28982 4688 29034
rect 4736 28982 4768 29034
rect 4768 28982 4792 29034
rect 4840 28982 4892 29034
rect 4892 28982 4896 29034
rect 4632 28980 4688 28982
rect 4736 28980 4792 28982
rect 4840 28980 4896 28982
rect 4944 28980 5000 29036
rect 5048 29034 5104 29036
rect 5152 29034 5208 29036
rect 5048 28982 5068 29034
rect 5068 28982 5104 29034
rect 5152 28982 5192 29034
rect 5192 28982 5208 29034
rect 5048 28980 5104 28982
rect 5152 28980 5208 28982
rect 3836 28588 3892 28644
rect 3948 28530 4004 28532
rect 3948 28478 3950 28530
rect 3950 28478 4002 28530
rect 4002 28478 4004 28530
rect 3948 28476 4004 28478
rect 3836 28364 3892 28420
rect 4172 28812 4228 28868
rect 4732 28812 4788 28868
rect 4508 28642 4564 28644
rect 4508 28590 4510 28642
rect 4510 28590 4562 28642
rect 4562 28590 4564 28642
rect 4508 28588 4564 28590
rect 4844 28530 4900 28532
rect 4844 28478 4846 28530
rect 4846 28478 4898 28530
rect 4898 28478 4900 28530
rect 4844 28476 4900 28478
rect 5180 28476 5236 28532
rect 4956 27580 5012 27636
rect 5516 28364 5572 28420
rect 5516 28140 5572 28196
rect 4008 27466 4064 27468
rect 4112 27466 4168 27468
rect 4008 27414 4024 27466
rect 4024 27414 4064 27466
rect 4112 27414 4148 27466
rect 4148 27414 4168 27466
rect 4008 27412 4064 27414
rect 4112 27412 4168 27414
rect 4216 27412 4272 27468
rect 4320 27466 4376 27468
rect 4424 27466 4480 27468
rect 4528 27466 4584 27468
rect 4320 27414 4324 27466
rect 4324 27414 4376 27466
rect 4424 27414 4448 27466
rect 4448 27414 4480 27466
rect 4528 27414 4572 27466
rect 4572 27414 4584 27466
rect 4320 27412 4376 27414
rect 4424 27412 4480 27414
rect 4528 27412 4584 27414
rect 4632 27466 4688 27468
rect 4736 27466 4792 27468
rect 4840 27466 4896 27468
rect 4632 27414 4644 27466
rect 4644 27414 4688 27466
rect 4736 27414 4768 27466
rect 4768 27414 4792 27466
rect 4840 27414 4892 27466
rect 4892 27414 4896 27466
rect 4632 27412 4688 27414
rect 4736 27412 4792 27414
rect 4840 27412 4896 27414
rect 4944 27412 5000 27468
rect 5048 27466 5104 27468
rect 5152 27466 5208 27468
rect 5048 27414 5068 27466
rect 5068 27414 5104 27466
rect 5152 27414 5192 27466
rect 5192 27414 5208 27466
rect 5048 27412 5104 27414
rect 5152 27412 5208 27414
rect 2940 27020 2996 27076
rect 2604 26460 2660 26516
rect 3164 26796 3220 26852
rect 3052 26012 3108 26068
rect 2044 24556 2100 24612
rect 1708 22876 1764 22932
rect 1820 23436 1876 23492
rect 1708 22428 1764 22484
rect 1932 23266 1988 23268
rect 1932 23214 1934 23266
rect 1934 23214 1986 23266
rect 1986 23214 1988 23266
rect 1932 23212 1988 23214
rect 1708 21586 1764 21588
rect 1708 21534 1710 21586
rect 1710 21534 1762 21586
rect 1762 21534 1764 21586
rect 1708 21532 1764 21534
rect 1820 21308 1876 21364
rect 2492 24610 2548 24612
rect 2492 24558 2494 24610
rect 2494 24558 2546 24610
rect 2546 24558 2548 24610
rect 2492 24556 2548 24558
rect 2940 24668 2996 24724
rect 2716 23772 2772 23828
rect 2156 23548 2212 23604
rect 2268 23100 2324 23156
rect 2268 22876 2324 22932
rect 2380 22764 2436 22820
rect 2492 22540 2548 22596
rect 2828 23436 2884 23492
rect 2492 22316 2548 22372
rect 2828 22316 2884 22372
rect 2604 21308 2660 21364
rect 2492 20188 2548 20244
rect 2492 19180 2548 19236
rect 2828 19180 2884 19236
rect 4284 27244 4340 27300
rect 3948 26962 4004 26964
rect 3948 26910 3950 26962
rect 3950 26910 4002 26962
rect 4002 26910 4004 26962
rect 3948 26908 4004 26910
rect 3612 26572 3668 26628
rect 3164 25452 3220 25508
rect 3276 26236 3332 26292
rect 3164 24668 3220 24724
rect 3500 25676 3556 25732
rect 3388 23714 3444 23716
rect 3388 23662 3390 23714
rect 3390 23662 3442 23714
rect 3442 23662 3444 23714
rect 3388 23660 3444 23662
rect 3276 23492 3332 23548
rect 3388 23042 3444 23044
rect 3388 22990 3390 23042
rect 3390 22990 3442 23042
rect 3442 22990 3444 23042
rect 3388 22988 3444 22990
rect 3836 26514 3892 26516
rect 3836 26462 3838 26514
rect 3838 26462 3890 26514
rect 3890 26462 3892 26514
rect 3836 26460 3892 26462
rect 4732 27298 4788 27300
rect 4732 27246 4734 27298
rect 4734 27246 4786 27298
rect 4786 27246 4788 27298
rect 4732 27244 4788 27246
rect 5068 27186 5124 27188
rect 5068 27134 5070 27186
rect 5070 27134 5122 27186
rect 5122 27134 5124 27186
rect 5068 27132 5124 27134
rect 4508 26908 4564 26964
rect 4844 27020 4900 27076
rect 5292 27020 5348 27076
rect 4620 26290 4676 26292
rect 4620 26238 4622 26290
rect 4622 26238 4674 26290
rect 4674 26238 4676 26290
rect 4620 26236 4676 26238
rect 5292 26460 5348 26516
rect 3612 23212 3668 23268
rect 3164 20690 3220 20692
rect 3164 20638 3166 20690
rect 3166 20638 3218 20690
rect 3218 20638 3220 20690
rect 3164 20636 3220 20638
rect 3612 19234 3668 19236
rect 3612 19182 3614 19234
rect 3614 19182 3666 19234
rect 3666 19182 3668 19234
rect 3612 19180 3668 19182
rect 3276 17836 3332 17892
rect 2492 17106 2548 17108
rect 2492 17054 2494 17106
rect 2494 17054 2546 17106
rect 2546 17054 2548 17106
rect 2492 17052 2548 17054
rect 1932 16994 1988 16996
rect 1932 16942 1934 16994
rect 1934 16942 1986 16994
rect 1986 16942 1988 16994
rect 1932 16940 1988 16942
rect 1708 14588 1764 14644
rect 1820 15148 1876 15204
rect 2940 16940 2996 16996
rect 2604 16044 2660 16100
rect 3276 16716 3332 16772
rect 4956 26066 5012 26068
rect 4956 26014 4958 26066
rect 4958 26014 5010 26066
rect 5010 26014 5012 26066
rect 4956 26012 5012 26014
rect 4008 25898 4064 25900
rect 4112 25898 4168 25900
rect 4008 25846 4024 25898
rect 4024 25846 4064 25898
rect 4112 25846 4148 25898
rect 4148 25846 4168 25898
rect 4008 25844 4064 25846
rect 4112 25844 4168 25846
rect 4216 25844 4272 25900
rect 4320 25898 4376 25900
rect 4424 25898 4480 25900
rect 4528 25898 4584 25900
rect 4320 25846 4324 25898
rect 4324 25846 4376 25898
rect 4424 25846 4448 25898
rect 4448 25846 4480 25898
rect 4528 25846 4572 25898
rect 4572 25846 4584 25898
rect 4320 25844 4376 25846
rect 4424 25844 4480 25846
rect 4528 25844 4584 25846
rect 4632 25898 4688 25900
rect 4736 25898 4792 25900
rect 4840 25898 4896 25900
rect 4632 25846 4644 25898
rect 4644 25846 4688 25898
rect 4736 25846 4768 25898
rect 4768 25846 4792 25898
rect 4840 25846 4892 25898
rect 4892 25846 4896 25898
rect 4632 25844 4688 25846
rect 4736 25844 4792 25846
rect 4840 25844 4896 25846
rect 4944 25844 5000 25900
rect 5048 25898 5104 25900
rect 5152 25898 5208 25900
rect 5048 25846 5068 25898
rect 5068 25846 5104 25898
rect 5152 25846 5192 25898
rect 5192 25846 5208 25898
rect 5048 25844 5104 25846
rect 5152 25844 5208 25846
rect 5852 28476 5908 28532
rect 6412 35084 6468 35140
rect 6524 39004 6580 39060
rect 6412 34690 6468 34692
rect 6412 34638 6414 34690
rect 6414 34638 6466 34690
rect 6466 34638 6468 34690
rect 6412 34636 6468 34638
rect 6524 34412 6580 34468
rect 6636 35196 6692 35252
rect 6524 34188 6580 34244
rect 6524 33964 6580 34020
rect 6188 32450 6244 32452
rect 6188 32398 6190 32450
rect 6190 32398 6242 32450
rect 6242 32398 6244 32450
rect 6188 32396 6244 32398
rect 6076 31724 6132 31780
rect 6076 30322 6132 30324
rect 6076 30270 6078 30322
rect 6078 30270 6130 30322
rect 6130 30270 6132 30322
rect 6076 30268 6132 30270
rect 6076 28476 6132 28532
rect 6188 28418 6244 28420
rect 6188 28366 6190 28418
rect 6190 28366 6242 28418
rect 6242 28366 6244 28418
rect 6188 28364 6244 28366
rect 5740 27804 5796 27860
rect 5628 27746 5684 27748
rect 5628 27694 5630 27746
rect 5630 27694 5682 27746
rect 5682 27694 5684 27746
rect 5628 27692 5684 27694
rect 5516 27634 5572 27636
rect 5516 27582 5518 27634
rect 5518 27582 5570 27634
rect 5570 27582 5572 27634
rect 5516 27580 5572 27582
rect 5516 27244 5572 27300
rect 6076 27692 6132 27748
rect 5964 27356 6020 27412
rect 6188 27580 6244 27636
rect 6076 27186 6132 27188
rect 6076 27134 6078 27186
rect 6078 27134 6130 27186
rect 6130 27134 6132 27186
rect 6076 27132 6132 27134
rect 5740 27020 5796 27076
rect 5628 26012 5684 26068
rect 5740 26796 5796 26852
rect 4172 25618 4228 25620
rect 4172 25566 4174 25618
rect 4174 25566 4226 25618
rect 4226 25566 4228 25618
rect 4172 25564 4228 25566
rect 3836 24722 3892 24724
rect 3836 24670 3838 24722
rect 3838 24670 3890 24722
rect 3890 24670 3892 24722
rect 3836 24668 3892 24670
rect 5852 26460 5908 26516
rect 6076 26572 6132 26628
rect 5404 25564 5460 25620
rect 4732 25394 4788 25396
rect 4732 25342 4734 25394
rect 4734 25342 4786 25394
rect 4786 25342 4788 25394
rect 4732 25340 4788 25342
rect 5292 25228 5348 25284
rect 4008 24330 4064 24332
rect 4112 24330 4168 24332
rect 4008 24278 4024 24330
rect 4024 24278 4064 24330
rect 4112 24278 4148 24330
rect 4148 24278 4168 24330
rect 4008 24276 4064 24278
rect 4112 24276 4168 24278
rect 4216 24276 4272 24332
rect 4320 24330 4376 24332
rect 4424 24330 4480 24332
rect 4528 24330 4584 24332
rect 4320 24278 4324 24330
rect 4324 24278 4376 24330
rect 4424 24278 4448 24330
rect 4448 24278 4480 24330
rect 4528 24278 4572 24330
rect 4572 24278 4584 24330
rect 4320 24276 4376 24278
rect 4424 24276 4480 24278
rect 4528 24276 4584 24278
rect 4632 24330 4688 24332
rect 4736 24330 4792 24332
rect 4840 24330 4896 24332
rect 4632 24278 4644 24330
rect 4644 24278 4688 24330
rect 4736 24278 4768 24330
rect 4768 24278 4792 24330
rect 4840 24278 4892 24330
rect 4892 24278 4896 24330
rect 4632 24276 4688 24278
rect 4736 24276 4792 24278
rect 4840 24276 4896 24278
rect 4944 24276 5000 24332
rect 5048 24330 5104 24332
rect 5152 24330 5208 24332
rect 5048 24278 5068 24330
rect 5068 24278 5104 24330
rect 5152 24278 5192 24330
rect 5192 24278 5208 24330
rect 5048 24276 5104 24278
rect 5152 24276 5208 24278
rect 3836 23436 3892 23492
rect 4508 23826 4564 23828
rect 4508 23774 4510 23826
rect 4510 23774 4562 23826
rect 4562 23774 4564 23826
rect 4508 23772 4564 23774
rect 4508 23548 4564 23604
rect 3948 23212 4004 23268
rect 5180 23436 5236 23492
rect 3948 22876 4004 22932
rect 4508 22930 4564 22932
rect 4508 22878 4510 22930
rect 4510 22878 4562 22930
rect 4562 22878 4564 22930
rect 4508 22876 4564 22878
rect 4008 22762 4064 22764
rect 4112 22762 4168 22764
rect 4008 22710 4024 22762
rect 4024 22710 4064 22762
rect 4112 22710 4148 22762
rect 4148 22710 4168 22762
rect 4008 22708 4064 22710
rect 4112 22708 4168 22710
rect 4216 22708 4272 22764
rect 4320 22762 4376 22764
rect 4424 22762 4480 22764
rect 4528 22762 4584 22764
rect 4320 22710 4324 22762
rect 4324 22710 4376 22762
rect 4424 22710 4448 22762
rect 4448 22710 4480 22762
rect 4528 22710 4572 22762
rect 4572 22710 4584 22762
rect 4320 22708 4376 22710
rect 4424 22708 4480 22710
rect 4528 22708 4584 22710
rect 4632 22762 4688 22764
rect 4736 22762 4792 22764
rect 4840 22762 4896 22764
rect 4632 22710 4644 22762
rect 4644 22710 4688 22762
rect 4736 22710 4768 22762
rect 4768 22710 4792 22762
rect 4840 22710 4892 22762
rect 4892 22710 4896 22762
rect 4632 22708 4688 22710
rect 4736 22708 4792 22710
rect 4840 22708 4896 22710
rect 4944 22708 5000 22764
rect 5048 22762 5104 22764
rect 5152 22762 5208 22764
rect 5048 22710 5068 22762
rect 5068 22710 5104 22762
rect 5152 22710 5192 22762
rect 5192 22710 5208 22762
rect 5048 22708 5104 22710
rect 5152 22708 5208 22710
rect 4172 22594 4228 22596
rect 4172 22542 4174 22594
rect 4174 22542 4226 22594
rect 4226 22542 4228 22594
rect 4172 22540 4228 22542
rect 4844 22092 4900 22148
rect 4844 21810 4900 21812
rect 4844 21758 4846 21810
rect 4846 21758 4898 21810
rect 4898 21758 4900 21810
rect 4844 21756 4900 21758
rect 3836 21644 3892 21700
rect 5404 23266 5460 23268
rect 5404 23214 5406 23266
rect 5406 23214 5458 23266
rect 5458 23214 5460 23266
rect 5404 23212 5460 23214
rect 5964 26012 6020 26068
rect 7196 45388 7252 45444
rect 7308 45276 7364 45332
rect 7308 44716 7364 44772
rect 7308 44380 7364 44436
rect 7644 45106 7700 45108
rect 7644 45054 7646 45106
rect 7646 45054 7698 45106
rect 7698 45054 7700 45106
rect 7644 45052 7700 45054
rect 7644 44716 7700 44772
rect 8092 47234 8148 47236
rect 8092 47182 8094 47234
rect 8094 47182 8146 47234
rect 8146 47182 8148 47234
rect 8092 47180 8148 47182
rect 8204 45388 8260 45444
rect 7980 45052 8036 45108
rect 8988 48130 9044 48132
rect 8988 48078 8990 48130
rect 8990 48078 9042 48130
rect 9042 48078 9044 48130
rect 8988 48076 9044 48078
rect 8764 47628 8820 47684
rect 9100 47346 9156 47348
rect 9100 47294 9102 47346
rect 9102 47294 9154 47346
rect 9154 47294 9156 47346
rect 9100 47292 9156 47294
rect 9100 46562 9156 46564
rect 9100 46510 9102 46562
rect 9102 46510 9154 46562
rect 9154 46510 9156 46562
rect 9100 46508 9156 46510
rect 9660 56476 9716 56532
rect 9660 54012 9716 54068
rect 9772 53676 9828 53732
rect 9660 51884 9716 51940
rect 9660 50034 9716 50036
rect 9660 49982 9662 50034
rect 9662 49982 9714 50034
rect 9714 49982 9716 50034
rect 9660 49980 9716 49982
rect 9772 49644 9828 49700
rect 9436 48524 9492 48580
rect 9996 62188 10052 62244
rect 10668 65490 10724 65492
rect 10668 65438 10670 65490
rect 10670 65438 10722 65490
rect 10722 65438 10724 65490
rect 10668 65436 10724 65438
rect 10444 64818 10500 64820
rect 10444 64766 10446 64818
rect 10446 64766 10498 64818
rect 10498 64766 10500 64818
rect 10444 64764 10500 64766
rect 11004 66498 11060 66500
rect 11004 66446 11006 66498
rect 11006 66446 11058 66498
rect 11058 66446 11060 66498
rect 11004 66444 11060 66446
rect 12012 69634 12068 69636
rect 12012 69582 12014 69634
rect 12014 69582 12066 69634
rect 12066 69582 12068 69634
rect 12012 69580 12068 69582
rect 11900 69244 11956 69300
rect 11228 69186 11284 69188
rect 11228 69134 11230 69186
rect 11230 69134 11282 69186
rect 11282 69134 11284 69186
rect 11228 69132 11284 69134
rect 12236 69132 12292 69188
rect 13020 73724 13076 73780
rect 13132 74956 13188 75012
rect 11228 67618 11284 67620
rect 11228 67566 11230 67618
rect 11230 67566 11282 67618
rect 11282 67566 11284 67618
rect 11228 67564 11284 67566
rect 11900 68460 11956 68516
rect 11452 67228 11508 67284
rect 12908 69132 12964 69188
rect 12572 67564 12628 67620
rect 12236 67228 12292 67284
rect 12572 67116 12628 67172
rect 11228 66162 11284 66164
rect 11228 66110 11230 66162
rect 11230 66110 11282 66162
rect 11282 66110 11284 66162
rect 11228 66108 11284 66110
rect 11116 65436 11172 65492
rect 10444 63756 10500 63812
rect 10444 63308 10500 63364
rect 10220 62076 10276 62132
rect 10332 61570 10388 61572
rect 10332 61518 10334 61570
rect 10334 61518 10386 61570
rect 10386 61518 10388 61570
rect 10332 61516 10388 61518
rect 10108 60674 10164 60676
rect 10108 60622 10110 60674
rect 10110 60622 10162 60674
rect 10162 60622 10164 60674
rect 10108 60620 10164 60622
rect 10220 58492 10276 58548
rect 9996 56812 10052 56868
rect 10556 57762 10612 57764
rect 10556 57710 10558 57762
rect 10558 57710 10610 57762
rect 10610 57710 10612 57762
rect 10556 57708 10612 57710
rect 10444 56588 10500 56644
rect 10108 56252 10164 56308
rect 10556 56476 10612 56532
rect 11340 64930 11396 64932
rect 11340 64878 11342 64930
rect 11342 64878 11394 64930
rect 11394 64878 11396 64930
rect 11340 64876 11396 64878
rect 11004 63308 11060 63364
rect 10892 62860 10948 62916
rect 10892 62354 10948 62356
rect 10892 62302 10894 62354
rect 10894 62302 10946 62354
rect 10946 62302 10948 62354
rect 10892 62300 10948 62302
rect 10780 61346 10836 61348
rect 10780 61294 10782 61346
rect 10782 61294 10834 61346
rect 10834 61294 10836 61346
rect 10780 61292 10836 61294
rect 10444 55916 10500 55972
rect 10780 57484 10836 57540
rect 10780 57148 10836 57204
rect 10108 55468 10164 55524
rect 10668 55970 10724 55972
rect 10668 55918 10670 55970
rect 10670 55918 10722 55970
rect 10722 55918 10724 55970
rect 10668 55916 10724 55918
rect 10220 55132 10276 55188
rect 10108 54908 10164 54964
rect 9996 54684 10052 54740
rect 10108 53116 10164 53172
rect 10220 54348 10276 54404
rect 10108 52220 10164 52276
rect 10668 55132 10724 55188
rect 10332 53788 10388 53844
rect 11676 67004 11732 67060
rect 11676 66332 11732 66388
rect 11788 64876 11844 64932
rect 12236 64876 12292 64932
rect 11228 61852 11284 61908
rect 12012 64428 12068 64484
rect 11004 61516 11060 61572
rect 11116 61292 11172 61348
rect 11004 61180 11060 61236
rect 11116 57148 11172 57204
rect 11004 55020 11060 55076
rect 10780 54626 10836 54628
rect 10780 54574 10782 54626
rect 10782 54574 10834 54626
rect 10834 54574 10836 54626
rect 10780 54572 10836 54574
rect 10668 53564 10724 53620
rect 10892 53506 10948 53508
rect 10892 53454 10894 53506
rect 10894 53454 10946 53506
rect 10946 53454 10948 53506
rect 10892 53452 10948 53454
rect 10220 49980 10276 50036
rect 10332 49698 10388 49700
rect 10332 49646 10334 49698
rect 10334 49646 10386 49698
rect 10386 49646 10388 49698
rect 10332 49644 10388 49646
rect 9996 48242 10052 48244
rect 9996 48190 9998 48242
rect 9998 48190 10050 48242
rect 10050 48190 10052 48242
rect 9996 48188 10052 48190
rect 9884 48130 9940 48132
rect 9884 48078 9886 48130
rect 9886 48078 9938 48130
rect 9938 48078 9940 48130
rect 9884 48076 9940 48078
rect 9436 47068 9492 47124
rect 9436 46620 9492 46676
rect 9324 45948 9380 46004
rect 6972 43708 7028 43764
rect 6972 39394 7028 39396
rect 6972 39342 6974 39394
rect 6974 39342 7026 39394
rect 7026 39342 7028 39394
rect 6972 39340 7028 39342
rect 6972 39004 7028 39060
rect 6860 34076 6916 34132
rect 6972 36540 7028 36596
rect 7196 42588 7252 42644
rect 7196 40684 7252 40740
rect 7420 42866 7476 42868
rect 7420 42814 7422 42866
rect 7422 42814 7474 42866
rect 7474 42814 7476 42866
rect 7420 42812 7476 42814
rect 7420 40626 7476 40628
rect 7420 40574 7422 40626
rect 7422 40574 7474 40626
rect 7474 40574 7476 40626
rect 7420 40572 7476 40574
rect 7532 41132 7588 41188
rect 7532 40236 7588 40292
rect 7308 39618 7364 39620
rect 7308 39566 7310 39618
rect 7310 39566 7362 39618
rect 7362 39566 7364 39618
rect 7308 39564 7364 39566
rect 7308 37772 7364 37828
rect 7084 36428 7140 36484
rect 7420 37324 7476 37380
rect 7084 35980 7140 36036
rect 7532 39116 7588 39172
rect 7532 36540 7588 36596
rect 8092 44268 8148 44324
rect 8092 43708 8148 43764
rect 9660 45106 9716 45108
rect 9660 45054 9662 45106
rect 9662 45054 9714 45106
rect 9714 45054 9716 45106
rect 9660 45052 9716 45054
rect 8316 44322 8372 44324
rect 8316 44270 8318 44322
rect 8318 44270 8370 44322
rect 8370 44270 8372 44322
rect 8316 44268 8372 44270
rect 8204 43426 8260 43428
rect 8204 43374 8206 43426
rect 8206 43374 8258 43426
rect 8258 43374 8260 43426
rect 8204 43372 8260 43374
rect 9660 44268 9716 44324
rect 8540 43372 8596 43428
rect 8204 42588 8260 42644
rect 8540 42866 8596 42868
rect 8540 42814 8542 42866
rect 8542 42814 8594 42866
rect 8594 42814 8596 42866
rect 8540 42812 8596 42814
rect 9212 42924 9268 42980
rect 8876 42812 8932 42868
rect 8428 41970 8484 41972
rect 8428 41918 8430 41970
rect 8430 41918 8482 41970
rect 8482 41918 8484 41970
rect 8428 41916 8484 41918
rect 7980 41132 8036 41188
rect 8316 41804 8372 41860
rect 8652 42530 8708 42532
rect 8652 42478 8654 42530
rect 8654 42478 8706 42530
rect 8706 42478 8708 42530
rect 8652 42476 8708 42478
rect 9212 42140 9268 42196
rect 8204 41074 8260 41076
rect 8204 41022 8206 41074
rect 8206 41022 8258 41074
rect 8258 41022 8260 41074
rect 8204 41020 8260 41022
rect 7980 40962 8036 40964
rect 7980 40910 7982 40962
rect 7982 40910 8034 40962
rect 8034 40910 8036 40962
rect 7980 40908 8036 40910
rect 7980 40626 8036 40628
rect 7980 40574 7982 40626
rect 7982 40574 8034 40626
rect 8034 40574 8036 40626
rect 7980 40572 8036 40574
rect 9660 42812 9716 42868
rect 9660 42476 9716 42532
rect 9212 41916 9268 41972
rect 9884 47682 9940 47684
rect 9884 47630 9886 47682
rect 9886 47630 9938 47682
rect 9938 47630 9940 47682
rect 9884 47628 9940 47630
rect 9772 41804 9828 41860
rect 8764 40572 8820 40628
rect 7868 40460 7924 40516
rect 8316 40514 8372 40516
rect 8316 40462 8318 40514
rect 8318 40462 8370 40514
rect 8370 40462 8372 40514
rect 8316 40460 8372 40462
rect 7980 40012 8036 40068
rect 8092 39058 8148 39060
rect 8092 39006 8094 39058
rect 8094 39006 8146 39058
rect 8146 39006 8148 39058
rect 8092 39004 8148 39006
rect 8092 38556 8148 38612
rect 7532 36258 7588 36260
rect 7532 36206 7534 36258
rect 7534 36206 7586 36258
rect 7586 36206 7588 36258
rect 7532 36204 7588 36206
rect 7868 36316 7924 36372
rect 7196 34972 7252 35028
rect 7420 35532 7476 35588
rect 7308 34914 7364 34916
rect 7308 34862 7310 34914
rect 7310 34862 7362 34914
rect 7362 34862 7364 34914
rect 7308 34860 7364 34862
rect 7084 34748 7140 34804
rect 7308 34412 7364 34468
rect 6972 34188 7028 34244
rect 7196 34076 7252 34132
rect 6748 33404 6804 33460
rect 6636 33234 6692 33236
rect 6636 33182 6638 33234
rect 6638 33182 6690 33234
rect 6690 33182 6692 33234
rect 6636 33180 6692 33182
rect 6636 32396 6692 32452
rect 6524 31836 6580 31892
rect 6412 27858 6468 27860
rect 6412 27806 6414 27858
rect 6414 27806 6466 27858
rect 6466 27806 6468 27858
rect 6412 27804 6468 27806
rect 6412 27298 6468 27300
rect 6412 27246 6414 27298
rect 6414 27246 6466 27298
rect 6466 27246 6468 27298
rect 6412 27244 6468 27246
rect 6300 27020 6356 27076
rect 7084 33964 7140 34020
rect 6860 32956 6916 33012
rect 7644 34636 7700 34692
rect 7644 34412 7700 34468
rect 7532 34076 7588 34132
rect 7420 33180 7476 33236
rect 7644 34188 7700 34244
rect 7532 32450 7588 32452
rect 7532 32398 7534 32450
rect 7534 32398 7586 32450
rect 7586 32398 7588 32450
rect 7532 32396 7588 32398
rect 6748 28140 6804 28196
rect 6860 29484 6916 29540
rect 7532 31836 7588 31892
rect 7308 30940 7364 30996
rect 7868 34018 7924 34020
rect 7868 33966 7870 34018
rect 7870 33966 7922 34018
rect 7922 33966 7924 34018
rect 7868 33964 7924 33966
rect 8764 39564 8820 39620
rect 8652 39116 8708 39172
rect 8316 38780 8372 38836
rect 8428 36540 8484 36596
rect 8652 38220 8708 38276
rect 8316 36428 8372 36484
rect 8428 35644 8484 35700
rect 8204 34188 8260 34244
rect 8428 34300 8484 34356
rect 8988 39394 9044 39396
rect 8988 39342 8990 39394
rect 8990 39342 9042 39394
rect 9042 39342 9044 39394
rect 8988 39340 9044 39342
rect 8988 38668 9044 38724
rect 9324 40572 9380 40628
rect 9660 39564 9716 39620
rect 9548 39394 9604 39396
rect 9548 39342 9550 39394
rect 9550 39342 9602 39394
rect 9602 39342 9604 39394
rect 9548 39340 9604 39342
rect 9436 39004 9492 39060
rect 8876 37826 8932 37828
rect 8876 37774 8878 37826
rect 8878 37774 8930 37826
rect 8930 37774 8932 37826
rect 8876 37772 8932 37774
rect 8764 36370 8820 36372
rect 8764 36318 8766 36370
rect 8766 36318 8818 36370
rect 8818 36318 8820 36370
rect 8764 36316 8820 36318
rect 9996 46674 10052 46676
rect 9996 46622 9998 46674
rect 9998 46622 10050 46674
rect 10050 46622 10052 46674
rect 9996 46620 10052 46622
rect 9996 45164 10052 45220
rect 10780 52892 10836 52948
rect 10556 52668 10612 52724
rect 11004 52780 11060 52836
rect 11004 52274 11060 52276
rect 11004 52222 11006 52274
rect 11006 52222 11058 52274
rect 11058 52222 11060 52274
rect 11004 52220 11060 52222
rect 10892 52050 10948 52052
rect 10892 51998 10894 52050
rect 10894 51998 10946 52050
rect 10946 51998 10948 52050
rect 10892 51996 10948 51998
rect 11004 48466 11060 48468
rect 11004 48414 11006 48466
rect 11006 48414 11058 48466
rect 11058 48414 11060 48466
rect 11004 48412 11060 48414
rect 12236 64316 12292 64372
rect 12796 65212 12852 65268
rect 14476 82738 14532 82740
rect 14476 82686 14478 82738
rect 14478 82686 14530 82738
rect 14530 82686 14532 82738
rect 14476 82684 14532 82686
rect 15148 82236 15204 82292
rect 14476 82066 14532 82068
rect 14476 82014 14478 82066
rect 14478 82014 14530 82066
rect 14530 82014 14532 82066
rect 14476 82012 14532 82014
rect 14364 81900 14420 81956
rect 15260 82796 15316 82852
rect 15372 82684 15428 82740
rect 16492 84140 16548 84196
rect 15932 83468 15988 83524
rect 15708 82796 15764 82852
rect 15596 82460 15652 82516
rect 13692 81842 13748 81844
rect 13692 81790 13694 81842
rect 13694 81790 13746 81842
rect 13746 81790 13748 81842
rect 13692 81788 13748 81790
rect 14028 81788 14084 81844
rect 14812 81842 14868 81844
rect 14812 81790 14814 81842
rect 14814 81790 14866 81842
rect 14866 81790 14868 81842
rect 14812 81788 14868 81790
rect 14700 81730 14756 81732
rect 14700 81678 14702 81730
rect 14702 81678 14754 81730
rect 14754 81678 14756 81730
rect 14700 81676 14756 81678
rect 15260 81676 15316 81732
rect 15372 82124 15428 82180
rect 14008 81562 14064 81564
rect 14112 81562 14168 81564
rect 14008 81510 14024 81562
rect 14024 81510 14064 81562
rect 14112 81510 14148 81562
rect 14148 81510 14168 81562
rect 14008 81508 14064 81510
rect 14112 81508 14168 81510
rect 14216 81508 14272 81564
rect 14320 81562 14376 81564
rect 14424 81562 14480 81564
rect 14528 81562 14584 81564
rect 14320 81510 14324 81562
rect 14324 81510 14376 81562
rect 14424 81510 14448 81562
rect 14448 81510 14480 81562
rect 14528 81510 14572 81562
rect 14572 81510 14584 81562
rect 14320 81508 14376 81510
rect 14424 81508 14480 81510
rect 14528 81508 14584 81510
rect 14632 81562 14688 81564
rect 14736 81562 14792 81564
rect 14840 81562 14896 81564
rect 14632 81510 14644 81562
rect 14644 81510 14688 81562
rect 14736 81510 14768 81562
rect 14768 81510 14792 81562
rect 14840 81510 14892 81562
rect 14892 81510 14896 81562
rect 14632 81508 14688 81510
rect 14736 81508 14792 81510
rect 14840 81508 14896 81510
rect 14944 81508 15000 81564
rect 15048 81562 15104 81564
rect 15152 81562 15208 81564
rect 15048 81510 15068 81562
rect 15068 81510 15104 81562
rect 15152 81510 15192 81562
rect 15192 81510 15208 81562
rect 15048 81508 15104 81510
rect 15152 81508 15208 81510
rect 14700 81340 14756 81396
rect 14140 81116 14196 81172
rect 13916 81058 13972 81060
rect 13916 81006 13918 81058
rect 13918 81006 13970 81058
rect 13970 81006 13972 81058
rect 13916 81004 13972 81006
rect 13356 77196 13412 77252
rect 13916 80444 13972 80500
rect 14588 81004 14644 81060
rect 14364 80332 14420 80388
rect 14476 80556 14532 80612
rect 15484 81340 15540 81396
rect 15036 81228 15092 81284
rect 14700 80444 14756 80500
rect 13916 80162 13972 80164
rect 13916 80110 13918 80162
rect 13918 80110 13970 80162
rect 13970 80110 13972 80162
rect 13916 80108 13972 80110
rect 15260 81282 15316 81284
rect 15260 81230 15262 81282
rect 15262 81230 15314 81282
rect 15314 81230 15316 81282
rect 15260 81228 15316 81230
rect 14812 80108 14868 80164
rect 15372 80332 15428 80388
rect 14008 79994 14064 79996
rect 14112 79994 14168 79996
rect 14008 79942 14024 79994
rect 14024 79942 14064 79994
rect 14112 79942 14148 79994
rect 14148 79942 14168 79994
rect 14008 79940 14064 79942
rect 14112 79940 14168 79942
rect 14216 79940 14272 79996
rect 14320 79994 14376 79996
rect 14424 79994 14480 79996
rect 14528 79994 14584 79996
rect 14320 79942 14324 79994
rect 14324 79942 14376 79994
rect 14424 79942 14448 79994
rect 14448 79942 14480 79994
rect 14528 79942 14572 79994
rect 14572 79942 14584 79994
rect 14320 79940 14376 79942
rect 14424 79940 14480 79942
rect 14528 79940 14584 79942
rect 14632 79994 14688 79996
rect 14736 79994 14792 79996
rect 14840 79994 14896 79996
rect 14632 79942 14644 79994
rect 14644 79942 14688 79994
rect 14736 79942 14768 79994
rect 14768 79942 14792 79994
rect 14840 79942 14892 79994
rect 14892 79942 14896 79994
rect 14632 79940 14688 79942
rect 14736 79940 14792 79942
rect 14840 79940 14896 79942
rect 14944 79940 15000 79996
rect 15048 79994 15104 79996
rect 15152 79994 15208 79996
rect 15048 79942 15068 79994
rect 15068 79942 15104 79994
rect 15152 79942 15192 79994
rect 15192 79942 15208 79994
rect 15048 79940 15104 79942
rect 15152 79940 15208 79942
rect 15260 79772 15316 79828
rect 13804 79490 13860 79492
rect 13804 79438 13806 79490
rect 13806 79438 13858 79490
rect 13858 79438 13860 79490
rect 13804 79436 13860 79438
rect 14252 79548 14308 79604
rect 13692 78876 13748 78932
rect 13356 75740 13412 75796
rect 15148 79436 15204 79492
rect 15596 79772 15652 79828
rect 16268 83244 16324 83300
rect 16268 82850 16324 82852
rect 16268 82798 16270 82850
rect 16270 82798 16322 82850
rect 16322 82798 16324 82850
rect 16268 82796 16324 82798
rect 15932 82348 15988 82404
rect 16492 82236 16548 82292
rect 16268 81954 16324 81956
rect 16268 81902 16270 81954
rect 16270 81902 16322 81954
rect 16322 81902 16324 81954
rect 16268 81900 16324 81902
rect 16156 81788 16212 81844
rect 16940 87330 16996 87332
rect 16940 87278 16942 87330
rect 16942 87278 16994 87330
rect 16994 87278 16996 87330
rect 16940 87276 16996 87278
rect 20412 87666 20468 87668
rect 20412 87614 20414 87666
rect 20414 87614 20466 87666
rect 20466 87614 20468 87666
rect 20412 87612 20468 87614
rect 17388 87276 17444 87332
rect 19404 87388 19460 87444
rect 16828 85762 16884 85764
rect 16828 85710 16830 85762
rect 16830 85710 16882 85762
rect 16882 85710 16884 85762
rect 16828 85708 16884 85710
rect 18060 85932 18116 85988
rect 18284 86044 18340 86100
rect 16716 84140 16772 84196
rect 17052 83298 17108 83300
rect 17052 83246 17054 83298
rect 17054 83246 17106 83298
rect 17106 83246 17108 83298
rect 17052 83244 17108 83246
rect 16828 82738 16884 82740
rect 16828 82686 16830 82738
rect 16830 82686 16882 82738
rect 16882 82686 16884 82738
rect 16828 82684 16884 82686
rect 16716 82348 16772 82404
rect 16716 81900 16772 81956
rect 16492 81730 16548 81732
rect 16492 81678 16494 81730
rect 16494 81678 16546 81730
rect 16546 81678 16548 81730
rect 16492 81676 16548 81678
rect 16492 81452 16548 81508
rect 16044 81340 16100 81396
rect 16716 81340 16772 81396
rect 17052 81788 17108 81844
rect 17052 81228 17108 81284
rect 16492 81170 16548 81172
rect 16492 81118 16494 81170
rect 16494 81118 16546 81170
rect 16546 81118 16548 81170
rect 16492 81116 16548 81118
rect 16716 81170 16772 81172
rect 16716 81118 16718 81170
rect 16718 81118 16770 81170
rect 16770 81118 16772 81170
rect 16716 81116 16772 81118
rect 15820 80386 15876 80388
rect 15820 80334 15822 80386
rect 15822 80334 15874 80386
rect 15874 80334 15876 80386
rect 15820 80332 15876 80334
rect 16380 81004 16436 81060
rect 16380 79436 16436 79492
rect 16716 80892 16772 80948
rect 15372 78988 15428 79044
rect 13916 78652 13972 78708
rect 13580 78540 13636 78596
rect 14008 78426 14064 78428
rect 14112 78426 14168 78428
rect 14008 78374 14024 78426
rect 14024 78374 14064 78426
rect 14112 78374 14148 78426
rect 14148 78374 14168 78426
rect 14008 78372 14064 78374
rect 14112 78372 14168 78374
rect 14216 78372 14272 78428
rect 14320 78426 14376 78428
rect 14424 78426 14480 78428
rect 14528 78426 14584 78428
rect 14320 78374 14324 78426
rect 14324 78374 14376 78426
rect 14424 78374 14448 78426
rect 14448 78374 14480 78426
rect 14528 78374 14572 78426
rect 14572 78374 14584 78426
rect 14320 78372 14376 78374
rect 14424 78372 14480 78374
rect 14528 78372 14584 78374
rect 14632 78426 14688 78428
rect 14736 78426 14792 78428
rect 14840 78426 14896 78428
rect 14632 78374 14644 78426
rect 14644 78374 14688 78426
rect 14736 78374 14768 78426
rect 14768 78374 14792 78426
rect 14840 78374 14892 78426
rect 14892 78374 14896 78426
rect 14632 78372 14688 78374
rect 14736 78372 14792 78374
rect 14840 78372 14896 78374
rect 14944 78372 15000 78428
rect 15048 78426 15104 78428
rect 15152 78426 15208 78428
rect 15048 78374 15068 78426
rect 15068 78374 15104 78426
rect 15152 78374 15192 78426
rect 15192 78374 15208 78426
rect 15048 78372 15104 78374
rect 15152 78372 15208 78374
rect 14700 78204 14756 78260
rect 13580 78092 13636 78148
rect 14588 77308 14644 77364
rect 13804 77250 13860 77252
rect 13804 77198 13806 77250
rect 13806 77198 13858 77250
rect 13858 77198 13860 77250
rect 13804 77196 13860 77198
rect 14028 77196 14084 77252
rect 15372 78034 15428 78036
rect 15372 77982 15374 78034
rect 15374 77982 15426 78034
rect 15426 77982 15428 78034
rect 15372 77980 15428 77982
rect 15372 77138 15428 77140
rect 15372 77086 15374 77138
rect 15374 77086 15426 77138
rect 15426 77086 15428 77138
rect 15372 77084 15428 77086
rect 15148 77026 15204 77028
rect 15148 76974 15150 77026
rect 15150 76974 15202 77026
rect 15202 76974 15204 77026
rect 15148 76972 15204 76974
rect 14008 76858 14064 76860
rect 14112 76858 14168 76860
rect 14008 76806 14024 76858
rect 14024 76806 14064 76858
rect 14112 76806 14148 76858
rect 14148 76806 14168 76858
rect 14008 76804 14064 76806
rect 14112 76804 14168 76806
rect 14216 76804 14272 76860
rect 14320 76858 14376 76860
rect 14424 76858 14480 76860
rect 14528 76858 14584 76860
rect 14320 76806 14324 76858
rect 14324 76806 14376 76858
rect 14424 76806 14448 76858
rect 14448 76806 14480 76858
rect 14528 76806 14572 76858
rect 14572 76806 14584 76858
rect 14320 76804 14376 76806
rect 14424 76804 14480 76806
rect 14528 76804 14584 76806
rect 14632 76858 14688 76860
rect 14736 76858 14792 76860
rect 14840 76858 14896 76860
rect 14632 76806 14644 76858
rect 14644 76806 14688 76858
rect 14736 76806 14768 76858
rect 14768 76806 14792 76858
rect 14840 76806 14892 76858
rect 14892 76806 14896 76858
rect 14632 76804 14688 76806
rect 14736 76804 14792 76806
rect 14840 76804 14896 76806
rect 14944 76804 15000 76860
rect 15048 76858 15104 76860
rect 15152 76858 15208 76860
rect 15048 76806 15068 76858
rect 15068 76806 15104 76858
rect 15152 76806 15192 76858
rect 15192 76806 15208 76858
rect 15048 76804 15104 76806
rect 15152 76804 15208 76806
rect 15372 76860 15428 76916
rect 15596 76748 15652 76804
rect 13580 76412 13636 76468
rect 15820 78540 15876 78596
rect 15708 76636 15764 76692
rect 14588 76578 14644 76580
rect 14588 76526 14590 76578
rect 14590 76526 14642 76578
rect 14642 76526 14644 76578
rect 14588 76524 14644 76526
rect 15820 76578 15876 76580
rect 15820 76526 15822 76578
rect 15822 76526 15874 76578
rect 15874 76526 15876 76578
rect 15820 76524 15876 76526
rect 15372 76412 15428 76468
rect 14476 75516 14532 75572
rect 13804 75404 13860 75460
rect 13580 73724 13636 73780
rect 13580 70924 13636 70980
rect 13580 70418 13636 70420
rect 13580 70366 13582 70418
rect 13582 70366 13634 70418
rect 13634 70366 13636 70418
rect 13580 70364 13636 70366
rect 13580 69186 13636 69188
rect 13580 69134 13582 69186
rect 13582 69134 13634 69186
rect 13634 69134 13636 69186
rect 13580 69132 13636 69134
rect 13356 69020 13412 69076
rect 13580 68796 13636 68852
rect 13244 67564 13300 67620
rect 13468 67676 13524 67732
rect 13244 67116 13300 67172
rect 13020 65100 13076 65156
rect 13132 66444 13188 66500
rect 13468 67228 13524 67284
rect 13580 67004 13636 67060
rect 14924 75794 14980 75796
rect 14924 75742 14926 75794
rect 14926 75742 14978 75794
rect 14978 75742 14980 75794
rect 14924 75740 14980 75742
rect 16044 77084 16100 77140
rect 16380 77922 16436 77924
rect 16380 77870 16382 77922
rect 16382 77870 16434 77922
rect 16434 77870 16436 77922
rect 16380 77868 16436 77870
rect 16380 76748 16436 76804
rect 16380 76466 16436 76468
rect 16380 76414 16382 76466
rect 16382 76414 16434 76466
rect 16434 76414 16436 76466
rect 16380 76412 16436 76414
rect 16044 76300 16100 76356
rect 14700 75404 14756 75460
rect 14008 75290 14064 75292
rect 14112 75290 14168 75292
rect 14008 75238 14024 75290
rect 14024 75238 14064 75290
rect 14112 75238 14148 75290
rect 14148 75238 14168 75290
rect 14008 75236 14064 75238
rect 14112 75236 14168 75238
rect 14216 75236 14272 75292
rect 14320 75290 14376 75292
rect 14424 75290 14480 75292
rect 14528 75290 14584 75292
rect 14320 75238 14324 75290
rect 14324 75238 14376 75290
rect 14424 75238 14448 75290
rect 14448 75238 14480 75290
rect 14528 75238 14572 75290
rect 14572 75238 14584 75290
rect 14320 75236 14376 75238
rect 14424 75236 14480 75238
rect 14528 75236 14584 75238
rect 14632 75290 14688 75292
rect 14736 75290 14792 75292
rect 14840 75290 14896 75292
rect 14632 75238 14644 75290
rect 14644 75238 14688 75290
rect 14736 75238 14768 75290
rect 14768 75238 14792 75290
rect 14840 75238 14892 75290
rect 14892 75238 14896 75290
rect 14632 75236 14688 75238
rect 14736 75236 14792 75238
rect 14840 75236 14896 75238
rect 14944 75236 15000 75292
rect 15048 75290 15104 75292
rect 15152 75290 15208 75292
rect 15048 75238 15068 75290
rect 15068 75238 15104 75290
rect 15152 75238 15192 75290
rect 15192 75238 15208 75290
rect 15048 75236 15104 75238
rect 15152 75236 15208 75238
rect 14252 75122 14308 75124
rect 14252 75070 14254 75122
rect 14254 75070 14306 75122
rect 14306 75070 14308 75122
rect 14252 75068 14308 75070
rect 14364 73836 14420 73892
rect 15372 73836 15428 73892
rect 14008 73722 14064 73724
rect 14112 73722 14168 73724
rect 14008 73670 14024 73722
rect 14024 73670 14064 73722
rect 14112 73670 14148 73722
rect 14148 73670 14168 73722
rect 14008 73668 14064 73670
rect 14112 73668 14168 73670
rect 14216 73668 14272 73724
rect 14320 73722 14376 73724
rect 14424 73722 14480 73724
rect 14528 73722 14584 73724
rect 14320 73670 14324 73722
rect 14324 73670 14376 73722
rect 14424 73670 14448 73722
rect 14448 73670 14480 73722
rect 14528 73670 14572 73722
rect 14572 73670 14584 73722
rect 14320 73668 14376 73670
rect 14424 73668 14480 73670
rect 14528 73668 14584 73670
rect 14632 73722 14688 73724
rect 14736 73722 14792 73724
rect 14840 73722 14896 73724
rect 14632 73670 14644 73722
rect 14644 73670 14688 73722
rect 14736 73670 14768 73722
rect 14768 73670 14792 73722
rect 14840 73670 14892 73722
rect 14892 73670 14896 73722
rect 14632 73668 14688 73670
rect 14736 73668 14792 73670
rect 14840 73668 14896 73670
rect 14944 73668 15000 73724
rect 15048 73722 15104 73724
rect 15152 73722 15208 73724
rect 15048 73670 15068 73722
rect 15068 73670 15104 73722
rect 15152 73670 15192 73722
rect 15192 73670 15208 73722
rect 15048 73668 15104 73670
rect 15152 73668 15208 73670
rect 14364 73554 14420 73556
rect 14364 73502 14366 73554
rect 14366 73502 14418 73554
rect 14418 73502 14420 73554
rect 14364 73500 14420 73502
rect 15708 75682 15764 75684
rect 15708 75630 15710 75682
rect 15710 75630 15762 75682
rect 15762 75630 15764 75682
rect 15708 75628 15764 75630
rect 16156 75628 16212 75684
rect 15708 75122 15764 75124
rect 15708 75070 15710 75122
rect 15710 75070 15762 75122
rect 15762 75070 15764 75122
rect 15708 75068 15764 75070
rect 16492 75068 16548 75124
rect 18172 84866 18228 84868
rect 18172 84814 18174 84866
rect 18174 84814 18226 84866
rect 18226 84814 18228 84866
rect 18172 84812 18228 84814
rect 17500 84194 17556 84196
rect 17500 84142 17502 84194
rect 17502 84142 17554 84194
rect 17554 84142 17556 84194
rect 17500 84140 17556 84142
rect 18620 85762 18676 85764
rect 18620 85710 18622 85762
rect 18622 85710 18674 85762
rect 18674 85710 18676 85762
rect 18620 85708 18676 85710
rect 18956 85708 19012 85764
rect 20412 87276 20468 87332
rect 20524 87500 20580 87556
rect 19292 84812 19348 84868
rect 18284 84028 18340 84084
rect 19068 84082 19124 84084
rect 19068 84030 19070 84082
rect 19070 84030 19122 84082
rect 19122 84030 19124 84082
rect 19068 84028 19124 84030
rect 18732 83692 18788 83748
rect 17612 82738 17668 82740
rect 17612 82686 17614 82738
rect 17614 82686 17666 82738
rect 17666 82686 17668 82738
rect 17612 82684 17668 82686
rect 18284 83522 18340 83524
rect 18284 83470 18286 83522
rect 18286 83470 18338 83522
rect 18338 83470 18340 83522
rect 18284 83468 18340 83470
rect 18396 83410 18452 83412
rect 18396 83358 18398 83410
rect 18398 83358 18450 83410
rect 18450 83358 18452 83410
rect 18396 83356 18452 83358
rect 17836 82460 17892 82516
rect 18732 82460 18788 82516
rect 17724 81452 17780 81508
rect 18060 82236 18116 82292
rect 17388 81170 17444 81172
rect 17388 81118 17390 81170
rect 17390 81118 17442 81170
rect 17442 81118 17444 81170
rect 17388 81116 17444 81118
rect 18844 81676 18900 81732
rect 18060 81058 18116 81060
rect 18060 81006 18062 81058
rect 18062 81006 18114 81058
rect 18114 81006 18116 81058
rect 18060 81004 18116 81006
rect 18284 81228 18340 81284
rect 18844 80892 18900 80948
rect 18956 83522 19012 83524
rect 18956 83470 18958 83522
rect 18958 83470 19010 83522
rect 19010 83470 19012 83522
rect 18956 83468 19012 83470
rect 20076 85874 20132 85876
rect 20076 85822 20078 85874
rect 20078 85822 20130 85874
rect 20130 85822 20132 85874
rect 20076 85820 20132 85822
rect 20300 84812 20356 84868
rect 19628 83692 19684 83748
rect 20300 84252 20356 84308
rect 20972 87442 21028 87444
rect 20972 87390 20974 87442
rect 20974 87390 21026 87442
rect 21026 87390 21028 87442
rect 20972 87388 21028 87390
rect 21308 87276 21364 87332
rect 24008 87050 24064 87052
rect 24112 87050 24168 87052
rect 24008 86998 24024 87050
rect 24024 86998 24064 87050
rect 24112 86998 24148 87050
rect 24148 86998 24168 87050
rect 24008 86996 24064 86998
rect 24112 86996 24168 86998
rect 24216 86996 24272 87052
rect 24320 87050 24376 87052
rect 24424 87050 24480 87052
rect 24528 87050 24584 87052
rect 24320 86998 24324 87050
rect 24324 86998 24376 87050
rect 24424 86998 24448 87050
rect 24448 86998 24480 87050
rect 24528 86998 24572 87050
rect 24572 86998 24584 87050
rect 24320 86996 24376 86998
rect 24424 86996 24480 86998
rect 24528 86996 24584 86998
rect 24632 87050 24688 87052
rect 24736 87050 24792 87052
rect 24840 87050 24896 87052
rect 24632 86998 24644 87050
rect 24644 86998 24688 87050
rect 24736 86998 24768 87050
rect 24768 86998 24792 87050
rect 24840 86998 24892 87050
rect 24892 86998 24896 87050
rect 24632 86996 24688 86998
rect 24736 86996 24792 86998
rect 24840 86996 24896 86998
rect 24944 86996 25000 87052
rect 25048 87050 25104 87052
rect 25152 87050 25208 87052
rect 25048 86998 25068 87050
rect 25068 86998 25104 87050
rect 25152 86998 25192 87050
rect 25192 86998 25208 87050
rect 25048 86996 25104 86998
rect 25152 86996 25208 86998
rect 21308 86044 21364 86100
rect 23100 85932 23156 85988
rect 23996 85932 24052 85988
rect 20748 85484 20804 85540
rect 23884 85820 23940 85876
rect 22540 85708 22596 85764
rect 20748 84978 20804 84980
rect 20748 84926 20750 84978
rect 20750 84926 20802 84978
rect 20802 84926 20804 84978
rect 20748 84924 20804 84926
rect 21980 84978 22036 84980
rect 21980 84926 21982 84978
rect 21982 84926 22034 84978
rect 22034 84926 22036 84978
rect 21980 84924 22036 84926
rect 23660 85762 23716 85764
rect 23660 85710 23662 85762
rect 23662 85710 23714 85762
rect 23714 85710 23716 85762
rect 23660 85708 23716 85710
rect 20972 84306 21028 84308
rect 20972 84254 20974 84306
rect 20974 84254 21026 84306
rect 21026 84254 21028 84306
rect 20972 84252 21028 84254
rect 20636 84140 20692 84196
rect 19068 83410 19124 83412
rect 19068 83358 19070 83410
rect 19070 83358 19122 83410
rect 19122 83358 19124 83410
rect 19068 83356 19124 83358
rect 20636 82460 20692 82516
rect 18956 81900 19012 81956
rect 21084 82514 21140 82516
rect 21084 82462 21086 82514
rect 21086 82462 21138 82514
rect 21138 82462 21140 82514
rect 21084 82460 21140 82462
rect 21756 84140 21812 84196
rect 20076 82124 20132 82180
rect 19180 81058 19236 81060
rect 19180 81006 19182 81058
rect 19182 81006 19234 81058
rect 19234 81006 19236 81058
rect 19180 81004 19236 81006
rect 18284 80556 18340 80612
rect 17500 80444 17556 80500
rect 19292 80892 19348 80948
rect 19404 80610 19460 80612
rect 19404 80558 19406 80610
rect 19406 80558 19458 80610
rect 19458 80558 19460 80610
rect 19404 80556 19460 80558
rect 19180 80444 19236 80500
rect 20076 81058 20132 81060
rect 20076 81006 20078 81058
rect 20078 81006 20130 81058
rect 20130 81006 20132 81058
rect 20076 81004 20132 81006
rect 18844 80220 18900 80276
rect 19964 80220 20020 80276
rect 17276 77196 17332 77252
rect 21420 82124 21476 82180
rect 22316 83580 22372 83636
rect 22540 83298 22596 83300
rect 22540 83246 22542 83298
rect 22542 83246 22594 83298
rect 22594 83246 22596 83298
rect 22540 83244 22596 83246
rect 21868 82124 21924 82180
rect 22092 82460 22148 82516
rect 20524 80892 20580 80948
rect 20748 78706 20804 78708
rect 20748 78654 20750 78706
rect 20750 78654 20802 78706
rect 20802 78654 20804 78706
rect 20748 78652 20804 78654
rect 20188 78428 20244 78484
rect 20300 78258 20356 78260
rect 20300 78206 20302 78258
rect 20302 78206 20354 78258
rect 20354 78206 20356 78258
rect 20300 78204 20356 78206
rect 19964 77196 20020 77252
rect 16828 76860 16884 76916
rect 17388 76860 17444 76916
rect 17724 76636 17780 76692
rect 16828 75628 16884 75684
rect 18732 76690 18788 76692
rect 18732 76638 18734 76690
rect 18734 76638 18786 76690
rect 18786 76638 18788 76690
rect 18732 76636 18788 76638
rect 20300 76690 20356 76692
rect 20300 76638 20302 76690
rect 20302 76638 20354 76690
rect 20354 76638 20356 76690
rect 20300 76636 20356 76638
rect 18284 76354 18340 76356
rect 18284 76302 18286 76354
rect 18286 76302 18338 76354
rect 18338 76302 18340 76354
rect 18284 76300 18340 76302
rect 17948 74732 18004 74788
rect 18844 76466 18900 76468
rect 18844 76414 18846 76466
rect 18846 76414 18898 76466
rect 18898 76414 18900 76466
rect 18844 76412 18900 76414
rect 20188 76412 20244 76468
rect 20748 76354 20804 76356
rect 20748 76302 20750 76354
rect 20750 76302 20802 76354
rect 20802 76302 20804 76354
rect 20748 76300 20804 76302
rect 19404 75458 19460 75460
rect 19404 75406 19406 75458
rect 19406 75406 19458 75458
rect 19458 75406 19460 75458
rect 19404 75404 19460 75406
rect 18508 74786 18564 74788
rect 18508 74734 18510 74786
rect 18510 74734 18562 74786
rect 18562 74734 18564 74786
rect 18508 74732 18564 74734
rect 18396 74284 18452 74340
rect 17948 73948 18004 74004
rect 14008 72154 14064 72156
rect 14112 72154 14168 72156
rect 14008 72102 14024 72154
rect 14024 72102 14064 72154
rect 14112 72102 14148 72154
rect 14148 72102 14168 72154
rect 14008 72100 14064 72102
rect 14112 72100 14168 72102
rect 14216 72100 14272 72156
rect 14320 72154 14376 72156
rect 14424 72154 14480 72156
rect 14528 72154 14584 72156
rect 14320 72102 14324 72154
rect 14324 72102 14376 72154
rect 14424 72102 14448 72154
rect 14448 72102 14480 72154
rect 14528 72102 14572 72154
rect 14572 72102 14584 72154
rect 14320 72100 14376 72102
rect 14424 72100 14480 72102
rect 14528 72100 14584 72102
rect 14632 72154 14688 72156
rect 14736 72154 14792 72156
rect 14840 72154 14896 72156
rect 14632 72102 14644 72154
rect 14644 72102 14688 72154
rect 14736 72102 14768 72154
rect 14768 72102 14792 72154
rect 14840 72102 14892 72154
rect 14892 72102 14896 72154
rect 14632 72100 14688 72102
rect 14736 72100 14792 72102
rect 14840 72100 14896 72102
rect 14944 72100 15000 72156
rect 15048 72154 15104 72156
rect 15152 72154 15208 72156
rect 15048 72102 15068 72154
rect 15068 72102 15104 72154
rect 15152 72102 15192 72154
rect 15192 72102 15208 72154
rect 15048 72100 15104 72102
rect 15152 72100 15208 72102
rect 15932 73554 15988 73556
rect 15932 73502 15934 73554
rect 15934 73502 15986 73554
rect 15986 73502 15988 73554
rect 15932 73500 15988 73502
rect 15260 71090 15316 71092
rect 15260 71038 15262 71090
rect 15262 71038 15314 71090
rect 15314 71038 15316 71090
rect 15260 71036 15316 71038
rect 15932 71036 15988 71092
rect 15260 70812 15316 70868
rect 14008 70586 14064 70588
rect 14112 70586 14168 70588
rect 14008 70534 14024 70586
rect 14024 70534 14064 70586
rect 14112 70534 14148 70586
rect 14148 70534 14168 70586
rect 14008 70532 14064 70534
rect 14112 70532 14168 70534
rect 14216 70532 14272 70588
rect 14320 70586 14376 70588
rect 14424 70586 14480 70588
rect 14528 70586 14584 70588
rect 14320 70534 14324 70586
rect 14324 70534 14376 70586
rect 14424 70534 14448 70586
rect 14448 70534 14480 70586
rect 14528 70534 14572 70586
rect 14572 70534 14584 70586
rect 14320 70532 14376 70534
rect 14424 70532 14480 70534
rect 14528 70532 14584 70534
rect 14632 70586 14688 70588
rect 14736 70586 14792 70588
rect 14840 70586 14896 70588
rect 14632 70534 14644 70586
rect 14644 70534 14688 70586
rect 14736 70534 14768 70586
rect 14768 70534 14792 70586
rect 14840 70534 14892 70586
rect 14892 70534 14896 70586
rect 14632 70532 14688 70534
rect 14736 70532 14792 70534
rect 14840 70532 14896 70534
rect 14944 70532 15000 70588
rect 15048 70586 15104 70588
rect 15152 70586 15208 70588
rect 15048 70534 15068 70586
rect 15068 70534 15104 70586
rect 15152 70534 15192 70586
rect 15192 70534 15208 70586
rect 15048 70532 15104 70534
rect 15152 70532 15208 70534
rect 15036 70364 15092 70420
rect 18284 73500 18340 73556
rect 18732 73500 18788 73556
rect 20524 75458 20580 75460
rect 20524 75406 20526 75458
rect 20526 75406 20578 75458
rect 20578 75406 20580 75458
rect 20524 75404 20580 75406
rect 19516 74338 19572 74340
rect 19516 74286 19518 74338
rect 19518 74286 19570 74338
rect 19570 74286 19572 74338
rect 19516 74284 19572 74286
rect 21980 81730 22036 81732
rect 21980 81678 21982 81730
rect 21982 81678 22034 81730
rect 22034 81678 22036 81730
rect 21980 81676 22036 81678
rect 21980 80892 22036 80948
rect 22428 82460 22484 82516
rect 22876 83298 22932 83300
rect 22876 83246 22878 83298
rect 22878 83246 22930 83298
rect 22930 83246 22932 83298
rect 22876 83244 22932 83246
rect 24556 85874 24612 85876
rect 24556 85822 24558 85874
rect 24558 85822 24610 85874
rect 24610 85822 24612 85874
rect 24556 85820 24612 85822
rect 23996 85762 24052 85764
rect 23996 85710 23998 85762
rect 23998 85710 24050 85762
rect 24050 85710 24052 85762
rect 23996 85708 24052 85710
rect 25340 85708 25396 85764
rect 24008 85482 24064 85484
rect 24112 85482 24168 85484
rect 24008 85430 24024 85482
rect 24024 85430 24064 85482
rect 24112 85430 24148 85482
rect 24148 85430 24168 85482
rect 24008 85428 24064 85430
rect 24112 85428 24168 85430
rect 24216 85428 24272 85484
rect 24320 85482 24376 85484
rect 24424 85482 24480 85484
rect 24528 85482 24584 85484
rect 24320 85430 24324 85482
rect 24324 85430 24376 85482
rect 24424 85430 24448 85482
rect 24448 85430 24480 85482
rect 24528 85430 24572 85482
rect 24572 85430 24584 85482
rect 24320 85428 24376 85430
rect 24424 85428 24480 85430
rect 24528 85428 24584 85430
rect 24632 85482 24688 85484
rect 24736 85482 24792 85484
rect 24840 85482 24896 85484
rect 24632 85430 24644 85482
rect 24644 85430 24688 85482
rect 24736 85430 24768 85482
rect 24768 85430 24792 85482
rect 24840 85430 24892 85482
rect 24892 85430 24896 85482
rect 24632 85428 24688 85430
rect 24736 85428 24792 85430
rect 24840 85428 24896 85430
rect 24944 85428 25000 85484
rect 25048 85482 25104 85484
rect 25152 85482 25208 85484
rect 25048 85430 25068 85482
rect 25068 85430 25104 85482
rect 25152 85430 25192 85482
rect 25192 85430 25208 85482
rect 25048 85428 25104 85430
rect 25152 85428 25208 85430
rect 24008 83914 24064 83916
rect 24112 83914 24168 83916
rect 24008 83862 24024 83914
rect 24024 83862 24064 83914
rect 24112 83862 24148 83914
rect 24148 83862 24168 83914
rect 24008 83860 24064 83862
rect 24112 83860 24168 83862
rect 24216 83860 24272 83916
rect 24320 83914 24376 83916
rect 24424 83914 24480 83916
rect 24528 83914 24584 83916
rect 24320 83862 24324 83914
rect 24324 83862 24376 83914
rect 24424 83862 24448 83914
rect 24448 83862 24480 83914
rect 24528 83862 24572 83914
rect 24572 83862 24584 83914
rect 24320 83860 24376 83862
rect 24424 83860 24480 83862
rect 24528 83860 24584 83862
rect 24632 83914 24688 83916
rect 24736 83914 24792 83916
rect 24840 83914 24896 83916
rect 24632 83862 24644 83914
rect 24644 83862 24688 83914
rect 24736 83862 24768 83914
rect 24768 83862 24792 83914
rect 24840 83862 24892 83914
rect 24892 83862 24896 83914
rect 24632 83860 24688 83862
rect 24736 83860 24792 83862
rect 24840 83860 24896 83862
rect 24944 83860 25000 83916
rect 25048 83914 25104 83916
rect 25152 83914 25208 83916
rect 25048 83862 25068 83914
rect 25068 83862 25104 83914
rect 25152 83862 25192 83914
rect 25192 83862 25208 83914
rect 25048 83860 25104 83862
rect 25152 83860 25208 83862
rect 23884 82684 23940 82740
rect 22540 81730 22596 81732
rect 22540 81678 22542 81730
rect 22542 81678 22594 81730
rect 22594 81678 22596 81730
rect 22540 81676 22596 81678
rect 22316 81058 22372 81060
rect 22316 81006 22318 81058
rect 22318 81006 22370 81058
rect 22370 81006 22372 81058
rect 22316 81004 22372 81006
rect 23660 81058 23716 81060
rect 23660 81006 23662 81058
rect 23662 81006 23714 81058
rect 23714 81006 23716 81058
rect 23660 81004 23716 81006
rect 20972 78428 21028 78484
rect 21196 77250 21252 77252
rect 21196 77198 21198 77250
rect 21198 77198 21250 77250
rect 21250 77198 21252 77250
rect 21196 77196 21252 77198
rect 21308 76300 21364 76356
rect 21980 78428 22036 78484
rect 21756 76636 21812 76692
rect 21868 77196 21924 77252
rect 22988 78706 23044 78708
rect 22988 78654 22990 78706
rect 22990 78654 23042 78706
rect 23042 78654 23044 78706
rect 22988 78652 23044 78654
rect 22204 78204 22260 78260
rect 22316 77196 22372 77252
rect 24556 82738 24612 82740
rect 24556 82686 24558 82738
rect 24558 82686 24610 82738
rect 24610 82686 24612 82738
rect 24556 82684 24612 82686
rect 24108 82460 24164 82516
rect 24008 82346 24064 82348
rect 24112 82346 24168 82348
rect 24008 82294 24024 82346
rect 24024 82294 24064 82346
rect 24112 82294 24148 82346
rect 24148 82294 24168 82346
rect 24008 82292 24064 82294
rect 24112 82292 24168 82294
rect 24216 82292 24272 82348
rect 24320 82346 24376 82348
rect 24424 82346 24480 82348
rect 24528 82346 24584 82348
rect 24320 82294 24324 82346
rect 24324 82294 24376 82346
rect 24424 82294 24448 82346
rect 24448 82294 24480 82346
rect 24528 82294 24572 82346
rect 24572 82294 24584 82346
rect 24320 82292 24376 82294
rect 24424 82292 24480 82294
rect 24528 82292 24584 82294
rect 24632 82346 24688 82348
rect 24736 82346 24792 82348
rect 24840 82346 24896 82348
rect 24632 82294 24644 82346
rect 24644 82294 24688 82346
rect 24736 82294 24768 82346
rect 24768 82294 24792 82346
rect 24840 82294 24892 82346
rect 24892 82294 24896 82346
rect 24632 82292 24688 82294
rect 24736 82292 24792 82294
rect 24840 82292 24896 82294
rect 24944 82292 25000 82348
rect 25048 82346 25104 82348
rect 25152 82346 25208 82348
rect 25048 82294 25068 82346
rect 25068 82294 25104 82346
rect 25152 82294 25192 82346
rect 25192 82294 25208 82346
rect 25048 82292 25104 82294
rect 25152 82292 25208 82294
rect 25788 82738 25844 82740
rect 25788 82686 25790 82738
rect 25790 82686 25842 82738
rect 25842 82686 25844 82738
rect 25788 82684 25844 82686
rect 25340 82124 25396 82180
rect 24008 80778 24064 80780
rect 24112 80778 24168 80780
rect 24008 80726 24024 80778
rect 24024 80726 24064 80778
rect 24112 80726 24148 80778
rect 24148 80726 24168 80778
rect 24008 80724 24064 80726
rect 24112 80724 24168 80726
rect 24216 80724 24272 80780
rect 24320 80778 24376 80780
rect 24424 80778 24480 80780
rect 24528 80778 24584 80780
rect 24320 80726 24324 80778
rect 24324 80726 24376 80778
rect 24424 80726 24448 80778
rect 24448 80726 24480 80778
rect 24528 80726 24572 80778
rect 24572 80726 24584 80778
rect 24320 80724 24376 80726
rect 24424 80724 24480 80726
rect 24528 80724 24584 80726
rect 24632 80778 24688 80780
rect 24736 80778 24792 80780
rect 24840 80778 24896 80780
rect 24632 80726 24644 80778
rect 24644 80726 24688 80778
rect 24736 80726 24768 80778
rect 24768 80726 24792 80778
rect 24840 80726 24892 80778
rect 24892 80726 24896 80778
rect 24632 80724 24688 80726
rect 24736 80724 24792 80726
rect 24840 80724 24896 80726
rect 24944 80724 25000 80780
rect 25048 80778 25104 80780
rect 25152 80778 25208 80780
rect 25048 80726 25068 80778
rect 25068 80726 25104 80778
rect 25152 80726 25192 80778
rect 25192 80726 25208 80778
rect 25048 80724 25104 80726
rect 25152 80724 25208 80726
rect 24008 79210 24064 79212
rect 24112 79210 24168 79212
rect 24008 79158 24024 79210
rect 24024 79158 24064 79210
rect 24112 79158 24148 79210
rect 24148 79158 24168 79210
rect 24008 79156 24064 79158
rect 24112 79156 24168 79158
rect 24216 79156 24272 79212
rect 24320 79210 24376 79212
rect 24424 79210 24480 79212
rect 24528 79210 24584 79212
rect 24320 79158 24324 79210
rect 24324 79158 24376 79210
rect 24424 79158 24448 79210
rect 24448 79158 24480 79210
rect 24528 79158 24572 79210
rect 24572 79158 24584 79210
rect 24320 79156 24376 79158
rect 24424 79156 24480 79158
rect 24528 79156 24584 79158
rect 24632 79210 24688 79212
rect 24736 79210 24792 79212
rect 24840 79210 24896 79212
rect 24632 79158 24644 79210
rect 24644 79158 24688 79210
rect 24736 79158 24768 79210
rect 24768 79158 24792 79210
rect 24840 79158 24892 79210
rect 24892 79158 24896 79210
rect 24632 79156 24688 79158
rect 24736 79156 24792 79158
rect 24840 79156 24896 79158
rect 24944 79156 25000 79212
rect 25048 79210 25104 79212
rect 25152 79210 25208 79212
rect 25048 79158 25068 79210
rect 25068 79158 25104 79210
rect 25152 79158 25192 79210
rect 25192 79158 25208 79210
rect 25048 79156 25104 79158
rect 25152 79156 25208 79158
rect 34008 95674 34064 95676
rect 34112 95674 34168 95676
rect 34008 95622 34024 95674
rect 34024 95622 34064 95674
rect 34112 95622 34148 95674
rect 34148 95622 34168 95674
rect 34008 95620 34064 95622
rect 34112 95620 34168 95622
rect 34216 95620 34272 95676
rect 34320 95674 34376 95676
rect 34424 95674 34480 95676
rect 34528 95674 34584 95676
rect 34320 95622 34324 95674
rect 34324 95622 34376 95674
rect 34424 95622 34448 95674
rect 34448 95622 34480 95674
rect 34528 95622 34572 95674
rect 34572 95622 34584 95674
rect 34320 95620 34376 95622
rect 34424 95620 34480 95622
rect 34528 95620 34584 95622
rect 34632 95674 34688 95676
rect 34736 95674 34792 95676
rect 34840 95674 34896 95676
rect 34632 95622 34644 95674
rect 34644 95622 34688 95674
rect 34736 95622 34768 95674
rect 34768 95622 34792 95674
rect 34840 95622 34892 95674
rect 34892 95622 34896 95674
rect 34632 95620 34688 95622
rect 34736 95620 34792 95622
rect 34840 95620 34896 95622
rect 34944 95620 35000 95676
rect 35048 95674 35104 95676
rect 35152 95674 35208 95676
rect 35048 95622 35068 95674
rect 35068 95622 35104 95674
rect 35152 95622 35192 95674
rect 35192 95622 35208 95674
rect 35048 95620 35104 95622
rect 35152 95620 35208 95622
rect 34008 94106 34064 94108
rect 34112 94106 34168 94108
rect 34008 94054 34024 94106
rect 34024 94054 34064 94106
rect 34112 94054 34148 94106
rect 34148 94054 34168 94106
rect 34008 94052 34064 94054
rect 34112 94052 34168 94054
rect 34216 94052 34272 94108
rect 34320 94106 34376 94108
rect 34424 94106 34480 94108
rect 34528 94106 34584 94108
rect 34320 94054 34324 94106
rect 34324 94054 34376 94106
rect 34424 94054 34448 94106
rect 34448 94054 34480 94106
rect 34528 94054 34572 94106
rect 34572 94054 34584 94106
rect 34320 94052 34376 94054
rect 34424 94052 34480 94054
rect 34528 94052 34584 94054
rect 34632 94106 34688 94108
rect 34736 94106 34792 94108
rect 34840 94106 34896 94108
rect 34632 94054 34644 94106
rect 34644 94054 34688 94106
rect 34736 94054 34768 94106
rect 34768 94054 34792 94106
rect 34840 94054 34892 94106
rect 34892 94054 34896 94106
rect 34632 94052 34688 94054
rect 34736 94052 34792 94054
rect 34840 94052 34896 94054
rect 34944 94052 35000 94108
rect 35048 94106 35104 94108
rect 35152 94106 35208 94108
rect 35048 94054 35068 94106
rect 35068 94054 35104 94106
rect 35152 94054 35192 94106
rect 35192 94054 35208 94106
rect 35048 94052 35104 94054
rect 35152 94052 35208 94054
rect 34008 92538 34064 92540
rect 34112 92538 34168 92540
rect 34008 92486 34024 92538
rect 34024 92486 34064 92538
rect 34112 92486 34148 92538
rect 34148 92486 34168 92538
rect 34008 92484 34064 92486
rect 34112 92484 34168 92486
rect 34216 92484 34272 92540
rect 34320 92538 34376 92540
rect 34424 92538 34480 92540
rect 34528 92538 34584 92540
rect 34320 92486 34324 92538
rect 34324 92486 34376 92538
rect 34424 92486 34448 92538
rect 34448 92486 34480 92538
rect 34528 92486 34572 92538
rect 34572 92486 34584 92538
rect 34320 92484 34376 92486
rect 34424 92484 34480 92486
rect 34528 92484 34584 92486
rect 34632 92538 34688 92540
rect 34736 92538 34792 92540
rect 34840 92538 34896 92540
rect 34632 92486 34644 92538
rect 34644 92486 34688 92538
rect 34736 92486 34768 92538
rect 34768 92486 34792 92538
rect 34840 92486 34892 92538
rect 34892 92486 34896 92538
rect 34632 92484 34688 92486
rect 34736 92484 34792 92486
rect 34840 92484 34896 92486
rect 34944 92484 35000 92540
rect 35048 92538 35104 92540
rect 35152 92538 35208 92540
rect 35048 92486 35068 92538
rect 35068 92486 35104 92538
rect 35152 92486 35192 92538
rect 35192 92486 35208 92538
rect 35048 92484 35104 92486
rect 35152 92484 35208 92486
rect 34008 90970 34064 90972
rect 34112 90970 34168 90972
rect 34008 90918 34024 90970
rect 34024 90918 34064 90970
rect 34112 90918 34148 90970
rect 34148 90918 34168 90970
rect 34008 90916 34064 90918
rect 34112 90916 34168 90918
rect 34216 90916 34272 90972
rect 34320 90970 34376 90972
rect 34424 90970 34480 90972
rect 34528 90970 34584 90972
rect 34320 90918 34324 90970
rect 34324 90918 34376 90970
rect 34424 90918 34448 90970
rect 34448 90918 34480 90970
rect 34528 90918 34572 90970
rect 34572 90918 34584 90970
rect 34320 90916 34376 90918
rect 34424 90916 34480 90918
rect 34528 90916 34584 90918
rect 34632 90970 34688 90972
rect 34736 90970 34792 90972
rect 34840 90970 34896 90972
rect 34632 90918 34644 90970
rect 34644 90918 34688 90970
rect 34736 90918 34768 90970
rect 34768 90918 34792 90970
rect 34840 90918 34892 90970
rect 34892 90918 34896 90970
rect 34632 90916 34688 90918
rect 34736 90916 34792 90918
rect 34840 90916 34896 90918
rect 34944 90916 35000 90972
rect 35048 90970 35104 90972
rect 35152 90970 35208 90972
rect 35048 90918 35068 90970
rect 35068 90918 35104 90970
rect 35152 90918 35192 90970
rect 35192 90918 35208 90970
rect 35048 90916 35104 90918
rect 35152 90916 35208 90918
rect 34008 89402 34064 89404
rect 34112 89402 34168 89404
rect 34008 89350 34024 89402
rect 34024 89350 34064 89402
rect 34112 89350 34148 89402
rect 34148 89350 34168 89402
rect 34008 89348 34064 89350
rect 34112 89348 34168 89350
rect 34216 89348 34272 89404
rect 34320 89402 34376 89404
rect 34424 89402 34480 89404
rect 34528 89402 34584 89404
rect 34320 89350 34324 89402
rect 34324 89350 34376 89402
rect 34424 89350 34448 89402
rect 34448 89350 34480 89402
rect 34528 89350 34572 89402
rect 34572 89350 34584 89402
rect 34320 89348 34376 89350
rect 34424 89348 34480 89350
rect 34528 89348 34584 89350
rect 34632 89402 34688 89404
rect 34736 89402 34792 89404
rect 34840 89402 34896 89404
rect 34632 89350 34644 89402
rect 34644 89350 34688 89402
rect 34736 89350 34768 89402
rect 34768 89350 34792 89402
rect 34840 89350 34892 89402
rect 34892 89350 34896 89402
rect 34632 89348 34688 89350
rect 34736 89348 34792 89350
rect 34840 89348 34896 89350
rect 34944 89348 35000 89404
rect 35048 89402 35104 89404
rect 35152 89402 35208 89404
rect 35048 89350 35068 89402
rect 35068 89350 35104 89402
rect 35152 89350 35192 89402
rect 35192 89350 35208 89402
rect 35048 89348 35104 89350
rect 35152 89348 35208 89350
rect 34008 87834 34064 87836
rect 34112 87834 34168 87836
rect 34008 87782 34024 87834
rect 34024 87782 34064 87834
rect 34112 87782 34148 87834
rect 34148 87782 34168 87834
rect 34008 87780 34064 87782
rect 34112 87780 34168 87782
rect 34216 87780 34272 87836
rect 34320 87834 34376 87836
rect 34424 87834 34480 87836
rect 34528 87834 34584 87836
rect 34320 87782 34324 87834
rect 34324 87782 34376 87834
rect 34424 87782 34448 87834
rect 34448 87782 34480 87834
rect 34528 87782 34572 87834
rect 34572 87782 34584 87834
rect 34320 87780 34376 87782
rect 34424 87780 34480 87782
rect 34528 87780 34584 87782
rect 34632 87834 34688 87836
rect 34736 87834 34792 87836
rect 34840 87834 34896 87836
rect 34632 87782 34644 87834
rect 34644 87782 34688 87834
rect 34736 87782 34768 87834
rect 34768 87782 34792 87834
rect 34840 87782 34892 87834
rect 34892 87782 34896 87834
rect 34632 87780 34688 87782
rect 34736 87780 34792 87782
rect 34840 87780 34896 87782
rect 34944 87780 35000 87836
rect 35048 87834 35104 87836
rect 35152 87834 35208 87836
rect 35048 87782 35068 87834
rect 35068 87782 35104 87834
rect 35152 87782 35192 87834
rect 35192 87782 35208 87834
rect 35048 87780 35104 87782
rect 35152 87780 35208 87782
rect 34008 86266 34064 86268
rect 34112 86266 34168 86268
rect 34008 86214 34024 86266
rect 34024 86214 34064 86266
rect 34112 86214 34148 86266
rect 34148 86214 34168 86266
rect 34008 86212 34064 86214
rect 34112 86212 34168 86214
rect 34216 86212 34272 86268
rect 34320 86266 34376 86268
rect 34424 86266 34480 86268
rect 34528 86266 34584 86268
rect 34320 86214 34324 86266
rect 34324 86214 34376 86266
rect 34424 86214 34448 86266
rect 34448 86214 34480 86266
rect 34528 86214 34572 86266
rect 34572 86214 34584 86266
rect 34320 86212 34376 86214
rect 34424 86212 34480 86214
rect 34528 86212 34584 86214
rect 34632 86266 34688 86268
rect 34736 86266 34792 86268
rect 34840 86266 34896 86268
rect 34632 86214 34644 86266
rect 34644 86214 34688 86266
rect 34736 86214 34768 86266
rect 34768 86214 34792 86266
rect 34840 86214 34892 86266
rect 34892 86214 34896 86266
rect 34632 86212 34688 86214
rect 34736 86212 34792 86214
rect 34840 86212 34896 86214
rect 34944 86212 35000 86268
rect 35048 86266 35104 86268
rect 35152 86266 35208 86268
rect 35048 86214 35068 86266
rect 35068 86214 35104 86266
rect 35152 86214 35192 86266
rect 35192 86214 35208 86266
rect 35048 86212 35104 86214
rect 35152 86212 35208 86214
rect 34008 84698 34064 84700
rect 34112 84698 34168 84700
rect 34008 84646 34024 84698
rect 34024 84646 34064 84698
rect 34112 84646 34148 84698
rect 34148 84646 34168 84698
rect 34008 84644 34064 84646
rect 34112 84644 34168 84646
rect 34216 84644 34272 84700
rect 34320 84698 34376 84700
rect 34424 84698 34480 84700
rect 34528 84698 34584 84700
rect 34320 84646 34324 84698
rect 34324 84646 34376 84698
rect 34424 84646 34448 84698
rect 34448 84646 34480 84698
rect 34528 84646 34572 84698
rect 34572 84646 34584 84698
rect 34320 84644 34376 84646
rect 34424 84644 34480 84646
rect 34528 84644 34584 84646
rect 34632 84698 34688 84700
rect 34736 84698 34792 84700
rect 34840 84698 34896 84700
rect 34632 84646 34644 84698
rect 34644 84646 34688 84698
rect 34736 84646 34768 84698
rect 34768 84646 34792 84698
rect 34840 84646 34892 84698
rect 34892 84646 34896 84698
rect 34632 84644 34688 84646
rect 34736 84644 34792 84646
rect 34840 84644 34896 84646
rect 34944 84644 35000 84700
rect 35048 84698 35104 84700
rect 35152 84698 35208 84700
rect 35048 84646 35068 84698
rect 35068 84646 35104 84698
rect 35152 84646 35192 84698
rect 35192 84646 35208 84698
rect 35048 84644 35104 84646
rect 35152 84644 35208 84646
rect 34008 83130 34064 83132
rect 34112 83130 34168 83132
rect 34008 83078 34024 83130
rect 34024 83078 34064 83130
rect 34112 83078 34148 83130
rect 34148 83078 34168 83130
rect 34008 83076 34064 83078
rect 34112 83076 34168 83078
rect 34216 83076 34272 83132
rect 34320 83130 34376 83132
rect 34424 83130 34480 83132
rect 34528 83130 34584 83132
rect 34320 83078 34324 83130
rect 34324 83078 34376 83130
rect 34424 83078 34448 83130
rect 34448 83078 34480 83130
rect 34528 83078 34572 83130
rect 34572 83078 34584 83130
rect 34320 83076 34376 83078
rect 34424 83076 34480 83078
rect 34528 83076 34584 83078
rect 34632 83130 34688 83132
rect 34736 83130 34792 83132
rect 34840 83130 34896 83132
rect 34632 83078 34644 83130
rect 34644 83078 34688 83130
rect 34736 83078 34768 83130
rect 34768 83078 34792 83130
rect 34840 83078 34892 83130
rect 34892 83078 34896 83130
rect 34632 83076 34688 83078
rect 34736 83076 34792 83078
rect 34840 83076 34896 83078
rect 34944 83076 35000 83132
rect 35048 83130 35104 83132
rect 35152 83130 35208 83132
rect 35048 83078 35068 83130
rect 35068 83078 35104 83130
rect 35152 83078 35192 83130
rect 35192 83078 35208 83130
rect 35048 83076 35104 83078
rect 35152 83076 35208 83078
rect 34008 81562 34064 81564
rect 34112 81562 34168 81564
rect 34008 81510 34024 81562
rect 34024 81510 34064 81562
rect 34112 81510 34148 81562
rect 34148 81510 34168 81562
rect 34008 81508 34064 81510
rect 34112 81508 34168 81510
rect 34216 81508 34272 81564
rect 34320 81562 34376 81564
rect 34424 81562 34480 81564
rect 34528 81562 34584 81564
rect 34320 81510 34324 81562
rect 34324 81510 34376 81562
rect 34424 81510 34448 81562
rect 34448 81510 34480 81562
rect 34528 81510 34572 81562
rect 34572 81510 34584 81562
rect 34320 81508 34376 81510
rect 34424 81508 34480 81510
rect 34528 81508 34584 81510
rect 34632 81562 34688 81564
rect 34736 81562 34792 81564
rect 34840 81562 34896 81564
rect 34632 81510 34644 81562
rect 34644 81510 34688 81562
rect 34736 81510 34768 81562
rect 34768 81510 34792 81562
rect 34840 81510 34892 81562
rect 34892 81510 34896 81562
rect 34632 81508 34688 81510
rect 34736 81508 34792 81510
rect 34840 81508 34896 81510
rect 34944 81508 35000 81564
rect 35048 81562 35104 81564
rect 35152 81562 35208 81564
rect 35048 81510 35068 81562
rect 35068 81510 35104 81562
rect 35152 81510 35192 81562
rect 35192 81510 35208 81562
rect 35048 81508 35104 81510
rect 35152 81508 35208 81510
rect 34008 79994 34064 79996
rect 34112 79994 34168 79996
rect 34008 79942 34024 79994
rect 34024 79942 34064 79994
rect 34112 79942 34148 79994
rect 34148 79942 34168 79994
rect 34008 79940 34064 79942
rect 34112 79940 34168 79942
rect 34216 79940 34272 79996
rect 34320 79994 34376 79996
rect 34424 79994 34480 79996
rect 34528 79994 34584 79996
rect 34320 79942 34324 79994
rect 34324 79942 34376 79994
rect 34424 79942 34448 79994
rect 34448 79942 34480 79994
rect 34528 79942 34572 79994
rect 34572 79942 34584 79994
rect 34320 79940 34376 79942
rect 34424 79940 34480 79942
rect 34528 79940 34584 79942
rect 34632 79994 34688 79996
rect 34736 79994 34792 79996
rect 34840 79994 34896 79996
rect 34632 79942 34644 79994
rect 34644 79942 34688 79994
rect 34736 79942 34768 79994
rect 34768 79942 34792 79994
rect 34840 79942 34892 79994
rect 34892 79942 34896 79994
rect 34632 79940 34688 79942
rect 34736 79940 34792 79942
rect 34840 79940 34896 79942
rect 34944 79940 35000 79996
rect 35048 79994 35104 79996
rect 35152 79994 35208 79996
rect 35048 79942 35068 79994
rect 35068 79942 35104 79994
rect 35152 79942 35192 79994
rect 35192 79942 35208 79994
rect 35048 79940 35104 79942
rect 35152 79940 35208 79942
rect 23884 78204 23940 78260
rect 23436 76524 23492 76580
rect 24332 78428 24388 78484
rect 19404 73500 19460 73556
rect 20636 73442 20692 73444
rect 20636 73390 20638 73442
rect 20638 73390 20690 73442
rect 20690 73390 20692 73442
rect 20636 73388 20692 73390
rect 19852 71820 19908 71876
rect 19292 70978 19348 70980
rect 19292 70926 19294 70978
rect 19294 70926 19346 70978
rect 19346 70926 19348 70978
rect 19292 70924 19348 70926
rect 13804 69692 13860 69748
rect 14252 69580 14308 69636
rect 14812 69580 14868 69636
rect 14028 69298 14084 69300
rect 14028 69246 14030 69298
rect 14030 69246 14082 69298
rect 14082 69246 14084 69298
rect 14028 69244 14084 69246
rect 14924 69522 14980 69524
rect 14924 69470 14926 69522
rect 14926 69470 14978 69522
rect 14978 69470 14980 69522
rect 14924 69468 14980 69470
rect 13916 69132 13972 69188
rect 15036 69132 15092 69188
rect 14008 69018 14064 69020
rect 14112 69018 14168 69020
rect 14008 68966 14024 69018
rect 14024 68966 14064 69018
rect 14112 68966 14148 69018
rect 14148 68966 14168 69018
rect 14008 68964 14064 68966
rect 14112 68964 14168 68966
rect 14216 68964 14272 69020
rect 14320 69018 14376 69020
rect 14424 69018 14480 69020
rect 14528 69018 14584 69020
rect 14320 68966 14324 69018
rect 14324 68966 14376 69018
rect 14424 68966 14448 69018
rect 14448 68966 14480 69018
rect 14528 68966 14572 69018
rect 14572 68966 14584 69018
rect 14320 68964 14376 68966
rect 14424 68964 14480 68966
rect 14528 68964 14584 68966
rect 14632 69018 14688 69020
rect 14736 69018 14792 69020
rect 14840 69018 14896 69020
rect 14632 68966 14644 69018
rect 14644 68966 14688 69018
rect 14736 68966 14768 69018
rect 14768 68966 14792 69018
rect 14840 68966 14892 69018
rect 14892 68966 14896 69018
rect 14632 68964 14688 68966
rect 14736 68964 14792 68966
rect 14840 68964 14896 68966
rect 14944 68964 15000 69020
rect 15048 69018 15104 69020
rect 15152 69018 15208 69020
rect 15048 68966 15068 69018
rect 15068 68966 15104 69018
rect 15152 68966 15192 69018
rect 15192 68966 15208 69018
rect 15048 68964 15104 68966
rect 15152 68964 15208 68966
rect 15596 69468 15652 69524
rect 15708 69580 15764 69636
rect 15484 69356 15540 69412
rect 16044 70306 16100 70308
rect 16044 70254 16046 70306
rect 16046 70254 16098 70306
rect 16098 70254 16100 70306
rect 16044 70252 16100 70254
rect 15260 68684 15316 68740
rect 14476 67842 14532 67844
rect 14476 67790 14478 67842
rect 14478 67790 14530 67842
rect 14530 67790 14532 67842
rect 14476 67788 14532 67790
rect 14028 67730 14084 67732
rect 14028 67678 14030 67730
rect 14030 67678 14082 67730
rect 14082 67678 14084 67730
rect 14028 67676 14084 67678
rect 14588 67676 14644 67732
rect 14252 67564 14308 67620
rect 14812 67618 14868 67620
rect 14812 67566 14814 67618
rect 14814 67566 14866 67618
rect 14866 67566 14868 67618
rect 14812 67564 14868 67566
rect 14008 67450 14064 67452
rect 14112 67450 14168 67452
rect 14008 67398 14024 67450
rect 14024 67398 14064 67450
rect 14112 67398 14148 67450
rect 14148 67398 14168 67450
rect 14008 67396 14064 67398
rect 14112 67396 14168 67398
rect 14216 67396 14272 67452
rect 14320 67450 14376 67452
rect 14424 67450 14480 67452
rect 14528 67450 14584 67452
rect 14320 67398 14324 67450
rect 14324 67398 14376 67450
rect 14424 67398 14448 67450
rect 14448 67398 14480 67450
rect 14528 67398 14572 67450
rect 14572 67398 14584 67450
rect 14320 67396 14376 67398
rect 14424 67396 14480 67398
rect 14528 67396 14584 67398
rect 14632 67450 14688 67452
rect 14736 67450 14792 67452
rect 14840 67450 14896 67452
rect 14632 67398 14644 67450
rect 14644 67398 14688 67450
rect 14736 67398 14768 67450
rect 14768 67398 14792 67450
rect 14840 67398 14892 67450
rect 14892 67398 14896 67450
rect 14632 67396 14688 67398
rect 14736 67396 14792 67398
rect 14840 67396 14896 67398
rect 14944 67396 15000 67452
rect 15048 67450 15104 67452
rect 15152 67450 15208 67452
rect 15048 67398 15068 67450
rect 15068 67398 15104 67450
rect 15152 67398 15192 67450
rect 15192 67398 15208 67450
rect 15048 67396 15104 67398
rect 15152 67396 15208 67398
rect 14924 67228 14980 67284
rect 13916 67170 13972 67172
rect 13916 67118 13918 67170
rect 13918 67118 13970 67170
rect 13970 67118 13972 67170
rect 13916 67116 13972 67118
rect 15820 69186 15876 69188
rect 15820 69134 15822 69186
rect 15822 69134 15874 69186
rect 15874 69134 15876 69186
rect 15820 69132 15876 69134
rect 15596 67676 15652 67732
rect 15708 68908 15764 68964
rect 16044 68796 16100 68852
rect 16156 69468 16212 69524
rect 15820 68684 15876 68740
rect 16492 70140 16548 70196
rect 16492 69356 16548 69412
rect 16268 68572 16324 68628
rect 16492 68684 16548 68740
rect 16716 70194 16772 70196
rect 16716 70142 16718 70194
rect 16718 70142 16770 70194
rect 16770 70142 16772 70194
rect 16716 70140 16772 70142
rect 16604 69020 16660 69076
rect 16156 67564 16212 67620
rect 16268 68012 16324 68068
rect 15932 67116 15988 67172
rect 14008 65882 14064 65884
rect 14112 65882 14168 65884
rect 14008 65830 14024 65882
rect 14024 65830 14064 65882
rect 14112 65830 14148 65882
rect 14148 65830 14168 65882
rect 14008 65828 14064 65830
rect 14112 65828 14168 65830
rect 14216 65828 14272 65884
rect 14320 65882 14376 65884
rect 14424 65882 14480 65884
rect 14528 65882 14584 65884
rect 14320 65830 14324 65882
rect 14324 65830 14376 65882
rect 14424 65830 14448 65882
rect 14448 65830 14480 65882
rect 14528 65830 14572 65882
rect 14572 65830 14584 65882
rect 14320 65828 14376 65830
rect 14424 65828 14480 65830
rect 14528 65828 14584 65830
rect 14632 65882 14688 65884
rect 14736 65882 14792 65884
rect 14840 65882 14896 65884
rect 14632 65830 14644 65882
rect 14644 65830 14688 65882
rect 14736 65830 14768 65882
rect 14768 65830 14792 65882
rect 14840 65830 14892 65882
rect 14892 65830 14896 65882
rect 14632 65828 14688 65830
rect 14736 65828 14792 65830
rect 14840 65828 14896 65830
rect 14944 65828 15000 65884
rect 15048 65882 15104 65884
rect 15152 65882 15208 65884
rect 15048 65830 15068 65882
rect 15068 65830 15104 65882
rect 15152 65830 15192 65882
rect 15192 65830 15208 65882
rect 15048 65828 15104 65830
rect 15152 65828 15208 65830
rect 13580 65324 13636 65380
rect 13916 65212 13972 65268
rect 14028 65324 14084 65380
rect 13244 64876 13300 64932
rect 13132 64652 13188 64708
rect 12572 64428 12628 64484
rect 12460 62972 12516 63028
rect 12348 62860 12404 62916
rect 12124 61852 12180 61908
rect 12348 61292 12404 61348
rect 11340 61180 11396 61236
rect 12908 62524 12964 62580
rect 13132 63922 13188 63924
rect 13132 63870 13134 63922
rect 13134 63870 13186 63922
rect 13186 63870 13188 63922
rect 13132 63868 13188 63870
rect 12796 62412 12852 62468
rect 12796 62076 12852 62132
rect 13468 64594 13524 64596
rect 13468 64542 13470 64594
rect 13470 64542 13522 64594
rect 13522 64542 13524 64594
rect 13468 64540 13524 64542
rect 13804 65100 13860 65156
rect 13916 64876 13972 64932
rect 14140 65100 14196 65156
rect 14588 64652 14644 64708
rect 13244 62300 13300 62356
rect 13356 62412 13412 62468
rect 13132 61852 13188 61908
rect 12684 60620 12740 60676
rect 14812 64876 14868 64932
rect 14700 64540 14756 64596
rect 16492 67730 16548 67732
rect 16492 67678 16494 67730
rect 16494 67678 16546 67730
rect 16546 67678 16548 67730
rect 16492 67676 16548 67678
rect 16716 68514 16772 68516
rect 16716 68462 16718 68514
rect 16718 68462 16770 68514
rect 16770 68462 16772 68514
rect 16716 68460 16772 68462
rect 16716 67676 16772 67732
rect 16716 67058 16772 67060
rect 16716 67006 16718 67058
rect 16718 67006 16770 67058
rect 16770 67006 16772 67058
rect 16716 67004 16772 67006
rect 15820 65324 15876 65380
rect 15372 64540 15428 64596
rect 14476 64428 14532 64484
rect 14008 64314 14064 64316
rect 14112 64314 14168 64316
rect 14008 64262 14024 64314
rect 14024 64262 14064 64314
rect 14112 64262 14148 64314
rect 14148 64262 14168 64314
rect 14008 64260 14064 64262
rect 14112 64260 14168 64262
rect 14216 64260 14272 64316
rect 14320 64314 14376 64316
rect 14424 64314 14480 64316
rect 14528 64314 14584 64316
rect 14320 64262 14324 64314
rect 14324 64262 14376 64314
rect 14424 64262 14448 64314
rect 14448 64262 14480 64314
rect 14528 64262 14572 64314
rect 14572 64262 14584 64314
rect 14320 64260 14376 64262
rect 14424 64260 14480 64262
rect 14528 64260 14584 64262
rect 14632 64314 14688 64316
rect 14736 64314 14792 64316
rect 14840 64314 14896 64316
rect 14632 64262 14644 64314
rect 14644 64262 14688 64314
rect 14736 64262 14768 64314
rect 14768 64262 14792 64314
rect 14840 64262 14892 64314
rect 14892 64262 14896 64314
rect 14632 64260 14688 64262
rect 14736 64260 14792 64262
rect 14840 64260 14896 64262
rect 14944 64260 15000 64316
rect 15048 64314 15104 64316
rect 15152 64314 15208 64316
rect 15048 64262 15068 64314
rect 15068 64262 15104 64314
rect 15152 64262 15192 64314
rect 15192 64262 15208 64314
rect 15048 64260 15104 64262
rect 15152 64260 15208 64262
rect 15372 64204 15428 64260
rect 14700 64092 14756 64148
rect 15260 64092 15316 64148
rect 13804 63756 13860 63812
rect 13916 63868 13972 63924
rect 14924 63756 14980 63812
rect 13692 63644 13748 63700
rect 14252 63698 14308 63700
rect 14252 63646 14254 63698
rect 14254 63646 14306 63698
rect 14306 63646 14308 63698
rect 14252 63644 14308 63646
rect 13804 63532 13860 63588
rect 13580 63420 13636 63476
rect 13580 63250 13636 63252
rect 13580 63198 13582 63250
rect 13582 63198 13634 63250
rect 13634 63198 13636 63250
rect 13580 63196 13636 63198
rect 13580 62972 13636 63028
rect 13580 62076 13636 62132
rect 14476 63026 14532 63028
rect 14476 62974 14478 63026
rect 14478 62974 14530 63026
rect 14530 62974 14532 63026
rect 14476 62972 14532 62974
rect 15260 63026 15316 63028
rect 15260 62974 15262 63026
rect 15262 62974 15314 63026
rect 15314 62974 15316 63026
rect 15260 62972 15316 62974
rect 14028 62914 14084 62916
rect 14028 62862 14030 62914
rect 14030 62862 14082 62914
rect 14082 62862 14084 62914
rect 14028 62860 14084 62862
rect 14008 62746 14064 62748
rect 14112 62746 14168 62748
rect 13804 62636 13860 62692
rect 14008 62694 14024 62746
rect 14024 62694 14064 62746
rect 14112 62694 14148 62746
rect 14148 62694 14168 62746
rect 14008 62692 14064 62694
rect 14112 62692 14168 62694
rect 14216 62692 14272 62748
rect 14320 62746 14376 62748
rect 14424 62746 14480 62748
rect 14528 62746 14584 62748
rect 14320 62694 14324 62746
rect 14324 62694 14376 62746
rect 14424 62694 14448 62746
rect 14448 62694 14480 62746
rect 14528 62694 14572 62746
rect 14572 62694 14584 62746
rect 14320 62692 14376 62694
rect 14424 62692 14480 62694
rect 14528 62692 14584 62694
rect 14632 62746 14688 62748
rect 14736 62746 14792 62748
rect 14840 62746 14896 62748
rect 14632 62694 14644 62746
rect 14644 62694 14688 62746
rect 14736 62694 14768 62746
rect 14768 62694 14792 62746
rect 14840 62694 14892 62746
rect 14892 62694 14896 62746
rect 14632 62692 14688 62694
rect 14736 62692 14792 62694
rect 14840 62692 14896 62694
rect 14944 62692 15000 62748
rect 15048 62746 15104 62748
rect 15152 62746 15208 62748
rect 15048 62694 15068 62746
rect 15068 62694 15104 62746
rect 15152 62694 15192 62746
rect 15192 62694 15208 62746
rect 15048 62692 15104 62694
rect 15152 62692 15208 62694
rect 14364 62578 14420 62580
rect 14364 62526 14366 62578
rect 14366 62526 14418 62578
rect 14418 62526 14420 62578
rect 14364 62524 14420 62526
rect 14588 62412 14644 62468
rect 14924 62354 14980 62356
rect 14924 62302 14926 62354
rect 14926 62302 14978 62354
rect 14978 62302 14980 62354
rect 14924 62300 14980 62302
rect 13916 62188 13972 62244
rect 13804 61628 13860 61684
rect 15596 63922 15652 63924
rect 15596 63870 15598 63922
rect 15598 63870 15650 63922
rect 15650 63870 15652 63922
rect 15596 63868 15652 63870
rect 15372 62354 15428 62356
rect 15372 62302 15374 62354
rect 15374 62302 15426 62354
rect 15426 62302 15428 62354
rect 15372 62300 15428 62302
rect 16156 64930 16212 64932
rect 16156 64878 16158 64930
rect 16158 64878 16210 64930
rect 16210 64878 16212 64930
rect 16156 64876 16212 64878
rect 16716 64482 16772 64484
rect 16716 64430 16718 64482
rect 16718 64430 16770 64482
rect 16770 64430 16772 64482
rect 16716 64428 16772 64430
rect 16156 64034 16212 64036
rect 16156 63982 16158 64034
rect 16158 63982 16210 64034
rect 16210 63982 16212 64034
rect 16156 63980 16212 63982
rect 15820 63644 15876 63700
rect 14588 62242 14644 62244
rect 14588 62190 14590 62242
rect 14590 62190 14642 62242
rect 14642 62190 14644 62242
rect 14588 62188 14644 62190
rect 14588 61964 14644 62020
rect 15036 62188 15092 62244
rect 14924 61682 14980 61684
rect 14924 61630 14926 61682
rect 14926 61630 14978 61682
rect 14978 61630 14980 61682
rect 14924 61628 14980 61630
rect 15372 61964 15428 62020
rect 15708 62412 15764 62468
rect 16380 62972 16436 63028
rect 15932 62524 15988 62580
rect 16380 62412 16436 62468
rect 16044 62354 16100 62356
rect 16044 62302 16046 62354
rect 16046 62302 16098 62354
rect 16098 62302 16100 62354
rect 16044 62300 16100 62302
rect 15596 61852 15652 61908
rect 15484 61628 15540 61684
rect 13692 61292 13748 61348
rect 14008 61178 14064 61180
rect 14112 61178 14168 61180
rect 14008 61126 14024 61178
rect 14024 61126 14064 61178
rect 14112 61126 14148 61178
rect 14148 61126 14168 61178
rect 14008 61124 14064 61126
rect 14112 61124 14168 61126
rect 14216 61124 14272 61180
rect 14320 61178 14376 61180
rect 14424 61178 14480 61180
rect 14528 61178 14584 61180
rect 14320 61126 14324 61178
rect 14324 61126 14376 61178
rect 14424 61126 14448 61178
rect 14448 61126 14480 61178
rect 14528 61126 14572 61178
rect 14572 61126 14584 61178
rect 14320 61124 14376 61126
rect 14424 61124 14480 61126
rect 14528 61124 14584 61126
rect 14632 61178 14688 61180
rect 14736 61178 14792 61180
rect 14840 61178 14896 61180
rect 14632 61126 14644 61178
rect 14644 61126 14688 61178
rect 14736 61126 14768 61178
rect 14768 61126 14792 61178
rect 14840 61126 14892 61178
rect 14892 61126 14896 61178
rect 14632 61124 14688 61126
rect 14736 61124 14792 61126
rect 14840 61124 14896 61126
rect 14944 61124 15000 61180
rect 15048 61178 15104 61180
rect 15152 61178 15208 61180
rect 15048 61126 15068 61178
rect 15068 61126 15104 61178
rect 15152 61126 15192 61178
rect 15192 61126 15208 61178
rect 15048 61124 15104 61126
rect 15152 61124 15208 61126
rect 13580 60508 13636 60564
rect 11676 60060 11732 60116
rect 11340 57596 11396 57652
rect 11788 57650 11844 57652
rect 11788 57598 11790 57650
rect 11790 57598 11842 57650
rect 11842 57598 11844 57650
rect 11788 57596 11844 57598
rect 11564 57148 11620 57204
rect 11340 56866 11396 56868
rect 11340 56814 11342 56866
rect 11342 56814 11394 56866
rect 11394 56814 11396 56866
rect 11340 56812 11396 56814
rect 11676 56978 11732 56980
rect 11676 56926 11678 56978
rect 11678 56926 11730 56978
rect 11730 56926 11732 56978
rect 11676 56924 11732 56926
rect 11340 56588 11396 56644
rect 11900 57036 11956 57092
rect 11788 56140 11844 56196
rect 11676 56082 11732 56084
rect 11676 56030 11678 56082
rect 11678 56030 11730 56082
rect 11730 56030 11732 56082
rect 11676 56028 11732 56030
rect 11676 55468 11732 55524
rect 11452 55020 11508 55076
rect 13580 59388 13636 59444
rect 13020 59330 13076 59332
rect 13020 59278 13022 59330
rect 13022 59278 13074 59330
rect 13074 59278 13076 59330
rect 13020 59276 13076 59278
rect 12572 59164 12628 59220
rect 12460 58492 12516 58548
rect 12124 56924 12180 56980
rect 12236 56476 12292 56532
rect 11340 54572 11396 54628
rect 11564 54684 11620 54740
rect 11452 54402 11508 54404
rect 11452 54350 11454 54402
rect 11454 54350 11506 54402
rect 11506 54350 11508 54402
rect 11452 54348 11508 54350
rect 11452 53676 11508 53732
rect 12012 55074 12068 55076
rect 12012 55022 12014 55074
rect 12014 55022 12066 55074
rect 12066 55022 12068 55074
rect 12012 55020 12068 55022
rect 11228 53228 11284 53284
rect 11228 52444 11284 52500
rect 11228 49810 11284 49812
rect 11228 49758 11230 49810
rect 11230 49758 11282 49810
rect 11282 49758 11284 49810
rect 11228 49756 11284 49758
rect 11228 49308 11284 49364
rect 10108 44268 10164 44324
rect 10668 47404 10724 47460
rect 10108 43708 10164 43764
rect 9996 43036 10052 43092
rect 9996 42812 10052 42868
rect 9996 42028 10052 42084
rect 10108 42140 10164 42196
rect 10556 45052 10612 45108
rect 11564 53228 11620 53284
rect 11452 52220 11508 52276
rect 11788 52668 11844 52724
rect 11788 52274 11844 52276
rect 11788 52222 11790 52274
rect 11790 52222 11842 52274
rect 11842 52222 11844 52274
rect 11788 52220 11844 52222
rect 11676 51884 11732 51940
rect 11228 47346 11284 47348
rect 11228 47294 11230 47346
rect 11230 47294 11282 47346
rect 11282 47294 11284 47346
rect 11228 47292 11284 47294
rect 11676 49756 11732 49812
rect 11564 49308 11620 49364
rect 11788 49308 11844 49364
rect 11788 48802 11844 48804
rect 11788 48750 11790 48802
rect 11790 48750 11842 48802
rect 11842 48750 11844 48802
rect 11788 48748 11844 48750
rect 11004 46620 11060 46676
rect 11676 48242 11732 48244
rect 11676 48190 11678 48242
rect 11678 48190 11730 48242
rect 11730 48190 11732 48242
rect 11676 48188 11732 48190
rect 11452 46508 11508 46564
rect 10892 45388 10948 45444
rect 10780 45052 10836 45108
rect 10556 44156 10612 44212
rect 10668 43484 10724 43540
rect 11004 44380 11060 44436
rect 10220 41244 10276 41300
rect 11004 44098 11060 44100
rect 11004 44046 11006 44098
rect 11006 44046 11058 44098
rect 11058 44046 11060 44098
rect 11004 44044 11060 44046
rect 11340 45330 11396 45332
rect 11340 45278 11342 45330
rect 11342 45278 11394 45330
rect 11394 45278 11396 45330
rect 11340 45276 11396 45278
rect 11452 44210 11508 44212
rect 11452 44158 11454 44210
rect 11454 44158 11506 44210
rect 11506 44158 11508 44210
rect 11452 44156 11508 44158
rect 11340 44044 11396 44100
rect 11116 43596 11172 43652
rect 9996 40460 10052 40516
rect 9996 39676 10052 39732
rect 10668 41804 10724 41860
rect 10668 41186 10724 41188
rect 10668 41134 10670 41186
rect 10670 41134 10722 41186
rect 10722 41134 10724 41186
rect 10668 41132 10724 41134
rect 10556 41074 10612 41076
rect 10556 41022 10558 41074
rect 10558 41022 10610 41074
rect 10610 41022 10612 41074
rect 10556 41020 10612 41022
rect 10892 42028 10948 42084
rect 9884 38220 9940 38276
rect 11116 41410 11172 41412
rect 11116 41358 11118 41410
rect 11118 41358 11170 41410
rect 11170 41358 11172 41410
rect 11116 41356 11172 41358
rect 11452 43372 11508 43428
rect 12348 57596 12404 57652
rect 12460 57372 12516 57428
rect 12460 56978 12516 56980
rect 12460 56926 12462 56978
rect 12462 56926 12514 56978
rect 12514 56926 12516 56978
rect 12460 56924 12516 56926
rect 12460 56252 12516 56308
rect 12460 55804 12516 55860
rect 12572 56364 12628 56420
rect 12796 57650 12852 57652
rect 12796 57598 12798 57650
rect 12798 57598 12850 57650
rect 12850 57598 12852 57650
rect 12796 57596 12852 57598
rect 12796 57372 12852 57428
rect 12684 56252 12740 56308
rect 13580 58546 13636 58548
rect 13580 58494 13582 58546
rect 13582 58494 13634 58546
rect 13634 58494 13636 58546
rect 13580 58492 13636 58494
rect 12908 56028 12964 56084
rect 13580 57090 13636 57092
rect 13580 57038 13582 57090
rect 13582 57038 13634 57090
rect 13634 57038 13636 57090
rect 13580 57036 13636 57038
rect 14008 59610 14064 59612
rect 14112 59610 14168 59612
rect 14008 59558 14024 59610
rect 14024 59558 14064 59610
rect 14112 59558 14148 59610
rect 14148 59558 14168 59610
rect 14008 59556 14064 59558
rect 14112 59556 14168 59558
rect 14216 59556 14272 59612
rect 14320 59610 14376 59612
rect 14424 59610 14480 59612
rect 14528 59610 14584 59612
rect 14320 59558 14324 59610
rect 14324 59558 14376 59610
rect 14424 59558 14448 59610
rect 14448 59558 14480 59610
rect 14528 59558 14572 59610
rect 14572 59558 14584 59610
rect 14320 59556 14376 59558
rect 14424 59556 14480 59558
rect 14528 59556 14584 59558
rect 14632 59610 14688 59612
rect 14736 59610 14792 59612
rect 14840 59610 14896 59612
rect 14632 59558 14644 59610
rect 14644 59558 14688 59610
rect 14736 59558 14768 59610
rect 14768 59558 14792 59610
rect 14840 59558 14892 59610
rect 14892 59558 14896 59610
rect 14632 59556 14688 59558
rect 14736 59556 14792 59558
rect 14840 59556 14896 59558
rect 14944 59556 15000 59612
rect 15048 59610 15104 59612
rect 15152 59610 15208 59612
rect 15048 59558 15068 59610
rect 15068 59558 15104 59610
rect 15152 59558 15192 59610
rect 15192 59558 15208 59610
rect 15048 59556 15104 59558
rect 15152 59556 15208 59558
rect 13916 59388 13972 59444
rect 14924 59388 14980 59444
rect 14700 58994 14756 58996
rect 14700 58942 14702 58994
rect 14702 58942 14754 58994
rect 14754 58942 14756 58994
rect 14700 58940 14756 58942
rect 14028 58828 14084 58884
rect 13916 58380 13972 58436
rect 14812 58434 14868 58436
rect 14812 58382 14814 58434
rect 14814 58382 14866 58434
rect 14866 58382 14868 58434
rect 14812 58380 14868 58382
rect 15372 59388 15428 59444
rect 15372 59218 15428 59220
rect 15372 59166 15374 59218
rect 15374 59166 15426 59218
rect 15426 59166 15428 59218
rect 15372 59164 15428 59166
rect 15036 58268 15092 58324
rect 14924 58156 14980 58212
rect 14008 58042 14064 58044
rect 14112 58042 14168 58044
rect 14008 57990 14024 58042
rect 14024 57990 14064 58042
rect 14112 57990 14148 58042
rect 14148 57990 14168 58042
rect 14008 57988 14064 57990
rect 14112 57988 14168 57990
rect 14216 57988 14272 58044
rect 14320 58042 14376 58044
rect 14424 58042 14480 58044
rect 14528 58042 14584 58044
rect 14320 57990 14324 58042
rect 14324 57990 14376 58042
rect 14424 57990 14448 58042
rect 14448 57990 14480 58042
rect 14528 57990 14572 58042
rect 14572 57990 14584 58042
rect 14320 57988 14376 57990
rect 14424 57988 14480 57990
rect 14528 57988 14584 57990
rect 14632 58042 14688 58044
rect 14736 58042 14792 58044
rect 14840 58042 14896 58044
rect 14632 57990 14644 58042
rect 14644 57990 14688 58042
rect 14736 57990 14768 58042
rect 14768 57990 14792 58042
rect 14840 57990 14892 58042
rect 14892 57990 14896 58042
rect 14632 57988 14688 57990
rect 14736 57988 14792 57990
rect 14840 57988 14896 57990
rect 14944 57988 15000 58044
rect 15048 58042 15104 58044
rect 15152 58042 15208 58044
rect 15048 57990 15068 58042
rect 15068 57990 15104 58042
rect 15152 57990 15192 58042
rect 15192 57990 15208 58042
rect 15048 57988 15104 57990
rect 15152 57988 15208 57990
rect 15932 60956 15988 61012
rect 16268 60956 16324 61012
rect 17388 69410 17444 69412
rect 17388 69358 17390 69410
rect 17390 69358 17442 69410
rect 17442 69358 17444 69410
rect 17388 69356 17444 69358
rect 17836 70028 17892 70084
rect 17948 69356 18004 69412
rect 17724 68908 17780 68964
rect 17836 69244 17892 69300
rect 16940 68572 16996 68628
rect 17052 68796 17108 68852
rect 17500 68626 17556 68628
rect 17500 68574 17502 68626
rect 17502 68574 17554 68626
rect 17554 68574 17556 68626
rect 17500 68572 17556 68574
rect 18508 70194 18564 70196
rect 18508 70142 18510 70194
rect 18510 70142 18562 70194
rect 18562 70142 18564 70194
rect 18508 70140 18564 70142
rect 19404 70082 19460 70084
rect 19404 70030 19406 70082
rect 19406 70030 19458 70082
rect 19458 70030 19460 70082
rect 19404 70028 19460 70030
rect 18172 68908 18228 68964
rect 18956 69468 19012 69524
rect 18396 69410 18452 69412
rect 18396 69358 18398 69410
rect 18398 69358 18450 69410
rect 18450 69358 18452 69410
rect 18396 69356 18452 69358
rect 18508 69298 18564 69300
rect 18508 69246 18510 69298
rect 18510 69246 18562 69298
rect 18562 69246 18564 69298
rect 18508 69244 18564 69246
rect 19404 69186 19460 69188
rect 19404 69134 19406 69186
rect 19406 69134 19458 69186
rect 19458 69134 19460 69186
rect 19404 69132 19460 69134
rect 18732 69020 18788 69076
rect 19068 68850 19124 68852
rect 19068 68798 19070 68850
rect 19070 68798 19122 68850
rect 19122 68798 19124 68850
rect 19068 68796 19124 68798
rect 17948 68514 18004 68516
rect 17948 68462 17950 68514
rect 17950 68462 18002 68514
rect 18002 68462 18004 68514
rect 17948 68460 18004 68462
rect 18172 68626 18228 68628
rect 18172 68574 18174 68626
rect 18174 68574 18226 68626
rect 18226 68574 18228 68626
rect 18172 68572 18228 68574
rect 17164 67004 17220 67060
rect 17388 67564 17444 67620
rect 17164 66274 17220 66276
rect 17164 66222 17166 66274
rect 17166 66222 17218 66274
rect 17218 66222 17220 66274
rect 17164 66220 17220 66222
rect 17164 65996 17220 66052
rect 17164 65212 17220 65268
rect 17276 64652 17332 64708
rect 16828 63026 16884 63028
rect 16828 62974 16830 63026
rect 16830 62974 16882 63026
rect 16882 62974 16884 63026
rect 16828 62972 16884 62974
rect 16604 62860 16660 62916
rect 17276 63196 17332 63252
rect 17052 62300 17108 62356
rect 17164 62636 17220 62692
rect 16940 62188 16996 62244
rect 16828 62076 16884 62132
rect 16940 61682 16996 61684
rect 16940 61630 16942 61682
rect 16942 61630 16994 61682
rect 16994 61630 16996 61682
rect 16940 61628 16996 61630
rect 16492 60732 16548 60788
rect 16156 60562 16212 60564
rect 16156 60510 16158 60562
rect 16158 60510 16210 60562
rect 16210 60510 16212 60562
rect 16156 60508 16212 60510
rect 15708 58322 15764 58324
rect 15708 58270 15710 58322
rect 15710 58270 15762 58322
rect 15762 58270 15764 58322
rect 15708 58268 15764 58270
rect 15036 57820 15092 57876
rect 13132 56812 13188 56868
rect 13804 57372 13860 57428
rect 13468 56028 13524 56084
rect 13020 55692 13076 55748
rect 12572 55468 12628 55524
rect 12348 55356 12404 55412
rect 12460 55186 12516 55188
rect 12460 55134 12462 55186
rect 12462 55134 12514 55186
rect 12514 55134 12516 55186
rect 12460 55132 12516 55134
rect 12236 53730 12292 53732
rect 12236 53678 12238 53730
rect 12238 53678 12290 53730
rect 12290 53678 12292 53730
rect 12236 53676 12292 53678
rect 13468 54124 13524 54180
rect 13692 55692 13748 55748
rect 14364 57650 14420 57652
rect 14364 57598 14366 57650
rect 14366 57598 14418 57650
rect 14418 57598 14420 57650
rect 14364 57596 14420 57598
rect 14252 57372 14308 57428
rect 14252 56866 14308 56868
rect 14252 56814 14254 56866
rect 14254 56814 14306 56866
rect 14306 56814 14308 56866
rect 14252 56812 14308 56814
rect 14364 56754 14420 56756
rect 14364 56702 14366 56754
rect 14366 56702 14418 56754
rect 14418 56702 14420 56754
rect 14364 56700 14420 56702
rect 15372 57036 15428 57092
rect 14008 56474 14064 56476
rect 14112 56474 14168 56476
rect 14008 56422 14024 56474
rect 14024 56422 14064 56474
rect 14112 56422 14148 56474
rect 14148 56422 14168 56474
rect 14008 56420 14064 56422
rect 14112 56420 14168 56422
rect 14216 56420 14272 56476
rect 14320 56474 14376 56476
rect 14424 56474 14480 56476
rect 14528 56474 14584 56476
rect 14320 56422 14324 56474
rect 14324 56422 14376 56474
rect 14424 56422 14448 56474
rect 14448 56422 14480 56474
rect 14528 56422 14572 56474
rect 14572 56422 14584 56474
rect 14320 56420 14376 56422
rect 14424 56420 14480 56422
rect 14528 56420 14584 56422
rect 14632 56474 14688 56476
rect 14736 56474 14792 56476
rect 14840 56474 14896 56476
rect 14632 56422 14644 56474
rect 14644 56422 14688 56474
rect 14736 56422 14768 56474
rect 14768 56422 14792 56474
rect 14840 56422 14892 56474
rect 14892 56422 14896 56474
rect 14632 56420 14688 56422
rect 14736 56420 14792 56422
rect 14840 56420 14896 56422
rect 14944 56420 15000 56476
rect 15048 56474 15104 56476
rect 15152 56474 15208 56476
rect 15048 56422 15068 56474
rect 15068 56422 15104 56474
rect 15152 56422 15192 56474
rect 15192 56422 15208 56474
rect 15048 56420 15104 56422
rect 15152 56420 15208 56422
rect 14028 56252 14084 56308
rect 13916 56140 13972 56196
rect 15036 56140 15092 56196
rect 14252 55970 14308 55972
rect 14252 55918 14254 55970
rect 14254 55918 14306 55970
rect 14306 55918 14308 55970
rect 14252 55916 14308 55918
rect 14588 55970 14644 55972
rect 14588 55918 14590 55970
rect 14590 55918 14642 55970
rect 14642 55918 14644 55970
rect 14588 55916 14644 55918
rect 14588 55692 14644 55748
rect 15484 55692 15540 55748
rect 14252 55356 14308 55412
rect 14028 55132 14084 55188
rect 15036 55074 15092 55076
rect 15036 55022 15038 55074
rect 15038 55022 15090 55074
rect 15090 55022 15092 55074
rect 15036 55020 15092 55022
rect 15484 55074 15540 55076
rect 15484 55022 15486 55074
rect 15486 55022 15538 55074
rect 15538 55022 15540 55074
rect 15484 55020 15540 55022
rect 14008 54906 14064 54908
rect 14112 54906 14168 54908
rect 14008 54854 14024 54906
rect 14024 54854 14064 54906
rect 14112 54854 14148 54906
rect 14148 54854 14168 54906
rect 14008 54852 14064 54854
rect 14112 54852 14168 54854
rect 14216 54852 14272 54908
rect 14320 54906 14376 54908
rect 14424 54906 14480 54908
rect 14528 54906 14584 54908
rect 14320 54854 14324 54906
rect 14324 54854 14376 54906
rect 14424 54854 14448 54906
rect 14448 54854 14480 54906
rect 14528 54854 14572 54906
rect 14572 54854 14584 54906
rect 14320 54852 14376 54854
rect 14424 54852 14480 54854
rect 14528 54852 14584 54854
rect 14632 54906 14688 54908
rect 14736 54906 14792 54908
rect 14840 54906 14896 54908
rect 14632 54854 14644 54906
rect 14644 54854 14688 54906
rect 14736 54854 14768 54906
rect 14768 54854 14792 54906
rect 14840 54854 14892 54906
rect 14892 54854 14896 54906
rect 14632 54852 14688 54854
rect 14736 54852 14792 54854
rect 14840 54852 14896 54854
rect 14944 54852 15000 54908
rect 15048 54906 15104 54908
rect 15152 54906 15208 54908
rect 15048 54854 15068 54906
rect 15068 54854 15104 54906
rect 15152 54854 15192 54906
rect 15192 54854 15208 54906
rect 15048 54852 15104 54854
rect 15152 54852 15208 54854
rect 13692 54684 13748 54740
rect 14364 54684 14420 54740
rect 13692 54290 13748 54292
rect 13692 54238 13694 54290
rect 13694 54238 13746 54290
rect 13746 54238 13748 54290
rect 13692 54236 13748 54238
rect 12348 53452 12404 53508
rect 12572 53004 12628 53060
rect 13580 53004 13636 53060
rect 13468 52444 13524 52500
rect 12124 52162 12180 52164
rect 12124 52110 12126 52162
rect 12126 52110 12178 52162
rect 12178 52110 12180 52162
rect 12124 52108 12180 52110
rect 12572 52162 12628 52164
rect 12572 52110 12574 52162
rect 12574 52110 12626 52162
rect 12626 52110 12628 52162
rect 12572 52108 12628 52110
rect 13468 51996 13524 52052
rect 13580 50316 13636 50372
rect 12908 49196 12964 49252
rect 12796 48914 12852 48916
rect 12796 48862 12798 48914
rect 12798 48862 12850 48914
rect 12850 48862 12852 48914
rect 12796 48860 12852 48862
rect 12124 47516 12180 47572
rect 13468 49644 13524 49700
rect 13804 53900 13860 53956
rect 13916 54012 13972 54068
rect 15036 54514 15092 54516
rect 15036 54462 15038 54514
rect 15038 54462 15090 54514
rect 15090 54462 15092 54514
rect 15036 54460 15092 54462
rect 15036 54124 15092 54180
rect 14476 53900 14532 53956
rect 15036 53900 15092 53956
rect 15036 53618 15092 53620
rect 15036 53566 15038 53618
rect 15038 53566 15090 53618
rect 15090 53566 15092 53618
rect 15036 53564 15092 53566
rect 15372 54348 15428 54404
rect 16156 58322 16212 58324
rect 16156 58270 16158 58322
rect 16158 58270 16210 58322
rect 16210 58270 16212 58322
rect 16156 58268 16212 58270
rect 16044 57820 16100 57876
rect 15820 57036 15876 57092
rect 15932 55132 15988 55188
rect 16044 55020 16100 55076
rect 14008 53338 14064 53340
rect 14112 53338 14168 53340
rect 14008 53286 14024 53338
rect 14024 53286 14064 53338
rect 14112 53286 14148 53338
rect 14148 53286 14168 53338
rect 14008 53284 14064 53286
rect 14112 53284 14168 53286
rect 14216 53284 14272 53340
rect 14320 53338 14376 53340
rect 14424 53338 14480 53340
rect 14528 53338 14584 53340
rect 14320 53286 14324 53338
rect 14324 53286 14376 53338
rect 14424 53286 14448 53338
rect 14448 53286 14480 53338
rect 14528 53286 14572 53338
rect 14572 53286 14584 53338
rect 14320 53284 14376 53286
rect 14424 53284 14480 53286
rect 14528 53284 14584 53286
rect 14632 53338 14688 53340
rect 14736 53338 14792 53340
rect 14840 53338 14896 53340
rect 14632 53286 14644 53338
rect 14644 53286 14688 53338
rect 14736 53286 14768 53338
rect 14768 53286 14792 53338
rect 14840 53286 14892 53338
rect 14892 53286 14896 53338
rect 14632 53284 14688 53286
rect 14736 53284 14792 53286
rect 14840 53284 14896 53286
rect 14944 53284 15000 53340
rect 15048 53338 15104 53340
rect 15152 53338 15208 53340
rect 15048 53286 15068 53338
rect 15068 53286 15104 53338
rect 15152 53286 15192 53338
rect 15192 53286 15208 53338
rect 15048 53284 15104 53286
rect 15152 53284 15208 53286
rect 13916 52946 13972 52948
rect 13916 52894 13918 52946
rect 13918 52894 13970 52946
rect 13970 52894 13972 52946
rect 13916 52892 13972 52894
rect 14140 52892 14196 52948
rect 14140 52668 14196 52724
rect 14028 51996 14084 52052
rect 14364 51996 14420 52052
rect 15372 51996 15428 52052
rect 14008 51770 14064 51772
rect 14112 51770 14168 51772
rect 14008 51718 14024 51770
rect 14024 51718 14064 51770
rect 14112 51718 14148 51770
rect 14148 51718 14168 51770
rect 14008 51716 14064 51718
rect 14112 51716 14168 51718
rect 14216 51716 14272 51772
rect 14320 51770 14376 51772
rect 14424 51770 14480 51772
rect 14528 51770 14584 51772
rect 14320 51718 14324 51770
rect 14324 51718 14376 51770
rect 14424 51718 14448 51770
rect 14448 51718 14480 51770
rect 14528 51718 14572 51770
rect 14572 51718 14584 51770
rect 14320 51716 14376 51718
rect 14424 51716 14480 51718
rect 14528 51716 14584 51718
rect 14632 51770 14688 51772
rect 14736 51770 14792 51772
rect 14840 51770 14896 51772
rect 14632 51718 14644 51770
rect 14644 51718 14688 51770
rect 14736 51718 14768 51770
rect 14768 51718 14792 51770
rect 14840 51718 14892 51770
rect 14892 51718 14896 51770
rect 14632 51716 14688 51718
rect 14736 51716 14792 51718
rect 14840 51716 14896 51718
rect 14944 51716 15000 51772
rect 15048 51770 15104 51772
rect 15152 51770 15208 51772
rect 15048 51718 15068 51770
rect 15068 51718 15104 51770
rect 15152 51718 15192 51770
rect 15192 51718 15208 51770
rect 15048 51716 15104 51718
rect 15152 51716 15208 51718
rect 14252 51602 14308 51604
rect 14252 51550 14254 51602
rect 14254 51550 14306 51602
rect 14306 51550 14308 51602
rect 14252 51548 14308 51550
rect 13916 50370 13972 50372
rect 13916 50318 13918 50370
rect 13918 50318 13970 50370
rect 13970 50318 13972 50370
rect 13916 50316 13972 50318
rect 15484 51884 15540 51940
rect 16380 58268 16436 58324
rect 16380 56364 16436 56420
rect 16380 55298 16436 55300
rect 16380 55246 16382 55298
rect 16382 55246 16434 55298
rect 16434 55246 16436 55298
rect 16380 55244 16436 55246
rect 16268 51996 16324 52052
rect 15484 51100 15540 51156
rect 15148 50764 15204 50820
rect 14812 50428 14868 50484
rect 14364 50316 14420 50372
rect 14008 50202 14064 50204
rect 14112 50202 14168 50204
rect 14008 50150 14024 50202
rect 14024 50150 14064 50202
rect 14112 50150 14148 50202
rect 14148 50150 14168 50202
rect 14008 50148 14064 50150
rect 14112 50148 14168 50150
rect 14216 50148 14272 50204
rect 14320 50202 14376 50204
rect 14424 50202 14480 50204
rect 14528 50202 14584 50204
rect 14320 50150 14324 50202
rect 14324 50150 14376 50202
rect 14424 50150 14448 50202
rect 14448 50150 14480 50202
rect 14528 50150 14572 50202
rect 14572 50150 14584 50202
rect 14320 50148 14376 50150
rect 14424 50148 14480 50150
rect 14528 50148 14584 50150
rect 14632 50202 14688 50204
rect 14736 50202 14792 50204
rect 14840 50202 14896 50204
rect 14632 50150 14644 50202
rect 14644 50150 14688 50202
rect 14736 50150 14768 50202
rect 14768 50150 14792 50202
rect 14840 50150 14892 50202
rect 14892 50150 14896 50202
rect 14632 50148 14688 50150
rect 14736 50148 14792 50150
rect 14840 50148 14896 50150
rect 14944 50148 15000 50204
rect 15048 50202 15104 50204
rect 15152 50202 15208 50204
rect 15048 50150 15068 50202
rect 15068 50150 15104 50202
rect 15152 50150 15192 50202
rect 15192 50150 15208 50202
rect 15048 50148 15104 50150
rect 15152 50148 15208 50150
rect 15484 50540 15540 50596
rect 14252 49644 14308 49700
rect 13356 48076 13412 48132
rect 11788 46674 11844 46676
rect 11788 46622 11790 46674
rect 11790 46622 11842 46674
rect 11842 46622 11844 46674
rect 11788 46620 11844 46622
rect 11788 45890 11844 45892
rect 11788 45838 11790 45890
rect 11790 45838 11842 45890
rect 11842 45838 11844 45890
rect 11788 45836 11844 45838
rect 11788 45388 11844 45444
rect 11788 45218 11844 45220
rect 11788 45166 11790 45218
rect 11790 45166 11842 45218
rect 11842 45166 11844 45218
rect 11788 45164 11844 45166
rect 11676 44380 11732 44436
rect 11676 42924 11732 42980
rect 13244 46956 13300 47012
rect 13132 45836 13188 45892
rect 13132 45052 13188 45108
rect 12572 44044 12628 44100
rect 12348 43484 12404 43540
rect 12908 44434 12964 44436
rect 12908 44382 12910 44434
rect 12910 44382 12962 44434
rect 12962 44382 12964 44434
rect 12908 44380 12964 44382
rect 13692 48802 13748 48804
rect 13692 48750 13694 48802
rect 13694 48750 13746 48802
rect 13746 48750 13748 48802
rect 13692 48748 13748 48750
rect 13580 48636 13636 48692
rect 13580 47570 13636 47572
rect 13580 47518 13582 47570
rect 13582 47518 13634 47570
rect 13634 47518 13636 47570
rect 13580 47516 13636 47518
rect 13580 47292 13636 47348
rect 13916 49026 13972 49028
rect 13916 48974 13918 49026
rect 13918 48974 13970 49026
rect 13970 48974 13972 49026
rect 13916 48972 13972 48974
rect 15708 50316 15764 50372
rect 15932 50372 15988 50428
rect 15708 49698 15764 49700
rect 15708 49646 15710 49698
rect 15710 49646 15762 49698
rect 15762 49646 15764 49698
rect 15708 49644 15764 49646
rect 15932 49644 15988 49700
rect 14252 48860 14308 48916
rect 14700 48860 14756 48916
rect 15372 48972 15428 49028
rect 15372 48748 15428 48804
rect 14008 48634 14064 48636
rect 14112 48634 14168 48636
rect 14008 48582 14024 48634
rect 14024 48582 14064 48634
rect 14112 48582 14148 48634
rect 14148 48582 14168 48634
rect 14008 48580 14064 48582
rect 14112 48580 14168 48582
rect 14216 48580 14272 48636
rect 14320 48634 14376 48636
rect 14424 48634 14480 48636
rect 14528 48634 14584 48636
rect 14320 48582 14324 48634
rect 14324 48582 14376 48634
rect 14424 48582 14448 48634
rect 14448 48582 14480 48634
rect 14528 48582 14572 48634
rect 14572 48582 14584 48634
rect 14320 48580 14376 48582
rect 14424 48580 14480 48582
rect 14528 48580 14584 48582
rect 14632 48634 14688 48636
rect 14736 48634 14792 48636
rect 14840 48634 14896 48636
rect 14632 48582 14644 48634
rect 14644 48582 14688 48634
rect 14736 48582 14768 48634
rect 14768 48582 14792 48634
rect 14840 48582 14892 48634
rect 14892 48582 14896 48634
rect 14632 48580 14688 48582
rect 14736 48580 14792 48582
rect 14840 48580 14896 48582
rect 14944 48580 15000 48636
rect 15048 48634 15104 48636
rect 15152 48634 15208 48636
rect 15048 48582 15068 48634
rect 15068 48582 15104 48634
rect 15152 48582 15192 48634
rect 15192 48582 15208 48634
rect 15048 48580 15104 48582
rect 15152 48580 15208 48582
rect 15596 48748 15652 48804
rect 14588 48076 14644 48132
rect 15372 48076 15428 48132
rect 13916 47404 13972 47460
rect 14700 47180 14756 47236
rect 14008 47066 14064 47068
rect 14112 47066 14168 47068
rect 14008 47014 14024 47066
rect 14024 47014 14064 47066
rect 14112 47014 14148 47066
rect 14148 47014 14168 47066
rect 14008 47012 14064 47014
rect 14112 47012 14168 47014
rect 14216 47012 14272 47068
rect 14320 47066 14376 47068
rect 14424 47066 14480 47068
rect 14528 47066 14584 47068
rect 14320 47014 14324 47066
rect 14324 47014 14376 47066
rect 14424 47014 14448 47066
rect 14448 47014 14480 47066
rect 14528 47014 14572 47066
rect 14572 47014 14584 47066
rect 14320 47012 14376 47014
rect 14424 47012 14480 47014
rect 14528 47012 14584 47014
rect 14632 47066 14688 47068
rect 14736 47066 14792 47068
rect 14840 47066 14896 47068
rect 14632 47014 14644 47066
rect 14644 47014 14688 47066
rect 14736 47014 14768 47066
rect 14768 47014 14792 47066
rect 14840 47014 14892 47066
rect 14892 47014 14896 47066
rect 14632 47012 14688 47014
rect 14736 47012 14792 47014
rect 14840 47012 14896 47014
rect 14944 47012 15000 47068
rect 15048 47066 15104 47068
rect 15152 47066 15208 47068
rect 15048 47014 15068 47066
rect 15068 47014 15104 47066
rect 15152 47014 15192 47066
rect 15192 47014 15208 47066
rect 15048 47012 15104 47014
rect 15152 47012 15208 47014
rect 13916 46844 13972 46900
rect 13804 45890 13860 45892
rect 13804 45838 13806 45890
rect 13806 45838 13858 45890
rect 13858 45838 13860 45890
rect 13804 45836 13860 45838
rect 13692 45330 13748 45332
rect 13692 45278 13694 45330
rect 13694 45278 13746 45330
rect 13746 45278 13748 45330
rect 13692 45276 13748 45278
rect 14008 45498 14064 45500
rect 14112 45498 14168 45500
rect 14008 45446 14024 45498
rect 14024 45446 14064 45498
rect 14112 45446 14148 45498
rect 14148 45446 14168 45498
rect 14008 45444 14064 45446
rect 14112 45444 14168 45446
rect 14216 45444 14272 45500
rect 14320 45498 14376 45500
rect 14424 45498 14480 45500
rect 14528 45498 14584 45500
rect 14320 45446 14324 45498
rect 14324 45446 14376 45498
rect 14424 45446 14448 45498
rect 14448 45446 14480 45498
rect 14528 45446 14572 45498
rect 14572 45446 14584 45498
rect 14320 45444 14376 45446
rect 14424 45444 14480 45446
rect 14528 45444 14584 45446
rect 14632 45498 14688 45500
rect 14736 45498 14792 45500
rect 14840 45498 14896 45500
rect 14632 45446 14644 45498
rect 14644 45446 14688 45498
rect 14736 45446 14768 45498
rect 14768 45446 14792 45498
rect 14840 45446 14892 45498
rect 14892 45446 14896 45498
rect 14632 45444 14688 45446
rect 14736 45444 14792 45446
rect 14840 45444 14896 45446
rect 14944 45444 15000 45500
rect 15048 45498 15104 45500
rect 15152 45498 15208 45500
rect 15048 45446 15068 45498
rect 15068 45446 15104 45498
rect 15152 45446 15192 45498
rect 15192 45446 15208 45498
rect 15048 45444 15104 45446
rect 15152 45444 15208 45446
rect 13804 45106 13860 45108
rect 13804 45054 13806 45106
rect 13806 45054 13858 45106
rect 13858 45054 13860 45106
rect 13804 45052 13860 45054
rect 13692 44828 13748 44884
rect 13804 44716 13860 44772
rect 13468 44380 13524 44436
rect 12796 43372 12852 43428
rect 11564 41970 11620 41972
rect 11564 41918 11566 41970
rect 11566 41918 11618 41970
rect 11618 41918 11620 41970
rect 11564 41916 11620 41918
rect 10780 39730 10836 39732
rect 10780 39678 10782 39730
rect 10782 39678 10834 39730
rect 10834 39678 10836 39730
rect 10780 39676 10836 39678
rect 11228 39730 11284 39732
rect 11228 39678 11230 39730
rect 11230 39678 11282 39730
rect 11282 39678 11284 39730
rect 11228 39676 11284 39678
rect 11228 39004 11284 39060
rect 11340 38834 11396 38836
rect 11340 38782 11342 38834
rect 11342 38782 11394 38834
rect 11394 38782 11396 38834
rect 11340 38780 11396 38782
rect 8988 36482 9044 36484
rect 8988 36430 8990 36482
rect 8990 36430 9042 36482
rect 9042 36430 9044 36482
rect 8988 36428 9044 36430
rect 8652 35810 8708 35812
rect 8652 35758 8654 35810
rect 8654 35758 8706 35810
rect 8706 35758 8708 35810
rect 8652 35756 8708 35758
rect 8652 35586 8708 35588
rect 8652 35534 8654 35586
rect 8654 35534 8706 35586
rect 8706 35534 8708 35586
rect 8652 35532 8708 35534
rect 9548 36370 9604 36372
rect 9548 36318 9550 36370
rect 9550 36318 9602 36370
rect 9602 36318 9604 36370
rect 9548 36316 9604 36318
rect 9100 35868 9156 35924
rect 8764 35308 8820 35364
rect 9660 35810 9716 35812
rect 9660 35758 9662 35810
rect 9662 35758 9714 35810
rect 9714 35758 9716 35810
rect 9660 35756 9716 35758
rect 9548 35420 9604 35476
rect 8988 34748 9044 34804
rect 9436 35196 9492 35252
rect 10444 37100 10500 37156
rect 10332 36482 10388 36484
rect 10332 36430 10334 36482
rect 10334 36430 10386 36482
rect 10386 36430 10388 36482
rect 10332 36428 10388 36430
rect 10332 35420 10388 35476
rect 9996 35308 10052 35364
rect 9884 35084 9940 35140
rect 9772 34860 9828 34916
rect 8316 33292 8372 33348
rect 8652 33852 8708 33908
rect 8316 33122 8372 33124
rect 8316 33070 8318 33122
rect 8318 33070 8370 33122
rect 8370 33070 8372 33122
rect 8316 33068 8372 33070
rect 7980 32562 8036 32564
rect 7980 32510 7982 32562
rect 7982 32510 8034 32562
rect 8034 32510 8036 32562
rect 7980 32508 8036 32510
rect 7980 31836 8036 31892
rect 7308 30210 7364 30212
rect 7308 30158 7310 30210
rect 7310 30158 7362 30210
rect 7362 30158 7364 30210
rect 7308 30156 7364 30158
rect 7532 30268 7588 30324
rect 7084 29596 7140 29652
rect 7420 29260 7476 29316
rect 6748 27580 6804 27636
rect 6636 26796 6692 26852
rect 6972 27244 7028 27300
rect 7084 28588 7140 28644
rect 6076 25506 6132 25508
rect 6076 25454 6078 25506
rect 6078 25454 6130 25506
rect 6130 25454 6132 25506
rect 6076 25452 6132 25454
rect 6300 25452 6356 25508
rect 6188 23436 6244 23492
rect 5404 22092 5460 22148
rect 4008 21194 4064 21196
rect 4112 21194 4168 21196
rect 4008 21142 4024 21194
rect 4024 21142 4064 21194
rect 4112 21142 4148 21194
rect 4148 21142 4168 21194
rect 4008 21140 4064 21142
rect 4112 21140 4168 21142
rect 4216 21140 4272 21196
rect 4320 21194 4376 21196
rect 4424 21194 4480 21196
rect 4528 21194 4584 21196
rect 4320 21142 4324 21194
rect 4324 21142 4376 21194
rect 4424 21142 4448 21194
rect 4448 21142 4480 21194
rect 4528 21142 4572 21194
rect 4572 21142 4584 21194
rect 4320 21140 4376 21142
rect 4424 21140 4480 21142
rect 4528 21140 4584 21142
rect 4632 21194 4688 21196
rect 4736 21194 4792 21196
rect 4840 21194 4896 21196
rect 4632 21142 4644 21194
rect 4644 21142 4688 21194
rect 4736 21142 4768 21194
rect 4768 21142 4792 21194
rect 4840 21142 4892 21194
rect 4892 21142 4896 21194
rect 4632 21140 4688 21142
rect 4736 21140 4792 21142
rect 4840 21140 4896 21142
rect 4944 21140 5000 21196
rect 5048 21194 5104 21196
rect 5152 21194 5208 21196
rect 5048 21142 5068 21194
rect 5068 21142 5104 21194
rect 5152 21142 5192 21194
rect 5192 21142 5208 21194
rect 5048 21140 5104 21142
rect 5152 21140 5208 21142
rect 4508 21026 4564 21028
rect 4508 20974 4510 21026
rect 4510 20974 4562 21026
rect 4562 20974 4564 21026
rect 4508 20972 4564 20974
rect 4620 20802 4676 20804
rect 4620 20750 4622 20802
rect 4622 20750 4674 20802
rect 4674 20750 4676 20802
rect 4620 20748 4676 20750
rect 5404 20748 5460 20804
rect 5516 20636 5572 20692
rect 6076 22092 6132 22148
rect 5628 21532 5684 21588
rect 5068 20578 5124 20580
rect 5068 20526 5070 20578
rect 5070 20526 5122 20578
rect 5122 20526 5124 20578
rect 5068 20524 5124 20526
rect 6188 21644 6244 21700
rect 7980 30268 8036 30324
rect 7868 30156 7924 30212
rect 7756 29986 7812 29988
rect 7756 29934 7758 29986
rect 7758 29934 7810 29986
rect 7810 29934 7812 29986
rect 7756 29932 7812 29934
rect 7868 28588 7924 28644
rect 7084 27020 7140 27076
rect 7308 26908 7364 26964
rect 7084 26796 7140 26852
rect 7196 26290 7252 26292
rect 7196 26238 7198 26290
rect 7198 26238 7250 26290
rect 7250 26238 7252 26290
rect 7196 26236 7252 26238
rect 7196 25900 7252 25956
rect 6636 24668 6692 24724
rect 6412 23548 6468 23604
rect 6412 23436 6468 23492
rect 6412 21532 6468 21588
rect 4008 19626 4064 19628
rect 4112 19626 4168 19628
rect 4008 19574 4024 19626
rect 4024 19574 4064 19626
rect 4112 19574 4148 19626
rect 4148 19574 4168 19626
rect 4008 19572 4064 19574
rect 4112 19572 4168 19574
rect 4216 19572 4272 19628
rect 4320 19626 4376 19628
rect 4424 19626 4480 19628
rect 4528 19626 4584 19628
rect 4320 19574 4324 19626
rect 4324 19574 4376 19626
rect 4424 19574 4448 19626
rect 4448 19574 4480 19626
rect 4528 19574 4572 19626
rect 4572 19574 4584 19626
rect 4320 19572 4376 19574
rect 4424 19572 4480 19574
rect 4528 19572 4584 19574
rect 4632 19626 4688 19628
rect 4736 19626 4792 19628
rect 4840 19626 4896 19628
rect 4632 19574 4644 19626
rect 4644 19574 4688 19626
rect 4736 19574 4768 19626
rect 4768 19574 4792 19626
rect 4840 19574 4892 19626
rect 4892 19574 4896 19626
rect 4632 19572 4688 19574
rect 4736 19572 4792 19574
rect 4840 19572 4896 19574
rect 4944 19572 5000 19628
rect 5048 19626 5104 19628
rect 5152 19626 5208 19628
rect 5048 19574 5068 19626
rect 5068 19574 5104 19626
rect 5152 19574 5192 19626
rect 5192 19574 5208 19626
rect 5048 19572 5104 19574
rect 5152 19572 5208 19574
rect 4008 18058 4064 18060
rect 4112 18058 4168 18060
rect 4008 18006 4024 18058
rect 4024 18006 4064 18058
rect 4112 18006 4148 18058
rect 4148 18006 4168 18058
rect 4008 18004 4064 18006
rect 4112 18004 4168 18006
rect 4216 18004 4272 18060
rect 4320 18058 4376 18060
rect 4424 18058 4480 18060
rect 4528 18058 4584 18060
rect 4320 18006 4324 18058
rect 4324 18006 4376 18058
rect 4424 18006 4448 18058
rect 4448 18006 4480 18058
rect 4528 18006 4572 18058
rect 4572 18006 4584 18058
rect 4320 18004 4376 18006
rect 4424 18004 4480 18006
rect 4528 18004 4584 18006
rect 4632 18058 4688 18060
rect 4736 18058 4792 18060
rect 4840 18058 4896 18060
rect 4632 18006 4644 18058
rect 4644 18006 4688 18058
rect 4736 18006 4768 18058
rect 4768 18006 4792 18058
rect 4840 18006 4892 18058
rect 4892 18006 4896 18058
rect 4632 18004 4688 18006
rect 4736 18004 4792 18006
rect 4840 18004 4896 18006
rect 4944 18004 5000 18060
rect 5048 18058 5104 18060
rect 5152 18058 5208 18060
rect 5048 18006 5068 18058
rect 5068 18006 5104 18058
rect 5152 18006 5192 18058
rect 5192 18006 5208 18058
rect 5048 18004 5104 18006
rect 5152 18004 5208 18006
rect 4172 17890 4228 17892
rect 4172 17838 4174 17890
rect 4174 17838 4226 17890
rect 4226 17838 4228 17890
rect 4172 17836 4228 17838
rect 3836 17724 3892 17780
rect 3164 14700 3220 14756
rect 1932 13468 1988 13524
rect 3612 13916 3668 13972
rect 2380 11564 2436 11620
rect 3388 11618 3444 11620
rect 3388 11566 3390 11618
rect 3390 11566 3442 11618
rect 3442 11566 3444 11618
rect 3388 11564 3444 11566
rect 3500 7980 3556 8036
rect 3500 6860 3556 6916
rect 4956 17554 5012 17556
rect 4956 17502 4958 17554
rect 4958 17502 5010 17554
rect 5010 17502 5012 17554
rect 4956 17500 5012 17502
rect 4620 16882 4676 16884
rect 4620 16830 4622 16882
rect 4622 16830 4674 16882
rect 4674 16830 4676 16882
rect 4620 16828 4676 16830
rect 3948 16770 4004 16772
rect 3948 16718 3950 16770
rect 3950 16718 4002 16770
rect 4002 16718 4004 16770
rect 3948 16716 4004 16718
rect 5404 16828 5460 16884
rect 4732 16604 4788 16660
rect 4008 16490 4064 16492
rect 4112 16490 4168 16492
rect 4008 16438 4024 16490
rect 4024 16438 4064 16490
rect 4112 16438 4148 16490
rect 4148 16438 4168 16490
rect 4008 16436 4064 16438
rect 4112 16436 4168 16438
rect 4216 16436 4272 16492
rect 4320 16490 4376 16492
rect 4424 16490 4480 16492
rect 4528 16490 4584 16492
rect 4320 16438 4324 16490
rect 4324 16438 4376 16490
rect 4424 16438 4448 16490
rect 4448 16438 4480 16490
rect 4528 16438 4572 16490
rect 4572 16438 4584 16490
rect 4320 16436 4376 16438
rect 4424 16436 4480 16438
rect 4528 16436 4584 16438
rect 4632 16490 4688 16492
rect 4736 16490 4792 16492
rect 4840 16490 4896 16492
rect 4632 16438 4644 16490
rect 4644 16438 4688 16490
rect 4736 16438 4768 16490
rect 4768 16438 4792 16490
rect 4840 16438 4892 16490
rect 4892 16438 4896 16490
rect 4632 16436 4688 16438
rect 4736 16436 4792 16438
rect 4840 16436 4896 16438
rect 4944 16436 5000 16492
rect 5048 16490 5104 16492
rect 5152 16490 5208 16492
rect 5048 16438 5068 16490
rect 5068 16438 5104 16490
rect 5152 16438 5192 16490
rect 5192 16438 5208 16490
rect 5048 16436 5104 16438
rect 5152 16436 5208 16438
rect 3948 16156 4004 16212
rect 4732 16210 4788 16212
rect 4732 16158 4734 16210
rect 4734 16158 4786 16210
rect 4786 16158 4788 16210
rect 4732 16156 4788 16158
rect 4172 15986 4228 15988
rect 4172 15934 4174 15986
rect 4174 15934 4226 15986
rect 4226 15934 4228 15986
rect 4172 15932 4228 15934
rect 5292 15932 5348 15988
rect 4732 15596 4788 15652
rect 5740 16882 5796 16884
rect 5740 16830 5742 16882
rect 5742 16830 5794 16882
rect 5794 16830 5796 16882
rect 5740 16828 5796 16830
rect 5852 16604 5908 16660
rect 6076 20802 6132 20804
rect 6076 20750 6078 20802
rect 6078 20750 6130 20802
rect 6130 20750 6132 20802
rect 6076 20748 6132 20750
rect 6188 20690 6244 20692
rect 6188 20638 6190 20690
rect 6190 20638 6242 20690
rect 6242 20638 6244 20690
rect 6188 20636 6244 20638
rect 6188 20242 6244 20244
rect 6188 20190 6190 20242
rect 6190 20190 6242 20242
rect 6242 20190 6244 20242
rect 6188 20188 6244 20190
rect 6412 18732 6468 18788
rect 6076 16716 6132 16772
rect 6188 16828 6244 16884
rect 5964 16268 6020 16324
rect 5740 15932 5796 15988
rect 5852 15538 5908 15540
rect 5852 15486 5854 15538
rect 5854 15486 5906 15538
rect 5906 15486 5908 15538
rect 5852 15484 5908 15486
rect 5628 15148 5684 15204
rect 4008 14922 4064 14924
rect 4112 14922 4168 14924
rect 4008 14870 4024 14922
rect 4024 14870 4064 14922
rect 4112 14870 4148 14922
rect 4148 14870 4168 14922
rect 4008 14868 4064 14870
rect 4112 14868 4168 14870
rect 4216 14868 4272 14924
rect 4320 14922 4376 14924
rect 4424 14922 4480 14924
rect 4528 14922 4584 14924
rect 4320 14870 4324 14922
rect 4324 14870 4376 14922
rect 4424 14870 4448 14922
rect 4448 14870 4480 14922
rect 4528 14870 4572 14922
rect 4572 14870 4584 14922
rect 4320 14868 4376 14870
rect 4424 14868 4480 14870
rect 4528 14868 4584 14870
rect 4632 14922 4688 14924
rect 4736 14922 4792 14924
rect 4840 14922 4896 14924
rect 4632 14870 4644 14922
rect 4644 14870 4688 14922
rect 4736 14870 4768 14922
rect 4768 14870 4792 14922
rect 4840 14870 4892 14922
rect 4892 14870 4896 14922
rect 4632 14868 4688 14870
rect 4736 14868 4792 14870
rect 4840 14868 4896 14870
rect 4944 14868 5000 14924
rect 5048 14922 5104 14924
rect 5152 14922 5208 14924
rect 5048 14870 5068 14922
rect 5068 14870 5104 14922
rect 5152 14870 5192 14922
rect 5192 14870 5208 14922
rect 5048 14868 5104 14870
rect 5152 14868 5208 14870
rect 4060 14754 4116 14756
rect 4060 14702 4062 14754
rect 4062 14702 4114 14754
rect 4114 14702 4116 14754
rect 4060 14700 4116 14702
rect 4732 14418 4788 14420
rect 4732 14366 4734 14418
rect 4734 14366 4786 14418
rect 4786 14366 4788 14418
rect 4732 14364 4788 14366
rect 6076 15426 6132 15428
rect 6076 15374 6078 15426
rect 6078 15374 6130 15426
rect 6130 15374 6132 15426
rect 6076 15372 6132 15374
rect 6412 15538 6468 15540
rect 6412 15486 6414 15538
rect 6414 15486 6466 15538
rect 6466 15486 6468 15538
rect 6412 15484 6468 15486
rect 5964 14476 6020 14532
rect 5740 14252 5796 14308
rect 4008 13354 4064 13356
rect 4112 13354 4168 13356
rect 4008 13302 4024 13354
rect 4024 13302 4064 13354
rect 4112 13302 4148 13354
rect 4148 13302 4168 13354
rect 4008 13300 4064 13302
rect 4112 13300 4168 13302
rect 4216 13300 4272 13356
rect 4320 13354 4376 13356
rect 4424 13354 4480 13356
rect 4528 13354 4584 13356
rect 4320 13302 4324 13354
rect 4324 13302 4376 13354
rect 4424 13302 4448 13354
rect 4448 13302 4480 13354
rect 4528 13302 4572 13354
rect 4572 13302 4584 13354
rect 4320 13300 4376 13302
rect 4424 13300 4480 13302
rect 4528 13300 4584 13302
rect 4632 13354 4688 13356
rect 4736 13354 4792 13356
rect 4840 13354 4896 13356
rect 4632 13302 4644 13354
rect 4644 13302 4688 13354
rect 4736 13302 4768 13354
rect 4768 13302 4792 13354
rect 4840 13302 4892 13354
rect 4892 13302 4896 13354
rect 4632 13300 4688 13302
rect 4736 13300 4792 13302
rect 4840 13300 4896 13302
rect 4944 13300 5000 13356
rect 5048 13354 5104 13356
rect 5152 13354 5208 13356
rect 5048 13302 5068 13354
rect 5068 13302 5104 13354
rect 5152 13302 5192 13354
rect 5192 13302 5208 13354
rect 5048 13300 5104 13302
rect 5152 13300 5208 13302
rect 4284 13020 4340 13076
rect 4844 13074 4900 13076
rect 4844 13022 4846 13074
rect 4846 13022 4898 13074
rect 4898 13022 4900 13074
rect 4844 13020 4900 13022
rect 6188 14306 6244 14308
rect 6188 14254 6190 14306
rect 6190 14254 6242 14306
rect 6242 14254 6244 14306
rect 6188 14252 6244 14254
rect 4844 12402 4900 12404
rect 4844 12350 4846 12402
rect 4846 12350 4898 12402
rect 4898 12350 4900 12402
rect 4844 12348 4900 12350
rect 6636 23436 6692 23492
rect 6860 25282 6916 25284
rect 6860 25230 6862 25282
rect 6862 25230 6914 25282
rect 6914 25230 6916 25282
rect 6860 25228 6916 25230
rect 7196 25228 7252 25284
rect 6636 23212 6692 23268
rect 8092 29538 8148 29540
rect 8092 29486 8094 29538
rect 8094 29486 8146 29538
rect 8146 29486 8148 29538
rect 8092 29484 8148 29486
rect 8092 27916 8148 27972
rect 7756 26514 7812 26516
rect 7756 26462 7758 26514
rect 7758 26462 7810 26514
rect 7810 26462 7812 26514
rect 7756 26460 7812 26462
rect 7644 25900 7700 25956
rect 8092 26460 8148 26516
rect 7644 25676 7700 25732
rect 8092 25618 8148 25620
rect 8092 25566 8094 25618
rect 8094 25566 8146 25618
rect 8146 25566 8148 25618
rect 8092 25564 8148 25566
rect 8316 32396 8372 32452
rect 8316 28364 8372 28420
rect 8540 27916 8596 27972
rect 9884 34354 9940 34356
rect 9884 34302 9886 34354
rect 9886 34302 9938 34354
rect 9938 34302 9940 34354
rect 9884 34300 9940 34302
rect 9548 34130 9604 34132
rect 9548 34078 9550 34130
rect 9550 34078 9602 34130
rect 9602 34078 9604 34130
rect 9548 34076 9604 34078
rect 9324 33068 9380 33124
rect 8876 31890 8932 31892
rect 8876 31838 8878 31890
rect 8878 31838 8930 31890
rect 8930 31838 8932 31890
rect 8876 31836 8932 31838
rect 9996 31836 10052 31892
rect 8988 30994 9044 30996
rect 8988 30942 8990 30994
rect 8990 30942 9042 30994
rect 9042 30942 9044 30994
rect 8988 30940 9044 30942
rect 9660 30940 9716 30996
rect 8876 29484 8932 29540
rect 9772 29932 9828 29988
rect 9996 29932 10052 29988
rect 9660 29314 9716 29316
rect 9660 29262 9662 29314
rect 9662 29262 9714 29314
rect 9714 29262 9716 29314
rect 9660 29260 9716 29262
rect 9884 28700 9940 28756
rect 9548 28642 9604 28644
rect 9548 28590 9550 28642
rect 9550 28590 9602 28642
rect 9602 28590 9604 28642
rect 9548 28588 9604 28590
rect 9548 27970 9604 27972
rect 9548 27918 9550 27970
rect 9550 27918 9602 27970
rect 9602 27918 9604 27970
rect 9548 27916 9604 27918
rect 8316 27020 8372 27076
rect 8652 27468 8708 27524
rect 9324 27244 9380 27300
rect 10556 34802 10612 34804
rect 10556 34750 10558 34802
rect 10558 34750 10610 34802
rect 10610 34750 10612 34802
rect 10556 34748 10612 34750
rect 10892 36594 10948 36596
rect 10892 36542 10894 36594
rect 10894 36542 10946 36594
rect 10946 36542 10948 36594
rect 10892 36540 10948 36542
rect 10892 35474 10948 35476
rect 10892 35422 10894 35474
rect 10894 35422 10946 35474
rect 10946 35422 10948 35474
rect 10892 35420 10948 35422
rect 10892 35138 10948 35140
rect 10892 35086 10894 35138
rect 10894 35086 10946 35138
rect 10946 35086 10948 35138
rect 10892 35084 10948 35086
rect 11116 34914 11172 34916
rect 11116 34862 11118 34914
rect 11118 34862 11170 34914
rect 11170 34862 11172 34914
rect 11116 34860 11172 34862
rect 10668 34300 10724 34356
rect 11788 40572 11844 40628
rect 11452 37154 11508 37156
rect 11452 37102 11454 37154
rect 11454 37102 11506 37154
rect 11506 37102 11508 37154
rect 11452 37100 11508 37102
rect 11564 38780 11620 38836
rect 11340 36370 11396 36372
rect 11340 36318 11342 36370
rect 11342 36318 11394 36370
rect 11394 36318 11396 36370
rect 11340 36316 11396 36318
rect 11228 34748 11284 34804
rect 10780 33964 10836 34020
rect 10556 33346 10612 33348
rect 10556 33294 10558 33346
rect 10558 33294 10610 33346
rect 10610 33294 10612 33346
rect 10556 33292 10612 33294
rect 10220 31724 10276 31780
rect 12012 41186 12068 41188
rect 12012 41134 12014 41186
rect 12014 41134 12066 41186
rect 12066 41134 12068 41186
rect 12012 41132 12068 41134
rect 12348 41410 12404 41412
rect 12348 41358 12350 41410
rect 12350 41358 12402 41410
rect 12402 41358 12404 41410
rect 12348 41356 12404 41358
rect 12796 42588 12852 42644
rect 13356 43426 13412 43428
rect 13356 43374 13358 43426
rect 13358 43374 13410 43426
rect 13410 43374 13412 43426
rect 13356 43372 13412 43374
rect 12236 37266 12292 37268
rect 12236 37214 12238 37266
rect 12238 37214 12290 37266
rect 12290 37214 12292 37266
rect 12236 37212 12292 37214
rect 12124 36316 12180 36372
rect 12012 35308 12068 35364
rect 11788 34914 11844 34916
rect 11788 34862 11790 34914
rect 11790 34862 11842 34914
rect 11842 34862 11844 34914
rect 11788 34860 11844 34862
rect 11676 34802 11732 34804
rect 11676 34750 11678 34802
rect 11678 34750 11730 34802
rect 11730 34750 11732 34802
rect 11676 34748 11732 34750
rect 11676 34018 11732 34020
rect 11676 33966 11678 34018
rect 11678 33966 11730 34018
rect 11730 33966 11732 34018
rect 11676 33964 11732 33966
rect 12124 34354 12180 34356
rect 12124 34302 12126 34354
rect 12126 34302 12178 34354
rect 12178 34302 12180 34354
rect 12124 34300 12180 34302
rect 12236 33852 12292 33908
rect 12572 37378 12628 37380
rect 12572 37326 12574 37378
rect 12574 37326 12626 37378
rect 12626 37326 12628 37378
rect 12572 37324 12628 37326
rect 12796 37100 12852 37156
rect 12012 33458 12068 33460
rect 12012 33406 12014 33458
rect 12014 33406 12066 33458
rect 12066 33406 12068 33458
rect 12012 33404 12068 33406
rect 10220 30268 10276 30324
rect 10332 30044 10388 30100
rect 11340 29986 11396 29988
rect 11340 29934 11342 29986
rect 11342 29934 11394 29986
rect 11394 29934 11396 29986
rect 11340 29932 11396 29934
rect 10780 29650 10836 29652
rect 10780 29598 10782 29650
rect 10782 29598 10834 29650
rect 10834 29598 10836 29650
rect 10780 29596 10836 29598
rect 11676 30210 11732 30212
rect 11676 30158 11678 30210
rect 11678 30158 11730 30210
rect 11730 30158 11732 30210
rect 11676 30156 11732 30158
rect 11900 29426 11956 29428
rect 11900 29374 11902 29426
rect 11902 29374 11954 29426
rect 11954 29374 11956 29426
rect 11900 29372 11956 29374
rect 11564 28588 11620 28644
rect 14140 45276 14196 45332
rect 14140 45106 14196 45108
rect 14140 45054 14142 45106
rect 14142 45054 14194 45106
rect 14194 45054 14196 45106
rect 14140 45052 14196 45054
rect 14364 45052 14420 45108
rect 13580 42978 13636 42980
rect 13580 42926 13582 42978
rect 13582 42926 13634 42978
rect 13634 42926 13636 42978
rect 13580 42924 13636 42926
rect 13468 40572 13524 40628
rect 13580 42642 13636 42644
rect 13580 42590 13582 42642
rect 13582 42590 13634 42642
rect 13634 42590 13636 42642
rect 13580 42588 13636 42590
rect 13580 40236 13636 40292
rect 13356 38668 13412 38724
rect 15148 45106 15204 45108
rect 15148 45054 15150 45106
rect 15150 45054 15202 45106
rect 15202 45054 15204 45106
rect 15148 45052 15204 45054
rect 15372 45052 15428 45108
rect 14364 44716 14420 44772
rect 15372 44716 15428 44772
rect 15484 44940 15540 44996
rect 14008 43930 14064 43932
rect 14112 43930 14168 43932
rect 14008 43878 14024 43930
rect 14024 43878 14064 43930
rect 14112 43878 14148 43930
rect 14148 43878 14168 43930
rect 14008 43876 14064 43878
rect 14112 43876 14168 43878
rect 14216 43876 14272 43932
rect 14320 43930 14376 43932
rect 14424 43930 14480 43932
rect 14528 43930 14584 43932
rect 14320 43878 14324 43930
rect 14324 43878 14376 43930
rect 14424 43878 14448 43930
rect 14448 43878 14480 43930
rect 14528 43878 14572 43930
rect 14572 43878 14584 43930
rect 14320 43876 14376 43878
rect 14424 43876 14480 43878
rect 14528 43876 14584 43878
rect 14632 43930 14688 43932
rect 14736 43930 14792 43932
rect 14840 43930 14896 43932
rect 14632 43878 14644 43930
rect 14644 43878 14688 43930
rect 14736 43878 14768 43930
rect 14768 43878 14792 43930
rect 14840 43878 14892 43930
rect 14892 43878 14896 43930
rect 14632 43876 14688 43878
rect 14736 43876 14792 43878
rect 14840 43876 14896 43878
rect 14944 43876 15000 43932
rect 15048 43930 15104 43932
rect 15152 43930 15208 43932
rect 15048 43878 15068 43930
rect 15068 43878 15104 43930
rect 15152 43878 15192 43930
rect 15192 43878 15208 43930
rect 15048 43876 15104 43878
rect 15152 43876 15208 43878
rect 13916 43650 13972 43652
rect 13916 43598 13918 43650
rect 13918 43598 13970 43650
rect 13970 43598 13972 43650
rect 13916 43596 13972 43598
rect 14252 43650 14308 43652
rect 14252 43598 14254 43650
rect 14254 43598 14306 43650
rect 14306 43598 14308 43650
rect 14252 43596 14308 43598
rect 15484 43650 15540 43652
rect 15484 43598 15486 43650
rect 15486 43598 15538 43650
rect 15538 43598 15540 43650
rect 15484 43596 15540 43598
rect 14476 43538 14532 43540
rect 14476 43486 14478 43538
rect 14478 43486 14530 43538
rect 14530 43486 14532 43538
rect 14476 43484 14532 43486
rect 14140 43372 14196 43428
rect 13804 42588 13860 42644
rect 14140 42588 14196 42644
rect 14008 42362 14064 42364
rect 14112 42362 14168 42364
rect 14008 42310 14024 42362
rect 14024 42310 14064 42362
rect 14112 42310 14148 42362
rect 14148 42310 14168 42362
rect 14008 42308 14064 42310
rect 14112 42308 14168 42310
rect 14216 42308 14272 42364
rect 14320 42362 14376 42364
rect 14424 42362 14480 42364
rect 14528 42362 14584 42364
rect 14320 42310 14324 42362
rect 14324 42310 14376 42362
rect 14424 42310 14448 42362
rect 14448 42310 14480 42362
rect 14528 42310 14572 42362
rect 14572 42310 14584 42362
rect 14320 42308 14376 42310
rect 14424 42308 14480 42310
rect 14528 42308 14584 42310
rect 14632 42362 14688 42364
rect 14736 42362 14792 42364
rect 14840 42362 14896 42364
rect 14632 42310 14644 42362
rect 14644 42310 14688 42362
rect 14736 42310 14768 42362
rect 14768 42310 14792 42362
rect 14840 42310 14892 42362
rect 14892 42310 14896 42362
rect 14632 42308 14688 42310
rect 14736 42308 14792 42310
rect 14840 42308 14896 42310
rect 14944 42308 15000 42364
rect 15048 42362 15104 42364
rect 15152 42362 15208 42364
rect 15048 42310 15068 42362
rect 15068 42310 15104 42362
rect 15152 42310 15192 42362
rect 15192 42310 15208 42362
rect 15048 42308 15104 42310
rect 15152 42308 15208 42310
rect 14008 40794 14064 40796
rect 14112 40794 14168 40796
rect 14008 40742 14024 40794
rect 14024 40742 14064 40794
rect 14112 40742 14148 40794
rect 14148 40742 14168 40794
rect 14008 40740 14064 40742
rect 14112 40740 14168 40742
rect 14216 40740 14272 40796
rect 14320 40794 14376 40796
rect 14424 40794 14480 40796
rect 14528 40794 14584 40796
rect 14320 40742 14324 40794
rect 14324 40742 14376 40794
rect 14424 40742 14448 40794
rect 14448 40742 14480 40794
rect 14528 40742 14572 40794
rect 14572 40742 14584 40794
rect 14320 40740 14376 40742
rect 14424 40740 14480 40742
rect 14528 40740 14584 40742
rect 14632 40794 14688 40796
rect 14736 40794 14792 40796
rect 14840 40794 14896 40796
rect 14632 40742 14644 40794
rect 14644 40742 14688 40794
rect 14736 40742 14768 40794
rect 14768 40742 14792 40794
rect 14840 40742 14892 40794
rect 14892 40742 14896 40794
rect 14632 40740 14688 40742
rect 14736 40740 14792 40742
rect 14840 40740 14896 40742
rect 14944 40740 15000 40796
rect 15048 40794 15104 40796
rect 15152 40794 15208 40796
rect 15048 40742 15068 40794
rect 15068 40742 15104 40794
rect 15152 40742 15192 40794
rect 15192 40742 15208 40794
rect 15048 40740 15104 40742
rect 15152 40740 15208 40742
rect 13804 40572 13860 40628
rect 14140 40626 14196 40628
rect 14140 40574 14142 40626
rect 14142 40574 14194 40626
rect 14194 40574 14196 40626
rect 14140 40572 14196 40574
rect 15148 40572 15204 40628
rect 14924 40348 14980 40404
rect 15036 40236 15092 40292
rect 14008 39226 14064 39228
rect 14112 39226 14168 39228
rect 14008 39174 14024 39226
rect 14024 39174 14064 39226
rect 14112 39174 14148 39226
rect 14148 39174 14168 39226
rect 14008 39172 14064 39174
rect 14112 39172 14168 39174
rect 14216 39172 14272 39228
rect 14320 39226 14376 39228
rect 14424 39226 14480 39228
rect 14528 39226 14584 39228
rect 14320 39174 14324 39226
rect 14324 39174 14376 39226
rect 14424 39174 14448 39226
rect 14448 39174 14480 39226
rect 14528 39174 14572 39226
rect 14572 39174 14584 39226
rect 14320 39172 14376 39174
rect 14424 39172 14480 39174
rect 14528 39172 14584 39174
rect 14632 39226 14688 39228
rect 14736 39226 14792 39228
rect 14840 39226 14896 39228
rect 14632 39174 14644 39226
rect 14644 39174 14688 39226
rect 14736 39174 14768 39226
rect 14768 39174 14792 39226
rect 14840 39174 14892 39226
rect 14892 39174 14896 39226
rect 14632 39172 14688 39174
rect 14736 39172 14792 39174
rect 14840 39172 14896 39174
rect 14944 39172 15000 39228
rect 15048 39226 15104 39228
rect 15152 39226 15208 39228
rect 15048 39174 15068 39226
rect 15068 39174 15104 39226
rect 15152 39174 15192 39226
rect 15192 39174 15208 39226
rect 15048 39172 15104 39174
rect 15152 39172 15208 39174
rect 14924 39058 14980 39060
rect 14924 39006 14926 39058
rect 14926 39006 14978 39058
rect 14978 39006 14980 39058
rect 14924 39004 14980 39006
rect 15484 38780 15540 38836
rect 15820 49026 15876 49028
rect 15820 48974 15822 49026
rect 15822 48974 15874 49026
rect 15874 48974 15876 49026
rect 15820 48972 15876 48974
rect 15932 48242 15988 48244
rect 15932 48190 15934 48242
rect 15934 48190 15986 48242
rect 15986 48190 15988 48242
rect 15932 48188 15988 48190
rect 16604 60508 16660 60564
rect 16604 58322 16660 58324
rect 16604 58270 16606 58322
rect 16606 58270 16658 58322
rect 16658 58270 16660 58322
rect 16604 58268 16660 58270
rect 17276 59388 17332 59444
rect 17612 67170 17668 67172
rect 17612 67118 17614 67170
rect 17614 67118 17666 67170
rect 17666 67118 17668 67170
rect 17612 67116 17668 67118
rect 17948 67004 18004 67060
rect 17836 66780 17892 66836
rect 17612 66050 17668 66052
rect 17612 65998 17614 66050
rect 17614 65998 17666 66050
rect 17666 65998 17668 66050
rect 17612 65996 17668 65998
rect 18172 66444 18228 66500
rect 18172 66220 18228 66276
rect 18508 66162 18564 66164
rect 18508 66110 18510 66162
rect 18510 66110 18562 66162
rect 18562 66110 18564 66162
rect 18508 66108 18564 66110
rect 18172 65212 18228 65268
rect 17612 63868 17668 63924
rect 18060 65100 18116 65156
rect 17724 61628 17780 61684
rect 17164 58434 17220 58436
rect 17164 58382 17166 58434
rect 17166 58382 17218 58434
rect 17218 58382 17220 58434
rect 17164 58380 17220 58382
rect 16828 57538 16884 57540
rect 16828 57486 16830 57538
rect 16830 57486 16882 57538
rect 16882 57486 16884 57538
rect 16828 57484 16884 57486
rect 16828 56812 16884 56868
rect 16828 56642 16884 56644
rect 16828 56590 16830 56642
rect 16830 56590 16882 56642
rect 16882 56590 16884 56642
rect 16828 56588 16884 56590
rect 17052 56028 17108 56084
rect 16828 55804 16884 55860
rect 18284 64706 18340 64708
rect 18284 64654 18286 64706
rect 18286 64654 18338 64706
rect 18338 64654 18340 64706
rect 18284 64652 18340 64654
rect 18284 64428 18340 64484
rect 18508 64428 18564 64484
rect 18284 63922 18340 63924
rect 18284 63870 18286 63922
rect 18286 63870 18338 63922
rect 18338 63870 18340 63922
rect 18284 63868 18340 63870
rect 18172 62636 18228 62692
rect 19180 68124 19236 68180
rect 18732 66892 18788 66948
rect 19740 68796 19796 68852
rect 19516 68572 19572 68628
rect 19404 67116 19460 67172
rect 18732 66220 18788 66276
rect 19180 67058 19236 67060
rect 19180 67006 19182 67058
rect 19182 67006 19234 67058
rect 19234 67006 19236 67058
rect 19180 67004 19236 67006
rect 19180 66780 19236 66836
rect 20748 68012 20804 68068
rect 20076 67618 20132 67620
rect 20076 67566 20078 67618
rect 20078 67566 20130 67618
rect 20130 67566 20132 67618
rect 20076 67564 20132 67566
rect 19180 66220 19236 66276
rect 19292 66444 19348 66500
rect 18956 65324 19012 65380
rect 19068 65212 19124 65268
rect 19180 65490 19236 65492
rect 19180 65438 19182 65490
rect 19182 65438 19234 65490
rect 19234 65438 19236 65490
rect 19180 65436 19236 65438
rect 19516 65996 19572 66052
rect 20188 66220 20244 66276
rect 19964 66108 20020 66164
rect 20636 66220 20692 66276
rect 20748 66162 20804 66164
rect 20748 66110 20750 66162
rect 20750 66110 20802 66162
rect 20802 66110 20804 66162
rect 20748 66108 20804 66110
rect 20300 65436 20356 65492
rect 20412 65660 20468 65716
rect 19740 65378 19796 65380
rect 19740 65326 19742 65378
rect 19742 65326 19794 65378
rect 19794 65326 19796 65378
rect 19740 65324 19796 65326
rect 20076 65324 20132 65380
rect 19516 65100 19572 65156
rect 18956 63868 19012 63924
rect 19068 62412 19124 62468
rect 17388 56588 17444 56644
rect 17388 56082 17444 56084
rect 17388 56030 17390 56082
rect 17390 56030 17442 56082
rect 17442 56030 17444 56082
rect 17388 56028 17444 56030
rect 16156 48972 16212 49028
rect 16828 53788 16884 53844
rect 17388 50540 17444 50596
rect 17276 50482 17332 50484
rect 17276 50430 17278 50482
rect 17278 50430 17330 50482
rect 17330 50430 17332 50482
rect 17276 50428 17332 50430
rect 17724 58156 17780 58212
rect 17612 57596 17668 57652
rect 17724 57148 17780 57204
rect 18172 58268 18228 58324
rect 18396 59442 18452 59444
rect 18396 59390 18398 59442
rect 18398 59390 18450 59442
rect 18450 59390 18452 59442
rect 18396 59388 18452 59390
rect 18508 58434 18564 58436
rect 18508 58382 18510 58434
rect 18510 58382 18562 58434
rect 18562 58382 18564 58434
rect 18508 58380 18564 58382
rect 18396 58322 18452 58324
rect 18396 58270 18398 58322
rect 18398 58270 18450 58322
rect 18450 58270 18452 58322
rect 18396 58268 18452 58270
rect 18732 59218 18788 59220
rect 18732 59166 18734 59218
rect 18734 59166 18786 59218
rect 18786 59166 18788 59218
rect 18732 59164 18788 59166
rect 18844 58604 18900 58660
rect 19068 59500 19124 59556
rect 18956 58828 19012 58884
rect 19068 58716 19124 58772
rect 18844 58156 18900 58212
rect 18396 58044 18452 58100
rect 18172 57538 18228 57540
rect 18172 57486 18174 57538
rect 18174 57486 18226 57538
rect 18226 57486 18228 57538
rect 18172 57484 18228 57486
rect 18060 56700 18116 56756
rect 18060 55858 18116 55860
rect 18060 55806 18062 55858
rect 18062 55806 18114 55858
rect 18114 55806 18116 55858
rect 18060 55804 18116 55806
rect 17836 55692 17892 55748
rect 19068 58044 19124 58100
rect 19964 64988 20020 65044
rect 19292 64482 19348 64484
rect 19292 64430 19294 64482
rect 19294 64430 19346 64482
rect 19346 64430 19348 64482
rect 19292 64428 19348 64430
rect 19964 63980 20020 64036
rect 19404 63026 19460 63028
rect 19404 62974 19406 63026
rect 19406 62974 19458 63026
rect 19458 62974 19460 63026
rect 19404 62972 19460 62974
rect 19404 62524 19460 62580
rect 19292 62466 19348 62468
rect 19292 62414 19294 62466
rect 19294 62414 19346 62466
rect 19346 62414 19348 62466
rect 19292 62412 19348 62414
rect 19292 58828 19348 58884
rect 19516 62300 19572 62356
rect 19628 62636 19684 62692
rect 20300 65266 20356 65268
rect 20300 65214 20302 65266
rect 20302 65214 20354 65266
rect 20354 65214 20356 65266
rect 20300 65212 20356 65214
rect 20524 65100 20580 65156
rect 25228 78428 25284 78484
rect 25340 78258 25396 78260
rect 25340 78206 25342 78258
rect 25342 78206 25394 78258
rect 25394 78206 25396 78258
rect 25340 78204 25396 78206
rect 20972 67228 21028 67284
rect 21196 71596 21252 71652
rect 21532 73500 21588 73556
rect 21756 73276 21812 73332
rect 22876 73330 22932 73332
rect 22876 73278 22878 73330
rect 22878 73278 22930 73330
rect 22930 73278 22932 73330
rect 22876 73276 22932 73278
rect 23436 73164 23492 73220
rect 22652 71874 22708 71876
rect 22652 71822 22654 71874
rect 22654 71822 22706 71874
rect 22706 71822 22708 71874
rect 22652 71820 22708 71822
rect 21420 70978 21476 70980
rect 21420 70926 21422 70978
rect 21422 70926 21474 70978
rect 21474 70926 21476 70978
rect 21420 70924 21476 70926
rect 24008 77642 24064 77644
rect 24112 77642 24168 77644
rect 24008 77590 24024 77642
rect 24024 77590 24064 77642
rect 24112 77590 24148 77642
rect 24148 77590 24168 77642
rect 24008 77588 24064 77590
rect 24112 77588 24168 77590
rect 24216 77588 24272 77644
rect 24320 77642 24376 77644
rect 24424 77642 24480 77644
rect 24528 77642 24584 77644
rect 24320 77590 24324 77642
rect 24324 77590 24376 77642
rect 24424 77590 24448 77642
rect 24448 77590 24480 77642
rect 24528 77590 24572 77642
rect 24572 77590 24584 77642
rect 24320 77588 24376 77590
rect 24424 77588 24480 77590
rect 24528 77588 24584 77590
rect 24632 77642 24688 77644
rect 24736 77642 24792 77644
rect 24840 77642 24896 77644
rect 24632 77590 24644 77642
rect 24644 77590 24688 77642
rect 24736 77590 24768 77642
rect 24768 77590 24792 77642
rect 24840 77590 24892 77642
rect 24892 77590 24896 77642
rect 24632 77588 24688 77590
rect 24736 77588 24792 77590
rect 24840 77588 24896 77590
rect 24944 77588 25000 77644
rect 25048 77642 25104 77644
rect 25152 77642 25208 77644
rect 25048 77590 25068 77642
rect 25068 77590 25104 77642
rect 25152 77590 25192 77642
rect 25192 77590 25208 77642
rect 25048 77588 25104 77590
rect 25152 77588 25208 77590
rect 24780 77308 24836 77364
rect 24220 77250 24276 77252
rect 24220 77198 24222 77250
rect 24222 77198 24274 77250
rect 24274 77198 24276 77250
rect 24220 77196 24276 77198
rect 25676 77362 25732 77364
rect 25676 77310 25678 77362
rect 25678 77310 25730 77362
rect 25730 77310 25732 77362
rect 25676 77308 25732 77310
rect 24008 76074 24064 76076
rect 24112 76074 24168 76076
rect 24008 76022 24024 76074
rect 24024 76022 24064 76074
rect 24112 76022 24148 76074
rect 24148 76022 24168 76074
rect 24008 76020 24064 76022
rect 24112 76020 24168 76022
rect 24216 76020 24272 76076
rect 24320 76074 24376 76076
rect 24424 76074 24480 76076
rect 24528 76074 24584 76076
rect 24320 76022 24324 76074
rect 24324 76022 24376 76074
rect 24424 76022 24448 76074
rect 24448 76022 24480 76074
rect 24528 76022 24572 76074
rect 24572 76022 24584 76074
rect 24320 76020 24376 76022
rect 24424 76020 24480 76022
rect 24528 76020 24584 76022
rect 24632 76074 24688 76076
rect 24736 76074 24792 76076
rect 24840 76074 24896 76076
rect 24632 76022 24644 76074
rect 24644 76022 24688 76074
rect 24736 76022 24768 76074
rect 24768 76022 24792 76074
rect 24840 76022 24892 76074
rect 24892 76022 24896 76074
rect 24632 76020 24688 76022
rect 24736 76020 24792 76022
rect 24840 76020 24896 76022
rect 24944 76020 25000 76076
rect 25048 76074 25104 76076
rect 25152 76074 25208 76076
rect 25048 76022 25068 76074
rect 25068 76022 25104 76074
rect 25152 76022 25192 76074
rect 25192 76022 25208 76074
rect 25048 76020 25104 76022
rect 25152 76020 25208 76022
rect 24008 74506 24064 74508
rect 24112 74506 24168 74508
rect 24008 74454 24024 74506
rect 24024 74454 24064 74506
rect 24112 74454 24148 74506
rect 24148 74454 24168 74506
rect 24008 74452 24064 74454
rect 24112 74452 24168 74454
rect 24216 74452 24272 74508
rect 24320 74506 24376 74508
rect 24424 74506 24480 74508
rect 24528 74506 24584 74508
rect 24320 74454 24324 74506
rect 24324 74454 24376 74506
rect 24424 74454 24448 74506
rect 24448 74454 24480 74506
rect 24528 74454 24572 74506
rect 24572 74454 24584 74506
rect 24320 74452 24376 74454
rect 24424 74452 24480 74454
rect 24528 74452 24584 74454
rect 24632 74506 24688 74508
rect 24736 74506 24792 74508
rect 24840 74506 24896 74508
rect 24632 74454 24644 74506
rect 24644 74454 24688 74506
rect 24736 74454 24768 74506
rect 24768 74454 24792 74506
rect 24840 74454 24892 74506
rect 24892 74454 24896 74506
rect 24632 74452 24688 74454
rect 24736 74452 24792 74454
rect 24840 74452 24896 74454
rect 24944 74452 25000 74508
rect 25048 74506 25104 74508
rect 25152 74506 25208 74508
rect 25048 74454 25068 74506
rect 25068 74454 25104 74506
rect 25152 74454 25192 74506
rect 25192 74454 25208 74506
rect 25048 74452 25104 74454
rect 25152 74452 25208 74454
rect 23884 73388 23940 73444
rect 23436 71650 23492 71652
rect 23436 71598 23438 71650
rect 23438 71598 23490 71650
rect 23490 71598 23492 71650
rect 23436 71596 23492 71598
rect 21420 68124 21476 68180
rect 21532 67564 21588 67620
rect 21532 67116 21588 67172
rect 21196 65436 21252 65492
rect 21308 66108 21364 66164
rect 21532 65660 21588 65716
rect 20860 65324 20916 65380
rect 21084 65266 21140 65268
rect 21084 65214 21086 65266
rect 21086 65214 21138 65266
rect 21138 65214 21140 65266
rect 21084 65212 21140 65214
rect 20188 64652 20244 64708
rect 20412 63922 20468 63924
rect 20412 63870 20414 63922
rect 20414 63870 20466 63922
rect 20466 63870 20468 63922
rect 20412 63868 20468 63870
rect 19852 62636 19908 62692
rect 20076 62860 20132 62916
rect 20300 62748 20356 62804
rect 20300 62412 20356 62468
rect 20188 62300 20244 62356
rect 20636 63026 20692 63028
rect 20636 62974 20638 63026
rect 20638 62974 20690 63026
rect 20690 62974 20692 63026
rect 20636 62972 20692 62974
rect 20748 62748 20804 62804
rect 20524 62412 20580 62468
rect 21420 61292 21476 61348
rect 20524 60114 20580 60116
rect 20524 60062 20526 60114
rect 20526 60062 20578 60114
rect 20578 60062 20580 60114
rect 20524 60060 20580 60062
rect 19740 59500 19796 59556
rect 20188 59500 20244 59556
rect 19852 59442 19908 59444
rect 19852 59390 19854 59442
rect 19854 59390 19906 59442
rect 19906 59390 19908 59442
rect 19852 59388 19908 59390
rect 19516 59106 19572 59108
rect 19516 59054 19518 59106
rect 19518 59054 19570 59106
rect 19570 59054 19572 59106
rect 19516 59052 19572 59054
rect 19740 58716 19796 58772
rect 19628 58604 19684 58660
rect 19404 58492 19460 58548
rect 20188 58940 20244 58996
rect 19852 58434 19908 58436
rect 19852 58382 19854 58434
rect 19854 58382 19906 58434
rect 19906 58382 19908 58434
rect 19852 58380 19908 58382
rect 20300 58380 20356 58436
rect 18620 57650 18676 57652
rect 18620 57598 18622 57650
rect 18622 57598 18674 57650
rect 18674 57598 18676 57650
rect 18620 57596 18676 57598
rect 18620 57372 18676 57428
rect 18508 56306 18564 56308
rect 18508 56254 18510 56306
rect 18510 56254 18562 56306
rect 18562 56254 18564 56306
rect 18508 56252 18564 56254
rect 18956 56306 19012 56308
rect 18956 56254 18958 56306
rect 18958 56254 19010 56306
rect 19010 56254 19012 56306
rect 18956 56252 19012 56254
rect 18396 55186 18452 55188
rect 18396 55134 18398 55186
rect 18398 55134 18450 55186
rect 18450 55134 18452 55186
rect 18396 55132 18452 55134
rect 18172 54124 18228 54180
rect 18284 54012 18340 54068
rect 18284 53004 18340 53060
rect 17612 51266 17668 51268
rect 17612 51214 17614 51266
rect 17614 51214 17666 51266
rect 17666 51214 17668 51266
rect 17612 51212 17668 51214
rect 16492 49756 16548 49812
rect 18172 51266 18228 51268
rect 18172 51214 18174 51266
rect 18174 51214 18226 51266
rect 18226 51214 18228 51266
rect 18172 51212 18228 51214
rect 18844 55244 18900 55300
rect 18732 55186 18788 55188
rect 18732 55134 18734 55186
rect 18734 55134 18786 55186
rect 18786 55134 18788 55186
rect 18732 55132 18788 55134
rect 18956 53564 19012 53620
rect 18956 52780 19012 52836
rect 18620 50706 18676 50708
rect 18620 50654 18622 50706
rect 18622 50654 18674 50706
rect 18674 50654 18676 50706
rect 18620 50652 18676 50654
rect 19404 57650 19460 57652
rect 19404 57598 19406 57650
rect 19406 57598 19458 57650
rect 19458 57598 19460 57650
rect 19404 57596 19460 57598
rect 19180 57484 19236 57540
rect 19964 57708 20020 57764
rect 20524 59164 20580 59220
rect 20636 59052 20692 59108
rect 20748 58940 20804 58996
rect 20860 58828 20916 58884
rect 19740 57372 19796 57428
rect 19740 56754 19796 56756
rect 19740 56702 19742 56754
rect 19742 56702 19794 56754
rect 19794 56702 19796 56754
rect 19740 56700 19796 56702
rect 19852 56364 19908 56420
rect 20076 56252 20132 56308
rect 19516 55244 19572 55300
rect 19628 55132 19684 55188
rect 19628 53954 19684 53956
rect 19628 53902 19630 53954
rect 19630 53902 19682 53954
rect 19682 53902 19684 53954
rect 19628 53900 19684 53902
rect 19964 54012 20020 54068
rect 19404 53618 19460 53620
rect 19404 53566 19406 53618
rect 19406 53566 19458 53618
rect 19458 53566 19460 53618
rect 19404 53564 19460 53566
rect 19852 52556 19908 52612
rect 20076 53900 20132 53956
rect 20300 57148 20356 57204
rect 20748 57650 20804 57652
rect 20748 57598 20750 57650
rect 20750 57598 20802 57650
rect 20802 57598 20804 57650
rect 20748 57596 20804 57598
rect 20524 57538 20580 57540
rect 20524 57486 20526 57538
rect 20526 57486 20578 57538
rect 20578 57486 20580 57538
rect 20524 57484 20580 57486
rect 20748 56194 20804 56196
rect 20748 56142 20750 56194
rect 20750 56142 20802 56194
rect 20802 56142 20804 56194
rect 20748 56140 20804 56142
rect 20300 56082 20356 56084
rect 20300 56030 20302 56082
rect 20302 56030 20354 56082
rect 20354 56030 20356 56082
rect 20300 56028 20356 56030
rect 20860 55916 20916 55972
rect 21980 61292 22036 61348
rect 22204 70476 22260 70532
rect 24332 73218 24388 73220
rect 24332 73166 24334 73218
rect 24334 73166 24386 73218
rect 24386 73166 24388 73218
rect 24332 73164 24388 73166
rect 24008 72938 24064 72940
rect 24112 72938 24168 72940
rect 24008 72886 24024 72938
rect 24024 72886 24064 72938
rect 24112 72886 24148 72938
rect 24148 72886 24168 72938
rect 24008 72884 24064 72886
rect 24112 72884 24168 72886
rect 24216 72884 24272 72940
rect 24320 72938 24376 72940
rect 24424 72938 24480 72940
rect 24528 72938 24584 72940
rect 24320 72886 24324 72938
rect 24324 72886 24376 72938
rect 24424 72886 24448 72938
rect 24448 72886 24480 72938
rect 24528 72886 24572 72938
rect 24572 72886 24584 72938
rect 24320 72884 24376 72886
rect 24424 72884 24480 72886
rect 24528 72884 24584 72886
rect 24632 72938 24688 72940
rect 24736 72938 24792 72940
rect 24840 72938 24896 72940
rect 24632 72886 24644 72938
rect 24644 72886 24688 72938
rect 24736 72886 24768 72938
rect 24768 72886 24792 72938
rect 24840 72886 24892 72938
rect 24892 72886 24896 72938
rect 24632 72884 24688 72886
rect 24736 72884 24792 72886
rect 24840 72884 24896 72886
rect 24944 72884 25000 72940
rect 25048 72938 25104 72940
rect 25152 72938 25208 72940
rect 25048 72886 25068 72938
rect 25068 72886 25104 72938
rect 25152 72886 25192 72938
rect 25192 72886 25208 72938
rect 25048 72884 25104 72886
rect 25152 72884 25208 72886
rect 23548 72268 23604 72324
rect 24332 72322 24388 72324
rect 24332 72270 24334 72322
rect 24334 72270 24386 72322
rect 24386 72270 24388 72322
rect 24332 72268 24388 72270
rect 24008 71370 24064 71372
rect 24112 71370 24168 71372
rect 24008 71318 24024 71370
rect 24024 71318 24064 71370
rect 24112 71318 24148 71370
rect 24148 71318 24168 71370
rect 24008 71316 24064 71318
rect 24112 71316 24168 71318
rect 24216 71316 24272 71372
rect 24320 71370 24376 71372
rect 24424 71370 24480 71372
rect 24528 71370 24584 71372
rect 24320 71318 24324 71370
rect 24324 71318 24376 71370
rect 24424 71318 24448 71370
rect 24448 71318 24480 71370
rect 24528 71318 24572 71370
rect 24572 71318 24584 71370
rect 24320 71316 24376 71318
rect 24424 71316 24480 71318
rect 24528 71316 24584 71318
rect 24632 71370 24688 71372
rect 24736 71370 24792 71372
rect 24840 71370 24896 71372
rect 24632 71318 24644 71370
rect 24644 71318 24688 71370
rect 24736 71318 24768 71370
rect 24768 71318 24792 71370
rect 24840 71318 24892 71370
rect 24892 71318 24896 71370
rect 24632 71316 24688 71318
rect 24736 71316 24792 71318
rect 24840 71316 24896 71318
rect 24944 71316 25000 71372
rect 25048 71370 25104 71372
rect 25152 71370 25208 71372
rect 25048 71318 25068 71370
rect 25068 71318 25104 71370
rect 25152 71318 25192 71370
rect 25192 71318 25208 71370
rect 25048 71316 25104 71318
rect 25152 71316 25208 71318
rect 24220 70978 24276 70980
rect 24220 70926 24222 70978
rect 24222 70926 24274 70978
rect 24274 70926 24276 70978
rect 24220 70924 24276 70926
rect 25116 70978 25172 70980
rect 25116 70926 25118 70978
rect 25118 70926 25170 70978
rect 25170 70926 25172 70978
rect 25116 70924 25172 70926
rect 23548 70700 23604 70756
rect 23884 70476 23940 70532
rect 23772 70028 23828 70084
rect 27356 70924 27412 70980
rect 25676 70476 25732 70532
rect 24668 70082 24724 70084
rect 24668 70030 24670 70082
rect 24670 70030 24722 70082
rect 24722 70030 24724 70082
rect 24668 70028 24724 70030
rect 25564 70194 25620 70196
rect 25564 70142 25566 70194
rect 25566 70142 25618 70194
rect 25618 70142 25620 70194
rect 25564 70140 25620 70142
rect 25116 70028 25172 70084
rect 24008 69802 24064 69804
rect 24112 69802 24168 69804
rect 24008 69750 24024 69802
rect 24024 69750 24064 69802
rect 24112 69750 24148 69802
rect 24148 69750 24168 69802
rect 24008 69748 24064 69750
rect 24112 69748 24168 69750
rect 24216 69748 24272 69804
rect 24320 69802 24376 69804
rect 24424 69802 24480 69804
rect 24528 69802 24584 69804
rect 24320 69750 24324 69802
rect 24324 69750 24376 69802
rect 24424 69750 24448 69802
rect 24448 69750 24480 69802
rect 24528 69750 24572 69802
rect 24572 69750 24584 69802
rect 24320 69748 24376 69750
rect 24424 69748 24480 69750
rect 24528 69748 24584 69750
rect 24632 69802 24688 69804
rect 24736 69802 24792 69804
rect 24840 69802 24896 69804
rect 24632 69750 24644 69802
rect 24644 69750 24688 69802
rect 24736 69750 24768 69802
rect 24768 69750 24792 69802
rect 24840 69750 24892 69802
rect 24892 69750 24896 69802
rect 24632 69748 24688 69750
rect 24736 69748 24792 69750
rect 24840 69748 24896 69750
rect 24944 69748 25000 69804
rect 25048 69802 25104 69804
rect 25152 69802 25208 69804
rect 25048 69750 25068 69802
rect 25068 69750 25104 69802
rect 25152 69750 25192 69802
rect 25192 69750 25208 69802
rect 25048 69748 25104 69750
rect 25152 69748 25208 69750
rect 24556 69580 24612 69636
rect 25340 69580 25396 69636
rect 27020 70364 27076 70420
rect 25900 69468 25956 69524
rect 24220 68626 24276 68628
rect 24220 68574 24222 68626
rect 24222 68574 24274 68626
rect 24274 68574 24276 68626
rect 24220 68572 24276 68574
rect 24668 68460 24724 68516
rect 24444 68348 24500 68404
rect 24008 68234 24064 68236
rect 24112 68234 24168 68236
rect 24008 68182 24024 68234
rect 24024 68182 24064 68234
rect 24112 68182 24148 68234
rect 24148 68182 24168 68234
rect 24008 68180 24064 68182
rect 24112 68180 24168 68182
rect 24216 68180 24272 68236
rect 24320 68234 24376 68236
rect 24424 68234 24480 68236
rect 24528 68234 24584 68236
rect 24320 68182 24324 68234
rect 24324 68182 24376 68234
rect 24424 68182 24448 68234
rect 24448 68182 24480 68234
rect 24528 68182 24572 68234
rect 24572 68182 24584 68234
rect 24320 68180 24376 68182
rect 24424 68180 24480 68182
rect 24528 68180 24584 68182
rect 24632 68234 24688 68236
rect 24736 68234 24792 68236
rect 24840 68234 24896 68236
rect 24632 68182 24644 68234
rect 24644 68182 24688 68234
rect 24736 68182 24768 68234
rect 24768 68182 24792 68234
rect 24840 68182 24892 68234
rect 24892 68182 24896 68234
rect 24632 68180 24688 68182
rect 24736 68180 24792 68182
rect 24840 68180 24896 68182
rect 24944 68180 25000 68236
rect 25048 68234 25104 68236
rect 25152 68234 25208 68236
rect 25048 68182 25068 68234
rect 25068 68182 25104 68234
rect 25152 68182 25192 68234
rect 25192 68182 25208 68234
rect 25048 68180 25104 68182
rect 25152 68180 25208 68182
rect 24444 68012 24500 68068
rect 23772 66892 23828 66948
rect 22540 66780 22596 66836
rect 22540 66162 22596 66164
rect 22540 66110 22542 66162
rect 22542 66110 22594 66162
rect 22594 66110 22596 66162
rect 22540 66108 22596 66110
rect 25564 68684 25620 68740
rect 25676 68626 25732 68628
rect 25676 68574 25678 68626
rect 25678 68574 25730 68626
rect 25730 68574 25732 68626
rect 25676 68572 25732 68574
rect 25340 67228 25396 67284
rect 25228 66946 25284 66948
rect 25228 66894 25230 66946
rect 25230 66894 25282 66946
rect 25282 66894 25284 66946
rect 25228 66892 25284 66894
rect 24444 66834 24500 66836
rect 24444 66782 24446 66834
rect 24446 66782 24498 66834
rect 24498 66782 24500 66834
rect 24444 66780 24500 66782
rect 24008 66666 24064 66668
rect 24112 66666 24168 66668
rect 24008 66614 24024 66666
rect 24024 66614 24064 66666
rect 24112 66614 24148 66666
rect 24148 66614 24168 66666
rect 24008 66612 24064 66614
rect 24112 66612 24168 66614
rect 24216 66612 24272 66668
rect 24320 66666 24376 66668
rect 24424 66666 24480 66668
rect 24528 66666 24584 66668
rect 24320 66614 24324 66666
rect 24324 66614 24376 66666
rect 24424 66614 24448 66666
rect 24448 66614 24480 66666
rect 24528 66614 24572 66666
rect 24572 66614 24584 66666
rect 24320 66612 24376 66614
rect 24424 66612 24480 66614
rect 24528 66612 24584 66614
rect 24632 66666 24688 66668
rect 24736 66666 24792 66668
rect 24840 66666 24896 66668
rect 24632 66614 24644 66666
rect 24644 66614 24688 66666
rect 24736 66614 24768 66666
rect 24768 66614 24792 66666
rect 24840 66614 24892 66666
rect 24892 66614 24896 66666
rect 24632 66612 24688 66614
rect 24736 66612 24792 66614
rect 24840 66612 24896 66614
rect 24944 66612 25000 66668
rect 25048 66666 25104 66668
rect 25152 66666 25208 66668
rect 25048 66614 25068 66666
rect 25068 66614 25104 66666
rect 25152 66614 25192 66666
rect 25192 66614 25208 66666
rect 25048 66612 25104 66614
rect 25152 66612 25208 66614
rect 23884 65996 23940 66052
rect 23436 63084 23492 63140
rect 22316 62412 22372 62468
rect 22092 59388 22148 59444
rect 23436 59778 23492 59780
rect 23436 59726 23438 59778
rect 23438 59726 23490 59778
rect 23490 59726 23492 59778
rect 23436 59724 23492 59726
rect 21532 59218 21588 59220
rect 21532 59166 21534 59218
rect 21534 59166 21586 59218
rect 21586 59166 21588 59218
rect 21532 59164 21588 59166
rect 21756 59052 21812 59108
rect 20300 55132 20356 55188
rect 21644 58434 21700 58436
rect 21644 58382 21646 58434
rect 21646 58382 21698 58434
rect 21698 58382 21700 58434
rect 21644 58380 21700 58382
rect 21532 57596 21588 57652
rect 21532 56812 21588 56868
rect 22204 59106 22260 59108
rect 22204 59054 22206 59106
rect 22206 59054 22258 59106
rect 22258 59054 22260 59106
rect 22204 59052 22260 59054
rect 23772 63138 23828 63140
rect 23772 63086 23774 63138
rect 23774 63086 23826 63138
rect 23826 63086 23828 63138
rect 23772 63084 23828 63086
rect 21420 56082 21476 56084
rect 21420 56030 21422 56082
rect 21422 56030 21474 56082
rect 21474 56030 21476 56082
rect 21420 56028 21476 56030
rect 21084 55132 21140 55188
rect 21196 54738 21252 54740
rect 21196 54686 21198 54738
rect 21198 54686 21250 54738
rect 21250 54686 21252 54738
rect 21196 54684 21252 54686
rect 20188 53788 20244 53844
rect 21644 55916 21700 55972
rect 22204 56140 22260 56196
rect 23100 56700 23156 56756
rect 22428 56140 22484 56196
rect 22092 55916 22148 55972
rect 22316 56082 22372 56084
rect 22316 56030 22318 56082
rect 22318 56030 22370 56082
rect 22370 56030 22372 56082
rect 22316 56028 22372 56030
rect 22764 56306 22820 56308
rect 22764 56254 22766 56306
rect 22766 56254 22818 56306
rect 22818 56254 22820 56306
rect 22764 56252 22820 56254
rect 21756 55244 21812 55300
rect 22092 54738 22148 54740
rect 22092 54686 22094 54738
rect 22094 54686 22146 54738
rect 22146 54686 22148 54738
rect 22092 54684 22148 54686
rect 21532 53564 21588 53620
rect 21644 53676 21700 53732
rect 20412 52556 20468 52612
rect 19964 52108 20020 52164
rect 19404 52050 19460 52052
rect 19404 51998 19406 52050
rect 19406 51998 19458 52050
rect 19458 51998 19460 52050
rect 19404 51996 19460 51998
rect 20188 52050 20244 52052
rect 20188 51998 20190 52050
rect 20190 51998 20242 52050
rect 20242 51998 20244 52050
rect 20188 51996 20244 51998
rect 19852 50706 19908 50708
rect 19852 50654 19854 50706
rect 19854 50654 19906 50706
rect 19906 50654 19908 50706
rect 19852 50652 19908 50654
rect 18844 50540 18900 50596
rect 17500 49698 17556 49700
rect 17500 49646 17502 49698
rect 17502 49646 17554 49698
rect 17554 49646 17556 49698
rect 17500 49644 17556 49646
rect 17052 49026 17108 49028
rect 17052 48974 17054 49026
rect 17054 48974 17106 49026
rect 17106 48974 17108 49026
rect 17052 48972 17108 48974
rect 16716 48748 16772 48804
rect 17948 48914 18004 48916
rect 17948 48862 17950 48914
rect 17950 48862 18002 48914
rect 18002 48862 18004 48914
rect 17948 48860 18004 48862
rect 17724 48748 17780 48804
rect 19292 50482 19348 50484
rect 19292 50430 19294 50482
rect 19294 50430 19346 50482
rect 19346 50430 19348 50482
rect 19292 50428 19348 50430
rect 18956 49810 19012 49812
rect 18956 49758 18958 49810
rect 18958 49758 19010 49810
rect 19010 49758 19012 49810
rect 18956 49756 19012 49758
rect 18620 48914 18676 48916
rect 18620 48862 18622 48914
rect 18622 48862 18674 48914
rect 18674 48862 18676 48914
rect 18620 48860 18676 48862
rect 17612 47458 17668 47460
rect 17612 47406 17614 47458
rect 17614 47406 17666 47458
rect 17666 47406 17668 47458
rect 17612 47404 17668 47406
rect 16380 45836 16436 45892
rect 17276 46956 17332 47012
rect 18396 46956 18452 47012
rect 17612 46508 17668 46564
rect 18284 46732 18340 46788
rect 16604 45724 16660 45780
rect 15932 45276 15988 45332
rect 15820 45164 15876 45220
rect 15932 44828 15988 44884
rect 16380 45330 16436 45332
rect 16380 45278 16382 45330
rect 16382 45278 16434 45330
rect 16434 45278 16436 45330
rect 16380 45276 16436 45278
rect 16604 45276 16660 45332
rect 16156 43260 16212 43316
rect 15932 40402 15988 40404
rect 15932 40350 15934 40402
rect 15934 40350 15986 40402
rect 15986 40350 15988 40402
rect 15932 40348 15988 40350
rect 13244 37212 13300 37268
rect 12572 36428 12628 36484
rect 12460 35420 12516 35476
rect 12460 34748 12516 34804
rect 12460 34300 12516 34356
rect 12460 30044 12516 30100
rect 12348 29596 12404 29652
rect 12460 29484 12516 29540
rect 9884 27692 9940 27748
rect 9772 27634 9828 27636
rect 9772 27582 9774 27634
rect 9774 27582 9826 27634
rect 9826 27582 9828 27634
rect 9772 27580 9828 27582
rect 8876 27020 8932 27076
rect 8876 25676 8932 25732
rect 11564 27804 11620 27860
rect 12348 27746 12404 27748
rect 12348 27694 12350 27746
rect 12350 27694 12402 27746
rect 12402 27694 12404 27746
rect 12348 27692 12404 27694
rect 15260 38556 15316 38612
rect 14008 37658 14064 37660
rect 14112 37658 14168 37660
rect 14008 37606 14024 37658
rect 14024 37606 14064 37658
rect 14112 37606 14148 37658
rect 14148 37606 14168 37658
rect 14008 37604 14064 37606
rect 14112 37604 14168 37606
rect 14216 37604 14272 37660
rect 14320 37658 14376 37660
rect 14424 37658 14480 37660
rect 14528 37658 14584 37660
rect 14320 37606 14324 37658
rect 14324 37606 14376 37658
rect 14424 37606 14448 37658
rect 14448 37606 14480 37658
rect 14528 37606 14572 37658
rect 14572 37606 14584 37658
rect 14320 37604 14376 37606
rect 14424 37604 14480 37606
rect 14528 37604 14584 37606
rect 14632 37658 14688 37660
rect 14736 37658 14792 37660
rect 14840 37658 14896 37660
rect 14632 37606 14644 37658
rect 14644 37606 14688 37658
rect 14736 37606 14768 37658
rect 14768 37606 14792 37658
rect 14840 37606 14892 37658
rect 14892 37606 14896 37658
rect 14632 37604 14688 37606
rect 14736 37604 14792 37606
rect 14840 37604 14896 37606
rect 14944 37604 15000 37660
rect 15048 37658 15104 37660
rect 15152 37658 15208 37660
rect 15048 37606 15068 37658
rect 15068 37606 15104 37658
rect 15152 37606 15192 37658
rect 15192 37606 15208 37658
rect 15048 37604 15104 37606
rect 15152 37604 15208 37606
rect 14812 37490 14868 37492
rect 14812 37438 14814 37490
rect 14814 37438 14866 37490
rect 14866 37438 14868 37490
rect 14812 37436 14868 37438
rect 15708 37436 15764 37492
rect 14028 37378 14084 37380
rect 14028 37326 14030 37378
rect 14030 37326 14082 37378
rect 14082 37326 14084 37378
rect 14028 37324 14084 37326
rect 13692 36876 13748 36932
rect 14252 37212 14308 37268
rect 15036 36876 15092 36932
rect 13580 36482 13636 36484
rect 13580 36430 13582 36482
rect 13582 36430 13634 36482
rect 13634 36430 13636 36482
rect 13580 36428 13636 36430
rect 12908 36258 12964 36260
rect 12908 36206 12910 36258
rect 12910 36206 12962 36258
rect 12962 36206 12964 36258
rect 12908 36204 12964 36206
rect 14812 36370 14868 36372
rect 14812 36318 14814 36370
rect 14814 36318 14866 36370
rect 14866 36318 14868 36370
rect 14812 36316 14868 36318
rect 13692 36204 13748 36260
rect 13580 35756 13636 35812
rect 12796 35644 12852 35700
rect 14008 36090 14064 36092
rect 14112 36090 14168 36092
rect 14008 36038 14024 36090
rect 14024 36038 14064 36090
rect 14112 36038 14148 36090
rect 14148 36038 14168 36090
rect 14008 36036 14064 36038
rect 14112 36036 14168 36038
rect 14216 36036 14272 36092
rect 14320 36090 14376 36092
rect 14424 36090 14480 36092
rect 14528 36090 14584 36092
rect 14320 36038 14324 36090
rect 14324 36038 14376 36090
rect 14424 36038 14448 36090
rect 14448 36038 14480 36090
rect 14528 36038 14572 36090
rect 14572 36038 14584 36090
rect 14320 36036 14376 36038
rect 14424 36036 14480 36038
rect 14528 36036 14584 36038
rect 14632 36090 14688 36092
rect 14736 36090 14792 36092
rect 14840 36090 14896 36092
rect 14632 36038 14644 36090
rect 14644 36038 14688 36090
rect 14736 36038 14768 36090
rect 14768 36038 14792 36090
rect 14840 36038 14892 36090
rect 14892 36038 14896 36090
rect 14632 36036 14688 36038
rect 14736 36036 14792 36038
rect 14840 36036 14896 36038
rect 14944 36036 15000 36092
rect 15048 36090 15104 36092
rect 15152 36090 15208 36092
rect 15048 36038 15068 36090
rect 15068 36038 15104 36090
rect 15152 36038 15192 36090
rect 15192 36038 15208 36090
rect 15048 36036 15104 36038
rect 15152 36036 15208 36038
rect 14924 35810 14980 35812
rect 14924 35758 14926 35810
rect 14926 35758 14978 35810
rect 14978 35758 14980 35810
rect 14924 35756 14980 35758
rect 14028 35698 14084 35700
rect 14028 35646 14030 35698
rect 14030 35646 14082 35698
rect 14082 35646 14084 35698
rect 14028 35644 14084 35646
rect 14588 35644 14644 35700
rect 13692 34972 13748 35028
rect 15148 35698 15204 35700
rect 15148 35646 15150 35698
rect 15150 35646 15202 35698
rect 15202 35646 15204 35698
rect 15148 35644 15204 35646
rect 14700 35196 14756 35252
rect 15036 35196 15092 35252
rect 14588 35084 14644 35140
rect 13020 34524 13076 34580
rect 12908 33852 12964 33908
rect 12908 32562 12964 32564
rect 12908 32510 12910 32562
rect 12910 32510 12962 32562
rect 12962 32510 12964 32562
rect 12908 32508 12964 32510
rect 12684 31890 12740 31892
rect 12684 31838 12686 31890
rect 12686 31838 12738 31890
rect 12738 31838 12740 31890
rect 12684 31836 12740 31838
rect 13580 34524 13636 34580
rect 13804 34524 13860 34580
rect 14008 34522 14064 34524
rect 14112 34522 14168 34524
rect 14008 34470 14024 34522
rect 14024 34470 14064 34522
rect 14112 34470 14148 34522
rect 14148 34470 14168 34522
rect 14008 34468 14064 34470
rect 14112 34468 14168 34470
rect 14216 34468 14272 34524
rect 14320 34522 14376 34524
rect 14424 34522 14480 34524
rect 14528 34522 14584 34524
rect 14320 34470 14324 34522
rect 14324 34470 14376 34522
rect 14424 34470 14448 34522
rect 14448 34470 14480 34522
rect 14528 34470 14572 34522
rect 14572 34470 14584 34522
rect 14320 34468 14376 34470
rect 14424 34468 14480 34470
rect 14528 34468 14584 34470
rect 14632 34522 14688 34524
rect 14736 34522 14792 34524
rect 14840 34522 14896 34524
rect 14632 34470 14644 34522
rect 14644 34470 14688 34522
rect 14736 34470 14768 34522
rect 14768 34470 14792 34522
rect 14840 34470 14892 34522
rect 14892 34470 14896 34522
rect 14632 34468 14688 34470
rect 14736 34468 14792 34470
rect 14840 34468 14896 34470
rect 14944 34468 15000 34524
rect 15048 34522 15104 34524
rect 15152 34522 15208 34524
rect 15048 34470 15068 34522
rect 15068 34470 15104 34522
rect 15152 34470 15192 34522
rect 15192 34470 15208 34522
rect 15048 34468 15104 34470
rect 15152 34468 15208 34470
rect 16044 37772 16100 37828
rect 16156 38892 16212 38948
rect 16044 36540 16100 36596
rect 15820 34354 15876 34356
rect 15820 34302 15822 34354
rect 15822 34302 15874 34354
rect 15874 34302 15876 34354
rect 15820 34300 15876 34302
rect 17500 45890 17556 45892
rect 17500 45838 17502 45890
rect 17502 45838 17554 45890
rect 17554 45838 17556 45890
rect 17500 45836 17556 45838
rect 17724 45276 17780 45332
rect 18284 45276 18340 45332
rect 16828 44994 16884 44996
rect 16828 44942 16830 44994
rect 16830 44942 16882 44994
rect 16882 44942 16884 44994
rect 16828 44940 16884 44942
rect 17388 45218 17444 45220
rect 17388 45166 17390 45218
rect 17390 45166 17442 45218
rect 17442 45166 17444 45218
rect 17388 45164 17444 45166
rect 17388 44828 17444 44884
rect 17388 43596 17444 43652
rect 16604 43372 16660 43428
rect 16716 43148 16772 43204
rect 17612 44492 17668 44548
rect 17724 44380 17780 44436
rect 17612 44210 17668 44212
rect 17612 44158 17614 44210
rect 17614 44158 17666 44210
rect 17666 44158 17668 44210
rect 17612 44156 17668 44158
rect 17500 43148 17556 43204
rect 16492 41356 16548 41412
rect 17500 41410 17556 41412
rect 17500 41358 17502 41410
rect 17502 41358 17554 41410
rect 17554 41358 17556 41410
rect 17500 41356 17556 41358
rect 16716 38946 16772 38948
rect 16716 38894 16718 38946
rect 16718 38894 16770 38946
rect 16770 38894 16772 38946
rect 16716 38892 16772 38894
rect 17836 42194 17892 42196
rect 17836 42142 17838 42194
rect 17838 42142 17890 42194
rect 17890 42142 17892 42194
rect 17836 42140 17892 42142
rect 17724 42082 17780 42084
rect 17724 42030 17726 42082
rect 17726 42030 17778 42082
rect 17778 42030 17780 42082
rect 17724 42028 17780 42030
rect 17612 40572 17668 40628
rect 18060 43596 18116 43652
rect 18060 42140 18116 42196
rect 18172 44156 18228 44212
rect 18620 47012 18676 47068
rect 18844 49084 18900 49140
rect 21644 52556 21700 52612
rect 21532 51996 21588 52052
rect 21420 51938 21476 51940
rect 21420 51886 21422 51938
rect 21422 51886 21474 51938
rect 21474 51886 21476 51938
rect 21420 51884 21476 51886
rect 20188 49196 20244 49252
rect 20076 49138 20132 49140
rect 20076 49086 20078 49138
rect 20078 49086 20130 49138
rect 20130 49086 20132 49138
rect 20076 49084 20132 49086
rect 19628 48802 19684 48804
rect 19628 48750 19630 48802
rect 19630 48750 19682 48802
rect 19682 48750 19684 48802
rect 19628 48748 19684 48750
rect 19852 47180 19908 47236
rect 18956 46898 19012 46900
rect 18956 46846 18958 46898
rect 18958 46846 19010 46898
rect 19010 46846 19012 46898
rect 18956 46844 19012 46846
rect 18732 45666 18788 45668
rect 18732 45614 18734 45666
rect 18734 45614 18786 45666
rect 18786 45614 18788 45666
rect 18732 45612 18788 45614
rect 18620 44882 18676 44884
rect 18620 44830 18622 44882
rect 18622 44830 18674 44882
rect 18674 44830 18676 44882
rect 18620 44828 18676 44830
rect 18508 44434 18564 44436
rect 18508 44382 18510 44434
rect 18510 44382 18562 44434
rect 18562 44382 18564 44434
rect 18508 44380 18564 44382
rect 18956 44492 19012 44548
rect 19292 45500 19348 45556
rect 19628 45612 19684 45668
rect 19068 44156 19124 44212
rect 19180 45276 19236 45332
rect 18620 43932 18676 43988
rect 18844 43820 18900 43876
rect 18396 43260 18452 43316
rect 18396 42028 18452 42084
rect 16492 38722 16548 38724
rect 16492 38670 16494 38722
rect 16494 38670 16546 38722
rect 16546 38670 16548 38722
rect 16492 38668 16548 38670
rect 16380 38556 16436 38612
rect 18956 43372 19012 43428
rect 19068 42194 19124 42196
rect 19068 42142 19070 42194
rect 19070 42142 19122 42194
rect 19122 42142 19124 42194
rect 19068 42140 19124 42142
rect 18732 41916 18788 41972
rect 19292 43538 19348 43540
rect 19292 43486 19294 43538
rect 19294 43486 19346 43538
rect 19346 43486 19348 43538
rect 19292 43484 19348 43486
rect 20972 48242 21028 48244
rect 20972 48190 20974 48242
rect 20974 48190 21026 48242
rect 21026 48190 21028 48242
rect 20972 48188 21028 48190
rect 21420 47516 21476 47572
rect 21644 47234 21700 47236
rect 21644 47182 21646 47234
rect 21646 47182 21698 47234
rect 21698 47182 21700 47234
rect 21644 47180 21700 47182
rect 21308 45890 21364 45892
rect 21308 45838 21310 45890
rect 21310 45838 21362 45890
rect 21362 45838 21364 45890
rect 21308 45836 21364 45838
rect 21532 45666 21588 45668
rect 21532 45614 21534 45666
rect 21534 45614 21586 45666
rect 21586 45614 21588 45666
rect 21532 45612 21588 45614
rect 19852 44828 19908 44884
rect 19964 44156 20020 44212
rect 19516 43820 19572 43876
rect 19740 43650 19796 43652
rect 19740 43598 19742 43650
rect 19742 43598 19794 43650
rect 19794 43598 19796 43650
rect 19740 43596 19796 43598
rect 19852 43426 19908 43428
rect 19852 43374 19854 43426
rect 19854 43374 19906 43426
rect 19906 43374 19908 43426
rect 19852 43372 19908 43374
rect 19292 42700 19348 42756
rect 22204 53228 22260 53284
rect 21868 52162 21924 52164
rect 21868 52110 21870 52162
rect 21870 52110 21922 52162
rect 21922 52110 21924 52162
rect 21868 52108 21924 52110
rect 21980 51884 22036 51940
rect 22316 52892 22372 52948
rect 22540 55132 22596 55188
rect 22988 56194 23044 56196
rect 22988 56142 22990 56194
rect 22990 56142 23042 56194
rect 23042 56142 23044 56194
rect 22988 56140 23044 56142
rect 22876 54684 22932 54740
rect 22876 53676 22932 53732
rect 22652 53228 22708 53284
rect 22540 52444 22596 52500
rect 22876 51602 22932 51604
rect 22876 51550 22878 51602
rect 22878 51550 22930 51602
rect 22930 51550 22932 51602
rect 22876 51548 22932 51550
rect 22428 50652 22484 50708
rect 23100 50706 23156 50708
rect 23100 50654 23102 50706
rect 23102 50654 23154 50706
rect 23154 50654 23156 50706
rect 23100 50652 23156 50654
rect 24556 66050 24612 66052
rect 24556 65998 24558 66050
rect 24558 65998 24610 66050
rect 24610 65998 24612 66050
rect 24556 65996 24612 65998
rect 26236 70140 26292 70196
rect 26460 70082 26516 70084
rect 26460 70030 26462 70082
rect 26462 70030 26514 70082
rect 26514 70030 26516 70082
rect 26460 70028 26516 70030
rect 27132 70194 27188 70196
rect 27132 70142 27134 70194
rect 27134 70142 27186 70194
rect 27186 70142 27188 70194
rect 27132 70140 27188 70142
rect 27020 69244 27076 69300
rect 26684 68572 26740 68628
rect 26348 68460 26404 68516
rect 26460 68348 26516 68404
rect 26460 67842 26516 67844
rect 26460 67790 26462 67842
rect 26462 67790 26514 67842
rect 26514 67790 26516 67842
rect 26460 67788 26516 67790
rect 25452 66220 25508 66276
rect 26236 66946 26292 66948
rect 26236 66894 26238 66946
rect 26238 66894 26290 66946
rect 26290 66894 26292 66946
rect 26236 66892 26292 66894
rect 26684 66946 26740 66948
rect 26684 66894 26686 66946
rect 26686 66894 26738 66946
rect 26738 66894 26740 66946
rect 26684 66892 26740 66894
rect 25004 65324 25060 65380
rect 24008 65098 24064 65100
rect 24112 65098 24168 65100
rect 24008 65046 24024 65098
rect 24024 65046 24064 65098
rect 24112 65046 24148 65098
rect 24148 65046 24168 65098
rect 24008 65044 24064 65046
rect 24112 65044 24168 65046
rect 24216 65044 24272 65100
rect 24320 65098 24376 65100
rect 24424 65098 24480 65100
rect 24528 65098 24584 65100
rect 24320 65046 24324 65098
rect 24324 65046 24376 65098
rect 24424 65046 24448 65098
rect 24448 65046 24480 65098
rect 24528 65046 24572 65098
rect 24572 65046 24584 65098
rect 24320 65044 24376 65046
rect 24424 65044 24480 65046
rect 24528 65044 24584 65046
rect 24632 65098 24688 65100
rect 24736 65098 24792 65100
rect 24840 65098 24896 65100
rect 24632 65046 24644 65098
rect 24644 65046 24688 65098
rect 24736 65046 24768 65098
rect 24768 65046 24792 65098
rect 24840 65046 24892 65098
rect 24892 65046 24896 65098
rect 24632 65044 24688 65046
rect 24736 65044 24792 65046
rect 24840 65044 24896 65046
rect 24944 65044 25000 65100
rect 25048 65098 25104 65100
rect 25152 65098 25208 65100
rect 25048 65046 25068 65098
rect 25068 65046 25104 65098
rect 25152 65046 25192 65098
rect 25192 65046 25208 65098
rect 25048 65044 25104 65046
rect 25152 65044 25208 65046
rect 24008 63530 24064 63532
rect 24112 63530 24168 63532
rect 24008 63478 24024 63530
rect 24024 63478 24064 63530
rect 24112 63478 24148 63530
rect 24148 63478 24168 63530
rect 24008 63476 24064 63478
rect 24112 63476 24168 63478
rect 24216 63476 24272 63532
rect 24320 63530 24376 63532
rect 24424 63530 24480 63532
rect 24528 63530 24584 63532
rect 24320 63478 24324 63530
rect 24324 63478 24376 63530
rect 24424 63478 24448 63530
rect 24448 63478 24480 63530
rect 24528 63478 24572 63530
rect 24572 63478 24584 63530
rect 24320 63476 24376 63478
rect 24424 63476 24480 63478
rect 24528 63476 24584 63478
rect 24632 63530 24688 63532
rect 24736 63530 24792 63532
rect 24840 63530 24896 63532
rect 24632 63478 24644 63530
rect 24644 63478 24688 63530
rect 24736 63478 24768 63530
rect 24768 63478 24792 63530
rect 24840 63478 24892 63530
rect 24892 63478 24896 63530
rect 24632 63476 24688 63478
rect 24736 63476 24792 63478
rect 24840 63476 24896 63478
rect 24944 63476 25000 63532
rect 25048 63530 25104 63532
rect 25152 63530 25208 63532
rect 25048 63478 25068 63530
rect 25068 63478 25104 63530
rect 25152 63478 25192 63530
rect 25192 63478 25208 63530
rect 25048 63476 25104 63478
rect 25152 63476 25208 63478
rect 24780 63250 24836 63252
rect 24780 63198 24782 63250
rect 24782 63198 24834 63250
rect 24834 63198 24836 63250
rect 24780 63196 24836 63198
rect 24892 63138 24948 63140
rect 24892 63086 24894 63138
rect 24894 63086 24946 63138
rect 24946 63086 24948 63138
rect 24892 63084 24948 63086
rect 24108 63026 24164 63028
rect 24108 62974 24110 63026
rect 24110 62974 24162 63026
rect 24162 62974 24164 63026
rect 24108 62972 24164 62974
rect 24668 63026 24724 63028
rect 24668 62974 24670 63026
rect 24670 62974 24722 63026
rect 24722 62974 24724 63026
rect 24668 62972 24724 62974
rect 25228 62860 25284 62916
rect 24108 62578 24164 62580
rect 24108 62526 24110 62578
rect 24110 62526 24162 62578
rect 24162 62526 24164 62578
rect 24108 62524 24164 62526
rect 24668 62466 24724 62468
rect 24668 62414 24670 62466
rect 24670 62414 24722 62466
rect 24722 62414 24724 62466
rect 24668 62412 24724 62414
rect 25676 63196 25732 63252
rect 25676 62412 25732 62468
rect 25340 62354 25396 62356
rect 25340 62302 25342 62354
rect 25342 62302 25394 62354
rect 25394 62302 25396 62354
rect 25340 62300 25396 62302
rect 23772 59724 23828 59780
rect 24008 61962 24064 61964
rect 24112 61962 24168 61964
rect 24008 61910 24024 61962
rect 24024 61910 24064 61962
rect 24112 61910 24148 61962
rect 24148 61910 24168 61962
rect 24008 61908 24064 61910
rect 24112 61908 24168 61910
rect 24216 61908 24272 61964
rect 24320 61962 24376 61964
rect 24424 61962 24480 61964
rect 24528 61962 24584 61964
rect 24320 61910 24324 61962
rect 24324 61910 24376 61962
rect 24424 61910 24448 61962
rect 24448 61910 24480 61962
rect 24528 61910 24572 61962
rect 24572 61910 24584 61962
rect 24320 61908 24376 61910
rect 24424 61908 24480 61910
rect 24528 61908 24584 61910
rect 24632 61962 24688 61964
rect 24736 61962 24792 61964
rect 24840 61962 24896 61964
rect 24632 61910 24644 61962
rect 24644 61910 24688 61962
rect 24736 61910 24768 61962
rect 24768 61910 24792 61962
rect 24840 61910 24892 61962
rect 24892 61910 24896 61962
rect 24632 61908 24688 61910
rect 24736 61908 24792 61910
rect 24840 61908 24896 61910
rect 24944 61908 25000 61964
rect 25048 61962 25104 61964
rect 25152 61962 25208 61964
rect 25048 61910 25068 61962
rect 25068 61910 25104 61962
rect 25152 61910 25192 61962
rect 25192 61910 25208 61962
rect 25048 61908 25104 61910
rect 25152 61908 25208 61910
rect 25788 61852 25844 61908
rect 24220 61740 24276 61796
rect 25228 61740 25284 61796
rect 24556 61458 24612 61460
rect 24556 61406 24558 61458
rect 24558 61406 24610 61458
rect 24610 61406 24612 61458
rect 24556 61404 24612 61406
rect 25788 61458 25844 61460
rect 25788 61406 25790 61458
rect 25790 61406 25842 61458
rect 25842 61406 25844 61458
rect 25788 61404 25844 61406
rect 26012 65490 26068 65492
rect 26012 65438 26014 65490
rect 26014 65438 26066 65490
rect 26066 65438 26068 65490
rect 26012 65436 26068 65438
rect 26012 62076 26068 62132
rect 26124 61852 26180 61908
rect 25340 60674 25396 60676
rect 25340 60622 25342 60674
rect 25342 60622 25394 60674
rect 25394 60622 25396 60674
rect 25340 60620 25396 60622
rect 26012 60620 26068 60676
rect 24008 60394 24064 60396
rect 24112 60394 24168 60396
rect 24008 60342 24024 60394
rect 24024 60342 24064 60394
rect 24112 60342 24148 60394
rect 24148 60342 24168 60394
rect 24008 60340 24064 60342
rect 24112 60340 24168 60342
rect 24216 60340 24272 60396
rect 24320 60394 24376 60396
rect 24424 60394 24480 60396
rect 24528 60394 24584 60396
rect 24320 60342 24324 60394
rect 24324 60342 24376 60394
rect 24424 60342 24448 60394
rect 24448 60342 24480 60394
rect 24528 60342 24572 60394
rect 24572 60342 24584 60394
rect 24320 60340 24376 60342
rect 24424 60340 24480 60342
rect 24528 60340 24584 60342
rect 24632 60394 24688 60396
rect 24736 60394 24792 60396
rect 24840 60394 24896 60396
rect 24632 60342 24644 60394
rect 24644 60342 24688 60394
rect 24736 60342 24768 60394
rect 24768 60342 24792 60394
rect 24840 60342 24892 60394
rect 24892 60342 24896 60394
rect 24632 60340 24688 60342
rect 24736 60340 24792 60342
rect 24840 60340 24896 60342
rect 24944 60340 25000 60396
rect 25048 60394 25104 60396
rect 25152 60394 25208 60396
rect 25048 60342 25068 60394
rect 25068 60342 25104 60394
rect 25152 60342 25192 60394
rect 25192 60342 25208 60394
rect 25048 60340 25104 60342
rect 25152 60340 25208 60342
rect 23884 59388 23940 59444
rect 23660 58210 23716 58212
rect 23660 58158 23662 58210
rect 23662 58158 23714 58210
rect 23714 58158 23716 58210
rect 23660 58156 23716 58158
rect 25340 59442 25396 59444
rect 25340 59390 25342 59442
rect 25342 59390 25394 59442
rect 25394 59390 25396 59442
rect 25340 59388 25396 59390
rect 24008 58826 24064 58828
rect 24112 58826 24168 58828
rect 24008 58774 24024 58826
rect 24024 58774 24064 58826
rect 24112 58774 24148 58826
rect 24148 58774 24168 58826
rect 24008 58772 24064 58774
rect 24112 58772 24168 58774
rect 24216 58772 24272 58828
rect 24320 58826 24376 58828
rect 24424 58826 24480 58828
rect 24528 58826 24584 58828
rect 24320 58774 24324 58826
rect 24324 58774 24376 58826
rect 24424 58774 24448 58826
rect 24448 58774 24480 58826
rect 24528 58774 24572 58826
rect 24572 58774 24584 58826
rect 24320 58772 24376 58774
rect 24424 58772 24480 58774
rect 24528 58772 24584 58774
rect 24632 58826 24688 58828
rect 24736 58826 24792 58828
rect 24840 58826 24896 58828
rect 24632 58774 24644 58826
rect 24644 58774 24688 58826
rect 24736 58774 24768 58826
rect 24768 58774 24792 58826
rect 24840 58774 24892 58826
rect 24892 58774 24896 58826
rect 24632 58772 24688 58774
rect 24736 58772 24792 58774
rect 24840 58772 24896 58774
rect 24944 58772 25000 58828
rect 25048 58826 25104 58828
rect 25152 58826 25208 58828
rect 25048 58774 25068 58826
rect 25068 58774 25104 58826
rect 25152 58774 25192 58826
rect 25192 58774 25208 58826
rect 25048 58772 25104 58774
rect 25152 58772 25208 58774
rect 23660 57596 23716 57652
rect 26012 58380 26068 58436
rect 25676 58268 25732 58324
rect 25452 57932 25508 57988
rect 26236 57932 26292 57988
rect 24780 57762 24836 57764
rect 24780 57710 24782 57762
rect 24782 57710 24834 57762
rect 24834 57710 24836 57762
rect 24780 57708 24836 57710
rect 24008 57258 24064 57260
rect 24112 57258 24168 57260
rect 24008 57206 24024 57258
rect 24024 57206 24064 57258
rect 24112 57206 24148 57258
rect 24148 57206 24168 57258
rect 24008 57204 24064 57206
rect 24112 57204 24168 57206
rect 24216 57204 24272 57260
rect 24320 57258 24376 57260
rect 24424 57258 24480 57260
rect 24528 57258 24584 57260
rect 24320 57206 24324 57258
rect 24324 57206 24376 57258
rect 24424 57206 24448 57258
rect 24448 57206 24480 57258
rect 24528 57206 24572 57258
rect 24572 57206 24584 57258
rect 24320 57204 24376 57206
rect 24424 57204 24480 57206
rect 24528 57204 24584 57206
rect 24632 57258 24688 57260
rect 24736 57258 24792 57260
rect 24840 57258 24896 57260
rect 24632 57206 24644 57258
rect 24644 57206 24688 57258
rect 24736 57206 24768 57258
rect 24768 57206 24792 57258
rect 24840 57206 24892 57258
rect 24892 57206 24896 57258
rect 24632 57204 24688 57206
rect 24736 57204 24792 57206
rect 24840 57204 24896 57206
rect 24944 57204 25000 57260
rect 25048 57258 25104 57260
rect 25152 57258 25208 57260
rect 25048 57206 25068 57258
rect 25068 57206 25104 57258
rect 25152 57206 25192 57258
rect 25192 57206 25208 57258
rect 25048 57204 25104 57206
rect 25152 57204 25208 57206
rect 25340 57260 25396 57316
rect 23996 56588 24052 56644
rect 25116 56866 25172 56868
rect 25116 56814 25118 56866
rect 25118 56814 25170 56866
rect 25170 56814 25172 56866
rect 25116 56812 25172 56814
rect 25676 57650 25732 57652
rect 25676 57598 25678 57650
rect 25678 57598 25730 57650
rect 25730 57598 25732 57650
rect 25676 57596 25732 57598
rect 26796 64876 26852 64932
rect 27020 63868 27076 63924
rect 26572 63026 26628 63028
rect 26572 62974 26574 63026
rect 26574 62974 26626 63026
rect 26626 62974 26628 63026
rect 26572 62972 26628 62974
rect 27132 63026 27188 63028
rect 27132 62974 27134 63026
rect 27134 62974 27186 63026
rect 27186 62974 27188 63026
rect 27132 62972 27188 62974
rect 26796 62914 26852 62916
rect 26796 62862 26798 62914
rect 26798 62862 26850 62914
rect 26850 62862 26852 62914
rect 26796 62860 26852 62862
rect 26908 61404 26964 61460
rect 26684 60956 26740 61012
rect 26684 59724 26740 59780
rect 25900 57260 25956 57316
rect 26572 58380 26628 58436
rect 24668 56140 24724 56196
rect 24008 55690 24064 55692
rect 24112 55690 24168 55692
rect 24008 55638 24024 55690
rect 24024 55638 24064 55690
rect 24112 55638 24148 55690
rect 24148 55638 24168 55690
rect 24008 55636 24064 55638
rect 24112 55636 24168 55638
rect 24216 55636 24272 55692
rect 24320 55690 24376 55692
rect 24424 55690 24480 55692
rect 24528 55690 24584 55692
rect 24320 55638 24324 55690
rect 24324 55638 24376 55690
rect 24424 55638 24448 55690
rect 24448 55638 24480 55690
rect 24528 55638 24572 55690
rect 24572 55638 24584 55690
rect 24320 55636 24376 55638
rect 24424 55636 24480 55638
rect 24528 55636 24584 55638
rect 24632 55690 24688 55692
rect 24736 55690 24792 55692
rect 24840 55690 24896 55692
rect 24632 55638 24644 55690
rect 24644 55638 24688 55690
rect 24736 55638 24768 55690
rect 24768 55638 24792 55690
rect 24840 55638 24892 55690
rect 24892 55638 24896 55690
rect 24632 55636 24688 55638
rect 24736 55636 24792 55638
rect 24840 55636 24896 55638
rect 24944 55636 25000 55692
rect 25048 55690 25104 55692
rect 25152 55690 25208 55692
rect 25048 55638 25068 55690
rect 25068 55638 25104 55690
rect 25152 55638 25192 55690
rect 25192 55638 25208 55690
rect 25048 55636 25104 55638
rect 25152 55636 25208 55638
rect 23548 54572 23604 54628
rect 23548 53788 23604 53844
rect 24008 54122 24064 54124
rect 24112 54122 24168 54124
rect 24008 54070 24024 54122
rect 24024 54070 24064 54122
rect 24112 54070 24148 54122
rect 24148 54070 24168 54122
rect 24008 54068 24064 54070
rect 24112 54068 24168 54070
rect 24216 54068 24272 54124
rect 24320 54122 24376 54124
rect 24424 54122 24480 54124
rect 24528 54122 24584 54124
rect 24320 54070 24324 54122
rect 24324 54070 24376 54122
rect 24424 54070 24448 54122
rect 24448 54070 24480 54122
rect 24528 54070 24572 54122
rect 24572 54070 24584 54122
rect 24320 54068 24376 54070
rect 24424 54068 24480 54070
rect 24528 54068 24584 54070
rect 24632 54122 24688 54124
rect 24736 54122 24792 54124
rect 24840 54122 24896 54124
rect 24632 54070 24644 54122
rect 24644 54070 24688 54122
rect 24736 54070 24768 54122
rect 24768 54070 24792 54122
rect 24840 54070 24892 54122
rect 24892 54070 24896 54122
rect 24632 54068 24688 54070
rect 24736 54068 24792 54070
rect 24840 54068 24896 54070
rect 24944 54068 25000 54124
rect 25048 54122 25104 54124
rect 25152 54122 25208 54124
rect 25048 54070 25068 54122
rect 25068 54070 25104 54122
rect 25152 54070 25192 54122
rect 25192 54070 25208 54122
rect 25048 54068 25104 54070
rect 25152 54068 25208 54070
rect 23660 53676 23716 53732
rect 24668 53788 24724 53844
rect 25116 53506 25172 53508
rect 25116 53454 25118 53506
rect 25118 53454 25170 53506
rect 25170 53454 25172 53506
rect 25116 53452 25172 53454
rect 23772 53228 23828 53284
rect 23660 53058 23716 53060
rect 23660 53006 23662 53058
rect 23662 53006 23714 53058
rect 23714 53006 23716 53058
rect 23660 53004 23716 53006
rect 24220 53228 24276 53284
rect 25340 53170 25396 53172
rect 25340 53118 25342 53170
rect 25342 53118 25394 53170
rect 25394 53118 25396 53170
rect 25340 53116 25396 53118
rect 24008 52554 24064 52556
rect 24112 52554 24168 52556
rect 24008 52502 24024 52554
rect 24024 52502 24064 52554
rect 24112 52502 24148 52554
rect 24148 52502 24168 52554
rect 24008 52500 24064 52502
rect 24112 52500 24168 52502
rect 24216 52500 24272 52556
rect 24320 52554 24376 52556
rect 24424 52554 24480 52556
rect 24528 52554 24584 52556
rect 24320 52502 24324 52554
rect 24324 52502 24376 52554
rect 24424 52502 24448 52554
rect 24448 52502 24480 52554
rect 24528 52502 24572 52554
rect 24572 52502 24584 52554
rect 24320 52500 24376 52502
rect 24424 52500 24480 52502
rect 24528 52500 24584 52502
rect 24632 52554 24688 52556
rect 24736 52554 24792 52556
rect 24840 52554 24896 52556
rect 24632 52502 24644 52554
rect 24644 52502 24688 52554
rect 24736 52502 24768 52554
rect 24768 52502 24792 52554
rect 24840 52502 24892 52554
rect 24892 52502 24896 52554
rect 24632 52500 24688 52502
rect 24736 52500 24792 52502
rect 24840 52500 24896 52502
rect 24944 52500 25000 52556
rect 25048 52554 25104 52556
rect 25152 52554 25208 52556
rect 25048 52502 25068 52554
rect 25068 52502 25104 52554
rect 25152 52502 25192 52554
rect 25192 52502 25208 52554
rect 25048 52500 25104 52502
rect 25152 52500 25208 52502
rect 26124 56642 26180 56644
rect 26124 56590 26126 56642
rect 26126 56590 26178 56642
rect 26178 56590 26180 56642
rect 26124 56588 26180 56590
rect 26684 58268 26740 58324
rect 26796 57820 26852 57876
rect 27916 70194 27972 70196
rect 27916 70142 27918 70194
rect 27918 70142 27970 70194
rect 27970 70142 27972 70194
rect 27916 70140 27972 70142
rect 28700 70140 28756 70196
rect 27580 70028 27636 70084
rect 27580 69244 27636 69300
rect 27916 68796 27972 68852
rect 28364 69298 28420 69300
rect 28364 69246 28366 69298
rect 28366 69246 28418 69298
rect 28418 69246 28420 69298
rect 28364 69244 28420 69246
rect 27804 67788 27860 67844
rect 29260 69522 29316 69524
rect 29260 69470 29262 69522
rect 29262 69470 29314 69522
rect 29314 69470 29316 69522
rect 29260 69468 29316 69470
rect 29148 69244 29204 69300
rect 28812 68850 28868 68852
rect 28812 68798 28814 68850
rect 28814 68798 28866 68850
rect 28866 68798 28868 68850
rect 28812 68796 28868 68798
rect 34008 78426 34064 78428
rect 34112 78426 34168 78428
rect 34008 78374 34024 78426
rect 34024 78374 34064 78426
rect 34112 78374 34148 78426
rect 34148 78374 34168 78426
rect 34008 78372 34064 78374
rect 34112 78372 34168 78374
rect 34216 78372 34272 78428
rect 34320 78426 34376 78428
rect 34424 78426 34480 78428
rect 34528 78426 34584 78428
rect 34320 78374 34324 78426
rect 34324 78374 34376 78426
rect 34424 78374 34448 78426
rect 34448 78374 34480 78426
rect 34528 78374 34572 78426
rect 34572 78374 34584 78426
rect 34320 78372 34376 78374
rect 34424 78372 34480 78374
rect 34528 78372 34584 78374
rect 34632 78426 34688 78428
rect 34736 78426 34792 78428
rect 34840 78426 34896 78428
rect 34632 78374 34644 78426
rect 34644 78374 34688 78426
rect 34736 78374 34768 78426
rect 34768 78374 34792 78426
rect 34840 78374 34892 78426
rect 34892 78374 34896 78426
rect 34632 78372 34688 78374
rect 34736 78372 34792 78374
rect 34840 78372 34896 78374
rect 34944 78372 35000 78428
rect 35048 78426 35104 78428
rect 35152 78426 35208 78428
rect 35048 78374 35068 78426
rect 35068 78374 35104 78426
rect 35152 78374 35192 78426
rect 35192 78374 35208 78426
rect 35048 78372 35104 78374
rect 35152 78372 35208 78374
rect 34008 76858 34064 76860
rect 34112 76858 34168 76860
rect 34008 76806 34024 76858
rect 34024 76806 34064 76858
rect 34112 76806 34148 76858
rect 34148 76806 34168 76858
rect 34008 76804 34064 76806
rect 34112 76804 34168 76806
rect 34216 76804 34272 76860
rect 34320 76858 34376 76860
rect 34424 76858 34480 76860
rect 34528 76858 34584 76860
rect 34320 76806 34324 76858
rect 34324 76806 34376 76858
rect 34424 76806 34448 76858
rect 34448 76806 34480 76858
rect 34528 76806 34572 76858
rect 34572 76806 34584 76858
rect 34320 76804 34376 76806
rect 34424 76804 34480 76806
rect 34528 76804 34584 76806
rect 34632 76858 34688 76860
rect 34736 76858 34792 76860
rect 34840 76858 34896 76860
rect 34632 76806 34644 76858
rect 34644 76806 34688 76858
rect 34736 76806 34768 76858
rect 34768 76806 34792 76858
rect 34840 76806 34892 76858
rect 34892 76806 34896 76858
rect 34632 76804 34688 76806
rect 34736 76804 34792 76806
rect 34840 76804 34896 76806
rect 34944 76804 35000 76860
rect 35048 76858 35104 76860
rect 35152 76858 35208 76860
rect 35048 76806 35068 76858
rect 35068 76806 35104 76858
rect 35152 76806 35192 76858
rect 35192 76806 35208 76858
rect 35048 76804 35104 76806
rect 35152 76804 35208 76806
rect 34008 75290 34064 75292
rect 34112 75290 34168 75292
rect 34008 75238 34024 75290
rect 34024 75238 34064 75290
rect 34112 75238 34148 75290
rect 34148 75238 34168 75290
rect 34008 75236 34064 75238
rect 34112 75236 34168 75238
rect 34216 75236 34272 75292
rect 34320 75290 34376 75292
rect 34424 75290 34480 75292
rect 34528 75290 34584 75292
rect 34320 75238 34324 75290
rect 34324 75238 34376 75290
rect 34424 75238 34448 75290
rect 34448 75238 34480 75290
rect 34528 75238 34572 75290
rect 34572 75238 34584 75290
rect 34320 75236 34376 75238
rect 34424 75236 34480 75238
rect 34528 75236 34584 75238
rect 34632 75290 34688 75292
rect 34736 75290 34792 75292
rect 34840 75290 34896 75292
rect 34632 75238 34644 75290
rect 34644 75238 34688 75290
rect 34736 75238 34768 75290
rect 34768 75238 34792 75290
rect 34840 75238 34892 75290
rect 34892 75238 34896 75290
rect 34632 75236 34688 75238
rect 34736 75236 34792 75238
rect 34840 75236 34896 75238
rect 34944 75236 35000 75292
rect 35048 75290 35104 75292
rect 35152 75290 35208 75292
rect 35048 75238 35068 75290
rect 35068 75238 35104 75290
rect 35152 75238 35192 75290
rect 35192 75238 35208 75290
rect 35048 75236 35104 75238
rect 35152 75236 35208 75238
rect 34008 73722 34064 73724
rect 34112 73722 34168 73724
rect 34008 73670 34024 73722
rect 34024 73670 34064 73722
rect 34112 73670 34148 73722
rect 34148 73670 34168 73722
rect 34008 73668 34064 73670
rect 34112 73668 34168 73670
rect 34216 73668 34272 73724
rect 34320 73722 34376 73724
rect 34424 73722 34480 73724
rect 34528 73722 34584 73724
rect 34320 73670 34324 73722
rect 34324 73670 34376 73722
rect 34424 73670 34448 73722
rect 34448 73670 34480 73722
rect 34528 73670 34572 73722
rect 34572 73670 34584 73722
rect 34320 73668 34376 73670
rect 34424 73668 34480 73670
rect 34528 73668 34584 73670
rect 34632 73722 34688 73724
rect 34736 73722 34792 73724
rect 34840 73722 34896 73724
rect 34632 73670 34644 73722
rect 34644 73670 34688 73722
rect 34736 73670 34768 73722
rect 34768 73670 34792 73722
rect 34840 73670 34892 73722
rect 34892 73670 34896 73722
rect 34632 73668 34688 73670
rect 34736 73668 34792 73670
rect 34840 73668 34896 73670
rect 34944 73668 35000 73724
rect 35048 73722 35104 73724
rect 35152 73722 35208 73724
rect 35048 73670 35068 73722
rect 35068 73670 35104 73722
rect 35152 73670 35192 73722
rect 35192 73670 35208 73722
rect 35048 73668 35104 73670
rect 35152 73668 35208 73670
rect 34008 72154 34064 72156
rect 34112 72154 34168 72156
rect 34008 72102 34024 72154
rect 34024 72102 34064 72154
rect 34112 72102 34148 72154
rect 34148 72102 34168 72154
rect 34008 72100 34064 72102
rect 34112 72100 34168 72102
rect 34216 72100 34272 72156
rect 34320 72154 34376 72156
rect 34424 72154 34480 72156
rect 34528 72154 34584 72156
rect 34320 72102 34324 72154
rect 34324 72102 34376 72154
rect 34424 72102 34448 72154
rect 34448 72102 34480 72154
rect 34528 72102 34572 72154
rect 34572 72102 34584 72154
rect 34320 72100 34376 72102
rect 34424 72100 34480 72102
rect 34528 72100 34584 72102
rect 34632 72154 34688 72156
rect 34736 72154 34792 72156
rect 34840 72154 34896 72156
rect 34632 72102 34644 72154
rect 34644 72102 34688 72154
rect 34736 72102 34768 72154
rect 34768 72102 34792 72154
rect 34840 72102 34892 72154
rect 34892 72102 34896 72154
rect 34632 72100 34688 72102
rect 34736 72100 34792 72102
rect 34840 72100 34896 72102
rect 34944 72100 35000 72156
rect 35048 72154 35104 72156
rect 35152 72154 35208 72156
rect 35048 72102 35068 72154
rect 35068 72102 35104 72154
rect 35152 72102 35192 72154
rect 35192 72102 35208 72154
rect 35048 72100 35104 72102
rect 35152 72100 35208 72102
rect 34972 71538 35028 71540
rect 34972 71486 34974 71538
rect 34974 71486 35026 71538
rect 35026 71486 35028 71538
rect 34972 71484 35028 71486
rect 30156 70924 30212 70980
rect 29820 70082 29876 70084
rect 29820 70030 29822 70082
rect 29822 70030 29874 70082
rect 29874 70030 29876 70082
rect 29820 70028 29876 70030
rect 29596 68572 29652 68628
rect 31836 70754 31892 70756
rect 31836 70702 31838 70754
rect 31838 70702 31890 70754
rect 31890 70702 31892 70754
rect 31836 70700 31892 70702
rect 31836 70140 31892 70196
rect 29036 68348 29092 68404
rect 32396 70476 32452 70532
rect 33068 70978 33124 70980
rect 33068 70926 33070 70978
rect 33070 70926 33122 70978
rect 33122 70926 33124 70978
rect 33068 70924 33124 70926
rect 33404 70476 33460 70532
rect 33180 70418 33236 70420
rect 33180 70366 33182 70418
rect 33182 70366 33234 70418
rect 33234 70366 33236 70418
rect 33180 70364 33236 70366
rect 32508 70082 32564 70084
rect 32508 70030 32510 70082
rect 32510 70030 32562 70082
rect 32562 70030 32564 70082
rect 32508 70028 32564 70030
rect 33292 70252 33348 70308
rect 30604 68796 30660 68852
rect 30156 68348 30212 68404
rect 29036 67228 29092 67284
rect 28588 66050 28644 66052
rect 28588 65998 28590 66050
rect 28590 65998 28642 66050
rect 28642 65998 28644 66050
rect 28588 65996 28644 65998
rect 28364 65714 28420 65716
rect 28364 65662 28366 65714
rect 28366 65662 28418 65714
rect 28418 65662 28420 65714
rect 28364 65660 28420 65662
rect 28812 63922 28868 63924
rect 28812 63870 28814 63922
rect 28814 63870 28866 63922
rect 28866 63870 28868 63922
rect 28812 63868 28868 63870
rect 28588 62748 28644 62804
rect 28252 62578 28308 62580
rect 28252 62526 28254 62578
rect 28254 62526 28306 62578
rect 28306 62526 28308 62578
rect 28252 62524 28308 62526
rect 28812 62242 28868 62244
rect 28812 62190 28814 62242
rect 28814 62190 28866 62242
rect 28866 62190 28868 62242
rect 28812 62188 28868 62190
rect 28476 61458 28532 61460
rect 28476 61406 28478 61458
rect 28478 61406 28530 61458
rect 28530 61406 28532 61458
rect 28476 61404 28532 61406
rect 28588 61346 28644 61348
rect 28588 61294 28590 61346
rect 28590 61294 28642 61346
rect 28642 61294 28644 61346
rect 28588 61292 28644 61294
rect 27020 60786 27076 60788
rect 27020 60734 27022 60786
rect 27022 60734 27074 60786
rect 27074 60734 27076 60786
rect 27020 60732 27076 60734
rect 28588 60956 28644 61012
rect 28364 59778 28420 59780
rect 28364 59726 28366 59778
rect 28366 59726 28418 59778
rect 28418 59726 28420 59778
rect 28364 59724 28420 59726
rect 27244 59052 27300 59108
rect 27804 58828 27860 58884
rect 27356 58434 27412 58436
rect 27356 58382 27358 58434
rect 27358 58382 27410 58434
rect 27410 58382 27412 58434
rect 27356 58380 27412 58382
rect 26348 56252 26404 56308
rect 26460 56140 26516 56196
rect 25676 53618 25732 53620
rect 25676 53566 25678 53618
rect 25678 53566 25730 53618
rect 25730 53566 25732 53618
rect 25676 53564 25732 53566
rect 23884 52220 23940 52276
rect 23772 52108 23828 52164
rect 23324 51996 23380 52052
rect 22316 48636 22372 48692
rect 22092 47570 22148 47572
rect 22092 47518 22094 47570
rect 22094 47518 22146 47570
rect 22146 47518 22148 47570
rect 22092 47516 22148 47518
rect 21980 47234 22036 47236
rect 21980 47182 21982 47234
rect 21982 47182 22034 47234
rect 22034 47182 22036 47234
rect 21980 47180 22036 47182
rect 22204 45890 22260 45892
rect 22204 45838 22206 45890
rect 22206 45838 22258 45890
rect 22258 45838 22260 45890
rect 22204 45836 22260 45838
rect 21868 45612 21924 45668
rect 22316 45276 22372 45332
rect 20412 44210 20468 44212
rect 20412 44158 20414 44210
rect 20414 44158 20466 44210
rect 20466 44158 20468 44210
rect 20412 44156 20468 44158
rect 21756 45052 21812 45108
rect 22316 44940 22372 44996
rect 21980 44322 22036 44324
rect 21980 44270 21982 44322
rect 21982 44270 22034 44322
rect 22034 44270 22036 44322
rect 21980 44268 22036 44270
rect 20972 43762 21028 43764
rect 20972 43710 20974 43762
rect 20974 43710 21026 43762
rect 21026 43710 21028 43762
rect 20972 43708 21028 43710
rect 20188 43484 20244 43540
rect 20748 42754 20804 42756
rect 20748 42702 20750 42754
rect 20750 42702 20802 42754
rect 20802 42702 20804 42754
rect 20748 42700 20804 42702
rect 20188 42530 20244 42532
rect 20188 42478 20190 42530
rect 20190 42478 20242 42530
rect 20242 42478 20244 42530
rect 20188 42476 20244 42478
rect 20972 42476 21028 42532
rect 19964 42140 20020 42196
rect 20748 42140 20804 42196
rect 16828 38780 16884 38836
rect 17388 38834 17444 38836
rect 17388 38782 17390 38834
rect 17390 38782 17442 38834
rect 17442 38782 17444 38834
rect 17388 38780 17444 38782
rect 17948 38668 18004 38724
rect 17612 38444 17668 38500
rect 16828 37324 16884 37380
rect 16492 37266 16548 37268
rect 16492 37214 16494 37266
rect 16494 37214 16546 37266
rect 16546 37214 16548 37266
rect 16492 37212 16548 37214
rect 16828 37154 16884 37156
rect 16828 37102 16830 37154
rect 16830 37102 16882 37154
rect 16882 37102 16884 37154
rect 16828 37100 16884 37102
rect 17500 37100 17556 37156
rect 16380 35810 16436 35812
rect 16380 35758 16382 35810
rect 16382 35758 16434 35810
rect 16434 35758 16436 35810
rect 16380 35756 16436 35758
rect 17052 35308 17108 35364
rect 16940 34748 16996 34804
rect 16716 34690 16772 34692
rect 16716 34638 16718 34690
rect 16718 34638 16770 34690
rect 16770 34638 16772 34690
rect 16716 34636 16772 34638
rect 16716 34354 16772 34356
rect 16716 34302 16718 34354
rect 16718 34302 16770 34354
rect 16770 34302 16772 34354
rect 16716 34300 16772 34302
rect 16492 34076 16548 34132
rect 13468 33852 13524 33908
rect 16380 33852 16436 33908
rect 15372 33404 15428 33460
rect 13916 33346 13972 33348
rect 13916 33294 13918 33346
rect 13918 33294 13970 33346
rect 13970 33294 13972 33346
rect 13916 33292 13972 33294
rect 13580 32508 13636 32564
rect 14476 33068 14532 33124
rect 14008 32954 14064 32956
rect 14112 32954 14168 32956
rect 14008 32902 14024 32954
rect 14024 32902 14064 32954
rect 14112 32902 14148 32954
rect 14148 32902 14168 32954
rect 14008 32900 14064 32902
rect 14112 32900 14168 32902
rect 14216 32900 14272 32956
rect 14320 32954 14376 32956
rect 14424 32954 14480 32956
rect 14528 32954 14584 32956
rect 14320 32902 14324 32954
rect 14324 32902 14376 32954
rect 14424 32902 14448 32954
rect 14448 32902 14480 32954
rect 14528 32902 14572 32954
rect 14572 32902 14584 32954
rect 14320 32900 14376 32902
rect 14424 32900 14480 32902
rect 14528 32900 14584 32902
rect 14632 32954 14688 32956
rect 14736 32954 14792 32956
rect 14840 32954 14896 32956
rect 14632 32902 14644 32954
rect 14644 32902 14688 32954
rect 14736 32902 14768 32954
rect 14768 32902 14792 32954
rect 14840 32902 14892 32954
rect 14892 32902 14896 32954
rect 14632 32900 14688 32902
rect 14736 32900 14792 32902
rect 14840 32900 14896 32902
rect 14944 32900 15000 32956
rect 15048 32954 15104 32956
rect 15152 32954 15208 32956
rect 15048 32902 15068 32954
rect 15068 32902 15104 32954
rect 15152 32902 15192 32954
rect 15192 32902 15208 32954
rect 15048 32900 15104 32902
rect 15152 32900 15208 32902
rect 14476 32732 14532 32788
rect 16268 33346 16324 33348
rect 16268 33294 16270 33346
rect 16270 33294 16322 33346
rect 16322 33294 16324 33346
rect 16268 33292 16324 33294
rect 15372 32786 15428 32788
rect 15372 32734 15374 32786
rect 15374 32734 15426 32786
rect 15426 32734 15428 32786
rect 15372 32732 15428 32734
rect 15932 32956 15988 33012
rect 16380 32956 16436 33012
rect 16268 32786 16324 32788
rect 16268 32734 16270 32786
rect 16270 32734 16322 32786
rect 16322 32734 16324 32786
rect 16268 32732 16324 32734
rect 15820 32396 15876 32452
rect 13020 31724 13076 31780
rect 13356 30882 13412 30884
rect 13356 30830 13358 30882
rect 13358 30830 13410 30882
rect 13410 30830 13412 30882
rect 13356 30828 13412 30830
rect 13020 30156 13076 30212
rect 13356 30156 13412 30212
rect 13692 31666 13748 31668
rect 13692 31614 13694 31666
rect 13694 31614 13746 31666
rect 13746 31614 13748 31666
rect 13692 31612 13748 31614
rect 14140 31612 14196 31668
rect 14924 31612 14980 31668
rect 15596 31666 15652 31668
rect 15596 31614 15598 31666
rect 15598 31614 15650 31666
rect 15650 31614 15652 31666
rect 15596 31612 15652 31614
rect 14008 31386 14064 31388
rect 14112 31386 14168 31388
rect 14008 31334 14024 31386
rect 14024 31334 14064 31386
rect 14112 31334 14148 31386
rect 14148 31334 14168 31386
rect 14008 31332 14064 31334
rect 14112 31332 14168 31334
rect 14216 31332 14272 31388
rect 14320 31386 14376 31388
rect 14424 31386 14480 31388
rect 14528 31386 14584 31388
rect 14320 31334 14324 31386
rect 14324 31334 14376 31386
rect 14424 31334 14448 31386
rect 14448 31334 14480 31386
rect 14528 31334 14572 31386
rect 14572 31334 14584 31386
rect 14320 31332 14376 31334
rect 14424 31332 14480 31334
rect 14528 31332 14584 31334
rect 14632 31386 14688 31388
rect 14736 31386 14792 31388
rect 14840 31386 14896 31388
rect 14632 31334 14644 31386
rect 14644 31334 14688 31386
rect 14736 31334 14768 31386
rect 14768 31334 14792 31386
rect 14840 31334 14892 31386
rect 14892 31334 14896 31386
rect 14632 31332 14688 31334
rect 14736 31332 14792 31334
rect 14840 31332 14896 31334
rect 14944 31332 15000 31388
rect 15048 31386 15104 31388
rect 15152 31386 15208 31388
rect 15048 31334 15068 31386
rect 15068 31334 15104 31386
rect 15152 31334 15192 31386
rect 15192 31334 15208 31386
rect 15048 31332 15104 31334
rect 15152 31332 15208 31334
rect 15820 31500 15876 31556
rect 13692 31052 13748 31108
rect 14364 30716 14420 30772
rect 14252 30210 14308 30212
rect 14252 30158 14254 30210
rect 14254 30158 14306 30210
rect 14306 30158 14308 30210
rect 14252 30156 14308 30158
rect 13468 30044 13524 30100
rect 14700 30268 14756 30324
rect 14364 29932 14420 29988
rect 14008 29818 14064 29820
rect 14112 29818 14168 29820
rect 14008 29766 14024 29818
rect 14024 29766 14064 29818
rect 14112 29766 14148 29818
rect 14148 29766 14168 29818
rect 14008 29764 14064 29766
rect 14112 29764 14168 29766
rect 14216 29764 14272 29820
rect 14320 29818 14376 29820
rect 14424 29818 14480 29820
rect 14528 29818 14584 29820
rect 14320 29766 14324 29818
rect 14324 29766 14376 29818
rect 14424 29766 14448 29818
rect 14448 29766 14480 29818
rect 14528 29766 14572 29818
rect 14572 29766 14584 29818
rect 14320 29764 14376 29766
rect 14424 29764 14480 29766
rect 14528 29764 14584 29766
rect 14632 29818 14688 29820
rect 14736 29818 14792 29820
rect 14840 29818 14896 29820
rect 14632 29766 14644 29818
rect 14644 29766 14688 29818
rect 14736 29766 14768 29818
rect 14768 29766 14792 29818
rect 14840 29766 14892 29818
rect 14892 29766 14896 29818
rect 14632 29764 14688 29766
rect 14736 29764 14792 29766
rect 14840 29764 14896 29766
rect 14944 29764 15000 29820
rect 15048 29818 15104 29820
rect 15152 29818 15208 29820
rect 15048 29766 15068 29818
rect 15068 29766 15104 29818
rect 15152 29766 15192 29818
rect 15192 29766 15208 29818
rect 15048 29764 15104 29766
rect 15152 29764 15208 29766
rect 15596 30770 15652 30772
rect 15596 30718 15598 30770
rect 15598 30718 15650 30770
rect 15650 30718 15652 30770
rect 15596 30716 15652 30718
rect 15596 30268 15652 30324
rect 15708 29932 15764 29988
rect 14476 29650 14532 29652
rect 14476 29598 14478 29650
rect 14478 29598 14530 29650
rect 14530 29598 14532 29650
rect 14476 29596 14532 29598
rect 15596 29596 15652 29652
rect 13804 29484 13860 29540
rect 13468 28924 13524 28980
rect 13580 29372 13636 29428
rect 13132 28364 13188 28420
rect 12684 27804 12740 27860
rect 12460 27468 12516 27524
rect 11564 27132 11620 27188
rect 13468 28252 13524 28308
rect 12236 26908 12292 26964
rect 9212 25282 9268 25284
rect 9212 25230 9214 25282
rect 9214 25230 9266 25282
rect 9266 25230 9268 25282
rect 9212 25228 9268 25230
rect 7756 22988 7812 23044
rect 7308 22428 7364 22484
rect 6748 21756 6804 21812
rect 6972 21698 7028 21700
rect 6972 21646 6974 21698
rect 6974 21646 7026 21698
rect 7026 21646 7028 21698
rect 6972 21644 7028 21646
rect 6860 21586 6916 21588
rect 6860 21534 6862 21586
rect 6862 21534 6914 21586
rect 6914 21534 6916 21586
rect 6860 21532 6916 21534
rect 7532 21586 7588 21588
rect 7532 21534 7534 21586
rect 7534 21534 7586 21586
rect 7586 21534 7588 21586
rect 7532 21532 7588 21534
rect 6748 20636 6804 20692
rect 6636 20524 6692 20580
rect 7420 18732 7476 18788
rect 7084 17500 7140 17556
rect 6972 16882 7028 16884
rect 6972 16830 6974 16882
rect 6974 16830 7026 16882
rect 7026 16830 7028 16882
rect 6972 16828 7028 16830
rect 6860 16770 6916 16772
rect 6860 16718 6862 16770
rect 6862 16718 6914 16770
rect 6914 16718 6916 16770
rect 6860 16716 6916 16718
rect 7420 16380 7476 16436
rect 7308 15484 7364 15540
rect 7196 15426 7252 15428
rect 7196 15374 7198 15426
rect 7198 15374 7250 15426
rect 7250 15374 7252 15426
rect 7196 15372 7252 15374
rect 6972 15090 7028 15092
rect 6972 15038 6974 15090
rect 6974 15038 7026 15090
rect 7026 15038 7028 15090
rect 6972 15036 7028 15038
rect 6524 14700 6580 14756
rect 6412 14364 6468 14420
rect 7196 14364 7252 14420
rect 6972 13692 7028 13748
rect 6524 13020 6580 13076
rect 5740 12348 5796 12404
rect 4060 12124 4116 12180
rect 5292 12124 5348 12180
rect 4008 11786 4064 11788
rect 4112 11786 4168 11788
rect 4008 11734 4024 11786
rect 4024 11734 4064 11786
rect 4112 11734 4148 11786
rect 4148 11734 4168 11786
rect 4008 11732 4064 11734
rect 4112 11732 4168 11734
rect 4216 11732 4272 11788
rect 4320 11786 4376 11788
rect 4424 11786 4480 11788
rect 4528 11786 4584 11788
rect 4320 11734 4324 11786
rect 4324 11734 4376 11786
rect 4424 11734 4448 11786
rect 4448 11734 4480 11786
rect 4528 11734 4572 11786
rect 4572 11734 4584 11786
rect 4320 11732 4376 11734
rect 4424 11732 4480 11734
rect 4528 11732 4584 11734
rect 4632 11786 4688 11788
rect 4736 11786 4792 11788
rect 4840 11786 4896 11788
rect 4632 11734 4644 11786
rect 4644 11734 4688 11786
rect 4736 11734 4768 11786
rect 4768 11734 4792 11786
rect 4840 11734 4892 11786
rect 4892 11734 4896 11786
rect 4632 11732 4688 11734
rect 4736 11732 4792 11734
rect 4840 11732 4896 11734
rect 4944 11732 5000 11788
rect 5048 11786 5104 11788
rect 5152 11786 5208 11788
rect 5048 11734 5068 11786
rect 5068 11734 5104 11786
rect 5152 11734 5192 11786
rect 5192 11734 5208 11786
rect 5048 11732 5104 11734
rect 5152 11732 5208 11734
rect 4396 11452 4452 11508
rect 5068 11506 5124 11508
rect 5068 11454 5070 11506
rect 5070 11454 5122 11506
rect 5122 11454 5124 11506
rect 5068 11452 5124 11454
rect 4508 11340 4564 11396
rect 4732 10834 4788 10836
rect 4732 10782 4734 10834
rect 4734 10782 4786 10834
rect 4786 10782 4788 10834
rect 4732 10780 4788 10782
rect 5516 12012 5572 12068
rect 5404 11340 5460 11396
rect 6076 12402 6132 12404
rect 6076 12350 6078 12402
rect 6078 12350 6130 12402
rect 6130 12350 6132 12402
rect 6076 12348 6132 12350
rect 7196 13692 7252 13748
rect 7084 13580 7140 13636
rect 6748 12348 6804 12404
rect 7196 13020 7252 13076
rect 6860 12290 6916 12292
rect 6860 12238 6862 12290
rect 6862 12238 6914 12290
rect 6914 12238 6916 12290
rect 6860 12236 6916 12238
rect 7084 12012 7140 12068
rect 8988 24722 9044 24724
rect 8988 24670 8990 24722
rect 8990 24670 9042 24722
rect 9042 24670 9044 24722
rect 8988 24668 9044 24670
rect 10220 25228 10276 25284
rect 8316 24444 8372 24500
rect 9660 24498 9716 24500
rect 9660 24446 9662 24498
rect 9662 24446 9714 24498
rect 9714 24446 9716 24498
rect 9660 24444 9716 24446
rect 9660 23100 9716 23156
rect 8428 21810 8484 21812
rect 8428 21758 8430 21810
rect 8430 21758 8482 21810
rect 8482 21758 8484 21810
rect 8428 21756 8484 21758
rect 8428 20802 8484 20804
rect 8428 20750 8430 20802
rect 8430 20750 8482 20802
rect 8482 20750 8484 20802
rect 8428 20748 8484 20750
rect 8876 21810 8932 21812
rect 8876 21758 8878 21810
rect 8878 21758 8930 21810
rect 8930 21758 8932 21810
rect 8876 21756 8932 21758
rect 8764 21698 8820 21700
rect 8764 21646 8766 21698
rect 8766 21646 8818 21698
rect 8818 21646 8820 21698
rect 8764 21644 8820 21646
rect 8540 17612 8596 17668
rect 8764 20578 8820 20580
rect 8764 20526 8766 20578
rect 8766 20526 8818 20578
rect 8818 20526 8820 20578
rect 8764 20524 8820 20526
rect 8652 17388 8708 17444
rect 8428 16994 8484 16996
rect 8428 16942 8430 16994
rect 8430 16942 8482 16994
rect 8482 16942 8484 16994
rect 8428 16940 8484 16942
rect 8092 16716 8148 16772
rect 7756 16658 7812 16660
rect 7756 16606 7758 16658
rect 7758 16606 7810 16658
rect 7810 16606 7812 16658
rect 7756 16604 7812 16606
rect 8316 16658 8372 16660
rect 8316 16606 8318 16658
rect 8318 16606 8370 16658
rect 8370 16606 8372 16658
rect 8316 16604 8372 16606
rect 7868 16380 7924 16436
rect 7532 15484 7588 15540
rect 8204 14418 8260 14420
rect 8204 14366 8206 14418
rect 8206 14366 8258 14418
rect 8258 14366 8260 14418
rect 8204 14364 8260 14366
rect 7756 13746 7812 13748
rect 7756 13694 7758 13746
rect 7758 13694 7810 13746
rect 7810 13694 7812 13746
rect 7756 13692 7812 13694
rect 8204 13634 8260 13636
rect 8204 13582 8206 13634
rect 8206 13582 8258 13634
rect 8258 13582 8260 13634
rect 8204 13580 8260 13582
rect 9100 20802 9156 20804
rect 9100 20750 9102 20802
rect 9102 20750 9154 20802
rect 9154 20750 9156 20802
rect 9100 20748 9156 20750
rect 9772 20748 9828 20804
rect 9324 20690 9380 20692
rect 9324 20638 9326 20690
rect 9326 20638 9378 20690
rect 9378 20638 9380 20690
rect 9324 20636 9380 20638
rect 8876 19964 8932 20020
rect 9548 20578 9604 20580
rect 9548 20526 9550 20578
rect 9550 20526 9602 20578
rect 9602 20526 9604 20578
rect 9548 20524 9604 20526
rect 9660 20076 9716 20132
rect 9212 17554 9268 17556
rect 9212 17502 9214 17554
rect 9214 17502 9266 17554
rect 9266 17502 9268 17554
rect 9212 17500 9268 17502
rect 8652 16156 8708 16212
rect 8428 14530 8484 14532
rect 8428 14478 8430 14530
rect 8430 14478 8482 14530
rect 8482 14478 8484 14530
rect 8428 14476 8484 14478
rect 8764 15090 8820 15092
rect 8764 15038 8766 15090
rect 8766 15038 8818 15090
rect 8818 15038 8820 15090
rect 8764 15036 8820 15038
rect 8876 14924 8932 14980
rect 8764 14418 8820 14420
rect 8764 14366 8766 14418
rect 8766 14366 8818 14418
rect 8818 14366 8820 14418
rect 8764 14364 8820 14366
rect 9100 14924 9156 14980
rect 9660 17500 9716 17556
rect 9548 16882 9604 16884
rect 9548 16830 9550 16882
rect 9550 16830 9602 16882
rect 9602 16830 9604 16882
rect 9548 16828 9604 16830
rect 9100 13916 9156 13972
rect 8540 13580 8596 13636
rect 7420 12236 7476 12292
rect 8204 12684 8260 12740
rect 7308 12066 7364 12068
rect 7308 12014 7310 12066
rect 7310 12014 7362 12066
rect 7362 12014 7364 12066
rect 7308 12012 7364 12014
rect 6972 11900 7028 11956
rect 5740 11170 5796 11172
rect 5740 11118 5742 11170
rect 5742 11118 5794 11170
rect 5794 11118 5796 11170
rect 5740 11116 5796 11118
rect 4008 10218 4064 10220
rect 4112 10218 4168 10220
rect 4008 10166 4024 10218
rect 4024 10166 4064 10218
rect 4112 10166 4148 10218
rect 4148 10166 4168 10218
rect 4008 10164 4064 10166
rect 4112 10164 4168 10166
rect 4216 10164 4272 10220
rect 4320 10218 4376 10220
rect 4424 10218 4480 10220
rect 4528 10218 4584 10220
rect 4320 10166 4324 10218
rect 4324 10166 4376 10218
rect 4424 10166 4448 10218
rect 4448 10166 4480 10218
rect 4528 10166 4572 10218
rect 4572 10166 4584 10218
rect 4320 10164 4376 10166
rect 4424 10164 4480 10166
rect 4528 10164 4584 10166
rect 4632 10218 4688 10220
rect 4736 10218 4792 10220
rect 4840 10218 4896 10220
rect 4632 10166 4644 10218
rect 4644 10166 4688 10218
rect 4736 10166 4768 10218
rect 4768 10166 4792 10218
rect 4840 10166 4892 10218
rect 4892 10166 4896 10218
rect 4632 10164 4688 10166
rect 4736 10164 4792 10166
rect 4840 10164 4896 10166
rect 4944 10164 5000 10220
rect 5048 10218 5104 10220
rect 5152 10218 5208 10220
rect 5048 10166 5068 10218
rect 5068 10166 5104 10218
rect 5152 10166 5192 10218
rect 5192 10166 5208 10218
rect 5048 10164 5104 10166
rect 5152 10164 5208 10166
rect 8316 11900 8372 11956
rect 6860 11394 6916 11396
rect 6860 11342 6862 11394
rect 6862 11342 6914 11394
rect 6914 11342 6916 11394
rect 6860 11340 6916 11342
rect 7980 11116 8036 11172
rect 5964 10834 6020 10836
rect 5964 10782 5966 10834
rect 5966 10782 6018 10834
rect 6018 10782 6020 10834
rect 5964 10780 6020 10782
rect 9212 13580 9268 13636
rect 8764 12850 8820 12852
rect 8764 12798 8766 12850
rect 8766 12798 8818 12850
rect 8818 12798 8820 12850
rect 8764 12796 8820 12798
rect 9100 12738 9156 12740
rect 9100 12686 9102 12738
rect 9102 12686 9154 12738
rect 9154 12686 9156 12738
rect 9100 12684 9156 12686
rect 8988 12402 9044 12404
rect 8988 12350 8990 12402
rect 8990 12350 9042 12402
rect 9042 12350 9044 12402
rect 8988 12348 9044 12350
rect 8988 12012 9044 12068
rect 8876 11116 8932 11172
rect 9660 15538 9716 15540
rect 9660 15486 9662 15538
rect 9662 15486 9714 15538
rect 9714 15486 9716 15538
rect 9660 15484 9716 15486
rect 9884 20018 9940 20020
rect 9884 19966 9886 20018
rect 9886 19966 9938 20018
rect 9938 19966 9940 20018
rect 9884 19964 9940 19966
rect 10556 24722 10612 24724
rect 10556 24670 10558 24722
rect 10558 24670 10610 24722
rect 10610 24670 10612 24722
rect 10556 24668 10612 24670
rect 10780 24332 10836 24388
rect 11564 24332 11620 24388
rect 11676 23826 11732 23828
rect 11676 23774 11678 23826
rect 11678 23774 11730 23826
rect 11730 23774 11732 23826
rect 11676 23772 11732 23774
rect 12572 25228 12628 25284
rect 13580 27916 13636 27972
rect 13692 28476 13748 28532
rect 13692 27692 13748 27748
rect 14700 29148 14756 29204
rect 13916 29036 13972 29092
rect 14364 28642 14420 28644
rect 14364 28590 14366 28642
rect 14366 28590 14418 28642
rect 14418 28590 14420 28642
rect 14364 28588 14420 28590
rect 15372 29202 15428 29204
rect 15372 29150 15374 29202
rect 15374 29150 15426 29202
rect 15426 29150 15428 29202
rect 15372 29148 15428 29150
rect 14924 29036 14980 29092
rect 15484 28588 15540 28644
rect 15260 28418 15316 28420
rect 15260 28366 15262 28418
rect 15262 28366 15314 28418
rect 15314 28366 15316 28418
rect 15260 28364 15316 28366
rect 14008 28250 14064 28252
rect 14112 28250 14168 28252
rect 14008 28198 14024 28250
rect 14024 28198 14064 28250
rect 14112 28198 14148 28250
rect 14148 28198 14168 28250
rect 14008 28196 14064 28198
rect 14112 28196 14168 28198
rect 14216 28196 14272 28252
rect 14320 28250 14376 28252
rect 14424 28250 14480 28252
rect 14528 28250 14584 28252
rect 14320 28198 14324 28250
rect 14324 28198 14376 28250
rect 14424 28198 14448 28250
rect 14448 28198 14480 28250
rect 14528 28198 14572 28250
rect 14572 28198 14584 28250
rect 14320 28196 14376 28198
rect 14424 28196 14480 28198
rect 14528 28196 14584 28198
rect 14632 28250 14688 28252
rect 14736 28250 14792 28252
rect 14840 28250 14896 28252
rect 14632 28198 14644 28250
rect 14644 28198 14688 28250
rect 14736 28198 14768 28250
rect 14768 28198 14792 28250
rect 14840 28198 14892 28250
rect 14892 28198 14896 28250
rect 14632 28196 14688 28198
rect 14736 28196 14792 28198
rect 14840 28196 14896 28198
rect 14944 28196 15000 28252
rect 15048 28250 15104 28252
rect 15152 28250 15208 28252
rect 15048 28198 15068 28250
rect 15068 28198 15104 28250
rect 15152 28198 15192 28250
rect 15192 28198 15208 28250
rect 15048 28196 15104 28198
rect 15152 28196 15208 28198
rect 16380 31164 16436 31220
rect 16044 30322 16100 30324
rect 16044 30270 16046 30322
rect 16046 30270 16098 30322
rect 16098 30270 16100 30322
rect 16044 30268 16100 30270
rect 16044 29372 16100 29428
rect 14028 27916 14084 27972
rect 13916 27858 13972 27860
rect 13916 27806 13918 27858
rect 13918 27806 13970 27858
rect 13970 27806 13972 27858
rect 13916 27804 13972 27806
rect 14028 27186 14084 27188
rect 14028 27134 14030 27186
rect 14030 27134 14082 27186
rect 14082 27134 14084 27186
rect 14028 27132 14084 27134
rect 14588 27970 14644 27972
rect 14588 27918 14590 27970
rect 14590 27918 14642 27970
rect 14642 27918 14644 27970
rect 14588 27916 14644 27918
rect 15708 27970 15764 27972
rect 15708 27918 15710 27970
rect 15710 27918 15762 27970
rect 15762 27918 15764 27970
rect 15708 27916 15764 27918
rect 15820 27858 15876 27860
rect 15820 27806 15822 27858
rect 15822 27806 15874 27858
rect 15874 27806 15876 27858
rect 15820 27804 15876 27806
rect 15260 27746 15316 27748
rect 15260 27694 15262 27746
rect 15262 27694 15314 27746
rect 15314 27694 15316 27746
rect 15260 27692 15316 27694
rect 17500 35196 17556 35252
rect 18284 38220 18340 38276
rect 18620 38556 18676 38612
rect 17948 37826 18004 37828
rect 17948 37774 17950 37826
rect 17950 37774 18002 37826
rect 18002 37774 18004 37826
rect 17948 37772 18004 37774
rect 17836 37490 17892 37492
rect 17836 37438 17838 37490
rect 17838 37438 17890 37490
rect 17890 37438 17892 37490
rect 17836 37436 17892 37438
rect 18060 37266 18116 37268
rect 18060 37214 18062 37266
rect 18062 37214 18114 37266
rect 18114 37214 18116 37266
rect 18060 37212 18116 37214
rect 18732 38274 18788 38276
rect 18732 38222 18734 38274
rect 18734 38222 18786 38274
rect 18786 38222 18788 38274
rect 18732 38220 18788 38222
rect 19180 39730 19236 39732
rect 19180 39678 19182 39730
rect 19182 39678 19234 39730
rect 19234 39678 19236 39730
rect 19180 39676 19236 39678
rect 19068 38556 19124 38612
rect 18956 37772 19012 37828
rect 18620 35532 18676 35588
rect 17164 33852 17220 33908
rect 17612 34802 17668 34804
rect 17612 34750 17614 34802
rect 17614 34750 17666 34802
rect 17666 34750 17668 34802
rect 17612 34748 17668 34750
rect 17836 34690 17892 34692
rect 17836 34638 17838 34690
rect 17838 34638 17890 34690
rect 17890 34638 17892 34690
rect 17836 34636 17892 34638
rect 17836 34300 17892 34356
rect 18620 35196 18676 35252
rect 18732 37324 18788 37380
rect 17052 33068 17108 33124
rect 18060 33628 18116 33684
rect 18172 34300 18228 34356
rect 17612 33068 17668 33124
rect 18508 33122 18564 33124
rect 18508 33070 18510 33122
rect 18510 33070 18562 33122
rect 18562 33070 18564 33122
rect 18508 33068 18564 33070
rect 18844 36258 18900 36260
rect 18844 36206 18846 36258
rect 18846 36206 18898 36258
rect 18898 36206 18900 36258
rect 18844 36204 18900 36206
rect 20748 41132 20804 41188
rect 20972 39676 21028 39732
rect 19516 39340 19572 39396
rect 19068 34802 19124 34804
rect 19068 34750 19070 34802
rect 19070 34750 19122 34802
rect 19122 34750 19124 34802
rect 19068 34748 19124 34750
rect 18956 33628 19012 33684
rect 19404 35532 19460 35588
rect 19852 38668 19908 38724
rect 19628 38050 19684 38052
rect 19628 37998 19630 38050
rect 19630 37998 19682 38050
rect 19682 37998 19684 38050
rect 19628 37996 19684 37998
rect 21532 43708 21588 43764
rect 21420 43260 21476 43316
rect 21756 43372 21812 43428
rect 22540 47458 22596 47460
rect 22540 47406 22542 47458
rect 22542 47406 22594 47458
rect 22594 47406 22596 47458
rect 22540 47404 22596 47406
rect 22876 48412 22932 48468
rect 23436 51884 23492 51940
rect 23772 51602 23828 51604
rect 23772 51550 23774 51602
rect 23774 51550 23826 51602
rect 23826 51550 23828 51602
rect 23772 51548 23828 51550
rect 24220 52108 24276 52164
rect 24892 51548 24948 51604
rect 25452 52274 25508 52276
rect 25452 52222 25454 52274
rect 25454 52222 25506 52274
rect 25506 52222 25508 52274
rect 25452 52220 25508 52222
rect 24008 50986 24064 50988
rect 24112 50986 24168 50988
rect 24008 50934 24024 50986
rect 24024 50934 24064 50986
rect 24112 50934 24148 50986
rect 24148 50934 24168 50986
rect 24008 50932 24064 50934
rect 24112 50932 24168 50934
rect 24216 50932 24272 50988
rect 24320 50986 24376 50988
rect 24424 50986 24480 50988
rect 24528 50986 24584 50988
rect 24320 50934 24324 50986
rect 24324 50934 24376 50986
rect 24424 50934 24448 50986
rect 24448 50934 24480 50986
rect 24528 50934 24572 50986
rect 24572 50934 24584 50986
rect 24320 50932 24376 50934
rect 24424 50932 24480 50934
rect 24528 50932 24584 50934
rect 24632 50986 24688 50988
rect 24736 50986 24792 50988
rect 24840 50986 24896 50988
rect 24632 50934 24644 50986
rect 24644 50934 24688 50986
rect 24736 50934 24768 50986
rect 24768 50934 24792 50986
rect 24840 50934 24892 50986
rect 24892 50934 24896 50986
rect 24632 50932 24688 50934
rect 24736 50932 24792 50934
rect 24840 50932 24896 50934
rect 24944 50932 25000 50988
rect 25048 50986 25104 50988
rect 25152 50986 25208 50988
rect 25048 50934 25068 50986
rect 25068 50934 25104 50986
rect 25152 50934 25192 50986
rect 25192 50934 25208 50986
rect 25048 50932 25104 50934
rect 25152 50932 25208 50934
rect 24332 50706 24388 50708
rect 24332 50654 24334 50706
rect 24334 50654 24386 50706
rect 24386 50654 24388 50706
rect 24332 50652 24388 50654
rect 24892 50706 24948 50708
rect 24892 50654 24894 50706
rect 24894 50654 24946 50706
rect 24946 50654 24948 50706
rect 24892 50652 24948 50654
rect 23996 50428 24052 50484
rect 23324 48636 23380 48692
rect 22764 46844 22820 46900
rect 22876 46732 22932 46788
rect 22988 44044 23044 44100
rect 23660 48354 23716 48356
rect 23660 48302 23662 48354
rect 23662 48302 23714 48354
rect 23714 48302 23716 48354
rect 23660 48300 23716 48302
rect 24008 49418 24064 49420
rect 24112 49418 24168 49420
rect 24008 49366 24024 49418
rect 24024 49366 24064 49418
rect 24112 49366 24148 49418
rect 24148 49366 24168 49418
rect 24008 49364 24064 49366
rect 24112 49364 24168 49366
rect 24216 49364 24272 49420
rect 24320 49418 24376 49420
rect 24424 49418 24480 49420
rect 24528 49418 24584 49420
rect 24320 49366 24324 49418
rect 24324 49366 24376 49418
rect 24424 49366 24448 49418
rect 24448 49366 24480 49418
rect 24528 49366 24572 49418
rect 24572 49366 24584 49418
rect 24320 49364 24376 49366
rect 24424 49364 24480 49366
rect 24528 49364 24584 49366
rect 24632 49418 24688 49420
rect 24736 49418 24792 49420
rect 24840 49418 24896 49420
rect 24632 49366 24644 49418
rect 24644 49366 24688 49418
rect 24736 49366 24768 49418
rect 24768 49366 24792 49418
rect 24840 49366 24892 49418
rect 24892 49366 24896 49418
rect 24632 49364 24688 49366
rect 24736 49364 24792 49366
rect 24840 49364 24896 49366
rect 24944 49364 25000 49420
rect 25048 49418 25104 49420
rect 25152 49418 25208 49420
rect 25048 49366 25068 49418
rect 25068 49366 25104 49418
rect 25152 49366 25192 49418
rect 25192 49366 25208 49418
rect 25048 49364 25104 49366
rect 25152 49364 25208 49366
rect 24332 49026 24388 49028
rect 24332 48974 24334 49026
rect 24334 48974 24386 49026
rect 24386 48974 24388 49026
rect 24332 48972 24388 48974
rect 25900 53452 25956 53508
rect 25676 52108 25732 52164
rect 26460 53954 26516 53956
rect 26460 53902 26462 53954
rect 26462 53902 26514 53954
rect 26514 53902 26516 53954
rect 26460 53900 26516 53902
rect 26796 53900 26852 53956
rect 26572 53788 26628 53844
rect 25788 52050 25844 52052
rect 25788 51998 25790 52050
rect 25790 51998 25842 52050
rect 25842 51998 25844 52050
rect 25788 51996 25844 51998
rect 25788 51602 25844 51604
rect 25788 51550 25790 51602
rect 25790 51550 25842 51602
rect 25842 51550 25844 51602
rect 25788 51548 25844 51550
rect 26460 53116 26516 53172
rect 26236 51548 26292 51604
rect 25564 50652 25620 50708
rect 25340 48860 25396 48916
rect 25452 49196 25508 49252
rect 23772 48188 23828 48244
rect 23772 47516 23828 47572
rect 23884 48412 23940 48468
rect 23660 47458 23716 47460
rect 23660 47406 23662 47458
rect 23662 47406 23714 47458
rect 23714 47406 23716 47458
rect 23660 47404 23716 47406
rect 24444 48466 24500 48468
rect 24444 48414 24446 48466
rect 24446 48414 24498 48466
rect 24498 48414 24500 48466
rect 24444 48412 24500 48414
rect 25340 48300 25396 48356
rect 24008 47850 24064 47852
rect 24112 47850 24168 47852
rect 24008 47798 24024 47850
rect 24024 47798 24064 47850
rect 24112 47798 24148 47850
rect 24148 47798 24168 47850
rect 24008 47796 24064 47798
rect 24112 47796 24168 47798
rect 24216 47796 24272 47852
rect 24320 47850 24376 47852
rect 24424 47850 24480 47852
rect 24528 47850 24584 47852
rect 24320 47798 24324 47850
rect 24324 47798 24376 47850
rect 24424 47798 24448 47850
rect 24448 47798 24480 47850
rect 24528 47798 24572 47850
rect 24572 47798 24584 47850
rect 24320 47796 24376 47798
rect 24424 47796 24480 47798
rect 24528 47796 24584 47798
rect 24632 47850 24688 47852
rect 24736 47850 24792 47852
rect 24840 47850 24896 47852
rect 24632 47798 24644 47850
rect 24644 47798 24688 47850
rect 24736 47798 24768 47850
rect 24768 47798 24792 47850
rect 24840 47798 24892 47850
rect 24892 47798 24896 47850
rect 24632 47796 24688 47798
rect 24736 47796 24792 47798
rect 24840 47796 24896 47798
rect 24944 47796 25000 47852
rect 25048 47850 25104 47852
rect 25152 47850 25208 47852
rect 25048 47798 25068 47850
rect 25068 47798 25104 47850
rect 25152 47798 25192 47850
rect 25192 47798 25208 47850
rect 25048 47796 25104 47798
rect 25152 47796 25208 47798
rect 24444 47516 24500 47572
rect 23996 47180 24052 47236
rect 23772 46844 23828 46900
rect 23548 45330 23604 45332
rect 23548 45278 23550 45330
rect 23550 45278 23602 45330
rect 23602 45278 23604 45330
rect 23548 45276 23604 45278
rect 23436 45164 23492 45220
rect 22540 42812 22596 42868
rect 22316 42754 22372 42756
rect 22316 42702 22318 42754
rect 22318 42702 22370 42754
rect 22370 42702 22372 42754
rect 22316 42700 22372 42702
rect 21532 41298 21588 41300
rect 21532 41246 21534 41298
rect 21534 41246 21586 41298
rect 21586 41246 21588 41298
rect 21532 41244 21588 41246
rect 21868 41186 21924 41188
rect 21868 41134 21870 41186
rect 21870 41134 21922 41186
rect 21922 41134 21924 41186
rect 21868 41132 21924 41134
rect 21532 40348 21588 40404
rect 21084 37324 21140 37380
rect 19628 37212 19684 37268
rect 20188 36204 20244 36260
rect 19852 35084 19908 35140
rect 20300 35868 20356 35924
rect 19516 34802 19572 34804
rect 19516 34750 19518 34802
rect 19518 34750 19570 34802
rect 19570 34750 19572 34802
rect 19516 34748 19572 34750
rect 19292 33404 19348 33460
rect 20636 35138 20692 35140
rect 20636 35086 20638 35138
rect 20638 35086 20690 35138
rect 20690 35086 20692 35138
rect 20636 35084 20692 35086
rect 20076 33964 20132 34020
rect 16604 31724 16660 31780
rect 17052 31778 17108 31780
rect 17052 31726 17054 31778
rect 17054 31726 17106 31778
rect 17106 31726 17108 31778
rect 17052 31724 17108 31726
rect 18172 31778 18228 31780
rect 18172 31726 18174 31778
rect 18174 31726 18226 31778
rect 18226 31726 18228 31778
rect 18172 31724 18228 31726
rect 17276 31612 17332 31668
rect 17388 31500 17444 31556
rect 17500 31164 17556 31220
rect 17388 30770 17444 30772
rect 17388 30718 17390 30770
rect 17390 30718 17442 30770
rect 17442 30718 17444 30770
rect 17388 30716 17444 30718
rect 17164 30156 17220 30212
rect 18732 31500 18788 31556
rect 17836 30156 17892 30212
rect 16380 28476 16436 28532
rect 16828 28476 16884 28532
rect 15148 27186 15204 27188
rect 15148 27134 15150 27186
rect 15150 27134 15202 27186
rect 15202 27134 15204 27186
rect 15148 27132 15204 27134
rect 15484 27020 15540 27076
rect 14364 26908 14420 26964
rect 14700 26962 14756 26964
rect 14700 26910 14702 26962
rect 14702 26910 14754 26962
rect 14754 26910 14756 26962
rect 14700 26908 14756 26910
rect 14008 26682 14064 26684
rect 14112 26682 14168 26684
rect 14008 26630 14024 26682
rect 14024 26630 14064 26682
rect 14112 26630 14148 26682
rect 14148 26630 14168 26682
rect 14008 26628 14064 26630
rect 14112 26628 14168 26630
rect 14216 26628 14272 26684
rect 14320 26682 14376 26684
rect 14424 26682 14480 26684
rect 14528 26682 14584 26684
rect 14320 26630 14324 26682
rect 14324 26630 14376 26682
rect 14424 26630 14448 26682
rect 14448 26630 14480 26682
rect 14528 26630 14572 26682
rect 14572 26630 14584 26682
rect 14320 26628 14376 26630
rect 14424 26628 14480 26630
rect 14528 26628 14584 26630
rect 14632 26682 14688 26684
rect 14736 26682 14792 26684
rect 14840 26682 14896 26684
rect 14632 26630 14644 26682
rect 14644 26630 14688 26682
rect 14736 26630 14768 26682
rect 14768 26630 14792 26682
rect 14840 26630 14892 26682
rect 14892 26630 14896 26682
rect 14632 26628 14688 26630
rect 14736 26628 14792 26630
rect 14840 26628 14896 26630
rect 14944 26628 15000 26684
rect 15048 26682 15104 26684
rect 15152 26682 15208 26684
rect 15048 26630 15068 26682
rect 15068 26630 15104 26682
rect 15152 26630 15192 26682
rect 15192 26630 15208 26682
rect 15048 26628 15104 26630
rect 15152 26628 15208 26630
rect 14028 25618 14084 25620
rect 14028 25566 14030 25618
rect 14030 25566 14082 25618
rect 14082 25566 14084 25618
rect 14028 25564 14084 25566
rect 14476 25564 14532 25620
rect 13580 25282 13636 25284
rect 13580 25230 13582 25282
rect 13582 25230 13634 25282
rect 13634 25230 13636 25282
rect 13580 25228 13636 25230
rect 15036 25282 15092 25284
rect 15036 25230 15038 25282
rect 15038 25230 15090 25282
rect 15090 25230 15092 25282
rect 15036 25228 15092 25230
rect 16380 26908 16436 26964
rect 14008 25114 14064 25116
rect 14112 25114 14168 25116
rect 14008 25062 14024 25114
rect 14024 25062 14064 25114
rect 14112 25062 14148 25114
rect 14148 25062 14168 25114
rect 14008 25060 14064 25062
rect 14112 25060 14168 25062
rect 14216 25060 14272 25116
rect 14320 25114 14376 25116
rect 14424 25114 14480 25116
rect 14528 25114 14584 25116
rect 14320 25062 14324 25114
rect 14324 25062 14376 25114
rect 14424 25062 14448 25114
rect 14448 25062 14480 25114
rect 14528 25062 14572 25114
rect 14572 25062 14584 25114
rect 14320 25060 14376 25062
rect 14424 25060 14480 25062
rect 14528 25060 14584 25062
rect 14632 25114 14688 25116
rect 14736 25114 14792 25116
rect 14840 25114 14896 25116
rect 14632 25062 14644 25114
rect 14644 25062 14688 25114
rect 14736 25062 14768 25114
rect 14768 25062 14792 25114
rect 14840 25062 14892 25114
rect 14892 25062 14896 25114
rect 14632 25060 14688 25062
rect 14736 25060 14792 25062
rect 14840 25060 14896 25062
rect 14944 25060 15000 25116
rect 15048 25114 15104 25116
rect 15152 25114 15208 25116
rect 15048 25062 15068 25114
rect 15068 25062 15104 25114
rect 15152 25062 15192 25114
rect 15192 25062 15208 25114
rect 15048 25060 15104 25062
rect 15152 25060 15208 25062
rect 12572 24780 12628 24836
rect 14028 24834 14084 24836
rect 14028 24782 14030 24834
rect 14030 24782 14082 24834
rect 14082 24782 14084 24834
rect 14028 24780 14084 24782
rect 12236 23772 12292 23828
rect 11228 23660 11284 23716
rect 11116 23154 11172 23156
rect 11116 23102 11118 23154
rect 11118 23102 11170 23154
rect 11170 23102 11172 23154
rect 11116 23100 11172 23102
rect 10556 22540 10612 22596
rect 11900 23714 11956 23716
rect 11900 23662 11902 23714
rect 11902 23662 11954 23714
rect 11954 23662 11956 23714
rect 11900 23660 11956 23662
rect 12460 22988 12516 23044
rect 11788 22316 11844 22372
rect 11564 22258 11620 22260
rect 11564 22206 11566 22258
rect 11566 22206 11618 22258
rect 11618 22206 11620 22258
rect 11564 22204 11620 22206
rect 10332 21308 10388 21364
rect 10332 20636 10388 20692
rect 10332 20130 10388 20132
rect 10332 20078 10334 20130
rect 10334 20078 10386 20130
rect 10386 20078 10388 20130
rect 10332 20076 10388 20078
rect 12460 22370 12516 22372
rect 12460 22318 12462 22370
rect 12462 22318 12514 22370
rect 12514 22318 12516 22370
rect 12460 22316 12516 22318
rect 12124 22258 12180 22260
rect 12124 22206 12126 22258
rect 12126 22206 12178 22258
rect 12178 22206 12180 22258
rect 12124 22204 12180 22206
rect 12236 22146 12292 22148
rect 12236 22094 12238 22146
rect 12238 22094 12290 22146
rect 12290 22094 12292 22146
rect 12236 22092 12292 22094
rect 10556 20076 10612 20132
rect 11564 20076 11620 20132
rect 11788 20076 11844 20132
rect 13356 23212 13412 23268
rect 12572 21420 12628 21476
rect 12908 20748 12964 20804
rect 13132 21362 13188 21364
rect 13132 21310 13134 21362
rect 13134 21310 13186 21362
rect 13186 21310 13188 21362
rect 13132 21308 13188 21310
rect 12348 20524 12404 20580
rect 13132 20188 13188 20244
rect 9996 17666 10052 17668
rect 9996 17614 9998 17666
rect 9998 17614 10050 17666
rect 10050 17614 10052 17666
rect 9996 17612 10052 17614
rect 10892 17612 10948 17668
rect 10780 17442 10836 17444
rect 10780 17390 10782 17442
rect 10782 17390 10834 17442
rect 10834 17390 10836 17442
rect 10780 17388 10836 17390
rect 10444 16994 10500 16996
rect 10444 16942 10446 16994
rect 10446 16942 10498 16994
rect 10498 16942 10500 16994
rect 10444 16940 10500 16942
rect 9548 15426 9604 15428
rect 9548 15374 9550 15426
rect 9550 15374 9602 15426
rect 9602 15374 9604 15426
rect 9548 15372 9604 15374
rect 11116 17388 11172 17444
rect 11228 17276 11284 17332
rect 11004 16994 11060 16996
rect 11004 16942 11006 16994
rect 11006 16942 11058 16994
rect 11058 16942 11060 16994
rect 11004 16940 11060 16942
rect 11228 16716 11284 16772
rect 11228 16210 11284 16212
rect 11228 16158 11230 16210
rect 11230 16158 11282 16210
rect 11282 16158 11284 16210
rect 11228 16156 11284 16158
rect 9996 14476 10052 14532
rect 9548 14364 9604 14420
rect 10556 14924 10612 14980
rect 10556 14476 10612 14532
rect 9548 13858 9604 13860
rect 9548 13806 9550 13858
rect 9550 13806 9602 13858
rect 9602 13806 9604 13858
rect 9548 13804 9604 13806
rect 9548 13580 9604 13636
rect 9884 13916 9940 13972
rect 10108 13468 10164 13524
rect 9772 12796 9828 12852
rect 11564 17388 11620 17444
rect 12572 20130 12628 20132
rect 12572 20078 12574 20130
rect 12574 20078 12626 20130
rect 12626 20078 12628 20130
rect 12572 20076 12628 20078
rect 12236 18562 12292 18564
rect 12236 18510 12238 18562
rect 12238 18510 12290 18562
rect 12290 18510 12292 18562
rect 12236 18508 12292 18510
rect 12012 17948 12068 18004
rect 12572 18284 12628 18340
rect 11900 17666 11956 17668
rect 11900 17614 11902 17666
rect 11902 17614 11954 17666
rect 11954 17614 11956 17666
rect 11900 17612 11956 17614
rect 12348 17442 12404 17444
rect 12348 17390 12350 17442
rect 12350 17390 12402 17442
rect 12402 17390 12404 17442
rect 12348 17388 12404 17390
rect 12572 17276 12628 17332
rect 13020 18284 13076 18340
rect 12684 17948 12740 18004
rect 11788 16940 11844 16996
rect 12348 16940 12404 16996
rect 12124 16716 12180 16772
rect 12908 17388 12964 17444
rect 12684 16604 12740 16660
rect 11564 15372 11620 15428
rect 12236 15820 12292 15876
rect 11452 14924 11508 14980
rect 11116 14530 11172 14532
rect 11116 14478 11118 14530
rect 11118 14478 11170 14530
rect 11170 14478 11172 14530
rect 11116 14476 11172 14478
rect 11452 14642 11508 14644
rect 11452 14590 11454 14642
rect 11454 14590 11506 14642
rect 11506 14590 11508 14642
rect 11452 14588 11508 14590
rect 10780 13804 10836 13860
rect 10444 13020 10500 13076
rect 11900 14530 11956 14532
rect 11900 14478 11902 14530
rect 11902 14478 11954 14530
rect 11954 14478 11956 14530
rect 11900 14476 11956 14478
rect 11228 13916 11284 13972
rect 12348 14924 12404 14980
rect 11452 13580 11508 13636
rect 10332 12402 10388 12404
rect 10332 12350 10334 12402
rect 10334 12350 10386 12402
rect 10386 12350 10388 12402
rect 10332 12348 10388 12350
rect 12348 14530 12404 14532
rect 12348 14478 12350 14530
rect 12350 14478 12402 14530
rect 12402 14478 12404 14530
rect 12348 14476 12404 14478
rect 12348 13970 12404 13972
rect 12348 13918 12350 13970
rect 12350 13918 12402 13970
rect 12402 13918 12404 13970
rect 12348 13916 12404 13918
rect 13468 23100 13524 23156
rect 13580 23660 13636 23716
rect 15484 25228 15540 25284
rect 14364 23772 14420 23828
rect 15372 24444 15428 24500
rect 13916 23660 13972 23716
rect 16492 24332 16548 24388
rect 16492 23714 16548 23716
rect 16492 23662 16494 23714
rect 16494 23662 16546 23714
rect 16546 23662 16548 23714
rect 16492 23660 16548 23662
rect 16604 23772 16660 23828
rect 13692 23436 13748 23492
rect 14008 23546 14064 23548
rect 14112 23546 14168 23548
rect 14008 23494 14024 23546
rect 14024 23494 14064 23546
rect 14112 23494 14148 23546
rect 14148 23494 14168 23546
rect 14008 23492 14064 23494
rect 14112 23492 14168 23494
rect 14216 23492 14272 23548
rect 14320 23546 14376 23548
rect 14424 23546 14480 23548
rect 14528 23546 14584 23548
rect 14320 23494 14324 23546
rect 14324 23494 14376 23546
rect 14424 23494 14448 23546
rect 14448 23494 14480 23546
rect 14528 23494 14572 23546
rect 14572 23494 14584 23546
rect 14320 23492 14376 23494
rect 14424 23492 14480 23494
rect 14528 23492 14584 23494
rect 14632 23546 14688 23548
rect 14736 23546 14792 23548
rect 14840 23546 14896 23548
rect 14632 23494 14644 23546
rect 14644 23494 14688 23546
rect 14736 23494 14768 23546
rect 14768 23494 14792 23546
rect 14840 23494 14892 23546
rect 14892 23494 14896 23546
rect 14632 23492 14688 23494
rect 14736 23492 14792 23494
rect 14840 23492 14896 23494
rect 14944 23492 15000 23548
rect 15048 23546 15104 23548
rect 15152 23546 15208 23548
rect 15048 23494 15068 23546
rect 15068 23494 15104 23546
rect 15152 23494 15192 23546
rect 15192 23494 15208 23546
rect 15048 23492 15104 23494
rect 15152 23492 15208 23494
rect 15484 23548 15540 23604
rect 16268 23548 16324 23604
rect 15932 23324 15988 23380
rect 14588 23154 14644 23156
rect 14588 23102 14590 23154
rect 14590 23102 14642 23154
rect 14642 23102 14644 23154
rect 14588 23100 14644 23102
rect 13804 22652 13860 22708
rect 13916 22876 13972 22932
rect 15372 22370 15428 22372
rect 15372 22318 15374 22370
rect 15374 22318 15426 22370
rect 15426 22318 15428 22370
rect 15372 22316 15428 22318
rect 14140 22258 14196 22260
rect 14140 22206 14142 22258
rect 14142 22206 14194 22258
rect 14194 22206 14196 22258
rect 14140 22204 14196 22206
rect 14700 22258 14756 22260
rect 14700 22206 14702 22258
rect 14702 22206 14754 22258
rect 14754 22206 14756 22258
rect 14700 22204 14756 22206
rect 13692 22092 13748 22148
rect 14008 21978 14064 21980
rect 14112 21978 14168 21980
rect 14008 21926 14024 21978
rect 14024 21926 14064 21978
rect 14112 21926 14148 21978
rect 14148 21926 14168 21978
rect 14008 21924 14064 21926
rect 14112 21924 14168 21926
rect 14216 21924 14272 21980
rect 14320 21978 14376 21980
rect 14424 21978 14480 21980
rect 14528 21978 14584 21980
rect 14320 21926 14324 21978
rect 14324 21926 14376 21978
rect 14424 21926 14448 21978
rect 14448 21926 14480 21978
rect 14528 21926 14572 21978
rect 14572 21926 14584 21978
rect 14320 21924 14376 21926
rect 14424 21924 14480 21926
rect 14528 21924 14584 21926
rect 14632 21978 14688 21980
rect 14736 21978 14792 21980
rect 14840 21978 14896 21980
rect 14632 21926 14644 21978
rect 14644 21926 14688 21978
rect 14736 21926 14768 21978
rect 14768 21926 14792 21978
rect 14840 21926 14892 21978
rect 14892 21926 14896 21978
rect 14632 21924 14688 21926
rect 14736 21924 14792 21926
rect 14840 21924 14896 21926
rect 14944 21924 15000 21980
rect 15048 21978 15104 21980
rect 15152 21978 15208 21980
rect 15048 21926 15068 21978
rect 15068 21926 15104 21978
rect 15152 21926 15192 21978
rect 15192 21926 15208 21978
rect 15048 21924 15104 21926
rect 15152 21924 15208 21926
rect 15260 21756 15316 21812
rect 13692 21196 13748 21252
rect 14140 20972 14196 21028
rect 13692 20860 13748 20916
rect 14140 20578 14196 20580
rect 14140 20526 14142 20578
rect 14142 20526 14194 20578
rect 14194 20526 14196 20578
rect 14140 20524 14196 20526
rect 14588 20524 14644 20580
rect 15148 21308 15204 21364
rect 15148 20914 15204 20916
rect 15148 20862 15150 20914
rect 15150 20862 15202 20914
rect 15202 20862 15204 20914
rect 15148 20860 15204 20862
rect 15596 21308 15652 21364
rect 14008 20410 14064 20412
rect 14112 20410 14168 20412
rect 14008 20358 14024 20410
rect 14024 20358 14064 20410
rect 14112 20358 14148 20410
rect 14148 20358 14168 20410
rect 14008 20356 14064 20358
rect 14112 20356 14168 20358
rect 14216 20356 14272 20412
rect 14320 20410 14376 20412
rect 14424 20410 14480 20412
rect 14528 20410 14584 20412
rect 14320 20358 14324 20410
rect 14324 20358 14376 20410
rect 14424 20358 14448 20410
rect 14448 20358 14480 20410
rect 14528 20358 14572 20410
rect 14572 20358 14584 20410
rect 14320 20356 14376 20358
rect 14424 20356 14480 20358
rect 14528 20356 14584 20358
rect 14632 20410 14688 20412
rect 14736 20410 14792 20412
rect 14840 20410 14896 20412
rect 14632 20358 14644 20410
rect 14644 20358 14688 20410
rect 14736 20358 14768 20410
rect 14768 20358 14792 20410
rect 14840 20358 14892 20410
rect 14892 20358 14896 20410
rect 14632 20356 14688 20358
rect 14736 20356 14792 20358
rect 14840 20356 14896 20358
rect 14944 20356 15000 20412
rect 15048 20410 15104 20412
rect 15152 20410 15208 20412
rect 15048 20358 15068 20410
rect 15068 20358 15104 20410
rect 15152 20358 15192 20410
rect 15192 20358 15208 20410
rect 15048 20356 15104 20358
rect 15152 20356 15208 20358
rect 14028 20188 14084 20244
rect 13692 20076 13748 20132
rect 13916 19964 13972 20020
rect 14252 19906 14308 19908
rect 14252 19854 14254 19906
rect 14254 19854 14306 19906
rect 14306 19854 14308 19906
rect 14252 19852 14308 19854
rect 13692 19068 13748 19124
rect 14812 20018 14868 20020
rect 14812 19966 14814 20018
rect 14814 19966 14866 20018
rect 14866 19966 14868 20018
rect 14812 19964 14868 19966
rect 14588 19346 14644 19348
rect 14588 19294 14590 19346
rect 14590 19294 14642 19346
rect 14642 19294 14644 19346
rect 14588 19292 14644 19294
rect 14700 19234 14756 19236
rect 14700 19182 14702 19234
rect 14702 19182 14754 19234
rect 14754 19182 14756 19234
rect 14700 19180 14756 19182
rect 15596 20076 15652 20132
rect 16044 20076 16100 20132
rect 15708 19852 15764 19908
rect 14364 19068 14420 19124
rect 14252 19010 14308 19012
rect 14252 18958 14254 19010
rect 14254 18958 14306 19010
rect 14306 18958 14308 19010
rect 14252 18956 14308 18958
rect 14008 18842 14064 18844
rect 14112 18842 14168 18844
rect 14008 18790 14024 18842
rect 14024 18790 14064 18842
rect 14112 18790 14148 18842
rect 14148 18790 14168 18842
rect 14008 18788 14064 18790
rect 14112 18788 14168 18790
rect 14216 18788 14272 18844
rect 14320 18842 14376 18844
rect 14424 18842 14480 18844
rect 14528 18842 14584 18844
rect 14320 18790 14324 18842
rect 14324 18790 14376 18842
rect 14424 18790 14448 18842
rect 14448 18790 14480 18842
rect 14528 18790 14572 18842
rect 14572 18790 14584 18842
rect 14320 18788 14376 18790
rect 14424 18788 14480 18790
rect 14528 18788 14584 18790
rect 14632 18842 14688 18844
rect 14736 18842 14792 18844
rect 14840 18842 14896 18844
rect 14632 18790 14644 18842
rect 14644 18790 14688 18842
rect 14736 18790 14768 18842
rect 14768 18790 14792 18842
rect 14840 18790 14892 18842
rect 14892 18790 14896 18842
rect 14632 18788 14688 18790
rect 14736 18788 14792 18790
rect 14840 18788 14896 18790
rect 14944 18788 15000 18844
rect 15048 18842 15104 18844
rect 15152 18842 15208 18844
rect 15048 18790 15068 18842
rect 15068 18790 15104 18842
rect 15152 18790 15192 18842
rect 15192 18790 15208 18842
rect 15048 18788 15104 18790
rect 15152 18788 15208 18790
rect 13916 18508 13972 18564
rect 15820 19292 15876 19348
rect 14812 18284 14868 18340
rect 15820 18284 15876 18340
rect 13804 17948 13860 18004
rect 13244 16716 13300 16772
rect 13580 16604 13636 16660
rect 13244 16156 13300 16212
rect 13356 16380 13412 16436
rect 13132 15820 13188 15876
rect 14364 17442 14420 17444
rect 14364 17390 14366 17442
rect 14366 17390 14418 17442
rect 14418 17390 14420 17442
rect 14364 17388 14420 17390
rect 14008 17274 14064 17276
rect 14112 17274 14168 17276
rect 14008 17222 14024 17274
rect 14024 17222 14064 17274
rect 14112 17222 14148 17274
rect 14148 17222 14168 17274
rect 14008 17220 14064 17222
rect 14112 17220 14168 17222
rect 14216 17220 14272 17276
rect 14320 17274 14376 17276
rect 14424 17274 14480 17276
rect 14528 17274 14584 17276
rect 14320 17222 14324 17274
rect 14324 17222 14376 17274
rect 14424 17222 14448 17274
rect 14448 17222 14480 17274
rect 14528 17222 14572 17274
rect 14572 17222 14584 17274
rect 14320 17220 14376 17222
rect 14424 17220 14480 17222
rect 14528 17220 14584 17222
rect 14632 17274 14688 17276
rect 14736 17274 14792 17276
rect 14840 17274 14896 17276
rect 14632 17222 14644 17274
rect 14644 17222 14688 17274
rect 14736 17222 14768 17274
rect 14768 17222 14792 17274
rect 14840 17222 14892 17274
rect 14892 17222 14896 17274
rect 14632 17220 14688 17222
rect 14736 17220 14792 17222
rect 14840 17220 14896 17222
rect 14944 17220 15000 17276
rect 15048 17274 15104 17276
rect 15152 17274 15208 17276
rect 15048 17222 15068 17274
rect 15068 17222 15104 17274
rect 15152 17222 15192 17274
rect 15192 17222 15208 17274
rect 15048 17220 15104 17222
rect 15152 17220 15208 17222
rect 15372 17164 15428 17220
rect 14924 17052 14980 17108
rect 14028 16268 14084 16324
rect 14028 15932 14084 15988
rect 14700 16210 14756 16212
rect 14700 16158 14702 16210
rect 14702 16158 14754 16210
rect 14754 16158 14756 16210
rect 14700 16156 14756 16158
rect 15484 16994 15540 16996
rect 15484 16942 15486 16994
rect 15486 16942 15538 16994
rect 15538 16942 15540 16994
rect 15484 16940 15540 16942
rect 15708 16940 15764 16996
rect 15596 16828 15652 16884
rect 14588 15932 14644 15988
rect 14140 15874 14196 15876
rect 14140 15822 14142 15874
rect 14142 15822 14194 15874
rect 14194 15822 14196 15874
rect 14140 15820 14196 15822
rect 12796 14924 12852 14980
rect 13356 14924 13412 14980
rect 13132 14588 13188 14644
rect 13468 13916 13524 13972
rect 12460 13692 12516 13748
rect 13244 13692 13300 13748
rect 11676 13020 11732 13076
rect 10892 12402 10948 12404
rect 10892 12350 10894 12402
rect 10894 12350 10946 12402
rect 10946 12350 10948 12402
rect 10892 12348 10948 12350
rect 10220 12178 10276 12180
rect 10220 12126 10222 12178
rect 10222 12126 10274 12178
rect 10274 12126 10276 12178
rect 10220 12124 10276 12126
rect 9660 11116 9716 11172
rect 10892 11004 10948 11060
rect 4008 8650 4064 8652
rect 4112 8650 4168 8652
rect 4008 8598 4024 8650
rect 4024 8598 4064 8650
rect 4112 8598 4148 8650
rect 4148 8598 4168 8650
rect 4008 8596 4064 8598
rect 4112 8596 4168 8598
rect 4216 8596 4272 8652
rect 4320 8650 4376 8652
rect 4424 8650 4480 8652
rect 4528 8650 4584 8652
rect 4320 8598 4324 8650
rect 4324 8598 4376 8650
rect 4424 8598 4448 8650
rect 4448 8598 4480 8650
rect 4528 8598 4572 8650
rect 4572 8598 4584 8650
rect 4320 8596 4376 8598
rect 4424 8596 4480 8598
rect 4528 8596 4584 8598
rect 4632 8650 4688 8652
rect 4736 8650 4792 8652
rect 4840 8650 4896 8652
rect 4632 8598 4644 8650
rect 4644 8598 4688 8650
rect 4736 8598 4768 8650
rect 4768 8598 4792 8650
rect 4840 8598 4892 8650
rect 4892 8598 4896 8650
rect 4632 8596 4688 8598
rect 4736 8596 4792 8598
rect 4840 8596 4896 8598
rect 4944 8596 5000 8652
rect 5048 8650 5104 8652
rect 5152 8650 5208 8652
rect 5048 8598 5068 8650
rect 5068 8598 5104 8650
rect 5152 8598 5192 8650
rect 5192 8598 5208 8650
rect 5048 8596 5104 8598
rect 5152 8596 5208 8598
rect 5404 7980 5460 8036
rect 4732 7698 4788 7700
rect 4732 7646 4734 7698
rect 4734 7646 4786 7698
rect 4786 7646 4788 7698
rect 4732 7644 4788 7646
rect 4008 7082 4064 7084
rect 4112 7082 4168 7084
rect 4008 7030 4024 7082
rect 4024 7030 4064 7082
rect 4112 7030 4148 7082
rect 4148 7030 4168 7082
rect 4008 7028 4064 7030
rect 4112 7028 4168 7030
rect 4216 7028 4272 7084
rect 4320 7082 4376 7084
rect 4424 7082 4480 7084
rect 4528 7082 4584 7084
rect 4320 7030 4324 7082
rect 4324 7030 4376 7082
rect 4424 7030 4448 7082
rect 4448 7030 4480 7082
rect 4528 7030 4572 7082
rect 4572 7030 4584 7082
rect 4320 7028 4376 7030
rect 4424 7028 4480 7030
rect 4528 7028 4584 7030
rect 4632 7082 4688 7084
rect 4736 7082 4792 7084
rect 4840 7082 4896 7084
rect 4632 7030 4644 7082
rect 4644 7030 4688 7082
rect 4736 7030 4768 7082
rect 4768 7030 4792 7082
rect 4840 7030 4892 7082
rect 4892 7030 4896 7082
rect 4632 7028 4688 7030
rect 4736 7028 4792 7030
rect 4840 7028 4896 7030
rect 4944 7028 5000 7084
rect 5048 7082 5104 7084
rect 5152 7082 5208 7084
rect 5048 7030 5068 7082
rect 5068 7030 5104 7082
rect 5152 7030 5192 7082
rect 5192 7030 5208 7082
rect 5048 7028 5104 7030
rect 5152 7028 5208 7030
rect 3612 6748 3668 6804
rect 4172 6860 4228 6916
rect 2492 6690 2548 6692
rect 2492 6638 2494 6690
rect 2494 6638 2546 6690
rect 2546 6638 2548 6690
rect 2492 6636 2548 6638
rect 4060 6690 4116 6692
rect 4060 6638 4062 6690
rect 4062 6638 4114 6690
rect 4114 6638 4116 6690
rect 4060 6636 4116 6638
rect 3052 6466 3108 6468
rect 3052 6414 3054 6466
rect 3054 6414 3106 6466
rect 3106 6414 3108 6466
rect 3052 6412 3108 6414
rect 2156 5964 2212 6020
rect 3500 6018 3556 6020
rect 3500 5966 3502 6018
rect 3502 5966 3554 6018
rect 3554 5966 3556 6018
rect 3500 5964 3556 5966
rect 2044 5628 2100 5684
rect 1932 4284 1988 4340
rect 4508 6802 4564 6804
rect 4508 6750 4510 6802
rect 4510 6750 4562 6802
rect 4562 6750 4564 6802
rect 4508 6748 4564 6750
rect 4732 6748 4788 6804
rect 5292 6636 5348 6692
rect 3612 5794 3668 5796
rect 3612 5742 3614 5794
rect 3614 5742 3666 5794
rect 3666 5742 3668 5794
rect 3612 5740 3668 5742
rect 2828 5628 2884 5684
rect 4008 5514 4064 5516
rect 4112 5514 4168 5516
rect 4008 5462 4024 5514
rect 4024 5462 4064 5514
rect 4112 5462 4148 5514
rect 4148 5462 4168 5514
rect 4008 5460 4064 5462
rect 4112 5460 4168 5462
rect 4216 5460 4272 5516
rect 4320 5514 4376 5516
rect 4424 5514 4480 5516
rect 4528 5514 4584 5516
rect 4320 5462 4324 5514
rect 4324 5462 4376 5514
rect 4424 5462 4448 5514
rect 4448 5462 4480 5514
rect 4528 5462 4572 5514
rect 4572 5462 4584 5514
rect 4320 5460 4376 5462
rect 4424 5460 4480 5462
rect 4528 5460 4584 5462
rect 4632 5514 4688 5516
rect 4736 5514 4792 5516
rect 4840 5514 4896 5516
rect 4632 5462 4644 5514
rect 4644 5462 4688 5514
rect 4736 5462 4768 5514
rect 4768 5462 4792 5514
rect 4840 5462 4892 5514
rect 4892 5462 4896 5514
rect 4632 5460 4688 5462
rect 4736 5460 4792 5462
rect 4840 5460 4896 5462
rect 4944 5460 5000 5516
rect 5048 5514 5104 5516
rect 5152 5514 5208 5516
rect 5048 5462 5068 5514
rect 5068 5462 5104 5514
rect 5152 5462 5192 5514
rect 5192 5462 5208 5514
rect 5048 5460 5104 5462
rect 5152 5460 5208 5462
rect 5292 5068 5348 5124
rect 4732 4956 4788 5012
rect 5516 7308 5572 7364
rect 9212 10108 9268 10164
rect 12908 12850 12964 12852
rect 12908 12798 12910 12850
rect 12910 12798 12962 12850
rect 12962 12798 12964 12850
rect 12908 12796 12964 12798
rect 14008 15706 14064 15708
rect 14112 15706 14168 15708
rect 14008 15654 14024 15706
rect 14024 15654 14064 15706
rect 14112 15654 14148 15706
rect 14148 15654 14168 15706
rect 14008 15652 14064 15654
rect 14112 15652 14168 15654
rect 14216 15652 14272 15708
rect 14320 15706 14376 15708
rect 14424 15706 14480 15708
rect 14528 15706 14584 15708
rect 14320 15654 14324 15706
rect 14324 15654 14376 15706
rect 14424 15654 14448 15706
rect 14448 15654 14480 15706
rect 14528 15654 14572 15706
rect 14572 15654 14584 15706
rect 14320 15652 14376 15654
rect 14424 15652 14480 15654
rect 14528 15652 14584 15654
rect 14632 15706 14688 15708
rect 14736 15706 14792 15708
rect 14840 15706 14896 15708
rect 14632 15654 14644 15706
rect 14644 15654 14688 15706
rect 14736 15654 14768 15706
rect 14768 15654 14792 15706
rect 14840 15654 14892 15706
rect 14892 15654 14896 15706
rect 14632 15652 14688 15654
rect 14736 15652 14792 15654
rect 14840 15652 14896 15654
rect 14944 15652 15000 15708
rect 15048 15706 15104 15708
rect 15152 15706 15208 15708
rect 15048 15654 15068 15706
rect 15068 15654 15104 15706
rect 15152 15654 15192 15706
rect 15192 15654 15208 15706
rect 15048 15652 15104 15654
rect 15152 15652 15208 15654
rect 13916 15426 13972 15428
rect 13916 15374 13918 15426
rect 13918 15374 13970 15426
rect 13970 15374 13972 15426
rect 13916 15372 13972 15374
rect 14364 15202 14420 15204
rect 14364 15150 14366 15202
rect 14366 15150 14418 15202
rect 14418 15150 14420 15202
rect 14364 15148 14420 15150
rect 15372 14476 15428 14532
rect 14008 14138 14064 14140
rect 14112 14138 14168 14140
rect 14008 14086 14024 14138
rect 14024 14086 14064 14138
rect 14112 14086 14148 14138
rect 14148 14086 14168 14138
rect 14008 14084 14064 14086
rect 14112 14084 14168 14086
rect 14216 14084 14272 14140
rect 14320 14138 14376 14140
rect 14424 14138 14480 14140
rect 14528 14138 14584 14140
rect 14320 14086 14324 14138
rect 14324 14086 14376 14138
rect 14424 14086 14448 14138
rect 14448 14086 14480 14138
rect 14528 14086 14572 14138
rect 14572 14086 14584 14138
rect 14320 14084 14376 14086
rect 14424 14084 14480 14086
rect 14528 14084 14584 14086
rect 14632 14138 14688 14140
rect 14736 14138 14792 14140
rect 14840 14138 14896 14140
rect 14632 14086 14644 14138
rect 14644 14086 14688 14138
rect 14736 14086 14768 14138
rect 14768 14086 14792 14138
rect 14840 14086 14892 14138
rect 14892 14086 14896 14138
rect 14632 14084 14688 14086
rect 14736 14084 14792 14086
rect 14840 14084 14896 14086
rect 14944 14084 15000 14140
rect 15048 14138 15104 14140
rect 15152 14138 15208 14140
rect 15048 14086 15068 14138
rect 15068 14086 15104 14138
rect 15152 14086 15192 14138
rect 15192 14086 15208 14138
rect 15048 14084 15104 14086
rect 15152 14084 15208 14086
rect 14252 13746 14308 13748
rect 14252 13694 14254 13746
rect 14254 13694 14306 13746
rect 14306 13694 14308 13746
rect 14252 13692 14308 13694
rect 14812 13746 14868 13748
rect 14812 13694 14814 13746
rect 14814 13694 14866 13746
rect 14866 13694 14868 13746
rect 14812 13692 14868 13694
rect 15372 13692 15428 13748
rect 15708 15372 15764 15428
rect 14924 13132 14980 13188
rect 15260 13468 15316 13524
rect 14364 12850 14420 12852
rect 14364 12798 14366 12850
rect 14366 12798 14418 12850
rect 14418 12798 14420 12850
rect 14364 12796 14420 12798
rect 13580 11788 13636 11844
rect 13244 11564 13300 11620
rect 12012 11170 12068 11172
rect 12012 11118 12014 11170
rect 12014 11118 12066 11170
rect 12066 11118 12068 11170
rect 12012 11116 12068 11118
rect 12460 11004 12516 11060
rect 13244 11004 13300 11060
rect 13244 10834 13300 10836
rect 13244 10782 13246 10834
rect 13246 10782 13298 10834
rect 13298 10782 13300 10834
rect 13244 10780 13300 10782
rect 10892 10108 10948 10164
rect 6076 8316 6132 8372
rect 5852 8034 5908 8036
rect 5852 7982 5854 8034
rect 5854 7982 5906 8034
rect 5906 7982 5908 8034
rect 5852 7980 5908 7982
rect 7308 8316 7364 8372
rect 6636 7980 6692 8036
rect 6076 7698 6132 7700
rect 6076 7646 6078 7698
rect 6078 7646 6130 7698
rect 6130 7646 6132 7698
rect 6076 7644 6132 7646
rect 6748 7420 6804 7476
rect 6636 7362 6692 7364
rect 6636 7310 6638 7362
rect 6638 7310 6690 7362
rect 6690 7310 6692 7362
rect 6636 7308 6692 7310
rect 5628 6860 5684 6916
rect 6860 7308 6916 7364
rect 6300 6748 6356 6804
rect 5740 6466 5796 6468
rect 5740 6414 5742 6466
rect 5742 6414 5794 6466
rect 5794 6414 5796 6466
rect 5740 6412 5796 6414
rect 6748 6636 6804 6692
rect 6412 6578 6468 6580
rect 6412 6526 6414 6578
rect 6414 6526 6466 6578
rect 6466 6526 6468 6578
rect 6412 6524 6468 6526
rect 6748 5852 6804 5908
rect 5964 5740 6020 5796
rect 7980 8370 8036 8372
rect 7980 8318 7982 8370
rect 7982 8318 8034 8370
rect 8034 8318 8036 8370
rect 7980 8316 8036 8318
rect 9212 8316 9268 8372
rect 7532 7474 7588 7476
rect 7532 7422 7534 7474
rect 7534 7422 7586 7474
rect 7586 7422 7588 7474
rect 7532 7420 7588 7422
rect 7980 7420 8036 7476
rect 7644 7308 7700 7364
rect 7756 6690 7812 6692
rect 7756 6638 7758 6690
rect 7758 6638 7810 6690
rect 7810 6638 7812 6690
rect 7756 6636 7812 6638
rect 6076 5122 6132 5124
rect 6076 5070 6078 5122
rect 6078 5070 6130 5122
rect 6130 5070 6132 5122
rect 6076 5068 6132 5070
rect 6636 4956 6692 5012
rect 3836 4284 3892 4340
rect 7532 6412 7588 6468
rect 7980 7250 8036 7252
rect 7980 7198 7982 7250
rect 7982 7198 8034 7250
rect 8034 7198 8036 7250
rect 7980 7196 8036 7198
rect 8092 6914 8148 6916
rect 8092 6862 8094 6914
rect 8094 6862 8146 6914
rect 8146 6862 8148 6914
rect 8092 6860 8148 6862
rect 8428 7196 8484 7252
rect 7980 6578 8036 6580
rect 7980 6526 7982 6578
rect 7982 6526 8034 6578
rect 8034 6526 8036 6578
rect 7980 6524 8036 6526
rect 7532 5740 7588 5796
rect 7308 4956 7364 5012
rect 7532 4956 7588 5012
rect 5964 4284 6020 4340
rect 4008 3946 4064 3948
rect 4112 3946 4168 3948
rect 4008 3894 4024 3946
rect 4024 3894 4064 3946
rect 4112 3894 4148 3946
rect 4148 3894 4168 3946
rect 4008 3892 4064 3894
rect 4112 3892 4168 3894
rect 4216 3892 4272 3948
rect 4320 3946 4376 3948
rect 4424 3946 4480 3948
rect 4528 3946 4584 3948
rect 4320 3894 4324 3946
rect 4324 3894 4376 3946
rect 4424 3894 4448 3946
rect 4448 3894 4480 3946
rect 4528 3894 4572 3946
rect 4572 3894 4584 3946
rect 4320 3892 4376 3894
rect 4424 3892 4480 3894
rect 4528 3892 4584 3894
rect 4632 3946 4688 3948
rect 4736 3946 4792 3948
rect 4840 3946 4896 3948
rect 4632 3894 4644 3946
rect 4644 3894 4688 3946
rect 4736 3894 4768 3946
rect 4768 3894 4792 3946
rect 4840 3894 4892 3946
rect 4892 3894 4896 3946
rect 4632 3892 4688 3894
rect 4736 3892 4792 3894
rect 4840 3892 4896 3894
rect 4944 3892 5000 3948
rect 5048 3946 5104 3948
rect 5152 3946 5208 3948
rect 5048 3894 5068 3946
rect 5068 3894 5104 3946
rect 5152 3894 5192 3946
rect 5192 3894 5208 3946
rect 5048 3892 5104 3894
rect 5152 3892 5208 3894
rect 5964 3666 6020 3668
rect 5964 3614 5966 3666
rect 5966 3614 6018 3666
rect 6018 3614 6020 3666
rect 5964 3612 6020 3614
rect 8316 6524 8372 6580
rect 8540 6860 8596 6916
rect 8764 6860 8820 6916
rect 8540 6076 8596 6132
rect 8428 5906 8484 5908
rect 8428 5854 8430 5906
rect 8430 5854 8482 5906
rect 8482 5854 8484 5906
rect 8428 5852 8484 5854
rect 8316 5628 8372 5684
rect 8540 5740 8596 5796
rect 8764 5628 8820 5684
rect 8876 5852 8932 5908
rect 9100 5852 9156 5908
rect 9212 5628 9268 5684
rect 9772 6860 9828 6916
rect 9324 5068 9380 5124
rect 9996 6690 10052 6692
rect 9996 6638 9998 6690
rect 9998 6638 10050 6690
rect 10050 6638 10052 6690
rect 9996 6636 10052 6638
rect 9996 5906 10052 5908
rect 9996 5854 9998 5906
rect 9998 5854 10050 5906
rect 10050 5854 10052 5906
rect 9996 5852 10052 5854
rect 11116 5740 11172 5796
rect 14588 12684 14644 12740
rect 16380 21196 16436 21252
rect 17052 22204 17108 22260
rect 17276 29596 17332 29652
rect 17388 29426 17444 29428
rect 17388 29374 17390 29426
rect 17390 29374 17442 29426
rect 17442 29374 17444 29426
rect 17388 29372 17444 29374
rect 17612 28476 17668 28532
rect 18732 29426 18788 29428
rect 18732 29374 18734 29426
rect 18734 29374 18786 29426
rect 18786 29374 18788 29426
rect 18732 29372 18788 29374
rect 19740 30210 19796 30212
rect 19740 30158 19742 30210
rect 19742 30158 19794 30210
rect 19794 30158 19796 30210
rect 19740 30156 19796 30158
rect 20860 32508 20916 32564
rect 20076 30156 20132 30212
rect 19292 29650 19348 29652
rect 19292 29598 19294 29650
rect 19294 29598 19346 29650
rect 19346 29598 19348 29650
rect 19292 29596 19348 29598
rect 19740 29596 19796 29652
rect 18284 28642 18340 28644
rect 18284 28590 18286 28642
rect 18286 28590 18338 28642
rect 18338 28590 18340 28642
rect 18284 28588 18340 28590
rect 18396 28082 18452 28084
rect 18396 28030 18398 28082
rect 18398 28030 18450 28082
rect 18450 28030 18452 28082
rect 18396 28028 18452 28030
rect 17836 27858 17892 27860
rect 17836 27806 17838 27858
rect 17838 27806 17890 27858
rect 17890 27806 17892 27858
rect 17836 27804 17892 27806
rect 19292 27804 19348 27860
rect 21196 33628 21252 33684
rect 21308 33516 21364 33572
rect 21308 32562 21364 32564
rect 21308 32510 21310 32562
rect 21310 32510 21362 32562
rect 21362 32510 21364 32562
rect 21308 32508 21364 32510
rect 21756 39676 21812 39732
rect 22092 41132 22148 41188
rect 21980 40572 22036 40628
rect 22540 41916 22596 41972
rect 22652 41298 22708 41300
rect 22652 41246 22654 41298
rect 22654 41246 22706 41298
rect 22706 41246 22708 41298
rect 22652 41244 22708 41246
rect 22204 40626 22260 40628
rect 22204 40574 22206 40626
rect 22206 40574 22258 40626
rect 22258 40574 22260 40626
rect 22204 40572 22260 40574
rect 23324 42812 23380 42868
rect 23100 40572 23156 40628
rect 23660 44098 23716 44100
rect 23660 44046 23662 44098
rect 23662 44046 23714 44098
rect 23714 44046 23716 44098
rect 23660 44044 23716 44046
rect 23660 42588 23716 42644
rect 23660 40684 23716 40740
rect 23660 40236 23716 40292
rect 23548 39788 23604 39844
rect 22092 37996 22148 38052
rect 21868 37436 21924 37492
rect 22204 37660 22260 37716
rect 21532 37324 21588 37380
rect 22428 37378 22484 37380
rect 22428 37326 22430 37378
rect 22430 37326 22482 37378
rect 22482 37326 22484 37378
rect 22428 37324 22484 37326
rect 23100 36204 23156 36260
rect 22876 35922 22932 35924
rect 22876 35870 22878 35922
rect 22878 35870 22930 35922
rect 22930 35870 22932 35922
rect 22876 35868 22932 35870
rect 21532 35644 21588 35700
rect 23100 34914 23156 34916
rect 23100 34862 23102 34914
rect 23102 34862 23154 34914
rect 23154 34862 23156 34914
rect 23100 34860 23156 34862
rect 21532 31836 21588 31892
rect 21644 34748 21700 34804
rect 21420 31612 21476 31668
rect 21420 30210 21476 30212
rect 21420 30158 21422 30210
rect 21422 30158 21474 30210
rect 21474 30158 21476 30210
rect 21420 30156 21476 30158
rect 19852 29484 19908 29540
rect 21084 29372 21140 29428
rect 23436 36316 23492 36372
rect 23548 35868 23604 35924
rect 23660 37324 23716 37380
rect 25340 47180 25396 47236
rect 24008 46282 24064 46284
rect 24112 46282 24168 46284
rect 24008 46230 24024 46282
rect 24024 46230 24064 46282
rect 24112 46230 24148 46282
rect 24148 46230 24168 46282
rect 24008 46228 24064 46230
rect 24112 46228 24168 46230
rect 24216 46228 24272 46284
rect 24320 46282 24376 46284
rect 24424 46282 24480 46284
rect 24528 46282 24584 46284
rect 24320 46230 24324 46282
rect 24324 46230 24376 46282
rect 24424 46230 24448 46282
rect 24448 46230 24480 46282
rect 24528 46230 24572 46282
rect 24572 46230 24584 46282
rect 24320 46228 24376 46230
rect 24424 46228 24480 46230
rect 24528 46228 24584 46230
rect 24632 46282 24688 46284
rect 24736 46282 24792 46284
rect 24840 46282 24896 46284
rect 24632 46230 24644 46282
rect 24644 46230 24688 46282
rect 24736 46230 24768 46282
rect 24768 46230 24792 46282
rect 24840 46230 24892 46282
rect 24892 46230 24896 46282
rect 24632 46228 24688 46230
rect 24736 46228 24792 46230
rect 24840 46228 24896 46230
rect 24944 46228 25000 46284
rect 25048 46282 25104 46284
rect 25152 46282 25208 46284
rect 25048 46230 25068 46282
rect 25068 46230 25104 46282
rect 25152 46230 25192 46282
rect 25192 46230 25208 46282
rect 25048 46228 25104 46230
rect 25152 46228 25208 46230
rect 28140 58434 28196 58436
rect 28140 58382 28142 58434
rect 28142 58382 28194 58434
rect 28194 58382 28196 58434
rect 28140 58380 28196 58382
rect 28476 58380 28532 58436
rect 28140 57874 28196 57876
rect 28140 57822 28142 57874
rect 28142 57822 28194 57874
rect 28194 57822 28196 57874
rect 28140 57820 28196 57822
rect 28588 57820 28644 57876
rect 28700 60396 28756 60452
rect 29372 67730 29428 67732
rect 29372 67678 29374 67730
rect 29374 67678 29426 67730
rect 29426 67678 29428 67730
rect 29372 67676 29428 67678
rect 30716 67676 30772 67732
rect 29372 66220 29428 66276
rect 29372 65660 29428 65716
rect 29260 63922 29316 63924
rect 29260 63870 29262 63922
rect 29262 63870 29314 63922
rect 29314 63870 29316 63922
rect 29260 63868 29316 63870
rect 29148 62354 29204 62356
rect 29148 62302 29150 62354
rect 29150 62302 29202 62354
rect 29202 62302 29204 62354
rect 29148 62300 29204 62302
rect 29596 62578 29652 62580
rect 29596 62526 29598 62578
rect 29598 62526 29650 62578
rect 29650 62526 29652 62578
rect 29596 62524 29652 62526
rect 29932 63810 29988 63812
rect 29932 63758 29934 63810
rect 29934 63758 29986 63810
rect 29986 63758 29988 63810
rect 29932 63756 29988 63758
rect 31164 66780 31220 66836
rect 31276 67116 31332 67172
rect 30828 65490 30884 65492
rect 30828 65438 30830 65490
rect 30830 65438 30882 65490
rect 30882 65438 30884 65490
rect 30828 65436 30884 65438
rect 31388 66892 31444 66948
rect 33404 69804 33460 69860
rect 33852 70924 33908 70980
rect 33516 69580 33572 69636
rect 33740 70364 33796 70420
rect 34008 70586 34064 70588
rect 34112 70586 34168 70588
rect 34008 70534 34024 70586
rect 34024 70534 34064 70586
rect 34112 70534 34148 70586
rect 34148 70534 34168 70586
rect 34008 70532 34064 70534
rect 34112 70532 34168 70534
rect 34216 70532 34272 70588
rect 34320 70586 34376 70588
rect 34424 70586 34480 70588
rect 34528 70586 34584 70588
rect 34320 70534 34324 70586
rect 34324 70534 34376 70586
rect 34424 70534 34448 70586
rect 34448 70534 34480 70586
rect 34528 70534 34572 70586
rect 34572 70534 34584 70586
rect 34320 70532 34376 70534
rect 34424 70532 34480 70534
rect 34528 70532 34584 70534
rect 34632 70586 34688 70588
rect 34736 70586 34792 70588
rect 34840 70586 34896 70588
rect 34632 70534 34644 70586
rect 34644 70534 34688 70586
rect 34736 70534 34768 70586
rect 34768 70534 34792 70586
rect 34840 70534 34892 70586
rect 34892 70534 34896 70586
rect 34632 70532 34688 70534
rect 34736 70532 34792 70534
rect 34840 70532 34896 70534
rect 34944 70532 35000 70588
rect 35048 70586 35104 70588
rect 35152 70586 35208 70588
rect 35048 70534 35068 70586
rect 35068 70534 35104 70586
rect 35152 70534 35192 70586
rect 35192 70534 35208 70586
rect 35048 70532 35104 70534
rect 35152 70532 35208 70534
rect 35756 70754 35812 70756
rect 35756 70702 35758 70754
rect 35758 70702 35810 70754
rect 35810 70702 35812 70754
rect 35756 70700 35812 70702
rect 35308 70476 35364 70532
rect 35644 70476 35700 70532
rect 32060 67564 32116 67620
rect 30268 64540 30324 64596
rect 30492 63138 30548 63140
rect 30492 63086 30494 63138
rect 30494 63086 30546 63138
rect 30546 63086 30548 63138
rect 30492 63084 30548 63086
rect 30044 62354 30100 62356
rect 30044 62302 30046 62354
rect 30046 62302 30098 62354
rect 30098 62302 30100 62354
rect 30044 62300 30100 62302
rect 29596 61292 29652 61348
rect 29372 60396 29428 60452
rect 29596 60508 29652 60564
rect 31052 63138 31108 63140
rect 31052 63086 31054 63138
rect 31054 63086 31106 63138
rect 31106 63086 31108 63138
rect 31052 63084 31108 63086
rect 30716 62748 30772 62804
rect 31052 62860 31108 62916
rect 30492 62188 30548 62244
rect 31612 66780 31668 66836
rect 32172 67116 32228 67172
rect 32956 67618 33012 67620
rect 32956 67566 32958 67618
rect 32958 67566 33010 67618
rect 33010 67566 33012 67618
rect 32956 67564 33012 67566
rect 32396 66834 32452 66836
rect 32396 66782 32398 66834
rect 32398 66782 32450 66834
rect 32450 66782 32452 66834
rect 32396 66780 32452 66782
rect 31836 66220 31892 66276
rect 31948 66162 32004 66164
rect 31948 66110 31950 66162
rect 31950 66110 32002 66162
rect 32002 66110 32004 66162
rect 31948 66108 32004 66110
rect 31836 65996 31892 66052
rect 33292 67170 33348 67172
rect 33292 67118 33294 67170
rect 33294 67118 33346 67170
rect 33346 67118 33348 67170
rect 33292 67116 33348 67118
rect 34412 70364 34468 70420
rect 35196 70028 35252 70084
rect 34972 69804 35028 69860
rect 34636 69634 34692 69636
rect 34636 69582 34638 69634
rect 34638 69582 34690 69634
rect 34690 69582 34692 69634
rect 34636 69580 34692 69582
rect 35532 69804 35588 69860
rect 33964 69132 34020 69188
rect 35532 69244 35588 69300
rect 34008 69018 34064 69020
rect 34112 69018 34168 69020
rect 34008 68966 34024 69018
rect 34024 68966 34064 69018
rect 34112 68966 34148 69018
rect 34148 68966 34168 69018
rect 34008 68964 34064 68966
rect 34112 68964 34168 68966
rect 34216 68964 34272 69020
rect 34320 69018 34376 69020
rect 34424 69018 34480 69020
rect 34528 69018 34584 69020
rect 34320 68966 34324 69018
rect 34324 68966 34376 69018
rect 34424 68966 34448 69018
rect 34448 68966 34480 69018
rect 34528 68966 34572 69018
rect 34572 68966 34584 69018
rect 34320 68964 34376 68966
rect 34424 68964 34480 68966
rect 34528 68964 34584 68966
rect 34632 69018 34688 69020
rect 34736 69018 34792 69020
rect 34840 69018 34896 69020
rect 34632 68966 34644 69018
rect 34644 68966 34688 69018
rect 34736 68966 34768 69018
rect 34768 68966 34792 69018
rect 34840 68966 34892 69018
rect 34892 68966 34896 69018
rect 34632 68964 34688 68966
rect 34736 68964 34792 68966
rect 34840 68964 34896 68966
rect 34944 68964 35000 69020
rect 35048 69018 35104 69020
rect 35152 69018 35208 69020
rect 35048 68966 35068 69018
rect 35068 68966 35104 69018
rect 35152 68966 35192 69018
rect 35192 68966 35208 69018
rect 35048 68964 35104 68966
rect 35152 68964 35208 68966
rect 34972 68796 35028 68852
rect 35756 69244 35812 69300
rect 36092 69916 36148 69972
rect 35980 69298 36036 69300
rect 35980 69246 35982 69298
rect 35982 69246 36034 69298
rect 36034 69246 36036 69298
rect 35980 69244 36036 69246
rect 34008 67450 34064 67452
rect 34112 67450 34168 67452
rect 34008 67398 34024 67450
rect 34024 67398 34064 67450
rect 34112 67398 34148 67450
rect 34148 67398 34168 67450
rect 34008 67396 34064 67398
rect 34112 67396 34168 67398
rect 34216 67396 34272 67452
rect 34320 67450 34376 67452
rect 34424 67450 34480 67452
rect 34528 67450 34584 67452
rect 34320 67398 34324 67450
rect 34324 67398 34376 67450
rect 34424 67398 34448 67450
rect 34448 67398 34480 67450
rect 34528 67398 34572 67450
rect 34572 67398 34584 67450
rect 34320 67396 34376 67398
rect 34424 67396 34480 67398
rect 34528 67396 34584 67398
rect 34632 67450 34688 67452
rect 34736 67450 34792 67452
rect 34840 67450 34896 67452
rect 34632 67398 34644 67450
rect 34644 67398 34688 67450
rect 34736 67398 34768 67450
rect 34768 67398 34792 67450
rect 34840 67398 34892 67450
rect 34892 67398 34896 67450
rect 34632 67396 34688 67398
rect 34736 67396 34792 67398
rect 34840 67396 34896 67398
rect 34944 67396 35000 67452
rect 35048 67450 35104 67452
rect 35152 67450 35208 67452
rect 35048 67398 35068 67450
rect 35068 67398 35104 67450
rect 35152 67398 35192 67450
rect 35192 67398 35208 67450
rect 35048 67396 35104 67398
rect 35152 67396 35208 67398
rect 34524 67228 34580 67284
rect 33180 66892 33236 66948
rect 32732 66050 32788 66052
rect 32732 65998 32734 66050
rect 32734 65998 32786 66050
rect 32786 65998 32788 66050
rect 32732 65996 32788 65998
rect 33740 66108 33796 66164
rect 35308 67228 35364 67284
rect 36652 70306 36708 70308
rect 36652 70254 36654 70306
rect 36654 70254 36706 70306
rect 36706 70254 36708 70306
rect 36652 70252 36708 70254
rect 36316 70140 36372 70196
rect 37436 69970 37492 69972
rect 37436 69918 37438 69970
rect 37438 69918 37490 69970
rect 37490 69918 37492 69970
rect 37436 69916 37492 69918
rect 37772 70082 37828 70084
rect 37772 70030 37774 70082
rect 37774 70030 37826 70082
rect 37826 70030 37828 70082
rect 37772 70028 37828 70030
rect 38108 70194 38164 70196
rect 38108 70142 38110 70194
rect 38110 70142 38162 70194
rect 38162 70142 38164 70194
rect 38108 70140 38164 70142
rect 37884 69916 37940 69972
rect 37548 69244 37604 69300
rect 36204 68796 36260 68852
rect 35868 67842 35924 67844
rect 35868 67790 35870 67842
rect 35870 67790 35922 67842
rect 35922 67790 35924 67842
rect 35868 67788 35924 67790
rect 37100 67842 37156 67844
rect 37100 67790 37102 67842
rect 37102 67790 37154 67842
rect 37154 67790 37156 67842
rect 37100 67788 37156 67790
rect 35644 66332 35700 66388
rect 34008 65882 34064 65884
rect 34112 65882 34168 65884
rect 34008 65830 34024 65882
rect 34024 65830 34064 65882
rect 34112 65830 34148 65882
rect 34148 65830 34168 65882
rect 34008 65828 34064 65830
rect 34112 65828 34168 65830
rect 34216 65828 34272 65884
rect 34320 65882 34376 65884
rect 34424 65882 34480 65884
rect 34528 65882 34584 65884
rect 34320 65830 34324 65882
rect 34324 65830 34376 65882
rect 34424 65830 34448 65882
rect 34448 65830 34480 65882
rect 34528 65830 34572 65882
rect 34572 65830 34584 65882
rect 34320 65828 34376 65830
rect 34424 65828 34480 65830
rect 34528 65828 34584 65830
rect 34632 65882 34688 65884
rect 34736 65882 34792 65884
rect 34840 65882 34896 65884
rect 34632 65830 34644 65882
rect 34644 65830 34688 65882
rect 34736 65830 34768 65882
rect 34768 65830 34792 65882
rect 34840 65830 34892 65882
rect 34892 65830 34896 65882
rect 34632 65828 34688 65830
rect 34736 65828 34792 65830
rect 34840 65828 34896 65830
rect 34944 65828 35000 65884
rect 35048 65882 35104 65884
rect 35152 65882 35208 65884
rect 35048 65830 35068 65882
rect 35068 65830 35104 65882
rect 35152 65830 35192 65882
rect 35192 65830 35208 65882
rect 35048 65828 35104 65830
rect 35152 65828 35208 65830
rect 34636 64876 34692 64932
rect 36988 66386 37044 66388
rect 36988 66334 36990 66386
rect 36990 66334 37042 66386
rect 37042 66334 37044 66386
rect 36988 66332 37044 66334
rect 36876 66108 36932 66164
rect 36092 64988 36148 65044
rect 35532 64930 35588 64932
rect 35532 64878 35534 64930
rect 35534 64878 35586 64930
rect 35586 64878 35588 64930
rect 35532 64876 35588 64878
rect 35868 64930 35924 64932
rect 35868 64878 35870 64930
rect 35870 64878 35922 64930
rect 35922 64878 35924 64930
rect 35868 64876 35924 64878
rect 34008 64314 34064 64316
rect 34112 64314 34168 64316
rect 34008 64262 34024 64314
rect 34024 64262 34064 64314
rect 34112 64262 34148 64314
rect 34148 64262 34168 64314
rect 34008 64260 34064 64262
rect 34112 64260 34168 64262
rect 34216 64260 34272 64316
rect 34320 64314 34376 64316
rect 34424 64314 34480 64316
rect 34528 64314 34584 64316
rect 34320 64262 34324 64314
rect 34324 64262 34376 64314
rect 34424 64262 34448 64314
rect 34448 64262 34480 64314
rect 34528 64262 34572 64314
rect 34572 64262 34584 64314
rect 34320 64260 34376 64262
rect 34424 64260 34480 64262
rect 34528 64260 34584 64262
rect 34632 64314 34688 64316
rect 34736 64314 34792 64316
rect 34840 64314 34896 64316
rect 34632 64262 34644 64314
rect 34644 64262 34688 64314
rect 34736 64262 34768 64314
rect 34768 64262 34792 64314
rect 34840 64262 34892 64314
rect 34892 64262 34896 64314
rect 34632 64260 34688 64262
rect 34736 64260 34792 64262
rect 34840 64260 34896 64262
rect 34944 64260 35000 64316
rect 35048 64314 35104 64316
rect 35152 64314 35208 64316
rect 35048 64262 35068 64314
rect 35068 64262 35104 64314
rect 35152 64262 35192 64314
rect 35192 64262 35208 64314
rect 35048 64260 35104 64262
rect 35152 64260 35208 64262
rect 31836 63756 31892 63812
rect 31500 62860 31556 62916
rect 31276 62748 31332 62804
rect 30156 61068 30212 61124
rect 29932 60956 29988 61012
rect 30044 60060 30100 60116
rect 30044 59890 30100 59892
rect 30044 59838 30046 59890
rect 30046 59838 30098 59890
rect 30098 59838 30100 59890
rect 30044 59836 30100 59838
rect 28812 59388 28868 59444
rect 29932 59388 29988 59444
rect 29708 58828 29764 58884
rect 29932 58434 29988 58436
rect 29932 58382 29934 58434
rect 29934 58382 29986 58434
rect 29986 58382 29988 58434
rect 29932 58380 29988 58382
rect 27692 56140 27748 56196
rect 28140 56140 28196 56196
rect 27356 54514 27412 54516
rect 27356 54462 27358 54514
rect 27358 54462 27410 54514
rect 27410 54462 27412 54514
rect 27356 54460 27412 54462
rect 27356 53788 27412 53844
rect 26908 51436 26964 51492
rect 27692 53954 27748 53956
rect 27692 53902 27694 53954
rect 27694 53902 27746 53954
rect 27746 53902 27748 53954
rect 27692 53900 27748 53902
rect 27580 52050 27636 52052
rect 27580 51998 27582 52050
rect 27582 51998 27634 52050
rect 27634 51998 27636 52050
rect 27580 51996 27636 51998
rect 27580 51436 27636 51492
rect 28476 53618 28532 53620
rect 28476 53566 28478 53618
rect 28478 53566 28530 53618
rect 28530 53566 28532 53618
rect 28476 53564 28532 53566
rect 29372 53506 29428 53508
rect 29372 53454 29374 53506
rect 29374 53454 29426 53506
rect 29426 53454 29428 53506
rect 29372 53452 29428 53454
rect 27132 50316 27188 50372
rect 26460 49922 26516 49924
rect 26460 49870 26462 49922
rect 26462 49870 26514 49922
rect 26514 49870 26516 49922
rect 26460 49868 26516 49870
rect 26236 49250 26292 49252
rect 26236 49198 26238 49250
rect 26238 49198 26290 49250
rect 26290 49198 26292 49250
rect 26236 49196 26292 49198
rect 25676 48972 25732 49028
rect 26684 48972 26740 49028
rect 26236 48860 26292 48916
rect 25788 47516 25844 47572
rect 24780 45890 24836 45892
rect 24780 45838 24782 45890
rect 24782 45838 24834 45890
rect 24834 45838 24836 45890
rect 24780 45836 24836 45838
rect 24108 45724 24164 45780
rect 24332 45666 24388 45668
rect 24332 45614 24334 45666
rect 24334 45614 24386 45666
rect 24386 45614 24388 45666
rect 24332 45612 24388 45614
rect 24332 45330 24388 45332
rect 24332 45278 24334 45330
rect 24334 45278 24386 45330
rect 24386 45278 24388 45330
rect 24332 45276 24388 45278
rect 25116 44828 25172 44884
rect 24008 44714 24064 44716
rect 24112 44714 24168 44716
rect 24008 44662 24024 44714
rect 24024 44662 24064 44714
rect 24112 44662 24148 44714
rect 24148 44662 24168 44714
rect 24008 44660 24064 44662
rect 24112 44660 24168 44662
rect 24216 44660 24272 44716
rect 24320 44714 24376 44716
rect 24424 44714 24480 44716
rect 24528 44714 24584 44716
rect 24320 44662 24324 44714
rect 24324 44662 24376 44714
rect 24424 44662 24448 44714
rect 24448 44662 24480 44714
rect 24528 44662 24572 44714
rect 24572 44662 24584 44714
rect 24320 44660 24376 44662
rect 24424 44660 24480 44662
rect 24528 44660 24584 44662
rect 24632 44714 24688 44716
rect 24736 44714 24792 44716
rect 24840 44714 24896 44716
rect 24632 44662 24644 44714
rect 24644 44662 24688 44714
rect 24736 44662 24768 44714
rect 24768 44662 24792 44714
rect 24840 44662 24892 44714
rect 24892 44662 24896 44714
rect 24632 44660 24688 44662
rect 24736 44660 24792 44662
rect 24840 44660 24896 44662
rect 24944 44660 25000 44716
rect 25048 44714 25104 44716
rect 25152 44714 25208 44716
rect 25048 44662 25068 44714
rect 25068 44662 25104 44714
rect 25152 44662 25192 44714
rect 25192 44662 25208 44714
rect 25048 44660 25104 44662
rect 25152 44660 25208 44662
rect 25788 45948 25844 46004
rect 26012 46562 26068 46564
rect 26012 46510 26014 46562
rect 26014 46510 26066 46562
rect 26066 46510 26068 46562
rect 26012 46508 26068 46510
rect 26012 45724 26068 45780
rect 27020 49026 27076 49028
rect 27020 48974 27022 49026
rect 27022 48974 27074 49026
rect 27074 48974 27076 49026
rect 27020 48972 27076 48974
rect 26908 48748 26964 48804
rect 27020 48300 27076 48356
rect 26460 46898 26516 46900
rect 26460 46846 26462 46898
rect 26462 46846 26514 46898
rect 26514 46846 26516 46898
rect 26460 46844 26516 46846
rect 27356 48242 27412 48244
rect 27356 48190 27358 48242
rect 27358 48190 27410 48242
rect 27410 48190 27412 48242
rect 27356 48188 27412 48190
rect 27132 47068 27188 47124
rect 26572 46732 26628 46788
rect 26572 46508 26628 46564
rect 26236 45836 26292 45892
rect 25788 45106 25844 45108
rect 25788 45054 25790 45106
rect 25790 45054 25842 45106
rect 25842 45054 25844 45106
rect 25788 45052 25844 45054
rect 25452 44994 25508 44996
rect 25452 44942 25454 44994
rect 25454 44942 25506 44994
rect 25506 44942 25508 44994
rect 25452 44940 25508 44942
rect 23884 44380 23940 44436
rect 24008 43146 24064 43148
rect 24112 43146 24168 43148
rect 24008 43094 24024 43146
rect 24024 43094 24064 43146
rect 24112 43094 24148 43146
rect 24148 43094 24168 43146
rect 24008 43092 24064 43094
rect 24112 43092 24168 43094
rect 24216 43092 24272 43148
rect 24320 43146 24376 43148
rect 24424 43146 24480 43148
rect 24528 43146 24584 43148
rect 24320 43094 24324 43146
rect 24324 43094 24376 43146
rect 24424 43094 24448 43146
rect 24448 43094 24480 43146
rect 24528 43094 24572 43146
rect 24572 43094 24584 43146
rect 24320 43092 24376 43094
rect 24424 43092 24480 43094
rect 24528 43092 24584 43094
rect 24632 43146 24688 43148
rect 24736 43146 24792 43148
rect 24840 43146 24896 43148
rect 24632 43094 24644 43146
rect 24644 43094 24688 43146
rect 24736 43094 24768 43146
rect 24768 43094 24792 43146
rect 24840 43094 24892 43146
rect 24892 43094 24896 43146
rect 24632 43092 24688 43094
rect 24736 43092 24792 43094
rect 24840 43092 24896 43094
rect 24944 43092 25000 43148
rect 25048 43146 25104 43148
rect 25152 43146 25208 43148
rect 25048 43094 25068 43146
rect 25068 43094 25104 43146
rect 25152 43094 25192 43146
rect 25192 43094 25208 43146
rect 25048 43092 25104 43094
rect 25152 43092 25208 43094
rect 23884 42812 23940 42868
rect 25004 42866 25060 42868
rect 25004 42814 25006 42866
rect 25006 42814 25058 42866
rect 25058 42814 25060 42866
rect 25004 42812 25060 42814
rect 24556 42642 24612 42644
rect 24556 42590 24558 42642
rect 24558 42590 24610 42642
rect 24610 42590 24612 42642
rect 24556 42588 24612 42590
rect 24444 41970 24500 41972
rect 24444 41918 24446 41970
rect 24446 41918 24498 41970
rect 24498 41918 24500 41970
rect 24444 41916 24500 41918
rect 25340 41970 25396 41972
rect 25340 41918 25342 41970
rect 25342 41918 25394 41970
rect 25394 41918 25396 41970
rect 25340 41916 25396 41918
rect 25452 41746 25508 41748
rect 25452 41694 25454 41746
rect 25454 41694 25506 41746
rect 25506 41694 25508 41746
rect 25452 41692 25508 41694
rect 24008 41578 24064 41580
rect 24112 41578 24168 41580
rect 24008 41526 24024 41578
rect 24024 41526 24064 41578
rect 24112 41526 24148 41578
rect 24148 41526 24168 41578
rect 24008 41524 24064 41526
rect 24112 41524 24168 41526
rect 24216 41524 24272 41580
rect 24320 41578 24376 41580
rect 24424 41578 24480 41580
rect 24528 41578 24584 41580
rect 24320 41526 24324 41578
rect 24324 41526 24376 41578
rect 24424 41526 24448 41578
rect 24448 41526 24480 41578
rect 24528 41526 24572 41578
rect 24572 41526 24584 41578
rect 24320 41524 24376 41526
rect 24424 41524 24480 41526
rect 24528 41524 24584 41526
rect 24632 41578 24688 41580
rect 24736 41578 24792 41580
rect 24840 41578 24896 41580
rect 24632 41526 24644 41578
rect 24644 41526 24688 41578
rect 24736 41526 24768 41578
rect 24768 41526 24792 41578
rect 24840 41526 24892 41578
rect 24892 41526 24896 41578
rect 24632 41524 24688 41526
rect 24736 41524 24792 41526
rect 24840 41524 24896 41526
rect 24944 41524 25000 41580
rect 25048 41578 25104 41580
rect 25152 41578 25208 41580
rect 25048 41526 25068 41578
rect 25068 41526 25104 41578
rect 25152 41526 25192 41578
rect 25192 41526 25208 41578
rect 25048 41524 25104 41526
rect 25152 41524 25208 41526
rect 25452 41356 25508 41412
rect 24668 41244 24724 41300
rect 24780 41186 24836 41188
rect 24780 41134 24782 41186
rect 24782 41134 24834 41186
rect 24834 41134 24836 41186
rect 24780 41132 24836 41134
rect 25452 41186 25508 41188
rect 25452 41134 25454 41186
rect 25454 41134 25506 41186
rect 25506 41134 25508 41186
rect 25452 41132 25508 41134
rect 24556 41074 24612 41076
rect 24556 41022 24558 41074
rect 24558 41022 24610 41074
rect 24610 41022 24612 41074
rect 24556 41020 24612 41022
rect 25228 41074 25284 41076
rect 25228 41022 25230 41074
rect 25230 41022 25282 41074
rect 25282 41022 25284 41074
rect 25228 41020 25284 41022
rect 23884 40962 23940 40964
rect 23884 40910 23886 40962
rect 23886 40910 23938 40962
rect 23938 40910 23940 40962
rect 23884 40908 23940 40910
rect 24444 40962 24500 40964
rect 24444 40910 24446 40962
rect 24446 40910 24498 40962
rect 24498 40910 24500 40962
rect 24444 40908 24500 40910
rect 25452 40572 25508 40628
rect 24332 40236 24388 40292
rect 25452 40236 25508 40292
rect 24008 40010 24064 40012
rect 24112 40010 24168 40012
rect 24008 39958 24024 40010
rect 24024 39958 24064 40010
rect 24112 39958 24148 40010
rect 24148 39958 24168 40010
rect 24008 39956 24064 39958
rect 24112 39956 24168 39958
rect 24216 39956 24272 40012
rect 24320 40010 24376 40012
rect 24424 40010 24480 40012
rect 24528 40010 24584 40012
rect 24320 39958 24324 40010
rect 24324 39958 24376 40010
rect 24424 39958 24448 40010
rect 24448 39958 24480 40010
rect 24528 39958 24572 40010
rect 24572 39958 24584 40010
rect 24320 39956 24376 39958
rect 24424 39956 24480 39958
rect 24528 39956 24584 39958
rect 24632 40010 24688 40012
rect 24736 40010 24792 40012
rect 24840 40010 24896 40012
rect 24632 39958 24644 40010
rect 24644 39958 24688 40010
rect 24736 39958 24768 40010
rect 24768 39958 24792 40010
rect 24840 39958 24892 40010
rect 24892 39958 24896 40010
rect 24632 39956 24688 39958
rect 24736 39956 24792 39958
rect 24840 39956 24896 39958
rect 24944 39956 25000 40012
rect 25048 40010 25104 40012
rect 25152 40010 25208 40012
rect 25048 39958 25068 40010
rect 25068 39958 25104 40010
rect 25152 39958 25192 40010
rect 25192 39958 25208 40010
rect 25048 39956 25104 39958
rect 25152 39956 25208 39958
rect 24108 39788 24164 39844
rect 24556 39564 24612 39620
rect 24008 38442 24064 38444
rect 24112 38442 24168 38444
rect 24008 38390 24024 38442
rect 24024 38390 24064 38442
rect 24112 38390 24148 38442
rect 24148 38390 24168 38442
rect 24008 38388 24064 38390
rect 24112 38388 24168 38390
rect 24216 38388 24272 38444
rect 24320 38442 24376 38444
rect 24424 38442 24480 38444
rect 24528 38442 24584 38444
rect 24320 38390 24324 38442
rect 24324 38390 24376 38442
rect 24424 38390 24448 38442
rect 24448 38390 24480 38442
rect 24528 38390 24572 38442
rect 24572 38390 24584 38442
rect 24320 38388 24376 38390
rect 24424 38388 24480 38390
rect 24528 38388 24584 38390
rect 24632 38442 24688 38444
rect 24736 38442 24792 38444
rect 24840 38442 24896 38444
rect 24632 38390 24644 38442
rect 24644 38390 24688 38442
rect 24736 38390 24768 38442
rect 24768 38390 24792 38442
rect 24840 38390 24892 38442
rect 24892 38390 24896 38442
rect 24632 38388 24688 38390
rect 24736 38388 24792 38390
rect 24840 38388 24896 38390
rect 24944 38388 25000 38444
rect 25048 38442 25104 38444
rect 25152 38442 25208 38444
rect 25048 38390 25068 38442
rect 25068 38390 25104 38442
rect 25152 38390 25192 38442
rect 25192 38390 25208 38442
rect 25048 38388 25104 38390
rect 25152 38388 25208 38390
rect 24892 38162 24948 38164
rect 24892 38110 24894 38162
rect 24894 38110 24946 38162
rect 24946 38110 24948 38162
rect 24892 38108 24948 38110
rect 26348 45106 26404 45108
rect 26348 45054 26350 45106
rect 26350 45054 26402 45106
rect 26402 45054 26404 45106
rect 26348 45052 26404 45054
rect 26124 44940 26180 44996
rect 28476 53116 28532 53172
rect 29372 51324 29428 51380
rect 28028 50316 28084 50372
rect 27692 49868 27748 49924
rect 28588 48802 28644 48804
rect 28588 48750 28590 48802
rect 28590 48750 28642 48802
rect 28642 48750 28644 48802
rect 28588 48748 28644 48750
rect 30268 60396 30324 60452
rect 30156 59276 30212 59332
rect 30604 61404 30660 61460
rect 30604 60844 30660 60900
rect 34860 63868 34916 63924
rect 34748 63250 34804 63252
rect 34748 63198 34750 63250
rect 34750 63198 34802 63250
rect 34802 63198 34804 63250
rect 34748 63196 34804 63198
rect 35084 63026 35140 63028
rect 35084 62974 35086 63026
rect 35086 62974 35138 63026
rect 35138 62974 35140 63026
rect 35084 62972 35140 62974
rect 34008 62746 34064 62748
rect 34112 62746 34168 62748
rect 34008 62694 34024 62746
rect 34024 62694 34064 62746
rect 34112 62694 34148 62746
rect 34148 62694 34168 62746
rect 34008 62692 34064 62694
rect 34112 62692 34168 62694
rect 34216 62692 34272 62748
rect 34320 62746 34376 62748
rect 34424 62746 34480 62748
rect 34528 62746 34584 62748
rect 34320 62694 34324 62746
rect 34324 62694 34376 62746
rect 34424 62694 34448 62746
rect 34448 62694 34480 62746
rect 34528 62694 34572 62746
rect 34572 62694 34584 62746
rect 34320 62692 34376 62694
rect 34424 62692 34480 62694
rect 34528 62692 34584 62694
rect 34632 62746 34688 62748
rect 34736 62746 34792 62748
rect 34840 62746 34896 62748
rect 34632 62694 34644 62746
rect 34644 62694 34688 62746
rect 34736 62694 34768 62746
rect 34768 62694 34792 62746
rect 34840 62694 34892 62746
rect 34892 62694 34896 62746
rect 34632 62692 34688 62694
rect 34736 62692 34792 62694
rect 34840 62692 34896 62694
rect 34944 62692 35000 62748
rect 35048 62746 35104 62748
rect 35152 62746 35208 62748
rect 35048 62694 35068 62746
rect 35068 62694 35104 62746
rect 35152 62694 35192 62746
rect 35192 62694 35208 62746
rect 35048 62692 35104 62694
rect 35152 62692 35208 62694
rect 33628 62524 33684 62580
rect 33404 62354 33460 62356
rect 33404 62302 33406 62354
rect 33406 62302 33458 62354
rect 33458 62302 33460 62354
rect 33404 62300 33460 62302
rect 30828 61068 30884 61124
rect 30716 59836 30772 59892
rect 30492 59442 30548 59444
rect 30492 59390 30494 59442
rect 30494 59390 30546 59442
rect 30546 59390 30548 59442
rect 30492 59388 30548 59390
rect 30380 58828 30436 58884
rect 31052 60620 31108 60676
rect 30380 58156 30436 58212
rect 30940 60002 30996 60004
rect 30940 59950 30942 60002
rect 30942 59950 30994 60002
rect 30994 59950 30996 60002
rect 30940 59948 30996 59950
rect 31052 59724 31108 59780
rect 31276 59276 31332 59332
rect 30940 58210 30996 58212
rect 30940 58158 30942 58210
rect 30942 58158 30994 58210
rect 30994 58158 30996 58210
rect 30940 58156 30996 58158
rect 31052 58828 31108 58884
rect 30828 57820 30884 57876
rect 31724 60844 31780 60900
rect 31500 60786 31556 60788
rect 31500 60734 31502 60786
rect 31502 60734 31554 60786
rect 31554 60734 31556 60786
rect 31500 60732 31556 60734
rect 32508 61346 32564 61348
rect 32508 61294 32510 61346
rect 32510 61294 32562 61346
rect 32562 61294 32564 61346
rect 32508 61292 32564 61294
rect 31724 59948 31780 60004
rect 31612 59724 31668 59780
rect 32060 60620 32116 60676
rect 32396 60172 32452 60228
rect 32284 60060 32340 60116
rect 31612 58492 31668 58548
rect 31388 58210 31444 58212
rect 31388 58158 31390 58210
rect 31390 58158 31442 58210
rect 31442 58158 31444 58210
rect 31388 58156 31444 58158
rect 31164 56588 31220 56644
rect 30268 56140 30324 56196
rect 31164 56028 31220 56084
rect 30380 54460 30436 54516
rect 30940 53676 30996 53732
rect 30268 53564 30324 53620
rect 30828 53618 30884 53620
rect 30828 53566 30830 53618
rect 30830 53566 30882 53618
rect 30882 53566 30884 53618
rect 30828 53564 30884 53566
rect 30268 52892 30324 52948
rect 30044 52274 30100 52276
rect 30044 52222 30046 52274
rect 30046 52222 30098 52274
rect 30098 52222 30100 52274
rect 30044 52220 30100 52222
rect 30268 52162 30324 52164
rect 30268 52110 30270 52162
rect 30270 52110 30322 52162
rect 30322 52110 30324 52162
rect 30268 52108 30324 52110
rect 29596 49196 29652 49252
rect 30156 50652 30212 50708
rect 28700 48412 28756 48468
rect 30380 48524 30436 48580
rect 29260 47570 29316 47572
rect 29260 47518 29262 47570
rect 29262 47518 29314 47570
rect 29314 47518 29316 47570
rect 29260 47516 29316 47518
rect 29484 47292 29540 47348
rect 27468 46732 27524 46788
rect 27916 46844 27972 46900
rect 28364 46956 28420 47012
rect 27244 44994 27300 44996
rect 27244 44942 27246 44994
rect 27246 44942 27298 44994
rect 27298 44942 27300 44994
rect 27244 44940 27300 44942
rect 26012 44268 26068 44324
rect 26236 44828 26292 44884
rect 26012 43260 26068 43316
rect 26124 42812 26180 42868
rect 26796 43260 26852 43316
rect 26572 42812 26628 42868
rect 26236 41916 26292 41972
rect 25788 41356 25844 41412
rect 25788 41186 25844 41188
rect 25788 41134 25790 41186
rect 25790 41134 25842 41186
rect 25842 41134 25844 41186
rect 25788 41132 25844 41134
rect 26012 41298 26068 41300
rect 26012 41246 26014 41298
rect 26014 41246 26066 41298
rect 26066 41246 26068 41298
rect 26012 41244 26068 41246
rect 27020 42754 27076 42756
rect 27020 42702 27022 42754
rect 27022 42702 27074 42754
rect 27074 42702 27076 42754
rect 27020 42700 27076 42702
rect 27020 41970 27076 41972
rect 27020 41918 27022 41970
rect 27022 41918 27074 41970
rect 27074 41918 27076 41970
rect 27020 41916 27076 41918
rect 26908 41186 26964 41188
rect 26908 41134 26910 41186
rect 26910 41134 26962 41186
rect 26962 41134 26964 41186
rect 26908 41132 26964 41134
rect 26796 40572 26852 40628
rect 27132 41692 27188 41748
rect 27356 41356 27412 41412
rect 27020 40348 27076 40404
rect 26124 39730 26180 39732
rect 26124 39678 26126 39730
rect 26126 39678 26178 39730
rect 26178 39678 26180 39730
rect 26124 39676 26180 39678
rect 25676 39618 25732 39620
rect 25676 39566 25678 39618
rect 25678 39566 25730 39618
rect 25730 39566 25732 39618
rect 25676 39564 25732 39566
rect 27804 45724 27860 45780
rect 28700 46956 28756 47012
rect 30828 52946 30884 52948
rect 30828 52894 30830 52946
rect 30830 52894 30882 52946
rect 30882 52894 30884 52946
rect 30828 52892 30884 52894
rect 31276 53676 31332 53732
rect 33180 61010 33236 61012
rect 33180 60958 33182 61010
rect 33182 60958 33234 61010
rect 33234 60958 33236 61010
rect 33180 60956 33236 60958
rect 33068 60844 33124 60900
rect 33292 60786 33348 60788
rect 33292 60734 33294 60786
rect 33294 60734 33346 60786
rect 33346 60734 33348 60786
rect 33292 60732 33348 60734
rect 34412 62412 34468 62468
rect 33628 61292 33684 61348
rect 33740 62300 33796 62356
rect 36316 65436 36372 65492
rect 37660 65490 37716 65492
rect 37660 65438 37662 65490
rect 37662 65438 37714 65490
rect 37714 65438 37716 65490
rect 37660 65436 37716 65438
rect 36988 64930 37044 64932
rect 36988 64878 36990 64930
rect 36990 64878 37042 64930
rect 37042 64878 37044 64930
rect 36988 64876 37044 64878
rect 37324 64988 37380 65044
rect 37324 63868 37380 63924
rect 35868 63026 35924 63028
rect 35868 62974 35870 63026
rect 35870 62974 35922 63026
rect 35922 62974 35924 63026
rect 35868 62972 35924 62974
rect 35532 62914 35588 62916
rect 35532 62862 35534 62914
rect 35534 62862 35586 62914
rect 35586 62862 35588 62914
rect 35532 62860 35588 62862
rect 35756 62914 35812 62916
rect 35756 62862 35758 62914
rect 35758 62862 35810 62914
rect 35810 62862 35812 62914
rect 35756 62860 35812 62862
rect 36764 62578 36820 62580
rect 36764 62526 36766 62578
rect 36766 62526 36818 62578
rect 36818 62526 36820 62578
rect 36764 62524 36820 62526
rect 36764 62076 36820 62132
rect 37548 62860 37604 62916
rect 37772 62076 37828 62132
rect 36204 61570 36260 61572
rect 36204 61518 36206 61570
rect 36206 61518 36258 61570
rect 36258 61518 36260 61570
rect 36204 61516 36260 61518
rect 33852 61346 33908 61348
rect 33852 61294 33854 61346
rect 33854 61294 33906 61346
rect 33906 61294 33908 61346
rect 33852 61292 33908 61294
rect 34412 61346 34468 61348
rect 34412 61294 34414 61346
rect 34414 61294 34466 61346
rect 34466 61294 34468 61346
rect 34412 61292 34468 61294
rect 34008 61178 34064 61180
rect 34112 61178 34168 61180
rect 34008 61126 34024 61178
rect 34024 61126 34064 61178
rect 34112 61126 34148 61178
rect 34148 61126 34168 61178
rect 34008 61124 34064 61126
rect 34112 61124 34168 61126
rect 34216 61124 34272 61180
rect 34320 61178 34376 61180
rect 34424 61178 34480 61180
rect 34528 61178 34584 61180
rect 34320 61126 34324 61178
rect 34324 61126 34376 61178
rect 34424 61126 34448 61178
rect 34448 61126 34480 61178
rect 34528 61126 34572 61178
rect 34572 61126 34584 61178
rect 34320 61124 34376 61126
rect 34424 61124 34480 61126
rect 34528 61124 34584 61126
rect 34632 61178 34688 61180
rect 34736 61178 34792 61180
rect 34840 61178 34896 61180
rect 34632 61126 34644 61178
rect 34644 61126 34688 61178
rect 34736 61126 34768 61178
rect 34768 61126 34792 61178
rect 34840 61126 34892 61178
rect 34892 61126 34896 61178
rect 34632 61124 34688 61126
rect 34736 61124 34792 61126
rect 34840 61124 34896 61126
rect 34944 61124 35000 61180
rect 35048 61178 35104 61180
rect 35152 61178 35208 61180
rect 35048 61126 35068 61178
rect 35068 61126 35104 61178
rect 35152 61126 35192 61178
rect 35192 61126 35208 61178
rect 35048 61124 35104 61126
rect 35152 61124 35208 61126
rect 33404 60620 33460 60676
rect 33740 60674 33796 60676
rect 33740 60622 33742 60674
rect 33742 60622 33794 60674
rect 33794 60622 33796 60674
rect 33740 60620 33796 60622
rect 33180 60562 33236 60564
rect 33180 60510 33182 60562
rect 33182 60510 33234 60562
rect 33234 60510 33236 60562
rect 33180 60508 33236 60510
rect 32508 59388 32564 59444
rect 33180 59778 33236 59780
rect 33180 59726 33182 59778
rect 33182 59726 33234 59778
rect 33234 59726 33236 59778
rect 33180 59724 33236 59726
rect 33180 59388 33236 59444
rect 33068 59330 33124 59332
rect 33068 59278 33070 59330
rect 33070 59278 33122 59330
rect 33122 59278 33124 59330
rect 33068 59276 33124 59278
rect 33292 58828 33348 58884
rect 32284 58546 32340 58548
rect 32284 58494 32286 58546
rect 32286 58494 32338 58546
rect 32338 58494 32340 58546
rect 32284 58492 32340 58494
rect 33404 58380 33460 58436
rect 32732 58210 32788 58212
rect 32732 58158 32734 58210
rect 32734 58158 32786 58210
rect 32786 58158 32788 58210
rect 32732 58156 32788 58158
rect 32060 56194 32116 56196
rect 32060 56142 32062 56194
rect 32062 56142 32114 56194
rect 32114 56142 32116 56194
rect 32060 56140 32116 56142
rect 33964 60226 34020 60228
rect 33964 60174 33966 60226
rect 33966 60174 34018 60226
rect 34018 60174 34020 60226
rect 33964 60172 34020 60174
rect 36204 60172 36260 60228
rect 37324 61570 37380 61572
rect 37324 61518 37326 61570
rect 37326 61518 37378 61570
rect 37378 61518 37380 61570
rect 37324 61516 37380 61518
rect 37548 60172 37604 60228
rect 38332 60172 38388 60228
rect 36428 60002 36484 60004
rect 36428 59950 36430 60002
rect 36430 59950 36482 60002
rect 36482 59950 36484 60002
rect 36428 59948 36484 59950
rect 37324 60002 37380 60004
rect 37324 59950 37326 60002
rect 37326 59950 37378 60002
rect 37378 59950 37380 60002
rect 37324 59948 37380 59950
rect 34300 59778 34356 59780
rect 34300 59726 34302 59778
rect 34302 59726 34354 59778
rect 34354 59726 34356 59778
rect 34300 59724 34356 59726
rect 34008 59610 34064 59612
rect 34112 59610 34168 59612
rect 34008 59558 34024 59610
rect 34024 59558 34064 59610
rect 34112 59558 34148 59610
rect 34148 59558 34168 59610
rect 34008 59556 34064 59558
rect 34112 59556 34168 59558
rect 34216 59556 34272 59612
rect 34320 59610 34376 59612
rect 34424 59610 34480 59612
rect 34528 59610 34584 59612
rect 34320 59558 34324 59610
rect 34324 59558 34376 59610
rect 34424 59558 34448 59610
rect 34448 59558 34480 59610
rect 34528 59558 34572 59610
rect 34572 59558 34584 59610
rect 34320 59556 34376 59558
rect 34424 59556 34480 59558
rect 34528 59556 34584 59558
rect 34632 59610 34688 59612
rect 34736 59610 34792 59612
rect 34840 59610 34896 59612
rect 34632 59558 34644 59610
rect 34644 59558 34688 59610
rect 34736 59558 34768 59610
rect 34768 59558 34792 59610
rect 34840 59558 34892 59610
rect 34892 59558 34896 59610
rect 34632 59556 34688 59558
rect 34736 59556 34792 59558
rect 34840 59556 34896 59558
rect 34944 59556 35000 59612
rect 35048 59610 35104 59612
rect 35152 59610 35208 59612
rect 35048 59558 35068 59610
rect 35068 59558 35104 59610
rect 35152 59558 35192 59610
rect 35192 59558 35208 59610
rect 35048 59556 35104 59558
rect 35152 59556 35208 59558
rect 34412 58268 34468 58324
rect 35196 58434 35252 58436
rect 35196 58382 35198 58434
rect 35198 58382 35250 58434
rect 35250 58382 35252 58434
rect 35196 58380 35252 58382
rect 34972 58156 35028 58212
rect 35084 58268 35140 58324
rect 35532 58322 35588 58324
rect 35532 58270 35534 58322
rect 35534 58270 35586 58322
rect 35586 58270 35588 58322
rect 35532 58268 35588 58270
rect 34008 58042 34064 58044
rect 34112 58042 34168 58044
rect 34008 57990 34024 58042
rect 34024 57990 34064 58042
rect 34112 57990 34148 58042
rect 34148 57990 34168 58042
rect 34008 57988 34064 57990
rect 34112 57988 34168 57990
rect 34216 57988 34272 58044
rect 34320 58042 34376 58044
rect 34424 58042 34480 58044
rect 34528 58042 34584 58044
rect 34320 57990 34324 58042
rect 34324 57990 34376 58042
rect 34424 57990 34448 58042
rect 34448 57990 34480 58042
rect 34528 57990 34572 58042
rect 34572 57990 34584 58042
rect 34320 57988 34376 57990
rect 34424 57988 34480 57990
rect 34528 57988 34584 57990
rect 34632 58042 34688 58044
rect 34736 58042 34792 58044
rect 34840 58042 34896 58044
rect 34632 57990 34644 58042
rect 34644 57990 34688 58042
rect 34736 57990 34768 58042
rect 34768 57990 34792 58042
rect 34840 57990 34892 58042
rect 34892 57990 34896 58042
rect 34632 57988 34688 57990
rect 34736 57988 34792 57990
rect 34840 57988 34896 57990
rect 34944 57988 35000 58044
rect 35048 58042 35104 58044
rect 35152 58042 35208 58044
rect 35048 57990 35068 58042
rect 35068 57990 35104 58042
rect 35152 57990 35192 58042
rect 35192 57990 35208 58042
rect 35048 57988 35104 57990
rect 35152 57988 35208 57990
rect 33404 57596 33460 57652
rect 32508 56082 32564 56084
rect 32508 56030 32510 56082
rect 32510 56030 32562 56082
rect 32562 56030 32564 56082
rect 32508 56028 32564 56030
rect 31388 53618 31444 53620
rect 31388 53566 31390 53618
rect 31390 53566 31442 53618
rect 31442 53566 31444 53618
rect 31388 53564 31444 53566
rect 31948 53618 32004 53620
rect 31948 53566 31950 53618
rect 31950 53566 32002 53618
rect 32002 53566 32004 53618
rect 31948 53564 32004 53566
rect 31276 53116 31332 53172
rect 31052 52220 31108 52276
rect 30716 52050 30772 52052
rect 30716 51998 30718 52050
rect 30718 51998 30770 52050
rect 30770 51998 30772 52050
rect 30716 51996 30772 51998
rect 30828 51938 30884 51940
rect 30828 51886 30830 51938
rect 30830 51886 30882 51938
rect 30882 51886 30884 51938
rect 30828 51884 30884 51886
rect 30940 51602 30996 51604
rect 30940 51550 30942 51602
rect 30942 51550 30994 51602
rect 30994 51550 30996 51602
rect 30940 51548 30996 51550
rect 30716 50706 30772 50708
rect 30716 50654 30718 50706
rect 30718 50654 30770 50706
rect 30770 50654 30772 50706
rect 30716 50652 30772 50654
rect 31052 49084 31108 49140
rect 31612 52108 31668 52164
rect 31724 51996 31780 52052
rect 32172 51884 32228 51940
rect 31164 49644 31220 49700
rect 30828 48466 30884 48468
rect 30828 48414 30830 48466
rect 30830 48414 30882 48466
rect 30882 48414 30884 48466
rect 30828 48412 30884 48414
rect 30492 48300 30548 48356
rect 30716 47404 30772 47460
rect 31724 49196 31780 49252
rect 31948 51378 32004 51380
rect 31948 51326 31950 51378
rect 31950 51326 32002 51378
rect 32002 51326 32004 51378
rect 31948 51324 32004 51326
rect 32620 51324 32676 51380
rect 31612 48914 31668 48916
rect 31612 48862 31614 48914
rect 31614 48862 31666 48914
rect 31666 48862 31668 48914
rect 31612 48860 31668 48862
rect 31276 48524 31332 48580
rect 31164 48242 31220 48244
rect 31164 48190 31166 48242
rect 31166 48190 31218 48242
rect 31218 48190 31220 48242
rect 31164 48188 31220 48190
rect 31276 48300 31332 48356
rect 32172 49138 32228 49140
rect 32172 49086 32174 49138
rect 32174 49086 32226 49138
rect 32226 49086 32228 49138
rect 32172 49084 32228 49086
rect 31836 48802 31892 48804
rect 31836 48750 31838 48802
rect 31838 48750 31890 48802
rect 31890 48750 31892 48802
rect 31836 48748 31892 48750
rect 31836 48242 31892 48244
rect 31836 48190 31838 48242
rect 31838 48190 31890 48242
rect 31890 48190 31892 48242
rect 31836 48188 31892 48190
rect 30380 47346 30436 47348
rect 30380 47294 30382 47346
rect 30382 47294 30434 47346
rect 30434 47294 30436 47346
rect 30380 47292 30436 47294
rect 31276 47180 31332 47236
rect 31500 47458 31556 47460
rect 31500 47406 31502 47458
rect 31502 47406 31554 47458
rect 31554 47406 31556 47458
rect 31500 47404 31556 47406
rect 29596 46956 29652 47012
rect 28700 45778 28756 45780
rect 28700 45726 28702 45778
rect 28702 45726 28754 45778
rect 28754 45726 28756 45778
rect 28700 45724 28756 45726
rect 28140 45666 28196 45668
rect 28140 45614 28142 45666
rect 28142 45614 28194 45666
rect 28194 45614 28196 45666
rect 28140 45612 28196 45614
rect 29260 45666 29316 45668
rect 29260 45614 29262 45666
rect 29262 45614 29314 45666
rect 29314 45614 29316 45666
rect 29260 45612 29316 45614
rect 27692 45106 27748 45108
rect 27692 45054 27694 45106
rect 27694 45054 27746 45106
rect 27746 45054 27748 45106
rect 27692 45052 27748 45054
rect 27580 44994 27636 44996
rect 27580 44942 27582 44994
rect 27582 44942 27634 44994
rect 27634 44942 27636 44994
rect 27580 44940 27636 44942
rect 29148 43650 29204 43652
rect 29148 43598 29150 43650
rect 29150 43598 29202 43650
rect 29202 43598 29204 43650
rect 29148 43596 29204 43598
rect 28140 42812 28196 42868
rect 27580 42754 27636 42756
rect 27580 42702 27582 42754
rect 27582 42702 27634 42754
rect 27634 42702 27636 42754
rect 27580 42700 27636 42702
rect 27804 41298 27860 41300
rect 27804 41246 27806 41298
rect 27806 41246 27858 41298
rect 27858 41246 27860 41298
rect 27804 41244 27860 41246
rect 29372 45500 29428 45556
rect 30156 46114 30212 46116
rect 30156 46062 30158 46114
rect 30158 46062 30210 46114
rect 30210 46062 30212 46114
rect 30156 46060 30212 46062
rect 30044 45778 30100 45780
rect 30044 45726 30046 45778
rect 30046 45726 30098 45778
rect 30098 45726 30100 45778
rect 30044 45724 30100 45726
rect 29820 45612 29876 45668
rect 29484 43484 29540 43540
rect 29372 43372 29428 43428
rect 29596 42812 29652 42868
rect 29260 41916 29316 41972
rect 28476 41186 28532 41188
rect 28476 41134 28478 41186
rect 28478 41134 28530 41186
rect 28530 41134 28532 41186
rect 28476 41132 28532 41134
rect 27916 40962 27972 40964
rect 27916 40910 27918 40962
rect 27918 40910 27970 40962
rect 27970 40910 27972 40962
rect 27916 40908 27972 40910
rect 29148 40908 29204 40964
rect 29036 40684 29092 40740
rect 25564 38108 25620 38164
rect 24668 37490 24724 37492
rect 24668 37438 24670 37490
rect 24670 37438 24722 37490
rect 24722 37438 24724 37490
rect 24668 37436 24724 37438
rect 23436 35532 23492 35588
rect 23212 34748 23268 34804
rect 21756 34018 21812 34020
rect 21756 33966 21758 34018
rect 21758 33966 21810 34018
rect 21810 33966 21812 34018
rect 21756 33964 21812 33966
rect 23212 33628 23268 33684
rect 22204 33516 22260 33572
rect 23548 35420 23604 35476
rect 27804 40348 27860 40404
rect 26460 37548 26516 37604
rect 25900 37436 25956 37492
rect 26684 37436 26740 37492
rect 27020 37378 27076 37380
rect 27020 37326 27022 37378
rect 27022 37326 27074 37378
rect 27074 37326 27076 37378
rect 27020 37324 27076 37326
rect 26684 37212 26740 37268
rect 24008 36874 24064 36876
rect 24112 36874 24168 36876
rect 24008 36822 24024 36874
rect 24024 36822 24064 36874
rect 24112 36822 24148 36874
rect 24148 36822 24168 36874
rect 24008 36820 24064 36822
rect 24112 36820 24168 36822
rect 24216 36820 24272 36876
rect 24320 36874 24376 36876
rect 24424 36874 24480 36876
rect 24528 36874 24584 36876
rect 24320 36822 24324 36874
rect 24324 36822 24376 36874
rect 24424 36822 24448 36874
rect 24448 36822 24480 36874
rect 24528 36822 24572 36874
rect 24572 36822 24584 36874
rect 24320 36820 24376 36822
rect 24424 36820 24480 36822
rect 24528 36820 24584 36822
rect 24632 36874 24688 36876
rect 24736 36874 24792 36876
rect 24840 36874 24896 36876
rect 24632 36822 24644 36874
rect 24644 36822 24688 36874
rect 24736 36822 24768 36874
rect 24768 36822 24792 36874
rect 24840 36822 24892 36874
rect 24892 36822 24896 36874
rect 24632 36820 24688 36822
rect 24736 36820 24792 36822
rect 24840 36820 24896 36822
rect 24944 36820 25000 36876
rect 25048 36874 25104 36876
rect 25152 36874 25208 36876
rect 25048 36822 25068 36874
rect 25068 36822 25104 36874
rect 25152 36822 25192 36874
rect 25192 36822 25208 36874
rect 25048 36820 25104 36822
rect 25152 36820 25208 36822
rect 25340 35756 25396 35812
rect 23660 35196 23716 35252
rect 23996 35698 24052 35700
rect 23996 35646 23998 35698
rect 23998 35646 24050 35698
rect 24050 35646 24052 35698
rect 23996 35644 24052 35646
rect 23436 33516 23492 33572
rect 22540 33458 22596 33460
rect 22540 33406 22542 33458
rect 22542 33406 22594 33458
rect 22594 33406 22596 33458
rect 22540 33404 22596 33406
rect 22428 33068 22484 33124
rect 21756 31836 21812 31892
rect 22316 29538 22372 29540
rect 22316 29486 22318 29538
rect 22318 29486 22370 29538
rect 22370 29486 22372 29538
rect 22316 29484 22372 29486
rect 21644 28812 21700 28868
rect 20076 28700 20132 28756
rect 21980 28754 22036 28756
rect 21980 28702 21982 28754
rect 21982 28702 22034 28754
rect 22034 28702 22036 28754
rect 21980 28700 22036 28702
rect 20076 28028 20132 28084
rect 17836 23714 17892 23716
rect 17836 23662 17838 23714
rect 17838 23662 17890 23714
rect 17890 23662 17892 23714
rect 17836 23660 17892 23662
rect 18732 24946 18788 24948
rect 18732 24894 18734 24946
rect 18734 24894 18786 24946
rect 18786 24894 18788 24946
rect 18732 24892 18788 24894
rect 19516 24892 19572 24948
rect 18284 24610 18340 24612
rect 18284 24558 18286 24610
rect 18286 24558 18338 24610
rect 18338 24558 18340 24610
rect 18284 24556 18340 24558
rect 19740 24556 19796 24612
rect 18844 23826 18900 23828
rect 18844 23774 18846 23826
rect 18846 23774 18898 23826
rect 18898 23774 18900 23826
rect 18844 23772 18900 23774
rect 20972 27858 21028 27860
rect 20972 27806 20974 27858
rect 20974 27806 21026 27858
rect 21026 27806 21028 27858
rect 20972 27804 21028 27806
rect 20972 27244 21028 27300
rect 20412 26460 20468 26516
rect 21196 26684 21252 26740
rect 22316 27244 22372 27300
rect 21420 26572 21476 26628
rect 21980 26684 22036 26740
rect 21756 26514 21812 26516
rect 21756 26462 21758 26514
rect 21758 26462 21810 26514
rect 21810 26462 21812 26514
rect 21756 26460 21812 26462
rect 20300 25676 20356 25732
rect 20748 25676 20804 25732
rect 19852 23826 19908 23828
rect 19852 23774 19854 23826
rect 19854 23774 19906 23826
rect 19906 23774 19908 23826
rect 19852 23772 19908 23774
rect 20188 24556 20244 24612
rect 18284 23548 18340 23604
rect 18396 22988 18452 23044
rect 17500 22316 17556 22372
rect 20412 23826 20468 23828
rect 20412 23774 20414 23826
rect 20414 23774 20466 23826
rect 20466 23774 20468 23826
rect 20412 23772 20468 23774
rect 20636 23660 20692 23716
rect 20412 22316 20468 22372
rect 20188 22204 20244 22260
rect 18508 22146 18564 22148
rect 18508 22094 18510 22146
rect 18510 22094 18562 22146
rect 18562 22094 18564 22146
rect 18508 22092 18564 22094
rect 16716 21698 16772 21700
rect 16716 21646 16718 21698
rect 16718 21646 16770 21698
rect 16770 21646 16772 21698
rect 16716 21644 16772 21646
rect 16604 21586 16660 21588
rect 16604 21534 16606 21586
rect 16606 21534 16658 21586
rect 16658 21534 16660 21586
rect 16604 21532 16660 21534
rect 16716 20860 16772 20916
rect 16492 19964 16548 20020
rect 16604 19852 16660 19908
rect 16268 16940 16324 16996
rect 16380 18956 16436 19012
rect 16716 18450 16772 18452
rect 16716 18398 16718 18450
rect 16718 18398 16770 18450
rect 16770 18398 16772 18450
rect 16716 18396 16772 18398
rect 16604 18284 16660 18340
rect 16492 17164 16548 17220
rect 16716 16044 16772 16100
rect 16716 14924 16772 14980
rect 19404 22146 19460 22148
rect 19404 22094 19406 22146
rect 19406 22094 19458 22146
rect 19458 22094 19460 22146
rect 19404 22092 19460 22094
rect 18620 21644 18676 21700
rect 17500 21586 17556 21588
rect 17500 21534 17502 21586
rect 17502 21534 17554 21586
rect 17554 21534 17556 21586
rect 17500 21532 17556 21534
rect 18284 20130 18340 20132
rect 18284 20078 18286 20130
rect 18286 20078 18338 20130
rect 18338 20078 18340 20130
rect 18284 20076 18340 20078
rect 18060 18956 18116 19012
rect 17052 16828 17108 16884
rect 17164 14700 17220 14756
rect 18732 20130 18788 20132
rect 18732 20078 18734 20130
rect 18734 20078 18786 20130
rect 18786 20078 18788 20130
rect 18732 20076 18788 20078
rect 20300 20076 20356 20132
rect 18956 19234 19012 19236
rect 18956 19182 18958 19234
rect 18958 19182 19010 19234
rect 19010 19182 19012 19234
rect 18956 19180 19012 19182
rect 18508 19068 18564 19124
rect 17948 17778 18004 17780
rect 17948 17726 17950 17778
rect 17950 17726 18002 17778
rect 18002 17726 18004 17778
rect 17948 17724 18004 17726
rect 17612 16882 17668 16884
rect 17612 16830 17614 16882
rect 17614 16830 17666 16882
rect 17666 16830 17668 16882
rect 17612 16828 17668 16830
rect 17612 16098 17668 16100
rect 17612 16046 17614 16098
rect 17614 16046 17666 16098
rect 17666 16046 17668 16098
rect 17612 16044 17668 16046
rect 17612 14364 17668 14420
rect 16828 13804 16884 13860
rect 18060 17388 18116 17444
rect 18060 15932 18116 15988
rect 18620 17554 18676 17556
rect 18620 17502 18622 17554
rect 18622 17502 18674 17554
rect 18674 17502 18676 17554
rect 18620 17500 18676 17502
rect 18508 17388 18564 17444
rect 19516 19122 19572 19124
rect 19516 19070 19518 19122
rect 19518 19070 19570 19122
rect 19570 19070 19572 19122
rect 19516 19068 19572 19070
rect 19628 19010 19684 19012
rect 19628 18958 19630 19010
rect 19630 18958 19682 19010
rect 19682 18958 19684 19010
rect 19628 18956 19684 18958
rect 19292 18172 19348 18228
rect 20524 19404 20580 19460
rect 20524 19234 20580 19236
rect 20524 19182 20526 19234
rect 20526 19182 20578 19234
rect 20578 19182 20580 19234
rect 20524 19180 20580 19182
rect 20300 19122 20356 19124
rect 20300 19070 20302 19122
rect 20302 19070 20354 19122
rect 20354 19070 20356 19122
rect 20300 19068 20356 19070
rect 19404 17666 19460 17668
rect 19404 17614 19406 17666
rect 19406 17614 19458 17666
rect 19458 17614 19460 17666
rect 19404 17612 19460 17614
rect 19292 17500 19348 17556
rect 18508 17164 18564 17220
rect 18172 16940 18228 16996
rect 19292 16716 19348 16772
rect 18732 15314 18788 15316
rect 18732 15262 18734 15314
rect 18734 15262 18786 15314
rect 18786 15262 18788 15314
rect 18732 15260 18788 15262
rect 22092 26460 22148 26516
rect 21420 25228 21476 25284
rect 23436 32732 23492 32788
rect 22988 32620 23044 32676
rect 23660 32620 23716 32676
rect 22988 31890 23044 31892
rect 22988 31838 22990 31890
rect 22990 31838 23042 31890
rect 23042 31838 23044 31890
rect 22988 31836 23044 31838
rect 22540 31778 22596 31780
rect 22540 31726 22542 31778
rect 22542 31726 22594 31778
rect 22594 31726 22596 31778
rect 22540 31724 22596 31726
rect 23212 30268 23268 30324
rect 22988 28866 23044 28868
rect 22988 28814 22990 28866
rect 22990 28814 23042 28866
rect 23042 28814 23044 28866
rect 22988 28812 23044 28814
rect 23324 29538 23380 29540
rect 23324 29486 23326 29538
rect 23326 29486 23378 29538
rect 23378 29486 23380 29538
rect 23324 29484 23380 29486
rect 23436 28700 23492 28756
rect 22652 26124 22708 26180
rect 22316 25282 22372 25284
rect 22316 25230 22318 25282
rect 22318 25230 22370 25282
rect 22370 25230 22372 25282
rect 22316 25228 22372 25230
rect 22876 23996 22932 24052
rect 20972 23324 21028 23380
rect 20860 22482 20916 22484
rect 20860 22430 20862 22482
rect 20862 22430 20914 22482
rect 20914 22430 20916 22482
rect 20860 22428 20916 22430
rect 20972 22092 21028 22148
rect 21756 23772 21812 23828
rect 22764 23826 22820 23828
rect 22764 23774 22766 23826
rect 22766 23774 22818 23826
rect 22818 23774 22820 23826
rect 22764 23772 22820 23774
rect 23548 27692 23604 27748
rect 23212 26572 23268 26628
rect 23436 25228 23492 25284
rect 23100 24444 23156 24500
rect 21868 23324 21924 23380
rect 23436 23324 23492 23380
rect 21980 23212 22036 23268
rect 21308 22988 21364 23044
rect 20748 20860 20804 20916
rect 21756 22482 21812 22484
rect 21756 22430 21758 22482
rect 21758 22430 21810 22482
rect 21810 22430 21812 22482
rect 21756 22428 21812 22430
rect 23100 22370 23156 22372
rect 23100 22318 23102 22370
rect 23102 22318 23154 22370
rect 23154 22318 23156 22370
rect 23100 22316 23156 22318
rect 21980 22258 22036 22260
rect 21980 22206 21982 22258
rect 21982 22206 22034 22258
rect 22034 22206 22036 22258
rect 21980 22204 22036 22206
rect 21420 20972 21476 21028
rect 21532 21532 21588 21588
rect 22204 21026 22260 21028
rect 22204 20974 22206 21026
rect 22206 20974 22258 21026
rect 22258 20974 22260 21026
rect 22204 20972 22260 20974
rect 21532 20748 21588 20804
rect 22428 20748 22484 20804
rect 22988 21308 23044 21364
rect 23324 22092 23380 22148
rect 23436 21980 23492 22036
rect 23660 28082 23716 28084
rect 23660 28030 23662 28082
rect 23662 28030 23714 28082
rect 23714 28030 23716 28082
rect 23660 28028 23716 28030
rect 24444 35586 24500 35588
rect 24444 35534 24446 35586
rect 24446 35534 24498 35586
rect 24498 35534 24500 35586
rect 24444 35532 24500 35534
rect 25340 35474 25396 35476
rect 25340 35422 25342 35474
rect 25342 35422 25394 35474
rect 25394 35422 25396 35474
rect 25340 35420 25396 35422
rect 24008 35306 24064 35308
rect 24112 35306 24168 35308
rect 24008 35254 24024 35306
rect 24024 35254 24064 35306
rect 24112 35254 24148 35306
rect 24148 35254 24168 35306
rect 24008 35252 24064 35254
rect 24112 35252 24168 35254
rect 24216 35252 24272 35308
rect 24320 35306 24376 35308
rect 24424 35306 24480 35308
rect 24528 35306 24584 35308
rect 24320 35254 24324 35306
rect 24324 35254 24376 35306
rect 24424 35254 24448 35306
rect 24448 35254 24480 35306
rect 24528 35254 24572 35306
rect 24572 35254 24584 35306
rect 24320 35252 24376 35254
rect 24424 35252 24480 35254
rect 24528 35252 24584 35254
rect 24632 35306 24688 35308
rect 24736 35306 24792 35308
rect 24840 35306 24896 35308
rect 24632 35254 24644 35306
rect 24644 35254 24688 35306
rect 24736 35254 24768 35306
rect 24768 35254 24792 35306
rect 24840 35254 24892 35306
rect 24892 35254 24896 35306
rect 24632 35252 24688 35254
rect 24736 35252 24792 35254
rect 24840 35252 24896 35254
rect 24944 35252 25000 35308
rect 25048 35306 25104 35308
rect 25152 35306 25208 35308
rect 25048 35254 25068 35306
rect 25068 35254 25104 35306
rect 25152 35254 25192 35306
rect 25192 35254 25208 35306
rect 25048 35252 25104 35254
rect 25152 35252 25208 35254
rect 26460 36988 26516 37044
rect 25900 35810 25956 35812
rect 25900 35758 25902 35810
rect 25902 35758 25954 35810
rect 25954 35758 25956 35810
rect 25900 35756 25956 35758
rect 26908 37212 26964 37268
rect 26684 35420 26740 35476
rect 26012 34860 26068 34916
rect 25788 34802 25844 34804
rect 25788 34750 25790 34802
rect 25790 34750 25842 34802
rect 25842 34750 25844 34802
rect 25788 34748 25844 34750
rect 24008 33738 24064 33740
rect 24112 33738 24168 33740
rect 24008 33686 24024 33738
rect 24024 33686 24064 33738
rect 24112 33686 24148 33738
rect 24148 33686 24168 33738
rect 24008 33684 24064 33686
rect 24112 33684 24168 33686
rect 24216 33684 24272 33740
rect 24320 33738 24376 33740
rect 24424 33738 24480 33740
rect 24528 33738 24584 33740
rect 24320 33686 24324 33738
rect 24324 33686 24376 33738
rect 24424 33686 24448 33738
rect 24448 33686 24480 33738
rect 24528 33686 24572 33738
rect 24572 33686 24584 33738
rect 24320 33684 24376 33686
rect 24424 33684 24480 33686
rect 24528 33684 24584 33686
rect 24632 33738 24688 33740
rect 24736 33738 24792 33740
rect 24840 33738 24896 33740
rect 24632 33686 24644 33738
rect 24644 33686 24688 33738
rect 24736 33686 24768 33738
rect 24768 33686 24792 33738
rect 24840 33686 24892 33738
rect 24892 33686 24896 33738
rect 24632 33684 24688 33686
rect 24736 33684 24792 33686
rect 24840 33684 24896 33686
rect 24944 33684 25000 33740
rect 25048 33738 25104 33740
rect 25152 33738 25208 33740
rect 25048 33686 25068 33738
rect 25068 33686 25104 33738
rect 25152 33686 25192 33738
rect 25192 33686 25208 33738
rect 25048 33684 25104 33686
rect 25152 33684 25208 33686
rect 23996 33516 24052 33572
rect 23884 33458 23940 33460
rect 23884 33406 23886 33458
rect 23886 33406 23938 33458
rect 23938 33406 23940 33458
rect 23884 33404 23940 33406
rect 23996 32844 24052 32900
rect 24668 33068 24724 33124
rect 25228 33122 25284 33124
rect 25228 33070 25230 33122
rect 25230 33070 25282 33122
rect 25282 33070 25284 33122
rect 25228 33068 25284 33070
rect 25452 34524 25508 34580
rect 25452 33404 25508 33460
rect 24444 32620 24500 32676
rect 25340 32844 25396 32900
rect 23884 32284 23940 32340
rect 24780 32338 24836 32340
rect 24780 32286 24782 32338
rect 24782 32286 24834 32338
rect 24834 32286 24836 32338
rect 24780 32284 24836 32286
rect 24008 32170 24064 32172
rect 24112 32170 24168 32172
rect 24008 32118 24024 32170
rect 24024 32118 24064 32170
rect 24112 32118 24148 32170
rect 24148 32118 24168 32170
rect 24008 32116 24064 32118
rect 24112 32116 24168 32118
rect 24216 32116 24272 32172
rect 24320 32170 24376 32172
rect 24424 32170 24480 32172
rect 24528 32170 24584 32172
rect 24320 32118 24324 32170
rect 24324 32118 24376 32170
rect 24424 32118 24448 32170
rect 24448 32118 24480 32170
rect 24528 32118 24572 32170
rect 24572 32118 24584 32170
rect 24320 32116 24376 32118
rect 24424 32116 24480 32118
rect 24528 32116 24584 32118
rect 24632 32170 24688 32172
rect 24736 32170 24792 32172
rect 24840 32170 24896 32172
rect 24632 32118 24644 32170
rect 24644 32118 24688 32170
rect 24736 32118 24768 32170
rect 24768 32118 24792 32170
rect 24840 32118 24892 32170
rect 24892 32118 24896 32170
rect 24632 32116 24688 32118
rect 24736 32116 24792 32118
rect 24840 32116 24896 32118
rect 24944 32116 25000 32172
rect 25048 32170 25104 32172
rect 25152 32170 25208 32172
rect 25048 32118 25068 32170
rect 25068 32118 25104 32170
rect 25152 32118 25192 32170
rect 25192 32118 25208 32170
rect 25048 32116 25104 32118
rect 25152 32116 25208 32118
rect 23996 31836 24052 31892
rect 24008 30602 24064 30604
rect 24112 30602 24168 30604
rect 24008 30550 24024 30602
rect 24024 30550 24064 30602
rect 24112 30550 24148 30602
rect 24148 30550 24168 30602
rect 24008 30548 24064 30550
rect 24112 30548 24168 30550
rect 24216 30548 24272 30604
rect 24320 30602 24376 30604
rect 24424 30602 24480 30604
rect 24528 30602 24584 30604
rect 24320 30550 24324 30602
rect 24324 30550 24376 30602
rect 24424 30550 24448 30602
rect 24448 30550 24480 30602
rect 24528 30550 24572 30602
rect 24572 30550 24584 30602
rect 24320 30548 24376 30550
rect 24424 30548 24480 30550
rect 24528 30548 24584 30550
rect 24632 30602 24688 30604
rect 24736 30602 24792 30604
rect 24840 30602 24896 30604
rect 24632 30550 24644 30602
rect 24644 30550 24688 30602
rect 24736 30550 24768 30602
rect 24768 30550 24792 30602
rect 24840 30550 24892 30602
rect 24892 30550 24896 30602
rect 24632 30548 24688 30550
rect 24736 30548 24792 30550
rect 24840 30548 24896 30550
rect 24944 30548 25000 30604
rect 25048 30602 25104 30604
rect 25152 30602 25208 30604
rect 25048 30550 25068 30602
rect 25068 30550 25104 30602
rect 25152 30550 25192 30602
rect 25192 30550 25208 30602
rect 25048 30548 25104 30550
rect 25152 30548 25208 30550
rect 25340 30156 25396 30212
rect 24008 29034 24064 29036
rect 24112 29034 24168 29036
rect 24008 28982 24024 29034
rect 24024 28982 24064 29034
rect 24112 28982 24148 29034
rect 24148 28982 24168 29034
rect 24008 28980 24064 28982
rect 24112 28980 24168 28982
rect 24216 28980 24272 29036
rect 24320 29034 24376 29036
rect 24424 29034 24480 29036
rect 24528 29034 24584 29036
rect 24320 28982 24324 29034
rect 24324 28982 24376 29034
rect 24424 28982 24448 29034
rect 24448 28982 24480 29034
rect 24528 28982 24572 29034
rect 24572 28982 24584 29034
rect 24320 28980 24376 28982
rect 24424 28980 24480 28982
rect 24528 28980 24584 28982
rect 24632 29034 24688 29036
rect 24736 29034 24792 29036
rect 24840 29034 24896 29036
rect 24632 28982 24644 29034
rect 24644 28982 24688 29034
rect 24736 28982 24768 29034
rect 24768 28982 24792 29034
rect 24840 28982 24892 29034
rect 24892 28982 24896 29034
rect 24632 28980 24688 28982
rect 24736 28980 24792 28982
rect 24840 28980 24896 28982
rect 24944 28980 25000 29036
rect 25048 29034 25104 29036
rect 25152 29034 25208 29036
rect 25048 28982 25068 29034
rect 25068 28982 25104 29034
rect 25152 28982 25192 29034
rect 25192 28982 25208 29034
rect 25048 28980 25104 28982
rect 25152 28980 25208 28982
rect 23884 27804 23940 27860
rect 25452 31836 25508 31892
rect 25564 31666 25620 31668
rect 25564 31614 25566 31666
rect 25566 31614 25618 31666
rect 25618 31614 25620 31666
rect 25564 31612 25620 31614
rect 27020 36428 27076 36484
rect 26908 34860 26964 34916
rect 27580 37772 27636 37828
rect 29708 41298 29764 41300
rect 29708 41246 29710 41298
rect 29710 41246 29762 41298
rect 29762 41246 29764 41298
rect 29708 41244 29764 41246
rect 29484 39730 29540 39732
rect 29484 39678 29486 39730
rect 29486 39678 29538 39730
rect 29538 39678 29540 39730
rect 29484 39676 29540 39678
rect 29932 41916 29988 41972
rect 29932 40684 29988 40740
rect 32284 48860 32340 48916
rect 31612 46844 31668 46900
rect 30940 46060 30996 46116
rect 31948 46508 32004 46564
rect 32060 48188 32116 48244
rect 30492 43596 30548 43652
rect 30156 43538 30212 43540
rect 30156 43486 30158 43538
rect 30158 43486 30210 43538
rect 30210 43486 30212 43538
rect 30156 43484 30212 43486
rect 30940 43426 30996 43428
rect 30940 43374 30942 43426
rect 30942 43374 30994 43426
rect 30994 43374 30996 43426
rect 30940 43372 30996 43374
rect 30268 42866 30324 42868
rect 30268 42814 30270 42866
rect 30270 42814 30322 42866
rect 30322 42814 30324 42866
rect 30268 42812 30324 42814
rect 30156 42476 30212 42532
rect 30492 42700 30548 42756
rect 30268 41916 30324 41972
rect 30828 42140 30884 42196
rect 31276 42476 31332 42532
rect 31052 41970 31108 41972
rect 31052 41918 31054 41970
rect 31054 41918 31106 41970
rect 31106 41918 31108 41970
rect 31052 41916 31108 41918
rect 30828 41356 30884 41412
rect 30268 41298 30324 41300
rect 30268 41246 30270 41298
rect 30270 41246 30322 41298
rect 30322 41246 30324 41298
rect 30268 41244 30324 41246
rect 30268 40572 30324 40628
rect 29932 40348 29988 40404
rect 30156 40460 30212 40516
rect 28252 39564 28308 39620
rect 27580 37378 27636 37380
rect 27580 37326 27582 37378
rect 27582 37326 27634 37378
rect 27634 37326 27636 37378
rect 27580 37324 27636 37326
rect 27356 36988 27412 37044
rect 28028 37548 28084 37604
rect 28252 37436 28308 37492
rect 27916 37212 27972 37268
rect 28252 37266 28308 37268
rect 28252 37214 28254 37266
rect 28254 37214 28306 37266
rect 28306 37214 28308 37266
rect 28252 37212 28308 37214
rect 27804 36988 27860 37044
rect 28028 37100 28084 37156
rect 27692 36652 27748 36708
rect 27692 36482 27748 36484
rect 27692 36430 27694 36482
rect 27694 36430 27746 36482
rect 27746 36430 27748 36482
rect 27692 36428 27748 36430
rect 29484 36988 29540 37044
rect 29036 36652 29092 36708
rect 30156 39676 30212 39732
rect 30604 41298 30660 41300
rect 30604 41246 30606 41298
rect 30606 41246 30658 41298
rect 30658 41246 30660 41298
rect 30604 41244 30660 41246
rect 30716 41186 30772 41188
rect 30716 41134 30718 41186
rect 30718 41134 30770 41186
rect 30770 41134 30772 41186
rect 30716 41132 30772 41134
rect 30604 40684 30660 40740
rect 29820 36988 29876 37044
rect 30492 39676 30548 39732
rect 30492 37772 30548 37828
rect 31724 42476 31780 42532
rect 32172 47404 32228 47460
rect 32172 47234 32228 47236
rect 32172 47182 32174 47234
rect 32174 47182 32226 47234
rect 32226 47182 32228 47234
rect 32172 47180 32228 47182
rect 32172 46898 32228 46900
rect 32172 46846 32174 46898
rect 32174 46846 32226 46898
rect 32226 46846 32228 46898
rect 32172 46844 32228 46846
rect 32508 48188 32564 48244
rect 32396 46732 32452 46788
rect 34076 57650 34132 57652
rect 34076 57598 34078 57650
rect 34078 57598 34130 57650
rect 34130 57598 34132 57650
rect 34076 57596 34132 57598
rect 34300 57874 34356 57876
rect 34300 57822 34302 57874
rect 34302 57822 34354 57874
rect 34354 57822 34356 57874
rect 34300 57820 34356 57822
rect 33292 56082 33348 56084
rect 33292 56030 33294 56082
rect 33294 56030 33346 56082
rect 33346 56030 33348 56082
rect 33292 56028 33348 56030
rect 33628 56028 33684 56084
rect 33852 56642 33908 56644
rect 33852 56590 33854 56642
rect 33854 56590 33906 56642
rect 33906 56590 33908 56642
rect 33852 56588 33908 56590
rect 34300 56642 34356 56644
rect 34300 56590 34302 56642
rect 34302 56590 34354 56642
rect 34354 56590 34356 56642
rect 34300 56588 34356 56590
rect 34860 57260 34916 57316
rect 34748 56924 34804 56980
rect 36876 58268 36932 58324
rect 35532 57260 35588 57316
rect 36428 58156 36484 58212
rect 36204 57090 36260 57092
rect 36204 57038 36206 57090
rect 36206 57038 36258 57090
rect 36258 57038 36260 57090
rect 36204 57036 36260 57038
rect 35084 56588 35140 56644
rect 34008 56474 34064 56476
rect 34112 56474 34168 56476
rect 34008 56422 34024 56474
rect 34024 56422 34064 56474
rect 34112 56422 34148 56474
rect 34148 56422 34168 56474
rect 34008 56420 34064 56422
rect 34112 56420 34168 56422
rect 34216 56420 34272 56476
rect 34320 56474 34376 56476
rect 34424 56474 34480 56476
rect 34528 56474 34584 56476
rect 34320 56422 34324 56474
rect 34324 56422 34376 56474
rect 34424 56422 34448 56474
rect 34448 56422 34480 56474
rect 34528 56422 34572 56474
rect 34572 56422 34584 56474
rect 34320 56420 34376 56422
rect 34424 56420 34480 56422
rect 34528 56420 34584 56422
rect 34632 56474 34688 56476
rect 34736 56474 34792 56476
rect 34840 56474 34896 56476
rect 34632 56422 34644 56474
rect 34644 56422 34688 56474
rect 34736 56422 34768 56474
rect 34768 56422 34792 56474
rect 34840 56422 34892 56474
rect 34892 56422 34896 56474
rect 34632 56420 34688 56422
rect 34736 56420 34792 56422
rect 34840 56420 34896 56422
rect 34944 56420 35000 56476
rect 35048 56474 35104 56476
rect 35152 56474 35208 56476
rect 35048 56422 35068 56474
rect 35068 56422 35104 56474
rect 35152 56422 35192 56474
rect 35192 56422 35208 56474
rect 35048 56420 35104 56422
rect 35152 56420 35208 56422
rect 36764 56924 36820 56980
rect 35980 56588 36036 56644
rect 36428 56588 36484 56644
rect 35308 56252 35364 56308
rect 36204 56306 36260 56308
rect 36204 56254 36206 56306
rect 36206 56254 36258 56306
rect 36258 56254 36260 56306
rect 36204 56252 36260 56254
rect 33852 55916 33908 55972
rect 35756 55916 35812 55972
rect 37100 58210 37156 58212
rect 37100 58158 37102 58210
rect 37102 58158 37154 58210
rect 37154 58158 37156 58210
rect 37100 58156 37156 58158
rect 36988 57090 37044 57092
rect 36988 57038 36990 57090
rect 36990 57038 37042 57090
rect 37042 57038 37044 57090
rect 36988 57036 37044 57038
rect 36988 56700 37044 56756
rect 37436 56754 37492 56756
rect 37436 56702 37438 56754
rect 37438 56702 37490 56754
rect 37490 56702 37492 56754
rect 37436 56700 37492 56702
rect 37100 55970 37156 55972
rect 37100 55918 37102 55970
rect 37102 55918 37154 55970
rect 37154 55918 37156 55970
rect 37100 55916 37156 55918
rect 36428 55244 36484 55300
rect 37100 55298 37156 55300
rect 37100 55246 37102 55298
rect 37102 55246 37154 55298
rect 37154 55246 37156 55298
rect 37100 55244 37156 55246
rect 37660 56252 37716 56308
rect 34008 54906 34064 54908
rect 34112 54906 34168 54908
rect 34008 54854 34024 54906
rect 34024 54854 34064 54906
rect 34112 54854 34148 54906
rect 34148 54854 34168 54906
rect 34008 54852 34064 54854
rect 34112 54852 34168 54854
rect 34216 54852 34272 54908
rect 34320 54906 34376 54908
rect 34424 54906 34480 54908
rect 34528 54906 34584 54908
rect 34320 54854 34324 54906
rect 34324 54854 34376 54906
rect 34424 54854 34448 54906
rect 34448 54854 34480 54906
rect 34528 54854 34572 54906
rect 34572 54854 34584 54906
rect 34320 54852 34376 54854
rect 34424 54852 34480 54854
rect 34528 54852 34584 54854
rect 34632 54906 34688 54908
rect 34736 54906 34792 54908
rect 34840 54906 34896 54908
rect 34632 54854 34644 54906
rect 34644 54854 34688 54906
rect 34736 54854 34768 54906
rect 34768 54854 34792 54906
rect 34840 54854 34892 54906
rect 34892 54854 34896 54906
rect 34632 54852 34688 54854
rect 34736 54852 34792 54854
rect 34840 54852 34896 54854
rect 34944 54852 35000 54908
rect 35048 54906 35104 54908
rect 35152 54906 35208 54908
rect 35048 54854 35068 54906
rect 35068 54854 35104 54906
rect 35152 54854 35192 54906
rect 35192 54854 35208 54906
rect 35048 54852 35104 54854
rect 35152 54852 35208 54854
rect 33180 51884 33236 51940
rect 34008 53338 34064 53340
rect 34112 53338 34168 53340
rect 34008 53286 34024 53338
rect 34024 53286 34064 53338
rect 34112 53286 34148 53338
rect 34148 53286 34168 53338
rect 34008 53284 34064 53286
rect 34112 53284 34168 53286
rect 34216 53284 34272 53340
rect 34320 53338 34376 53340
rect 34424 53338 34480 53340
rect 34528 53338 34584 53340
rect 34320 53286 34324 53338
rect 34324 53286 34376 53338
rect 34424 53286 34448 53338
rect 34448 53286 34480 53338
rect 34528 53286 34572 53338
rect 34572 53286 34584 53338
rect 34320 53284 34376 53286
rect 34424 53284 34480 53286
rect 34528 53284 34584 53286
rect 34632 53338 34688 53340
rect 34736 53338 34792 53340
rect 34840 53338 34896 53340
rect 34632 53286 34644 53338
rect 34644 53286 34688 53338
rect 34736 53286 34768 53338
rect 34768 53286 34792 53338
rect 34840 53286 34892 53338
rect 34892 53286 34896 53338
rect 34632 53284 34688 53286
rect 34736 53284 34792 53286
rect 34840 53284 34896 53286
rect 34944 53284 35000 53340
rect 35048 53338 35104 53340
rect 35152 53338 35208 53340
rect 35048 53286 35068 53338
rect 35068 53286 35104 53338
rect 35152 53286 35192 53338
rect 35192 53286 35208 53338
rect 35048 53284 35104 53286
rect 35152 53284 35208 53286
rect 33180 51378 33236 51380
rect 33180 51326 33182 51378
rect 33182 51326 33234 51378
rect 33234 51326 33236 51378
rect 33180 51324 33236 51326
rect 34860 51938 34916 51940
rect 34860 51886 34862 51938
rect 34862 51886 34914 51938
rect 34914 51886 34916 51938
rect 34860 51884 34916 51886
rect 34008 51770 34064 51772
rect 34112 51770 34168 51772
rect 34008 51718 34024 51770
rect 34024 51718 34064 51770
rect 34112 51718 34148 51770
rect 34148 51718 34168 51770
rect 34008 51716 34064 51718
rect 34112 51716 34168 51718
rect 34216 51716 34272 51772
rect 34320 51770 34376 51772
rect 34424 51770 34480 51772
rect 34528 51770 34584 51772
rect 34320 51718 34324 51770
rect 34324 51718 34376 51770
rect 34424 51718 34448 51770
rect 34448 51718 34480 51770
rect 34528 51718 34572 51770
rect 34572 51718 34584 51770
rect 34320 51716 34376 51718
rect 34424 51716 34480 51718
rect 34528 51716 34584 51718
rect 34632 51770 34688 51772
rect 34736 51770 34792 51772
rect 34840 51770 34896 51772
rect 34632 51718 34644 51770
rect 34644 51718 34688 51770
rect 34736 51718 34768 51770
rect 34768 51718 34792 51770
rect 34840 51718 34892 51770
rect 34892 51718 34896 51770
rect 34632 51716 34688 51718
rect 34736 51716 34792 51718
rect 34840 51716 34896 51718
rect 34944 51716 35000 51772
rect 35048 51770 35104 51772
rect 35152 51770 35208 51772
rect 35048 51718 35068 51770
rect 35068 51718 35104 51770
rect 35152 51718 35192 51770
rect 35192 51718 35208 51770
rect 35048 51716 35104 51718
rect 35152 51716 35208 51718
rect 33852 51548 33908 51604
rect 33852 50428 33908 50484
rect 34524 50482 34580 50484
rect 34524 50430 34526 50482
rect 34526 50430 34578 50482
rect 34578 50430 34580 50482
rect 34524 50428 34580 50430
rect 34008 50202 34064 50204
rect 34112 50202 34168 50204
rect 34008 50150 34024 50202
rect 34024 50150 34064 50202
rect 34112 50150 34148 50202
rect 34148 50150 34168 50202
rect 34008 50148 34064 50150
rect 34112 50148 34168 50150
rect 34216 50148 34272 50204
rect 34320 50202 34376 50204
rect 34424 50202 34480 50204
rect 34528 50202 34584 50204
rect 34320 50150 34324 50202
rect 34324 50150 34376 50202
rect 34424 50150 34448 50202
rect 34448 50150 34480 50202
rect 34528 50150 34572 50202
rect 34572 50150 34584 50202
rect 34320 50148 34376 50150
rect 34424 50148 34480 50150
rect 34528 50148 34584 50150
rect 34632 50202 34688 50204
rect 34736 50202 34792 50204
rect 34840 50202 34896 50204
rect 34632 50150 34644 50202
rect 34644 50150 34688 50202
rect 34736 50150 34768 50202
rect 34768 50150 34792 50202
rect 34840 50150 34892 50202
rect 34892 50150 34896 50202
rect 34632 50148 34688 50150
rect 34736 50148 34792 50150
rect 34840 50148 34896 50150
rect 34944 50148 35000 50204
rect 35048 50202 35104 50204
rect 35152 50202 35208 50204
rect 35048 50150 35068 50202
rect 35068 50150 35104 50202
rect 35152 50150 35192 50202
rect 35192 50150 35208 50202
rect 35048 50148 35104 50150
rect 35152 50148 35208 50150
rect 33180 49698 33236 49700
rect 33180 49646 33182 49698
rect 33182 49646 33234 49698
rect 33234 49646 33236 49698
rect 33180 49644 33236 49646
rect 33740 49644 33796 49700
rect 33516 49250 33572 49252
rect 33516 49198 33518 49250
rect 33518 49198 33570 49250
rect 33570 49198 33572 49250
rect 33516 49196 33572 49198
rect 33068 49026 33124 49028
rect 33068 48974 33070 49026
rect 33070 48974 33122 49026
rect 33122 48974 33124 49026
rect 33068 48972 33124 48974
rect 33628 49026 33684 49028
rect 33628 48974 33630 49026
rect 33630 48974 33682 49026
rect 33682 48974 33684 49026
rect 33628 48972 33684 48974
rect 32732 46956 32788 47012
rect 32620 46620 32676 46676
rect 33180 46562 33236 46564
rect 33180 46510 33182 46562
rect 33182 46510 33234 46562
rect 33234 46510 33236 46562
rect 33180 46508 33236 46510
rect 34300 48802 34356 48804
rect 34300 48750 34302 48802
rect 34302 48750 34354 48802
rect 34354 48750 34356 48802
rect 34300 48748 34356 48750
rect 34008 48634 34064 48636
rect 34112 48634 34168 48636
rect 34008 48582 34024 48634
rect 34024 48582 34064 48634
rect 34112 48582 34148 48634
rect 34148 48582 34168 48634
rect 34008 48580 34064 48582
rect 34112 48580 34168 48582
rect 34216 48580 34272 48636
rect 34320 48634 34376 48636
rect 34424 48634 34480 48636
rect 34528 48634 34584 48636
rect 34320 48582 34324 48634
rect 34324 48582 34376 48634
rect 34424 48582 34448 48634
rect 34448 48582 34480 48634
rect 34528 48582 34572 48634
rect 34572 48582 34584 48634
rect 34320 48580 34376 48582
rect 34424 48580 34480 48582
rect 34528 48580 34584 48582
rect 34632 48634 34688 48636
rect 34736 48634 34792 48636
rect 34840 48634 34896 48636
rect 34632 48582 34644 48634
rect 34644 48582 34688 48634
rect 34736 48582 34768 48634
rect 34768 48582 34792 48634
rect 34840 48582 34892 48634
rect 34892 48582 34896 48634
rect 34632 48580 34688 48582
rect 34736 48580 34792 48582
rect 34840 48580 34896 48582
rect 34944 48580 35000 48636
rect 35048 48634 35104 48636
rect 35152 48634 35208 48636
rect 35048 48582 35068 48634
rect 35068 48582 35104 48634
rect 35152 48582 35192 48634
rect 35192 48582 35208 48634
rect 35048 48580 35104 48582
rect 35152 48580 35208 48582
rect 34076 48242 34132 48244
rect 34076 48190 34078 48242
rect 34078 48190 34130 48242
rect 34130 48190 34132 48242
rect 34076 48188 34132 48190
rect 32284 46284 32340 46340
rect 33628 46396 33684 46452
rect 33180 45612 33236 45668
rect 33628 45388 33684 45444
rect 32508 44994 32564 44996
rect 32508 44942 32510 44994
rect 32510 44942 32562 44994
rect 32562 44942 32564 44994
rect 32508 44940 32564 44942
rect 34008 47066 34064 47068
rect 34112 47066 34168 47068
rect 34008 47014 34024 47066
rect 34024 47014 34064 47066
rect 34112 47014 34148 47066
rect 34148 47014 34168 47066
rect 34008 47012 34064 47014
rect 34112 47012 34168 47014
rect 34216 47012 34272 47068
rect 34320 47066 34376 47068
rect 34424 47066 34480 47068
rect 34528 47066 34584 47068
rect 34320 47014 34324 47066
rect 34324 47014 34376 47066
rect 34424 47014 34448 47066
rect 34448 47014 34480 47066
rect 34528 47014 34572 47066
rect 34572 47014 34584 47066
rect 34320 47012 34376 47014
rect 34424 47012 34480 47014
rect 34528 47012 34584 47014
rect 34632 47066 34688 47068
rect 34736 47066 34792 47068
rect 34840 47066 34896 47068
rect 34632 47014 34644 47066
rect 34644 47014 34688 47066
rect 34736 47014 34768 47066
rect 34768 47014 34792 47066
rect 34840 47014 34892 47066
rect 34892 47014 34896 47066
rect 34632 47012 34688 47014
rect 34736 47012 34792 47014
rect 34840 47012 34896 47014
rect 34944 47012 35000 47068
rect 35048 47066 35104 47068
rect 35152 47066 35208 47068
rect 35048 47014 35068 47066
rect 35068 47014 35104 47066
rect 35152 47014 35192 47066
rect 35192 47014 35208 47066
rect 35048 47012 35104 47014
rect 35152 47012 35208 47014
rect 34524 46786 34580 46788
rect 34524 46734 34526 46786
rect 34526 46734 34578 46786
rect 34578 46734 34580 46786
rect 34524 46732 34580 46734
rect 34188 46674 34244 46676
rect 34188 46622 34190 46674
rect 34190 46622 34242 46674
rect 34242 46622 34244 46674
rect 34188 46620 34244 46622
rect 34636 46284 34692 46340
rect 36428 48636 36484 48692
rect 36316 46844 36372 46900
rect 35756 46508 35812 46564
rect 35308 46396 35364 46452
rect 35644 46396 35700 46452
rect 35532 46284 35588 46340
rect 35420 45724 35476 45780
rect 34008 45498 34064 45500
rect 34112 45498 34168 45500
rect 34008 45446 34024 45498
rect 34024 45446 34064 45498
rect 34112 45446 34148 45498
rect 34148 45446 34168 45498
rect 34008 45444 34064 45446
rect 34112 45444 34168 45446
rect 34216 45444 34272 45500
rect 34320 45498 34376 45500
rect 34424 45498 34480 45500
rect 34528 45498 34584 45500
rect 34320 45446 34324 45498
rect 34324 45446 34376 45498
rect 34424 45446 34448 45498
rect 34448 45446 34480 45498
rect 34528 45446 34572 45498
rect 34572 45446 34584 45498
rect 34320 45444 34376 45446
rect 34424 45444 34480 45446
rect 34528 45444 34584 45446
rect 34632 45498 34688 45500
rect 34736 45498 34792 45500
rect 34840 45498 34896 45500
rect 34632 45446 34644 45498
rect 34644 45446 34688 45498
rect 34736 45446 34768 45498
rect 34768 45446 34792 45498
rect 34840 45446 34892 45498
rect 34892 45446 34896 45498
rect 34632 45444 34688 45446
rect 34736 45444 34792 45446
rect 34840 45444 34896 45446
rect 34944 45444 35000 45500
rect 35048 45498 35104 45500
rect 35152 45498 35208 45500
rect 35048 45446 35068 45498
rect 35068 45446 35104 45498
rect 35152 45446 35192 45498
rect 35192 45446 35208 45498
rect 35048 45444 35104 45446
rect 35152 45444 35208 45446
rect 34300 45276 34356 45332
rect 34860 45218 34916 45220
rect 34860 45166 34862 45218
rect 34862 45166 34914 45218
rect 34914 45166 34916 45218
rect 34860 45164 34916 45166
rect 33852 44994 33908 44996
rect 33852 44942 33854 44994
rect 33854 44942 33906 44994
rect 33906 44942 33908 44994
rect 33852 44940 33908 44942
rect 33740 44268 33796 44324
rect 34524 44322 34580 44324
rect 34524 44270 34526 44322
rect 34526 44270 34578 44322
rect 34578 44270 34580 44322
rect 34524 44268 34580 44270
rect 36204 46674 36260 46676
rect 36204 46622 36206 46674
rect 36206 46622 36258 46674
rect 36258 46622 36260 46674
rect 36204 46620 36260 46622
rect 35980 46396 36036 46452
rect 35756 45890 35812 45892
rect 35756 45838 35758 45890
rect 35758 45838 35810 45890
rect 35810 45838 35812 45890
rect 35756 45836 35812 45838
rect 36316 46284 36372 46340
rect 34748 44882 34804 44884
rect 34748 44830 34750 44882
rect 34750 44830 34802 44882
rect 34802 44830 34804 44882
rect 34748 44828 34804 44830
rect 34636 44210 34692 44212
rect 34636 44158 34638 44210
rect 34638 44158 34690 44210
rect 34690 44158 34692 44210
rect 34636 44156 34692 44158
rect 33852 44098 33908 44100
rect 33852 44046 33854 44098
rect 33854 44046 33906 44098
rect 33906 44046 33908 44098
rect 33852 44044 33908 44046
rect 32508 43372 32564 43428
rect 32172 42140 32228 42196
rect 31724 41580 31780 41636
rect 32172 41410 32228 41412
rect 32172 41358 32174 41410
rect 32174 41358 32226 41410
rect 32226 41358 32228 41410
rect 32172 41356 32228 41358
rect 32060 41186 32116 41188
rect 32060 41134 32062 41186
rect 32062 41134 32114 41186
rect 32114 41134 32116 41186
rect 32060 41132 32116 41134
rect 32396 41244 32452 41300
rect 32284 41132 32340 41188
rect 31612 40572 31668 40628
rect 30940 40348 30996 40404
rect 31500 40236 31556 40292
rect 32172 40402 32228 40404
rect 32172 40350 32174 40402
rect 32174 40350 32226 40402
rect 32226 40350 32228 40402
rect 32172 40348 32228 40350
rect 32396 40178 32452 40180
rect 32396 40126 32398 40178
rect 32398 40126 32450 40178
rect 32450 40126 32452 40178
rect 32396 40124 32452 40126
rect 30604 37436 30660 37492
rect 31836 38668 31892 38724
rect 30492 37212 30548 37268
rect 27356 35756 27412 35812
rect 27244 35474 27300 35476
rect 27244 35422 27246 35474
rect 27246 35422 27298 35474
rect 27298 35422 27300 35474
rect 27244 35420 27300 35422
rect 27804 35810 27860 35812
rect 27804 35758 27806 35810
rect 27806 35758 27858 35810
rect 27858 35758 27860 35810
rect 27804 35756 27860 35758
rect 27804 34802 27860 34804
rect 27804 34750 27806 34802
rect 27806 34750 27858 34802
rect 27858 34750 27860 34802
rect 27804 34748 27860 34750
rect 27132 34636 27188 34692
rect 26236 33458 26292 33460
rect 26236 33406 26238 33458
rect 26238 33406 26290 33458
rect 26290 33406 26292 33458
rect 26236 33404 26292 33406
rect 27020 33404 27076 33460
rect 25788 32786 25844 32788
rect 25788 32734 25790 32786
rect 25790 32734 25842 32786
rect 25842 32734 25844 32786
rect 25788 32732 25844 32734
rect 26236 32674 26292 32676
rect 26236 32622 26238 32674
rect 26238 32622 26290 32674
rect 26290 32622 26292 32674
rect 26236 32620 26292 32622
rect 27244 32674 27300 32676
rect 27244 32622 27246 32674
rect 27246 32622 27298 32674
rect 27298 32622 27300 32674
rect 27244 32620 27300 32622
rect 26236 32284 26292 32340
rect 26348 31836 26404 31892
rect 26572 31554 26628 31556
rect 26572 31502 26574 31554
rect 26574 31502 26626 31554
rect 26626 31502 26628 31554
rect 26572 31500 26628 31502
rect 27692 31778 27748 31780
rect 27692 31726 27694 31778
rect 27694 31726 27746 31778
rect 27746 31726 27748 31778
rect 27692 31724 27748 31726
rect 27132 31612 27188 31668
rect 27356 31554 27412 31556
rect 27356 31502 27358 31554
rect 27358 31502 27410 31554
rect 27410 31502 27412 31554
rect 27356 31500 27412 31502
rect 28252 34860 28308 34916
rect 31052 37826 31108 37828
rect 31052 37774 31054 37826
rect 31054 37774 31106 37826
rect 31106 37774 31108 37826
rect 31052 37772 31108 37774
rect 31164 37490 31220 37492
rect 31164 37438 31166 37490
rect 31166 37438 31218 37490
rect 31218 37438 31220 37490
rect 31164 37436 31220 37438
rect 31164 37100 31220 37156
rect 28476 35756 28532 35812
rect 28364 34300 28420 34356
rect 29708 34354 29764 34356
rect 29708 34302 29710 34354
rect 29710 34302 29762 34354
rect 29762 34302 29764 34354
rect 29708 34300 29764 34302
rect 28252 33628 28308 33684
rect 28028 31666 28084 31668
rect 28028 31614 28030 31666
rect 28030 31614 28082 31666
rect 28082 31614 28084 31666
rect 28028 31612 28084 31614
rect 28476 31724 28532 31780
rect 27804 31388 27860 31444
rect 27468 31052 27524 31108
rect 26012 30268 26068 30324
rect 25452 29932 25508 29988
rect 25340 28082 25396 28084
rect 25340 28030 25342 28082
rect 25342 28030 25394 28082
rect 25394 28030 25396 28082
rect 25340 28028 25396 28030
rect 24444 27746 24500 27748
rect 24444 27694 24446 27746
rect 24446 27694 24498 27746
rect 24498 27694 24500 27746
rect 24444 27692 24500 27694
rect 24008 27466 24064 27468
rect 24112 27466 24168 27468
rect 24008 27414 24024 27466
rect 24024 27414 24064 27466
rect 24112 27414 24148 27466
rect 24148 27414 24168 27466
rect 24008 27412 24064 27414
rect 24112 27412 24168 27414
rect 24216 27412 24272 27468
rect 24320 27466 24376 27468
rect 24424 27466 24480 27468
rect 24528 27466 24584 27468
rect 24320 27414 24324 27466
rect 24324 27414 24376 27466
rect 24424 27414 24448 27466
rect 24448 27414 24480 27466
rect 24528 27414 24572 27466
rect 24572 27414 24584 27466
rect 24320 27412 24376 27414
rect 24424 27412 24480 27414
rect 24528 27412 24584 27414
rect 24632 27466 24688 27468
rect 24736 27466 24792 27468
rect 24840 27466 24896 27468
rect 24632 27414 24644 27466
rect 24644 27414 24688 27466
rect 24736 27414 24768 27466
rect 24768 27414 24792 27466
rect 24840 27414 24892 27466
rect 24892 27414 24896 27466
rect 24632 27412 24688 27414
rect 24736 27412 24792 27414
rect 24840 27412 24896 27414
rect 24944 27412 25000 27468
rect 25048 27466 25104 27468
rect 25152 27466 25208 27468
rect 25048 27414 25068 27466
rect 25068 27414 25104 27466
rect 25152 27414 25192 27466
rect 25192 27414 25208 27466
rect 25048 27412 25104 27414
rect 25152 27412 25208 27414
rect 25452 29372 25508 29428
rect 25452 28642 25508 28644
rect 25452 28590 25454 28642
rect 25454 28590 25506 28642
rect 25506 28590 25508 28642
rect 25452 28588 25508 28590
rect 26684 30156 26740 30212
rect 26124 29986 26180 29988
rect 26124 29934 26126 29986
rect 26126 29934 26178 29986
rect 26178 29934 26180 29986
rect 26124 29932 26180 29934
rect 29036 31106 29092 31108
rect 29036 31054 29038 31106
rect 29038 31054 29090 31106
rect 29090 31054 29092 31106
rect 29036 31052 29092 31054
rect 28364 30828 28420 30884
rect 28364 30268 28420 30324
rect 30156 34300 30212 34356
rect 30268 33628 30324 33684
rect 30156 32732 30212 32788
rect 29820 31836 29876 31892
rect 29932 32620 29988 32676
rect 29372 30882 29428 30884
rect 29372 30830 29374 30882
rect 29374 30830 29426 30882
rect 29426 30830 29428 30882
rect 29372 30828 29428 30830
rect 27692 30044 27748 30100
rect 28588 30098 28644 30100
rect 28588 30046 28590 30098
rect 28590 30046 28642 30098
rect 28642 30046 28644 30098
rect 28588 30044 28644 30046
rect 27580 29932 27636 29988
rect 27132 29426 27188 29428
rect 27132 29374 27134 29426
rect 27134 29374 27186 29426
rect 27186 29374 27188 29426
rect 27132 29372 27188 29374
rect 29260 29986 29316 29988
rect 29260 29934 29262 29986
rect 29262 29934 29314 29986
rect 29314 29934 29316 29986
rect 29260 29932 29316 29934
rect 29596 31500 29652 31556
rect 29820 30268 29876 30324
rect 29820 30098 29876 30100
rect 29820 30046 29822 30098
rect 29822 30046 29874 30098
rect 29874 30046 29876 30098
rect 29820 30044 29876 30046
rect 28140 28642 28196 28644
rect 28140 28590 28142 28642
rect 28142 28590 28194 28642
rect 28194 28590 28196 28642
rect 28140 28588 28196 28590
rect 29708 28588 29764 28644
rect 26012 28028 26068 28084
rect 25676 27804 25732 27860
rect 25788 27244 25844 27300
rect 25676 27132 25732 27188
rect 23660 26684 23716 26740
rect 23772 26178 23828 26180
rect 23772 26126 23774 26178
rect 23774 26126 23826 26178
rect 23826 26126 23828 26178
rect 23772 26124 23828 26126
rect 23772 25730 23828 25732
rect 23772 25678 23774 25730
rect 23774 25678 23826 25730
rect 23826 25678 23828 25730
rect 23772 25676 23828 25678
rect 23772 23660 23828 23716
rect 24008 25898 24064 25900
rect 24112 25898 24168 25900
rect 24008 25846 24024 25898
rect 24024 25846 24064 25898
rect 24112 25846 24148 25898
rect 24148 25846 24168 25898
rect 24008 25844 24064 25846
rect 24112 25844 24168 25846
rect 24216 25844 24272 25900
rect 24320 25898 24376 25900
rect 24424 25898 24480 25900
rect 24528 25898 24584 25900
rect 24320 25846 24324 25898
rect 24324 25846 24376 25898
rect 24424 25846 24448 25898
rect 24448 25846 24480 25898
rect 24528 25846 24572 25898
rect 24572 25846 24584 25898
rect 24320 25844 24376 25846
rect 24424 25844 24480 25846
rect 24528 25844 24584 25846
rect 24632 25898 24688 25900
rect 24736 25898 24792 25900
rect 24840 25898 24896 25900
rect 24632 25846 24644 25898
rect 24644 25846 24688 25898
rect 24736 25846 24768 25898
rect 24768 25846 24792 25898
rect 24840 25846 24892 25898
rect 24892 25846 24896 25898
rect 24632 25844 24688 25846
rect 24736 25844 24792 25846
rect 24840 25844 24896 25846
rect 24944 25844 25000 25900
rect 25048 25898 25104 25900
rect 25152 25898 25208 25900
rect 25048 25846 25068 25898
rect 25068 25846 25104 25898
rect 25152 25846 25192 25898
rect 25192 25846 25208 25898
rect 25048 25844 25104 25846
rect 25152 25844 25208 25846
rect 24556 25282 24612 25284
rect 24556 25230 24558 25282
rect 24558 25230 24610 25282
rect 24610 25230 24612 25282
rect 24556 25228 24612 25230
rect 24668 24834 24724 24836
rect 24668 24782 24670 24834
rect 24670 24782 24722 24834
rect 24722 24782 24724 24834
rect 24668 24780 24724 24782
rect 25452 24834 25508 24836
rect 25452 24782 25454 24834
rect 25454 24782 25506 24834
rect 25506 24782 25508 24834
rect 25452 24780 25508 24782
rect 25228 24498 25284 24500
rect 25228 24446 25230 24498
rect 25230 24446 25282 24498
rect 25282 24446 25284 24498
rect 25228 24444 25284 24446
rect 24008 24330 24064 24332
rect 24112 24330 24168 24332
rect 24008 24278 24024 24330
rect 24024 24278 24064 24330
rect 24112 24278 24148 24330
rect 24148 24278 24168 24330
rect 24008 24276 24064 24278
rect 24112 24276 24168 24278
rect 24216 24276 24272 24332
rect 24320 24330 24376 24332
rect 24424 24330 24480 24332
rect 24528 24330 24584 24332
rect 24320 24278 24324 24330
rect 24324 24278 24376 24330
rect 24424 24278 24448 24330
rect 24448 24278 24480 24330
rect 24528 24278 24572 24330
rect 24572 24278 24584 24330
rect 24320 24276 24376 24278
rect 24424 24276 24480 24278
rect 24528 24276 24584 24278
rect 24632 24330 24688 24332
rect 24736 24330 24792 24332
rect 24840 24330 24896 24332
rect 24632 24278 24644 24330
rect 24644 24278 24688 24330
rect 24736 24278 24768 24330
rect 24768 24278 24792 24330
rect 24840 24278 24892 24330
rect 24892 24278 24896 24330
rect 24632 24276 24688 24278
rect 24736 24276 24792 24278
rect 24840 24276 24896 24278
rect 24944 24276 25000 24332
rect 25048 24330 25104 24332
rect 25152 24330 25208 24332
rect 25048 24278 25068 24330
rect 25068 24278 25104 24330
rect 25152 24278 25192 24330
rect 25192 24278 25208 24330
rect 25048 24276 25104 24278
rect 25152 24276 25208 24278
rect 24556 24050 24612 24052
rect 24556 23998 24558 24050
rect 24558 23998 24610 24050
rect 24610 23998 24612 24050
rect 24556 23996 24612 23998
rect 23660 23042 23716 23044
rect 23660 22990 23662 23042
rect 23662 22990 23714 23042
rect 23714 22990 23716 23042
rect 23660 22988 23716 22990
rect 24892 23938 24948 23940
rect 24892 23886 24894 23938
rect 24894 23886 24946 23938
rect 24946 23886 24948 23938
rect 24892 23884 24948 23886
rect 24444 23660 24500 23716
rect 24668 23714 24724 23716
rect 24668 23662 24670 23714
rect 24670 23662 24722 23714
rect 24722 23662 24724 23714
rect 24668 23660 24724 23662
rect 24108 23212 24164 23268
rect 25340 23266 25396 23268
rect 25340 23214 25342 23266
rect 25342 23214 25394 23266
rect 25394 23214 25396 23266
rect 25340 23212 25396 23214
rect 24008 22762 24064 22764
rect 24112 22762 24168 22764
rect 24008 22710 24024 22762
rect 24024 22710 24064 22762
rect 24112 22710 24148 22762
rect 24148 22710 24168 22762
rect 24008 22708 24064 22710
rect 24112 22708 24168 22710
rect 24216 22708 24272 22764
rect 24320 22762 24376 22764
rect 24424 22762 24480 22764
rect 24528 22762 24584 22764
rect 24320 22710 24324 22762
rect 24324 22710 24376 22762
rect 24424 22710 24448 22762
rect 24448 22710 24480 22762
rect 24528 22710 24572 22762
rect 24572 22710 24584 22762
rect 24320 22708 24376 22710
rect 24424 22708 24480 22710
rect 24528 22708 24584 22710
rect 24632 22762 24688 22764
rect 24736 22762 24792 22764
rect 24840 22762 24896 22764
rect 24632 22710 24644 22762
rect 24644 22710 24688 22762
rect 24736 22710 24768 22762
rect 24768 22710 24792 22762
rect 24840 22710 24892 22762
rect 24892 22710 24896 22762
rect 24632 22708 24688 22710
rect 24736 22708 24792 22710
rect 24840 22708 24896 22710
rect 24944 22708 25000 22764
rect 25048 22762 25104 22764
rect 25152 22762 25208 22764
rect 25048 22710 25068 22762
rect 25068 22710 25104 22762
rect 25152 22710 25192 22762
rect 25192 22710 25208 22762
rect 25048 22708 25104 22710
rect 25152 22708 25208 22710
rect 23996 22540 24052 22596
rect 23884 22482 23940 22484
rect 23884 22430 23886 22482
rect 23886 22430 23938 22482
rect 23938 22430 23940 22482
rect 23884 22428 23940 22430
rect 23548 21756 23604 21812
rect 23212 20748 23268 20804
rect 23996 22092 24052 22148
rect 24892 22258 24948 22260
rect 24892 22206 24894 22258
rect 24894 22206 24946 22258
rect 24946 22206 24948 22258
rect 24892 22204 24948 22206
rect 25228 22204 25284 22260
rect 25452 22428 25508 22484
rect 25452 22092 25508 22148
rect 24668 21756 24724 21812
rect 24780 21362 24836 21364
rect 24780 21310 24782 21362
rect 24782 21310 24834 21362
rect 24834 21310 24836 21362
rect 24780 21308 24836 21310
rect 24008 21194 24064 21196
rect 24112 21194 24168 21196
rect 24008 21142 24024 21194
rect 24024 21142 24064 21194
rect 24112 21142 24148 21194
rect 24148 21142 24168 21194
rect 24008 21140 24064 21142
rect 24112 21140 24168 21142
rect 24216 21140 24272 21196
rect 24320 21194 24376 21196
rect 24424 21194 24480 21196
rect 24528 21194 24584 21196
rect 24320 21142 24324 21194
rect 24324 21142 24376 21194
rect 24424 21142 24448 21194
rect 24448 21142 24480 21194
rect 24528 21142 24572 21194
rect 24572 21142 24584 21194
rect 24320 21140 24376 21142
rect 24424 21140 24480 21142
rect 24528 21140 24584 21142
rect 24632 21194 24688 21196
rect 24736 21194 24792 21196
rect 24840 21194 24896 21196
rect 24632 21142 24644 21194
rect 24644 21142 24688 21194
rect 24736 21142 24768 21194
rect 24768 21142 24792 21194
rect 24840 21142 24892 21194
rect 24892 21142 24896 21194
rect 24632 21140 24688 21142
rect 24736 21140 24792 21142
rect 24840 21140 24896 21142
rect 24944 21140 25000 21196
rect 25048 21194 25104 21196
rect 25152 21194 25208 21196
rect 25048 21142 25068 21194
rect 25068 21142 25104 21194
rect 25152 21142 25192 21194
rect 25192 21142 25208 21194
rect 25048 21140 25104 21142
rect 25152 21140 25208 21142
rect 24220 20972 24276 21028
rect 24108 20860 24164 20916
rect 23660 20578 23716 20580
rect 23660 20526 23662 20578
rect 23662 20526 23714 20578
rect 23714 20526 23716 20578
rect 23660 20524 23716 20526
rect 22540 19964 22596 20020
rect 23212 19964 23268 20020
rect 21420 19740 21476 19796
rect 21420 19404 21476 19460
rect 21196 18450 21252 18452
rect 21196 18398 21198 18450
rect 21198 18398 21250 18450
rect 21250 18398 21252 18450
rect 21196 18396 21252 18398
rect 21084 18226 21140 18228
rect 21084 18174 21086 18226
rect 21086 18174 21138 18226
rect 21138 18174 21140 18226
rect 21084 18172 21140 18174
rect 20412 17666 20468 17668
rect 20412 17614 20414 17666
rect 20414 17614 20466 17666
rect 20466 17614 20468 17666
rect 20412 17612 20468 17614
rect 20076 17052 20132 17108
rect 19516 16658 19572 16660
rect 19516 16606 19518 16658
rect 19518 16606 19570 16658
rect 19570 16606 19572 16658
rect 19516 16604 19572 16606
rect 20860 17106 20916 17108
rect 20860 17054 20862 17106
rect 20862 17054 20914 17106
rect 20914 17054 20916 17106
rect 20860 17052 20916 17054
rect 20412 16882 20468 16884
rect 20412 16830 20414 16882
rect 20414 16830 20466 16882
rect 20466 16830 20468 16882
rect 20412 16828 20468 16830
rect 21532 17612 21588 17668
rect 20188 16716 20244 16772
rect 21084 16716 21140 16772
rect 20748 16658 20804 16660
rect 20748 16606 20750 16658
rect 20750 16606 20802 16658
rect 20802 16606 20804 16658
rect 20748 16604 20804 16606
rect 18172 14700 18228 14756
rect 20524 15148 20580 15204
rect 18620 14642 18676 14644
rect 18620 14590 18622 14642
rect 18622 14590 18674 14642
rect 18674 14590 18676 14642
rect 18620 14588 18676 14590
rect 19852 14642 19908 14644
rect 19852 14590 19854 14642
rect 19854 14590 19906 14642
rect 19906 14590 19908 14642
rect 19852 14588 19908 14590
rect 18060 13858 18116 13860
rect 18060 13806 18062 13858
rect 18062 13806 18114 13858
rect 18114 13806 18116 13858
rect 18060 13804 18116 13806
rect 16044 13468 16100 13524
rect 15596 12908 15652 12964
rect 15260 12684 15316 12740
rect 14008 12570 14064 12572
rect 14112 12570 14168 12572
rect 14008 12518 14024 12570
rect 14024 12518 14064 12570
rect 14112 12518 14148 12570
rect 14148 12518 14168 12570
rect 14008 12516 14064 12518
rect 14112 12516 14168 12518
rect 14216 12516 14272 12572
rect 14320 12570 14376 12572
rect 14424 12570 14480 12572
rect 14528 12570 14584 12572
rect 14320 12518 14324 12570
rect 14324 12518 14376 12570
rect 14424 12518 14448 12570
rect 14448 12518 14480 12570
rect 14528 12518 14572 12570
rect 14572 12518 14584 12570
rect 14320 12516 14376 12518
rect 14424 12516 14480 12518
rect 14528 12516 14584 12518
rect 14632 12570 14688 12572
rect 14736 12570 14792 12572
rect 14840 12570 14896 12572
rect 14632 12518 14644 12570
rect 14644 12518 14688 12570
rect 14736 12518 14768 12570
rect 14768 12518 14792 12570
rect 14840 12518 14892 12570
rect 14892 12518 14896 12570
rect 14632 12516 14688 12518
rect 14736 12516 14792 12518
rect 14840 12516 14896 12518
rect 14944 12516 15000 12572
rect 15048 12570 15104 12572
rect 15152 12570 15208 12572
rect 15048 12518 15068 12570
rect 15068 12518 15104 12570
rect 15152 12518 15192 12570
rect 15192 12518 15208 12570
rect 15048 12516 15104 12518
rect 15152 12516 15208 12518
rect 13916 11564 13972 11620
rect 14588 12348 14644 12404
rect 14588 11116 14644 11172
rect 14008 11002 14064 11004
rect 14112 11002 14168 11004
rect 14008 10950 14024 11002
rect 14024 10950 14064 11002
rect 14112 10950 14148 11002
rect 14148 10950 14168 11002
rect 14008 10948 14064 10950
rect 14112 10948 14168 10950
rect 14216 10948 14272 11004
rect 14320 11002 14376 11004
rect 14424 11002 14480 11004
rect 14528 11002 14584 11004
rect 14320 10950 14324 11002
rect 14324 10950 14376 11002
rect 14424 10950 14448 11002
rect 14448 10950 14480 11002
rect 14528 10950 14572 11002
rect 14572 10950 14584 11002
rect 14320 10948 14376 10950
rect 14424 10948 14480 10950
rect 14528 10948 14584 10950
rect 14632 11002 14688 11004
rect 14736 11002 14792 11004
rect 14840 11002 14896 11004
rect 14632 10950 14644 11002
rect 14644 10950 14688 11002
rect 14736 10950 14768 11002
rect 14768 10950 14792 11002
rect 14840 10950 14892 11002
rect 14892 10950 14896 11002
rect 14632 10948 14688 10950
rect 14736 10948 14792 10950
rect 14840 10948 14896 10950
rect 14944 10948 15000 11004
rect 15048 11002 15104 11004
rect 15152 11002 15208 11004
rect 15048 10950 15068 11002
rect 15068 10950 15104 11002
rect 15152 10950 15192 11002
rect 15192 10950 15208 11002
rect 15048 10948 15104 10950
rect 15152 10948 15208 10950
rect 14588 10834 14644 10836
rect 14588 10782 14590 10834
rect 14590 10782 14642 10834
rect 14642 10782 14644 10834
rect 14588 10780 14644 10782
rect 15148 10780 15204 10836
rect 15820 13132 15876 13188
rect 16380 12962 16436 12964
rect 16380 12910 16382 12962
rect 16382 12910 16434 12962
rect 16434 12910 16436 12962
rect 16380 12908 16436 12910
rect 15484 11788 15540 11844
rect 15596 12738 15652 12740
rect 15596 12686 15598 12738
rect 15598 12686 15650 12738
rect 15650 12686 15652 12738
rect 15596 12684 15652 12686
rect 18956 14418 19012 14420
rect 18956 14366 18958 14418
rect 18958 14366 19010 14418
rect 19010 14366 19012 14418
rect 18956 14364 19012 14366
rect 20636 14588 20692 14644
rect 19516 14306 19572 14308
rect 19516 14254 19518 14306
rect 19518 14254 19570 14306
rect 19570 14254 19572 14306
rect 19516 14252 19572 14254
rect 20972 14252 21028 14308
rect 20188 13858 20244 13860
rect 20188 13806 20190 13858
rect 20190 13806 20242 13858
rect 20242 13806 20244 13858
rect 20188 13804 20244 13806
rect 21196 13858 21252 13860
rect 21196 13806 21198 13858
rect 21198 13806 21250 13858
rect 21250 13806 21252 13858
rect 21196 13804 21252 13806
rect 19180 12738 19236 12740
rect 19180 12686 19182 12738
rect 19182 12686 19234 12738
rect 19234 12686 19236 12738
rect 19180 12684 19236 12686
rect 16716 12348 16772 12404
rect 17500 12402 17556 12404
rect 17500 12350 17502 12402
rect 17502 12350 17554 12402
rect 17554 12350 17556 12402
rect 17500 12348 17556 12350
rect 17948 12066 18004 12068
rect 17948 12014 17950 12066
rect 17950 12014 18002 12066
rect 18002 12014 18004 12066
rect 17948 12012 18004 12014
rect 16380 11228 16436 11284
rect 20300 12738 20356 12740
rect 20300 12686 20302 12738
rect 20302 12686 20354 12738
rect 20354 12686 20356 12738
rect 20300 12684 20356 12686
rect 19852 12178 19908 12180
rect 19852 12126 19854 12178
rect 19854 12126 19906 12178
rect 19906 12126 19908 12178
rect 19852 12124 19908 12126
rect 19180 12012 19236 12068
rect 17836 11282 17892 11284
rect 17836 11230 17838 11282
rect 17838 11230 17890 11282
rect 17890 11230 17892 11282
rect 17836 11228 17892 11230
rect 15596 10332 15652 10388
rect 14008 9434 14064 9436
rect 14112 9434 14168 9436
rect 14008 9382 14024 9434
rect 14024 9382 14064 9434
rect 14112 9382 14148 9434
rect 14148 9382 14168 9434
rect 14008 9380 14064 9382
rect 14112 9380 14168 9382
rect 14216 9380 14272 9436
rect 14320 9434 14376 9436
rect 14424 9434 14480 9436
rect 14528 9434 14584 9436
rect 14320 9382 14324 9434
rect 14324 9382 14376 9434
rect 14424 9382 14448 9434
rect 14448 9382 14480 9434
rect 14528 9382 14572 9434
rect 14572 9382 14584 9434
rect 14320 9380 14376 9382
rect 14424 9380 14480 9382
rect 14528 9380 14584 9382
rect 14632 9434 14688 9436
rect 14736 9434 14792 9436
rect 14840 9434 14896 9436
rect 14632 9382 14644 9434
rect 14644 9382 14688 9434
rect 14736 9382 14768 9434
rect 14768 9382 14792 9434
rect 14840 9382 14892 9434
rect 14892 9382 14896 9434
rect 14632 9380 14688 9382
rect 14736 9380 14792 9382
rect 14840 9380 14896 9382
rect 14944 9380 15000 9436
rect 15048 9434 15104 9436
rect 15152 9434 15208 9436
rect 15048 9382 15068 9434
rect 15068 9382 15104 9434
rect 15152 9382 15192 9434
rect 15192 9382 15208 9434
rect 15048 9380 15104 9382
rect 15152 9380 15208 9382
rect 14008 7866 14064 7868
rect 14112 7866 14168 7868
rect 14008 7814 14024 7866
rect 14024 7814 14064 7866
rect 14112 7814 14148 7866
rect 14148 7814 14168 7866
rect 14008 7812 14064 7814
rect 14112 7812 14168 7814
rect 14216 7812 14272 7868
rect 14320 7866 14376 7868
rect 14424 7866 14480 7868
rect 14528 7866 14584 7868
rect 14320 7814 14324 7866
rect 14324 7814 14376 7866
rect 14424 7814 14448 7866
rect 14448 7814 14480 7866
rect 14528 7814 14572 7866
rect 14572 7814 14584 7866
rect 14320 7812 14376 7814
rect 14424 7812 14480 7814
rect 14528 7812 14584 7814
rect 14632 7866 14688 7868
rect 14736 7866 14792 7868
rect 14840 7866 14896 7868
rect 14632 7814 14644 7866
rect 14644 7814 14688 7866
rect 14736 7814 14768 7866
rect 14768 7814 14792 7866
rect 14840 7814 14892 7866
rect 14892 7814 14896 7866
rect 14632 7812 14688 7814
rect 14736 7812 14792 7814
rect 14840 7812 14896 7814
rect 14944 7812 15000 7868
rect 15048 7866 15104 7868
rect 15152 7866 15208 7868
rect 15048 7814 15068 7866
rect 15068 7814 15104 7866
rect 15152 7814 15192 7866
rect 15192 7814 15208 7866
rect 15048 7812 15104 7814
rect 15152 7812 15208 7814
rect 17052 11170 17108 11172
rect 17052 11118 17054 11170
rect 17054 11118 17106 11170
rect 17106 11118 17108 11170
rect 17052 11116 17108 11118
rect 19740 10668 19796 10724
rect 21420 17052 21476 17108
rect 22428 18060 22484 18116
rect 22316 17666 22372 17668
rect 22316 17614 22318 17666
rect 22318 17614 22370 17666
rect 22370 17614 22372 17666
rect 22316 17612 22372 17614
rect 21868 17500 21924 17556
rect 22204 17052 22260 17108
rect 22428 17276 22484 17332
rect 23660 20018 23716 20020
rect 23660 19966 23662 20018
rect 23662 19966 23714 20018
rect 23714 19966 23716 20018
rect 23660 19964 23716 19966
rect 23548 19906 23604 19908
rect 23548 19854 23550 19906
rect 23550 19854 23602 19906
rect 23602 19854 23604 19906
rect 23548 19852 23604 19854
rect 23772 19740 23828 19796
rect 24668 20860 24724 20916
rect 24556 20802 24612 20804
rect 24556 20750 24558 20802
rect 24558 20750 24610 20802
rect 24610 20750 24612 20802
rect 24556 20748 24612 20750
rect 25228 20860 25284 20916
rect 24780 20636 24836 20692
rect 25340 20188 25396 20244
rect 26348 27132 26404 27188
rect 25676 26124 25732 26180
rect 29708 27074 29764 27076
rect 29708 27022 29710 27074
rect 29710 27022 29762 27074
rect 29762 27022 29764 27074
rect 29708 27020 29764 27022
rect 31388 35644 31444 35700
rect 30828 35308 30884 35364
rect 31164 35420 31220 35476
rect 31724 38050 31780 38052
rect 31724 37998 31726 38050
rect 31726 37998 31778 38050
rect 31778 37998 31780 38050
rect 31724 37996 31780 37998
rect 31724 37212 31780 37268
rect 32284 39004 32340 39060
rect 32396 38946 32452 38948
rect 32396 38894 32398 38946
rect 32398 38894 32450 38946
rect 32450 38894 32452 38946
rect 32396 38892 32452 38894
rect 32060 38220 32116 38276
rect 31948 38108 32004 38164
rect 31948 37548 32004 37604
rect 32172 36540 32228 36596
rect 32620 38834 32676 38836
rect 32620 38782 32622 38834
rect 32622 38782 32674 38834
rect 32674 38782 32676 38834
rect 32620 38780 32676 38782
rect 32620 37996 32676 38052
rect 32508 37212 32564 37268
rect 32396 36876 32452 36932
rect 31724 36370 31780 36372
rect 31724 36318 31726 36370
rect 31726 36318 31778 36370
rect 31778 36318 31780 36370
rect 31724 36316 31780 36318
rect 31724 36092 31780 36148
rect 31724 35420 31780 35476
rect 31836 35756 31892 35812
rect 32172 36092 32228 36148
rect 32396 35868 32452 35924
rect 31612 35308 31668 35364
rect 31948 35420 32004 35476
rect 32172 35420 32228 35476
rect 30940 32956 30996 33012
rect 31388 33516 31444 33572
rect 31164 32786 31220 32788
rect 31164 32734 31166 32786
rect 31166 32734 31218 32786
rect 31218 32734 31220 32786
rect 31164 32732 31220 32734
rect 31388 32620 31444 32676
rect 30380 31388 30436 31444
rect 30492 31106 30548 31108
rect 30492 31054 30494 31106
rect 30494 31054 30546 31106
rect 30546 31054 30548 31106
rect 30492 31052 30548 31054
rect 31948 33516 32004 33572
rect 31612 32956 31668 33012
rect 31612 31500 31668 31556
rect 30268 30268 30324 30324
rect 30268 29372 30324 29428
rect 30044 27970 30100 27972
rect 30044 27918 30046 27970
rect 30046 27918 30098 27970
rect 30098 27918 30100 27970
rect 30044 27916 30100 27918
rect 30156 27634 30212 27636
rect 30156 27582 30158 27634
rect 30158 27582 30210 27634
rect 30210 27582 30212 27634
rect 30156 27580 30212 27582
rect 30156 27020 30212 27076
rect 29260 26178 29316 26180
rect 29260 26126 29262 26178
rect 29262 26126 29314 26178
rect 29314 26126 29316 26178
rect 29260 26124 29316 26126
rect 29820 26850 29876 26852
rect 29820 26798 29822 26850
rect 29822 26798 29874 26850
rect 29874 26798 29876 26850
rect 29820 26796 29876 26798
rect 29596 26236 29652 26292
rect 26796 25116 26852 25172
rect 26684 25004 26740 25060
rect 26012 24780 26068 24836
rect 25788 24610 25844 24612
rect 25788 24558 25790 24610
rect 25790 24558 25842 24610
rect 25842 24558 25844 24610
rect 25788 24556 25844 24558
rect 26012 24108 26068 24164
rect 26348 22092 26404 22148
rect 26684 24444 26740 24500
rect 26684 23660 26740 23716
rect 26460 21980 26516 22036
rect 27020 25116 27076 25172
rect 27356 25676 27412 25732
rect 27132 24892 27188 24948
rect 27244 24780 27300 24836
rect 29372 25564 29428 25620
rect 27468 25228 27524 25284
rect 27580 25340 27636 25396
rect 27244 23996 27300 24052
rect 27020 23884 27076 23940
rect 27020 23660 27076 23716
rect 27916 25394 27972 25396
rect 27916 25342 27918 25394
rect 27918 25342 27970 25394
rect 27970 25342 27972 25394
rect 27916 25340 27972 25342
rect 28252 25282 28308 25284
rect 28252 25230 28254 25282
rect 28254 25230 28306 25282
rect 28306 25230 28308 25282
rect 28252 25228 28308 25230
rect 27804 24722 27860 24724
rect 27804 24670 27806 24722
rect 27806 24670 27858 24722
rect 27858 24670 27860 24722
rect 27804 24668 27860 24670
rect 27916 24610 27972 24612
rect 27916 24558 27918 24610
rect 27918 24558 27970 24610
rect 27970 24558 27972 24610
rect 27916 24556 27972 24558
rect 27916 23996 27972 24052
rect 27580 23324 27636 23380
rect 27804 23548 27860 23604
rect 26908 22540 26964 22596
rect 27580 22540 27636 22596
rect 26796 21756 26852 21812
rect 27020 22092 27076 22148
rect 25788 20972 25844 21028
rect 25676 20860 25732 20916
rect 25452 20076 25508 20132
rect 25564 19964 25620 20020
rect 24008 19626 24064 19628
rect 24112 19626 24168 19628
rect 24008 19574 24024 19626
rect 24024 19574 24064 19626
rect 24112 19574 24148 19626
rect 24148 19574 24168 19626
rect 24008 19572 24064 19574
rect 24112 19572 24168 19574
rect 24216 19572 24272 19628
rect 24320 19626 24376 19628
rect 24424 19626 24480 19628
rect 24528 19626 24584 19628
rect 24320 19574 24324 19626
rect 24324 19574 24376 19626
rect 24424 19574 24448 19626
rect 24448 19574 24480 19626
rect 24528 19574 24572 19626
rect 24572 19574 24584 19626
rect 24320 19572 24376 19574
rect 24424 19572 24480 19574
rect 24528 19572 24584 19574
rect 24632 19626 24688 19628
rect 24736 19626 24792 19628
rect 24840 19626 24896 19628
rect 24632 19574 24644 19626
rect 24644 19574 24688 19626
rect 24736 19574 24768 19626
rect 24768 19574 24792 19626
rect 24840 19574 24892 19626
rect 24892 19574 24896 19626
rect 24632 19572 24688 19574
rect 24736 19572 24792 19574
rect 24840 19572 24896 19574
rect 24944 19572 25000 19628
rect 25048 19626 25104 19628
rect 25152 19626 25208 19628
rect 25048 19574 25068 19626
rect 25068 19574 25104 19626
rect 25152 19574 25192 19626
rect 25192 19574 25208 19626
rect 25048 19572 25104 19574
rect 25152 19572 25208 19574
rect 25676 19628 25732 19684
rect 25116 19234 25172 19236
rect 25116 19182 25118 19234
rect 25118 19182 25170 19234
rect 25170 19182 25172 19234
rect 25116 19180 25172 19182
rect 22652 18172 22708 18228
rect 23212 18060 23268 18116
rect 23772 18620 23828 18676
rect 23100 17612 23156 17668
rect 22764 17554 22820 17556
rect 22764 17502 22766 17554
rect 22766 17502 22818 17554
rect 22818 17502 22820 17554
rect 22764 17500 22820 17502
rect 23324 17164 23380 17220
rect 23548 17388 23604 17444
rect 22540 16940 22596 16996
rect 21644 16828 21700 16884
rect 21644 15932 21700 15988
rect 23212 16994 23268 16996
rect 23212 16942 23214 16994
rect 23214 16942 23266 16994
rect 23266 16942 23268 16994
rect 23212 16940 23268 16942
rect 22652 16828 22708 16884
rect 23324 16882 23380 16884
rect 23324 16830 23326 16882
rect 23326 16830 23378 16882
rect 23378 16830 23380 16882
rect 23324 16828 23380 16830
rect 22316 16770 22372 16772
rect 22316 16718 22318 16770
rect 22318 16718 22370 16770
rect 22370 16718 22372 16770
rect 22316 16716 22372 16718
rect 25788 18620 25844 18676
rect 24008 18058 24064 18060
rect 24112 18058 24168 18060
rect 24008 18006 24024 18058
rect 24024 18006 24064 18058
rect 24112 18006 24148 18058
rect 24148 18006 24168 18058
rect 24008 18004 24064 18006
rect 24112 18004 24168 18006
rect 24216 18004 24272 18060
rect 24320 18058 24376 18060
rect 24424 18058 24480 18060
rect 24528 18058 24584 18060
rect 24320 18006 24324 18058
rect 24324 18006 24376 18058
rect 24424 18006 24448 18058
rect 24448 18006 24480 18058
rect 24528 18006 24572 18058
rect 24572 18006 24584 18058
rect 24320 18004 24376 18006
rect 24424 18004 24480 18006
rect 24528 18004 24584 18006
rect 24632 18058 24688 18060
rect 24736 18058 24792 18060
rect 24840 18058 24896 18060
rect 24632 18006 24644 18058
rect 24644 18006 24688 18058
rect 24736 18006 24768 18058
rect 24768 18006 24792 18058
rect 24840 18006 24892 18058
rect 24892 18006 24896 18058
rect 24632 18004 24688 18006
rect 24736 18004 24792 18006
rect 24840 18004 24896 18006
rect 24944 18004 25000 18060
rect 25048 18058 25104 18060
rect 25152 18058 25208 18060
rect 25048 18006 25068 18058
rect 25068 18006 25104 18058
rect 25152 18006 25192 18058
rect 25192 18006 25208 18058
rect 25048 18004 25104 18006
rect 25152 18004 25208 18006
rect 23660 16994 23716 16996
rect 23660 16942 23662 16994
rect 23662 16942 23714 16994
rect 23714 16942 23716 16994
rect 23660 16940 23716 16942
rect 23884 17276 23940 17332
rect 24892 17442 24948 17444
rect 24892 17390 24894 17442
rect 24894 17390 24946 17442
rect 24946 17390 24948 17442
rect 24892 17388 24948 17390
rect 24220 17164 24276 17220
rect 24108 17106 24164 17108
rect 24108 17054 24110 17106
rect 24110 17054 24162 17106
rect 24162 17054 24164 17106
rect 24108 17052 24164 17054
rect 23772 16828 23828 16884
rect 25228 17164 25284 17220
rect 23772 16658 23828 16660
rect 23772 16606 23774 16658
rect 23774 16606 23826 16658
rect 23826 16606 23828 16658
rect 23772 16604 23828 16606
rect 22204 15484 22260 15540
rect 22652 15874 22708 15876
rect 22652 15822 22654 15874
rect 22654 15822 22706 15874
rect 22706 15822 22708 15874
rect 22652 15820 22708 15822
rect 22316 15260 22372 15316
rect 22988 15484 23044 15540
rect 21756 15148 21812 15204
rect 22204 15202 22260 15204
rect 22204 15150 22206 15202
rect 22206 15150 22258 15202
rect 22258 15150 22260 15202
rect 22204 15148 22260 15150
rect 21980 14642 22036 14644
rect 21980 14590 21982 14642
rect 21982 14590 22034 14642
rect 22034 14590 22036 14642
rect 21980 14588 22036 14590
rect 21756 12908 21812 12964
rect 21308 12684 21364 12740
rect 22428 13804 22484 13860
rect 22428 13074 22484 13076
rect 22428 13022 22430 13074
rect 22430 13022 22482 13074
rect 22482 13022 22484 13074
rect 22428 13020 22484 13022
rect 24008 16490 24064 16492
rect 24112 16490 24168 16492
rect 24008 16438 24024 16490
rect 24024 16438 24064 16490
rect 24112 16438 24148 16490
rect 24148 16438 24168 16490
rect 24008 16436 24064 16438
rect 24112 16436 24168 16438
rect 24216 16436 24272 16492
rect 24320 16490 24376 16492
rect 24424 16490 24480 16492
rect 24528 16490 24584 16492
rect 24320 16438 24324 16490
rect 24324 16438 24376 16490
rect 24424 16438 24448 16490
rect 24448 16438 24480 16490
rect 24528 16438 24572 16490
rect 24572 16438 24584 16490
rect 24320 16436 24376 16438
rect 24424 16436 24480 16438
rect 24528 16436 24584 16438
rect 24632 16490 24688 16492
rect 24736 16490 24792 16492
rect 24840 16490 24896 16492
rect 24632 16438 24644 16490
rect 24644 16438 24688 16490
rect 24736 16438 24768 16490
rect 24768 16438 24792 16490
rect 24840 16438 24892 16490
rect 24892 16438 24896 16490
rect 24632 16436 24688 16438
rect 24736 16436 24792 16438
rect 24840 16436 24896 16438
rect 24944 16436 25000 16492
rect 25048 16490 25104 16492
rect 25152 16490 25208 16492
rect 25048 16438 25068 16490
rect 25068 16438 25104 16490
rect 25152 16438 25192 16490
rect 25192 16438 25208 16490
rect 25048 16436 25104 16438
rect 25152 16436 25208 16438
rect 26908 19458 26964 19460
rect 26908 19406 26910 19458
rect 26910 19406 26962 19458
rect 26962 19406 26964 19458
rect 26908 19404 26964 19406
rect 26460 19122 26516 19124
rect 26460 19070 26462 19122
rect 26462 19070 26514 19122
rect 26514 19070 26516 19122
rect 26460 19068 26516 19070
rect 26348 18508 26404 18564
rect 26236 17500 26292 17556
rect 25452 16882 25508 16884
rect 25452 16830 25454 16882
rect 25454 16830 25506 16882
rect 25506 16830 25508 16882
rect 25452 16828 25508 16830
rect 25788 16268 25844 16324
rect 24556 16156 24612 16212
rect 23884 15820 23940 15876
rect 25116 15986 25172 15988
rect 25116 15934 25118 15986
rect 25118 15934 25170 15986
rect 25170 15934 25172 15986
rect 25116 15932 25172 15934
rect 23212 14588 23268 14644
rect 23772 14924 23828 14980
rect 24220 15036 24276 15092
rect 25340 15874 25396 15876
rect 25340 15822 25342 15874
rect 25342 15822 25394 15874
rect 25394 15822 25396 15874
rect 25340 15820 25396 15822
rect 25564 15314 25620 15316
rect 25564 15262 25566 15314
rect 25566 15262 25618 15314
rect 25618 15262 25620 15314
rect 25564 15260 25620 15262
rect 24444 15036 24500 15092
rect 24008 14922 24064 14924
rect 24112 14922 24168 14924
rect 24008 14870 24024 14922
rect 24024 14870 24064 14922
rect 24112 14870 24148 14922
rect 24148 14870 24168 14922
rect 24008 14868 24064 14870
rect 24112 14868 24168 14870
rect 24216 14868 24272 14924
rect 24320 14922 24376 14924
rect 24424 14922 24480 14924
rect 24528 14922 24584 14924
rect 24320 14870 24324 14922
rect 24324 14870 24376 14922
rect 24424 14870 24448 14922
rect 24448 14870 24480 14922
rect 24528 14870 24572 14922
rect 24572 14870 24584 14922
rect 24320 14868 24376 14870
rect 24424 14868 24480 14870
rect 24528 14868 24584 14870
rect 24632 14922 24688 14924
rect 24736 14922 24792 14924
rect 24840 14922 24896 14924
rect 24632 14870 24644 14922
rect 24644 14870 24688 14922
rect 24736 14870 24768 14922
rect 24768 14870 24792 14922
rect 24840 14870 24892 14922
rect 24892 14870 24896 14922
rect 24632 14868 24688 14870
rect 24736 14868 24792 14870
rect 24840 14868 24896 14870
rect 24944 14868 25000 14924
rect 25048 14922 25104 14924
rect 25152 14922 25208 14924
rect 25048 14870 25068 14922
rect 25068 14870 25104 14922
rect 25152 14870 25192 14922
rect 25192 14870 25208 14922
rect 25048 14868 25104 14870
rect 25152 14868 25208 14870
rect 24668 13692 24724 13748
rect 26124 13580 26180 13636
rect 24008 13354 24064 13356
rect 24112 13354 24168 13356
rect 24008 13302 24024 13354
rect 24024 13302 24064 13354
rect 24112 13302 24148 13354
rect 24148 13302 24168 13354
rect 24008 13300 24064 13302
rect 24112 13300 24168 13302
rect 24216 13300 24272 13356
rect 24320 13354 24376 13356
rect 24424 13354 24480 13356
rect 24528 13354 24584 13356
rect 24320 13302 24324 13354
rect 24324 13302 24376 13354
rect 24424 13302 24448 13354
rect 24448 13302 24480 13354
rect 24528 13302 24572 13354
rect 24572 13302 24584 13354
rect 24320 13300 24376 13302
rect 24424 13300 24480 13302
rect 24528 13300 24584 13302
rect 24632 13354 24688 13356
rect 24736 13354 24792 13356
rect 24840 13354 24896 13356
rect 24632 13302 24644 13354
rect 24644 13302 24688 13354
rect 24736 13302 24768 13354
rect 24768 13302 24792 13354
rect 24840 13302 24892 13354
rect 24892 13302 24896 13354
rect 24632 13300 24688 13302
rect 24736 13300 24792 13302
rect 24840 13300 24896 13302
rect 24944 13300 25000 13356
rect 25048 13354 25104 13356
rect 25152 13354 25208 13356
rect 25048 13302 25068 13354
rect 25068 13302 25104 13354
rect 25152 13302 25192 13354
rect 25192 13302 25208 13354
rect 25048 13300 25104 13302
rect 25152 13300 25208 13302
rect 23772 13132 23828 13188
rect 24556 13186 24612 13188
rect 24556 13134 24558 13186
rect 24558 13134 24610 13186
rect 24610 13134 24612 13186
rect 24556 13132 24612 13134
rect 23436 13020 23492 13076
rect 23212 12908 23268 12964
rect 22540 12124 22596 12180
rect 22540 10834 22596 10836
rect 22540 10782 22542 10834
rect 22542 10782 22594 10834
rect 22594 10782 22596 10834
rect 22540 10780 22596 10782
rect 24444 12962 24500 12964
rect 24444 12910 24446 12962
rect 24446 12910 24498 12962
rect 24498 12910 24500 12962
rect 24444 12908 24500 12910
rect 23996 12850 24052 12852
rect 23996 12798 23998 12850
rect 23998 12798 24050 12850
rect 24050 12798 24052 12850
rect 23996 12796 24052 12798
rect 26572 17164 26628 17220
rect 26796 18562 26852 18564
rect 26796 18510 26798 18562
rect 26798 18510 26850 18562
rect 26850 18510 26852 18562
rect 26796 18508 26852 18510
rect 26684 17052 26740 17108
rect 26796 17500 26852 17556
rect 27356 22428 27412 22484
rect 27356 22204 27412 22260
rect 27580 21980 27636 22036
rect 27692 21308 27748 21364
rect 27244 19628 27300 19684
rect 27356 20748 27412 20804
rect 27132 19234 27188 19236
rect 27132 19182 27134 19234
rect 27134 19182 27186 19234
rect 27186 19182 27188 19234
rect 27132 19180 27188 19182
rect 27468 19628 27524 19684
rect 27468 19180 27524 19236
rect 27804 19404 27860 19460
rect 28140 23884 28196 23940
rect 28812 25116 28868 25172
rect 28476 24946 28532 24948
rect 28476 24894 28478 24946
rect 28478 24894 28530 24946
rect 28530 24894 28532 24946
rect 28476 24892 28532 24894
rect 28812 24722 28868 24724
rect 28812 24670 28814 24722
rect 28814 24670 28866 24722
rect 28866 24670 28868 24722
rect 28812 24668 28868 24670
rect 29148 24892 29204 24948
rect 29708 25452 29764 25508
rect 29932 25004 29988 25060
rect 29484 24668 29540 24724
rect 29148 23884 29204 23940
rect 28140 23378 28196 23380
rect 28140 23326 28142 23378
rect 28142 23326 28194 23378
rect 28194 23326 28196 23378
rect 28140 23324 28196 23326
rect 28140 22594 28196 22596
rect 28140 22542 28142 22594
rect 28142 22542 28194 22594
rect 28194 22542 28196 22594
rect 28140 22540 28196 22542
rect 29596 24556 29652 24612
rect 29484 23996 29540 24052
rect 29372 23548 29428 23604
rect 29708 23714 29764 23716
rect 29708 23662 29710 23714
rect 29710 23662 29762 23714
rect 29762 23662 29764 23714
rect 29708 23660 29764 23662
rect 29596 23324 29652 23380
rect 29484 22482 29540 22484
rect 29484 22430 29486 22482
rect 29486 22430 29538 22482
rect 29538 22430 29540 22482
rect 29484 22428 29540 22430
rect 28588 21868 28644 21924
rect 28924 22316 28980 22372
rect 29708 22204 29764 22260
rect 29260 22146 29316 22148
rect 29260 22094 29262 22146
rect 29262 22094 29314 22146
rect 29314 22094 29316 22146
rect 29260 22092 29316 22094
rect 29148 21756 29204 21812
rect 28588 20860 28644 20916
rect 28252 20802 28308 20804
rect 28252 20750 28254 20802
rect 28254 20750 28306 20802
rect 28306 20750 28308 20802
rect 28252 20748 28308 20750
rect 28028 19964 28084 20020
rect 29708 21980 29764 22036
rect 30156 25618 30212 25620
rect 30156 25566 30158 25618
rect 30158 25566 30210 25618
rect 30210 25566 30212 25618
rect 30156 25564 30212 25566
rect 31500 30210 31556 30212
rect 31500 30158 31502 30210
rect 31502 30158 31554 30210
rect 31554 30158 31556 30210
rect 31500 30156 31556 30158
rect 31836 33068 31892 33124
rect 31724 30828 31780 30884
rect 31836 30210 31892 30212
rect 31836 30158 31838 30210
rect 31838 30158 31890 30210
rect 31890 30158 31892 30210
rect 31836 30156 31892 30158
rect 31612 29708 31668 29764
rect 30940 29426 30996 29428
rect 30940 29374 30942 29426
rect 30942 29374 30994 29426
rect 30994 29374 30996 29426
rect 30940 29372 30996 29374
rect 31612 28588 31668 28644
rect 31388 28476 31444 28532
rect 31724 28364 31780 28420
rect 30828 27580 30884 27636
rect 30940 26796 30996 26852
rect 30268 25452 30324 25508
rect 30716 26236 30772 26292
rect 30604 26124 30660 26180
rect 30268 24556 30324 24612
rect 30044 22652 30100 22708
rect 29708 21420 29764 21476
rect 29484 20802 29540 20804
rect 29484 20750 29486 20802
rect 29486 20750 29538 20802
rect 29538 20750 29540 20802
rect 29484 20748 29540 20750
rect 29596 20636 29652 20692
rect 28476 19740 28532 19796
rect 28364 19234 28420 19236
rect 28364 19182 28366 19234
rect 28366 19182 28418 19234
rect 28418 19182 28420 19234
rect 28364 19180 28420 19182
rect 29148 19234 29204 19236
rect 29148 19182 29150 19234
rect 29150 19182 29202 19234
rect 29202 19182 29204 19234
rect 29148 19180 29204 19182
rect 28476 19068 28532 19124
rect 27132 18620 27188 18676
rect 27916 18674 27972 18676
rect 27916 18622 27918 18674
rect 27918 18622 27970 18674
rect 27970 18622 27972 18674
rect 27916 18620 27972 18622
rect 28140 18620 28196 18676
rect 29708 20524 29764 20580
rect 29820 19906 29876 19908
rect 29820 19854 29822 19906
rect 29822 19854 29874 19906
rect 29874 19854 29876 19906
rect 29820 19852 29876 19854
rect 30492 24668 30548 24724
rect 30716 25506 30772 25508
rect 30716 25454 30718 25506
rect 30718 25454 30770 25506
rect 30770 25454 30772 25506
rect 30716 25452 30772 25454
rect 31388 25228 31444 25284
rect 30604 24162 30660 24164
rect 30604 24110 30606 24162
rect 30606 24110 30658 24162
rect 30658 24110 30660 24162
rect 30604 24108 30660 24110
rect 30268 23660 30324 23716
rect 30604 23324 30660 23380
rect 30492 22652 30548 22708
rect 30044 22258 30100 22260
rect 30044 22206 30046 22258
rect 30046 22206 30098 22258
rect 30098 22206 30100 22258
rect 30044 22204 30100 22206
rect 30156 22146 30212 22148
rect 30156 22094 30158 22146
rect 30158 22094 30210 22146
rect 30210 22094 30212 22146
rect 30156 22092 30212 22094
rect 29932 19740 29988 19796
rect 31052 24050 31108 24052
rect 31052 23998 31054 24050
rect 31054 23998 31106 24050
rect 31106 23998 31108 24050
rect 31052 23996 31108 23998
rect 32508 35308 32564 35364
rect 32396 34802 32452 34804
rect 32396 34750 32398 34802
rect 32398 34750 32450 34802
rect 32450 34750 32452 34802
rect 32396 34748 32452 34750
rect 35308 44044 35364 44100
rect 34008 43930 34064 43932
rect 34112 43930 34168 43932
rect 34008 43878 34024 43930
rect 34024 43878 34064 43930
rect 34112 43878 34148 43930
rect 34148 43878 34168 43930
rect 34008 43876 34064 43878
rect 34112 43876 34168 43878
rect 34216 43876 34272 43932
rect 34320 43930 34376 43932
rect 34424 43930 34480 43932
rect 34528 43930 34584 43932
rect 34320 43878 34324 43930
rect 34324 43878 34376 43930
rect 34424 43878 34448 43930
rect 34448 43878 34480 43930
rect 34528 43878 34572 43930
rect 34572 43878 34584 43930
rect 34320 43876 34376 43878
rect 34424 43876 34480 43878
rect 34528 43876 34584 43878
rect 34632 43930 34688 43932
rect 34736 43930 34792 43932
rect 34840 43930 34896 43932
rect 34632 43878 34644 43930
rect 34644 43878 34688 43930
rect 34736 43878 34768 43930
rect 34768 43878 34792 43930
rect 34840 43878 34892 43930
rect 34892 43878 34896 43930
rect 34632 43876 34688 43878
rect 34736 43876 34792 43878
rect 34840 43876 34896 43878
rect 34944 43876 35000 43932
rect 35048 43930 35104 43932
rect 35152 43930 35208 43932
rect 35048 43878 35068 43930
rect 35068 43878 35104 43930
rect 35152 43878 35192 43930
rect 35192 43878 35208 43930
rect 35048 43876 35104 43878
rect 35152 43876 35208 43878
rect 35980 45164 36036 45220
rect 37100 46674 37156 46676
rect 37100 46622 37102 46674
rect 37102 46622 37154 46674
rect 37154 46622 37156 46674
rect 37100 46620 37156 46622
rect 37884 46620 37940 46676
rect 37548 46396 37604 46452
rect 37996 46284 38052 46340
rect 37100 45890 37156 45892
rect 37100 45838 37102 45890
rect 37102 45838 37154 45890
rect 37154 45838 37156 45890
rect 37100 45836 37156 45838
rect 36988 45778 37044 45780
rect 36988 45726 36990 45778
rect 36990 45726 37042 45778
rect 37042 45726 37044 45778
rect 36988 45724 37044 45726
rect 35980 44828 36036 44884
rect 35868 44268 35924 44324
rect 34636 43426 34692 43428
rect 34636 43374 34638 43426
rect 34638 43374 34690 43426
rect 34690 43374 34692 43426
rect 34636 43372 34692 43374
rect 33852 43036 33908 43092
rect 34300 42812 34356 42868
rect 33740 42700 33796 42756
rect 33964 42700 34020 42756
rect 33628 42588 33684 42644
rect 33180 42140 33236 42196
rect 33516 42476 33572 42532
rect 33180 41580 33236 41636
rect 33292 41356 33348 41412
rect 32844 40572 32900 40628
rect 33180 40908 33236 40964
rect 33068 40402 33124 40404
rect 33068 40350 33070 40402
rect 33070 40350 33122 40402
rect 33122 40350 33124 40402
rect 33068 40348 33124 40350
rect 34972 42812 35028 42868
rect 34412 42754 34468 42756
rect 34412 42702 34414 42754
rect 34414 42702 34466 42754
rect 34466 42702 34468 42754
rect 34412 42700 34468 42702
rect 35084 42642 35140 42644
rect 35084 42590 35086 42642
rect 35086 42590 35138 42642
rect 35138 42590 35140 42642
rect 35084 42588 35140 42590
rect 36428 43650 36484 43652
rect 36428 43598 36430 43650
rect 36430 43598 36482 43650
rect 36482 43598 36484 43650
rect 36428 43596 36484 43598
rect 36316 42700 36372 42756
rect 36428 42642 36484 42644
rect 36428 42590 36430 42642
rect 36430 42590 36482 42642
rect 36482 42590 36484 42642
rect 36428 42588 36484 42590
rect 34008 42362 34064 42364
rect 34112 42362 34168 42364
rect 34008 42310 34024 42362
rect 34024 42310 34064 42362
rect 34112 42310 34148 42362
rect 34148 42310 34168 42362
rect 34008 42308 34064 42310
rect 34112 42308 34168 42310
rect 34216 42308 34272 42364
rect 34320 42362 34376 42364
rect 34424 42362 34480 42364
rect 34528 42362 34584 42364
rect 34320 42310 34324 42362
rect 34324 42310 34376 42362
rect 34424 42310 34448 42362
rect 34448 42310 34480 42362
rect 34528 42310 34572 42362
rect 34572 42310 34584 42362
rect 34320 42308 34376 42310
rect 34424 42308 34480 42310
rect 34528 42308 34584 42310
rect 34632 42362 34688 42364
rect 34736 42362 34792 42364
rect 34840 42362 34896 42364
rect 34632 42310 34644 42362
rect 34644 42310 34688 42362
rect 34736 42310 34768 42362
rect 34768 42310 34792 42362
rect 34840 42310 34892 42362
rect 34892 42310 34896 42362
rect 34632 42308 34688 42310
rect 34736 42308 34792 42310
rect 34840 42308 34896 42310
rect 34944 42308 35000 42364
rect 35048 42362 35104 42364
rect 35152 42362 35208 42364
rect 35048 42310 35068 42362
rect 35068 42310 35104 42362
rect 35152 42310 35192 42362
rect 35192 42310 35208 42362
rect 35048 42308 35104 42310
rect 35152 42308 35208 42310
rect 35196 42028 35252 42084
rect 33964 41916 34020 41972
rect 33852 41580 33908 41636
rect 35084 41970 35140 41972
rect 35084 41918 35086 41970
rect 35086 41918 35138 41970
rect 35138 41918 35140 41970
rect 35084 41916 35140 41918
rect 34748 41020 34804 41076
rect 36092 42476 36148 42532
rect 35532 42140 35588 42196
rect 35308 41916 35364 41972
rect 35756 41804 35812 41860
rect 35308 41186 35364 41188
rect 35308 41134 35310 41186
rect 35310 41134 35362 41186
rect 35362 41134 35364 41186
rect 35308 41132 35364 41134
rect 34008 40794 34064 40796
rect 34112 40794 34168 40796
rect 34008 40742 34024 40794
rect 34024 40742 34064 40794
rect 34112 40742 34148 40794
rect 34148 40742 34168 40794
rect 34008 40740 34064 40742
rect 34112 40740 34168 40742
rect 34216 40740 34272 40796
rect 34320 40794 34376 40796
rect 34424 40794 34480 40796
rect 34528 40794 34584 40796
rect 34320 40742 34324 40794
rect 34324 40742 34376 40794
rect 34424 40742 34448 40794
rect 34448 40742 34480 40794
rect 34528 40742 34572 40794
rect 34572 40742 34584 40794
rect 34320 40740 34376 40742
rect 34424 40740 34480 40742
rect 34528 40740 34584 40742
rect 34632 40794 34688 40796
rect 34736 40794 34792 40796
rect 34840 40794 34896 40796
rect 34632 40742 34644 40794
rect 34644 40742 34688 40794
rect 34736 40742 34768 40794
rect 34768 40742 34792 40794
rect 34840 40742 34892 40794
rect 34892 40742 34896 40794
rect 34632 40740 34688 40742
rect 34736 40740 34792 40742
rect 34840 40740 34896 40742
rect 34944 40740 35000 40796
rect 35048 40794 35104 40796
rect 35152 40794 35208 40796
rect 35048 40742 35068 40794
rect 35068 40742 35104 40794
rect 35152 40742 35192 40794
rect 35192 40742 35208 40794
rect 35048 40740 35104 40742
rect 35152 40740 35208 40742
rect 33292 40460 33348 40516
rect 33292 40290 33348 40292
rect 33292 40238 33294 40290
rect 33294 40238 33346 40290
rect 33346 40238 33348 40290
rect 33292 40236 33348 40238
rect 33404 40124 33460 40180
rect 33628 40626 33684 40628
rect 33628 40574 33630 40626
rect 33630 40574 33682 40626
rect 33682 40574 33684 40626
rect 33628 40572 33684 40574
rect 33964 40572 34020 40628
rect 33516 39788 33572 39844
rect 33516 38668 33572 38724
rect 34076 40514 34132 40516
rect 34076 40462 34078 40514
rect 34078 40462 34130 40514
rect 34130 40462 34132 40514
rect 34076 40460 34132 40462
rect 33964 39788 34020 39844
rect 34636 39730 34692 39732
rect 34636 39678 34638 39730
rect 34638 39678 34690 39730
rect 34690 39678 34692 39730
rect 34636 39676 34692 39678
rect 34008 39226 34064 39228
rect 34112 39226 34168 39228
rect 34008 39174 34024 39226
rect 34024 39174 34064 39226
rect 34112 39174 34148 39226
rect 34148 39174 34168 39226
rect 34008 39172 34064 39174
rect 34112 39172 34168 39174
rect 34216 39172 34272 39228
rect 34320 39226 34376 39228
rect 34424 39226 34480 39228
rect 34528 39226 34584 39228
rect 34320 39174 34324 39226
rect 34324 39174 34376 39226
rect 34424 39174 34448 39226
rect 34448 39174 34480 39226
rect 34528 39174 34572 39226
rect 34572 39174 34584 39226
rect 34320 39172 34376 39174
rect 34424 39172 34480 39174
rect 34528 39172 34584 39174
rect 34632 39226 34688 39228
rect 34736 39226 34792 39228
rect 34840 39226 34896 39228
rect 34632 39174 34644 39226
rect 34644 39174 34688 39226
rect 34736 39174 34768 39226
rect 34768 39174 34792 39226
rect 34840 39174 34892 39226
rect 34892 39174 34896 39226
rect 34632 39172 34688 39174
rect 34736 39172 34792 39174
rect 34840 39172 34896 39174
rect 34944 39172 35000 39228
rect 35048 39226 35104 39228
rect 35152 39226 35208 39228
rect 35048 39174 35068 39226
rect 35068 39174 35104 39226
rect 35152 39174 35192 39226
rect 35192 39174 35208 39226
rect 35048 39172 35104 39174
rect 35152 39172 35208 39174
rect 33740 39058 33796 39060
rect 33740 39006 33742 39058
rect 33742 39006 33794 39058
rect 33794 39006 33796 39058
rect 33740 39004 33796 39006
rect 34300 39058 34356 39060
rect 34300 39006 34302 39058
rect 34302 39006 34354 39058
rect 34354 39006 34356 39058
rect 34300 39004 34356 39006
rect 34188 38946 34244 38948
rect 34188 38894 34190 38946
rect 34190 38894 34242 38946
rect 34242 38894 34244 38946
rect 34188 38892 34244 38894
rect 34972 38892 35028 38948
rect 34748 38834 34804 38836
rect 34748 38782 34750 38834
rect 34750 38782 34802 38834
rect 34802 38782 34804 38834
rect 34748 38780 34804 38782
rect 33068 36876 33124 36932
rect 33516 37324 33572 37380
rect 33740 38162 33796 38164
rect 33740 38110 33742 38162
rect 33742 38110 33794 38162
rect 33794 38110 33796 38162
rect 33740 38108 33796 38110
rect 34076 38108 34132 38164
rect 35196 38668 35252 38724
rect 35868 40962 35924 40964
rect 35868 40910 35870 40962
rect 35870 40910 35922 40962
rect 35922 40910 35924 40962
rect 35868 40908 35924 40910
rect 35644 40348 35700 40404
rect 35868 38668 35924 38724
rect 36316 39788 36372 39844
rect 33628 37100 33684 37156
rect 33740 36876 33796 36932
rect 33852 37660 33908 37716
rect 33292 36594 33348 36596
rect 33292 36542 33294 36594
rect 33294 36542 33346 36594
rect 33346 36542 33348 36594
rect 33292 36540 33348 36542
rect 33068 36092 33124 36148
rect 33740 35868 33796 35924
rect 33068 35810 33124 35812
rect 33068 35758 33070 35810
rect 33070 35758 33122 35810
rect 33122 35758 33124 35810
rect 33068 35756 33124 35758
rect 32844 35420 32900 35476
rect 33628 35698 33684 35700
rect 33628 35646 33630 35698
rect 33630 35646 33682 35698
rect 33682 35646 33684 35698
rect 33628 35644 33684 35646
rect 33068 34636 33124 34692
rect 32508 34242 32564 34244
rect 32508 34190 32510 34242
rect 32510 34190 32562 34242
rect 32562 34190 32564 34242
rect 32508 34188 32564 34190
rect 32172 33068 32228 33124
rect 32956 33516 33012 33572
rect 32844 33292 32900 33348
rect 32732 33122 32788 33124
rect 32732 33070 32734 33122
rect 32734 33070 32786 33122
rect 32786 33070 32788 33122
rect 32732 33068 32788 33070
rect 32396 32786 32452 32788
rect 32396 32734 32398 32786
rect 32398 32734 32450 32786
rect 32450 32734 32452 32786
rect 32396 32732 32452 32734
rect 32396 32284 32452 32340
rect 32396 31554 32452 31556
rect 32396 31502 32398 31554
rect 32398 31502 32450 31554
rect 32450 31502 32452 31554
rect 32396 31500 32452 31502
rect 32284 31388 32340 31444
rect 33516 34972 33572 35028
rect 33516 33740 33572 33796
rect 33292 33628 33348 33684
rect 33740 35586 33796 35588
rect 33740 35534 33742 35586
rect 33742 35534 33794 35586
rect 33794 35534 33796 35586
rect 33740 35532 33796 35534
rect 34008 37658 34064 37660
rect 34112 37658 34168 37660
rect 34008 37606 34024 37658
rect 34024 37606 34064 37658
rect 34112 37606 34148 37658
rect 34148 37606 34168 37658
rect 34008 37604 34064 37606
rect 34112 37604 34168 37606
rect 34216 37604 34272 37660
rect 34320 37658 34376 37660
rect 34424 37658 34480 37660
rect 34528 37658 34584 37660
rect 34320 37606 34324 37658
rect 34324 37606 34376 37658
rect 34424 37606 34448 37658
rect 34448 37606 34480 37658
rect 34528 37606 34572 37658
rect 34572 37606 34584 37658
rect 34320 37604 34376 37606
rect 34424 37604 34480 37606
rect 34528 37604 34584 37606
rect 34632 37658 34688 37660
rect 34736 37658 34792 37660
rect 34840 37658 34896 37660
rect 34632 37606 34644 37658
rect 34644 37606 34688 37658
rect 34736 37606 34768 37658
rect 34768 37606 34792 37658
rect 34840 37606 34892 37658
rect 34892 37606 34896 37658
rect 34632 37604 34688 37606
rect 34736 37604 34792 37606
rect 34840 37604 34896 37606
rect 34944 37604 35000 37660
rect 35048 37658 35104 37660
rect 35152 37658 35208 37660
rect 35048 37606 35068 37658
rect 35068 37606 35104 37658
rect 35152 37606 35192 37658
rect 35192 37606 35208 37658
rect 35048 37604 35104 37606
rect 35152 37604 35208 37606
rect 34524 37436 34580 37492
rect 34188 36876 34244 36932
rect 35196 37266 35252 37268
rect 35196 37214 35198 37266
rect 35198 37214 35250 37266
rect 35250 37214 35252 37266
rect 35196 37212 35252 37214
rect 34188 36204 34244 36260
rect 35644 38220 35700 38276
rect 36092 38162 36148 38164
rect 36092 38110 36094 38162
rect 36094 38110 36146 38162
rect 36146 38110 36148 38162
rect 36092 38108 36148 38110
rect 36428 39116 36484 39172
rect 37548 44322 37604 44324
rect 37548 44270 37550 44322
rect 37550 44270 37602 44322
rect 37602 44270 37604 44322
rect 37548 44268 37604 44270
rect 36988 42754 37044 42756
rect 36988 42702 36990 42754
rect 36990 42702 37042 42754
rect 37042 42702 37044 42754
rect 36988 42700 37044 42702
rect 37100 42588 37156 42644
rect 36988 41916 37044 41972
rect 37660 43596 37716 43652
rect 37212 41916 37268 41972
rect 37660 42700 37716 42756
rect 37660 42530 37716 42532
rect 37660 42478 37662 42530
rect 37662 42478 37714 42530
rect 37714 42478 37716 42530
rect 37660 42476 37716 42478
rect 37548 42028 37604 42084
rect 37884 43596 37940 43652
rect 37884 42530 37940 42532
rect 37884 42478 37886 42530
rect 37886 42478 37938 42530
rect 37938 42478 37940 42530
rect 37884 42476 37940 42478
rect 37772 42364 37828 42420
rect 37884 41804 37940 41860
rect 37100 41356 37156 41412
rect 37212 41074 37268 41076
rect 37212 41022 37214 41074
rect 37214 41022 37266 41074
rect 37266 41022 37268 41074
rect 37212 41020 37268 41022
rect 34008 36090 34064 36092
rect 34112 36090 34168 36092
rect 34008 36038 34024 36090
rect 34024 36038 34064 36090
rect 34112 36038 34148 36090
rect 34148 36038 34168 36090
rect 34008 36036 34064 36038
rect 34112 36036 34168 36038
rect 34216 36036 34272 36092
rect 34320 36090 34376 36092
rect 34424 36090 34480 36092
rect 34528 36090 34584 36092
rect 34320 36038 34324 36090
rect 34324 36038 34376 36090
rect 34424 36038 34448 36090
rect 34448 36038 34480 36090
rect 34528 36038 34572 36090
rect 34572 36038 34584 36090
rect 34320 36036 34376 36038
rect 34424 36036 34480 36038
rect 34528 36036 34584 36038
rect 34632 36090 34688 36092
rect 34736 36090 34792 36092
rect 34840 36090 34896 36092
rect 34632 36038 34644 36090
rect 34644 36038 34688 36090
rect 34736 36038 34768 36090
rect 34768 36038 34792 36090
rect 34840 36038 34892 36090
rect 34892 36038 34896 36090
rect 34632 36036 34688 36038
rect 34736 36036 34792 36038
rect 34840 36036 34896 36038
rect 34944 36036 35000 36092
rect 35048 36090 35104 36092
rect 35152 36090 35208 36092
rect 35048 36038 35068 36090
rect 35068 36038 35104 36090
rect 35152 36038 35192 36090
rect 35192 36038 35208 36090
rect 35048 36036 35104 36038
rect 35152 36036 35208 36038
rect 34300 35868 34356 35924
rect 34636 35756 34692 35812
rect 34300 35420 34356 35476
rect 33180 33516 33236 33572
rect 33404 33068 33460 33124
rect 34524 34860 34580 34916
rect 35196 35868 35252 35924
rect 35420 35644 35476 35700
rect 36204 37378 36260 37380
rect 36204 37326 36206 37378
rect 36206 37326 36258 37378
rect 36258 37326 36260 37378
rect 36204 37324 36260 37326
rect 36316 37100 36372 37156
rect 35868 35026 35924 35028
rect 35868 34974 35870 35026
rect 35870 34974 35922 35026
rect 35922 34974 35924 35026
rect 35868 34972 35924 34974
rect 35084 34802 35140 34804
rect 35084 34750 35086 34802
rect 35086 34750 35138 34802
rect 35138 34750 35140 34802
rect 35084 34748 35140 34750
rect 37100 39116 37156 39172
rect 37660 41244 37716 41300
rect 37772 40572 37828 40628
rect 38220 42476 38276 42532
rect 37996 40908 38052 40964
rect 38220 40572 38276 40628
rect 38108 39788 38164 39844
rect 37212 39004 37268 39060
rect 37324 38332 37380 38388
rect 36988 37100 37044 37156
rect 36428 36204 36484 36260
rect 36204 35532 36260 35588
rect 36316 35644 36372 35700
rect 36988 36092 37044 36148
rect 38108 38892 38164 38948
rect 37884 38332 37940 38388
rect 37660 38108 37716 38164
rect 37324 37436 37380 37492
rect 37436 37324 37492 37380
rect 37324 36370 37380 36372
rect 37324 36318 37326 36370
rect 37326 36318 37378 36370
rect 37378 36318 37380 36370
rect 37324 36316 37380 36318
rect 37996 38162 38052 38164
rect 37996 38110 37998 38162
rect 37998 38110 38050 38162
rect 38050 38110 38052 38162
rect 37996 38108 38052 38110
rect 36540 35532 36596 35588
rect 37212 35698 37268 35700
rect 37212 35646 37214 35698
rect 37214 35646 37266 35698
rect 37266 35646 37268 35698
rect 37212 35644 37268 35646
rect 36988 35308 37044 35364
rect 37324 35138 37380 35140
rect 37324 35086 37326 35138
rect 37326 35086 37378 35138
rect 37378 35086 37380 35138
rect 37324 35084 37380 35086
rect 37772 35196 37828 35252
rect 37996 37324 38052 37380
rect 38108 36258 38164 36260
rect 38108 36206 38110 36258
rect 38110 36206 38162 36258
rect 38162 36206 38164 36258
rect 38108 36204 38164 36206
rect 37884 35084 37940 35140
rect 34860 34690 34916 34692
rect 34860 34638 34862 34690
rect 34862 34638 34914 34690
rect 34914 34638 34916 34690
rect 34860 34636 34916 34638
rect 34008 34522 34064 34524
rect 34112 34522 34168 34524
rect 34008 34470 34024 34522
rect 34024 34470 34064 34522
rect 34112 34470 34148 34522
rect 34148 34470 34168 34522
rect 34008 34468 34064 34470
rect 34112 34468 34168 34470
rect 34216 34468 34272 34524
rect 34320 34522 34376 34524
rect 34424 34522 34480 34524
rect 34528 34522 34584 34524
rect 34320 34470 34324 34522
rect 34324 34470 34376 34522
rect 34424 34470 34448 34522
rect 34448 34470 34480 34522
rect 34528 34470 34572 34522
rect 34572 34470 34584 34522
rect 34320 34468 34376 34470
rect 34424 34468 34480 34470
rect 34528 34468 34584 34470
rect 34632 34522 34688 34524
rect 34736 34522 34792 34524
rect 34840 34522 34896 34524
rect 34632 34470 34644 34522
rect 34644 34470 34688 34522
rect 34736 34470 34768 34522
rect 34768 34470 34792 34522
rect 34840 34470 34892 34522
rect 34892 34470 34896 34522
rect 34632 34468 34688 34470
rect 34736 34468 34792 34470
rect 34840 34468 34896 34470
rect 34944 34468 35000 34524
rect 35048 34522 35104 34524
rect 35152 34522 35208 34524
rect 35048 34470 35068 34522
rect 35068 34470 35104 34522
rect 35152 34470 35192 34522
rect 35192 34470 35208 34522
rect 35048 34468 35104 34470
rect 35152 34468 35208 34470
rect 33516 32732 33572 32788
rect 33516 32562 33572 32564
rect 33516 32510 33518 32562
rect 33518 32510 33570 32562
rect 33570 32510 33572 32562
rect 33516 32508 33572 32510
rect 32620 31778 32676 31780
rect 32620 31726 32622 31778
rect 32622 31726 32674 31778
rect 32674 31726 32676 31778
rect 32620 31724 32676 31726
rect 33404 32338 33460 32340
rect 33404 32286 33406 32338
rect 33406 32286 33458 32338
rect 33458 32286 33460 32338
rect 33404 32284 33460 32286
rect 32508 31052 32564 31108
rect 33516 31724 33572 31780
rect 32396 30940 32452 30996
rect 32508 30828 32564 30884
rect 32060 28364 32116 28420
rect 33068 29426 33124 29428
rect 33068 29374 33070 29426
rect 33070 29374 33122 29426
rect 33122 29374 33124 29426
rect 33068 29372 33124 29374
rect 32956 27916 33012 27972
rect 33068 28588 33124 28644
rect 33292 31388 33348 31444
rect 35868 34524 35924 34580
rect 34412 34188 34468 34244
rect 34188 33964 34244 34020
rect 34076 33628 34132 33684
rect 33964 33516 34020 33572
rect 33740 33234 33796 33236
rect 33740 33182 33742 33234
rect 33742 33182 33794 33234
rect 33794 33182 33796 33234
rect 33740 33180 33796 33182
rect 33740 32956 33796 33012
rect 33516 29372 33572 29428
rect 35084 33740 35140 33796
rect 35420 33516 35476 33572
rect 35084 33404 35140 33460
rect 34748 33346 34804 33348
rect 34748 33294 34750 33346
rect 34750 33294 34802 33346
rect 34802 33294 34804 33346
rect 34748 33292 34804 33294
rect 34076 33180 34132 33236
rect 34008 32954 34064 32956
rect 34112 32954 34168 32956
rect 34008 32902 34024 32954
rect 34024 32902 34064 32954
rect 34112 32902 34148 32954
rect 34148 32902 34168 32954
rect 34008 32900 34064 32902
rect 34112 32900 34168 32902
rect 34216 32900 34272 32956
rect 34320 32954 34376 32956
rect 34424 32954 34480 32956
rect 34528 32954 34584 32956
rect 34320 32902 34324 32954
rect 34324 32902 34376 32954
rect 34424 32902 34448 32954
rect 34448 32902 34480 32954
rect 34528 32902 34572 32954
rect 34572 32902 34584 32954
rect 34320 32900 34376 32902
rect 34424 32900 34480 32902
rect 34528 32900 34584 32902
rect 34632 32954 34688 32956
rect 34736 32954 34792 32956
rect 34840 32954 34896 32956
rect 34632 32902 34644 32954
rect 34644 32902 34688 32954
rect 34736 32902 34768 32954
rect 34768 32902 34792 32954
rect 34840 32902 34892 32954
rect 34892 32902 34896 32954
rect 34632 32900 34688 32902
rect 34736 32900 34792 32902
rect 34840 32900 34896 32902
rect 34944 32900 35000 32956
rect 35048 32954 35104 32956
rect 35152 32954 35208 32956
rect 35048 32902 35068 32954
rect 35068 32902 35104 32954
rect 35152 32902 35192 32954
rect 35192 32902 35208 32954
rect 35048 32900 35104 32902
rect 35152 32900 35208 32902
rect 34076 32786 34132 32788
rect 34076 32734 34078 32786
rect 34078 32734 34130 32786
rect 34130 32734 34132 32786
rect 34076 32732 34132 32734
rect 34524 32508 34580 32564
rect 34748 31836 34804 31892
rect 34188 31778 34244 31780
rect 34188 31726 34190 31778
rect 34190 31726 34242 31778
rect 34242 31726 34244 31778
rect 34188 31724 34244 31726
rect 36428 34860 36484 34916
rect 36876 34860 36932 34916
rect 37548 34860 37604 34916
rect 37212 34802 37268 34804
rect 37212 34750 37214 34802
rect 37214 34750 37266 34802
rect 37266 34750 37268 34802
rect 37212 34748 37268 34750
rect 37548 34690 37604 34692
rect 37548 34638 37550 34690
rect 37550 34638 37602 34690
rect 37602 34638 37604 34690
rect 37548 34636 37604 34638
rect 36988 34524 37044 34580
rect 37436 34354 37492 34356
rect 37436 34302 37438 34354
rect 37438 34302 37490 34354
rect 37490 34302 37492 34354
rect 37436 34300 37492 34302
rect 35532 33404 35588 33460
rect 36988 33740 37044 33796
rect 36092 32732 36148 32788
rect 36876 33516 36932 33572
rect 37212 33516 37268 33572
rect 37100 33404 37156 33460
rect 36988 32786 37044 32788
rect 36988 32734 36990 32786
rect 36990 32734 37042 32786
rect 37042 32734 37044 32786
rect 36988 32732 37044 32734
rect 35308 31948 35364 32004
rect 33964 31500 34020 31556
rect 34008 31386 34064 31388
rect 34112 31386 34168 31388
rect 34008 31334 34024 31386
rect 34024 31334 34064 31386
rect 34112 31334 34148 31386
rect 34148 31334 34168 31386
rect 34008 31332 34064 31334
rect 34112 31332 34168 31334
rect 34216 31332 34272 31388
rect 34320 31386 34376 31388
rect 34424 31386 34480 31388
rect 34528 31386 34584 31388
rect 34320 31334 34324 31386
rect 34324 31334 34376 31386
rect 34424 31334 34448 31386
rect 34448 31334 34480 31386
rect 34528 31334 34572 31386
rect 34572 31334 34584 31386
rect 34320 31332 34376 31334
rect 34424 31332 34480 31334
rect 34528 31332 34584 31334
rect 34632 31386 34688 31388
rect 34736 31386 34792 31388
rect 34840 31386 34896 31388
rect 34632 31334 34644 31386
rect 34644 31334 34688 31386
rect 34736 31334 34768 31386
rect 34768 31334 34792 31386
rect 34840 31334 34892 31386
rect 34892 31334 34896 31386
rect 34632 31332 34688 31334
rect 34736 31332 34792 31334
rect 34840 31332 34896 31334
rect 34944 31332 35000 31388
rect 35048 31386 35104 31388
rect 35152 31386 35208 31388
rect 35048 31334 35068 31386
rect 35068 31334 35104 31386
rect 35152 31334 35192 31386
rect 35192 31334 35208 31386
rect 35048 31332 35104 31334
rect 35152 31332 35208 31334
rect 37324 33292 37380 33348
rect 38108 35532 38164 35588
rect 37996 34860 38052 34916
rect 38108 35196 38164 35252
rect 37772 34300 37828 34356
rect 37884 34018 37940 34020
rect 37884 33966 37886 34018
rect 37886 33966 37938 34018
rect 37938 33966 37940 34018
rect 37884 33964 37940 33966
rect 34076 31106 34132 31108
rect 34076 31054 34078 31106
rect 34078 31054 34130 31106
rect 34130 31054 34132 31106
rect 34076 31052 34132 31054
rect 35196 30994 35252 30996
rect 35196 30942 35198 30994
rect 35198 30942 35250 30994
rect 35250 30942 35252 30994
rect 35196 30940 35252 30942
rect 36092 31948 36148 32004
rect 36204 31890 36260 31892
rect 36204 31838 36206 31890
rect 36206 31838 36258 31890
rect 36258 31838 36260 31890
rect 36204 31836 36260 31838
rect 34636 29932 34692 29988
rect 34008 29818 34064 29820
rect 34112 29818 34168 29820
rect 34008 29766 34024 29818
rect 34024 29766 34064 29818
rect 34112 29766 34148 29818
rect 34148 29766 34168 29818
rect 34008 29764 34064 29766
rect 34112 29764 34168 29766
rect 34216 29764 34272 29820
rect 34320 29818 34376 29820
rect 34424 29818 34480 29820
rect 34528 29818 34584 29820
rect 34320 29766 34324 29818
rect 34324 29766 34376 29818
rect 34424 29766 34448 29818
rect 34448 29766 34480 29818
rect 34528 29766 34572 29818
rect 34572 29766 34584 29818
rect 34320 29764 34376 29766
rect 34424 29764 34480 29766
rect 34528 29764 34584 29766
rect 34632 29818 34688 29820
rect 34736 29818 34792 29820
rect 34840 29818 34896 29820
rect 34632 29766 34644 29818
rect 34644 29766 34688 29818
rect 34736 29766 34768 29818
rect 34768 29766 34792 29818
rect 34840 29766 34892 29818
rect 34892 29766 34896 29818
rect 34632 29764 34688 29766
rect 34736 29764 34792 29766
rect 34840 29764 34896 29766
rect 34944 29764 35000 29820
rect 35048 29818 35104 29820
rect 35152 29818 35208 29820
rect 35048 29766 35068 29818
rect 35068 29766 35104 29818
rect 35152 29766 35192 29818
rect 35192 29766 35208 29818
rect 35048 29764 35104 29766
rect 35152 29764 35208 29766
rect 33292 28476 33348 28532
rect 32956 25676 33012 25732
rect 33740 25564 33796 25620
rect 33404 25282 33460 25284
rect 33404 25230 33406 25282
rect 33406 25230 33458 25282
rect 33458 25230 33460 25282
rect 33404 25228 33460 25230
rect 31388 23436 31444 23492
rect 31500 23714 31556 23716
rect 31500 23662 31502 23714
rect 31502 23662 31554 23714
rect 31554 23662 31556 23714
rect 31500 23660 31556 23662
rect 31948 23714 32004 23716
rect 31948 23662 31950 23714
rect 31950 23662 32002 23714
rect 32002 23662 32004 23714
rect 31948 23660 32004 23662
rect 30492 22092 30548 22148
rect 30044 21868 30100 21924
rect 30156 21420 30212 21476
rect 30380 20802 30436 20804
rect 30380 20750 30382 20802
rect 30382 20750 30434 20802
rect 30434 20750 30436 20802
rect 30380 20748 30436 20750
rect 30268 20076 30324 20132
rect 30156 20018 30212 20020
rect 30156 19966 30158 20018
rect 30158 19966 30210 20018
rect 30210 19966 30212 20018
rect 30156 19964 30212 19966
rect 31388 22652 31444 22708
rect 31052 21868 31108 21924
rect 30828 20076 30884 20132
rect 30268 19794 30324 19796
rect 30268 19742 30270 19794
rect 30270 19742 30322 19794
rect 30322 19742 30324 19794
rect 30268 19740 30324 19742
rect 30044 19180 30100 19236
rect 29036 18562 29092 18564
rect 29036 18510 29038 18562
rect 29038 18510 29090 18562
rect 29090 18510 29092 18562
rect 29036 18508 29092 18510
rect 28364 18284 28420 18340
rect 28252 17442 28308 17444
rect 28252 17390 28254 17442
rect 28254 17390 28306 17442
rect 28306 17390 28308 17442
rect 28252 17388 28308 17390
rect 27020 16940 27076 16996
rect 26796 16044 26852 16100
rect 26684 15932 26740 15988
rect 27580 15260 27636 15316
rect 26908 15036 26964 15092
rect 29596 18674 29652 18676
rect 29596 18622 29598 18674
rect 29598 18622 29650 18674
rect 29650 18622 29652 18674
rect 29596 18620 29652 18622
rect 29036 15820 29092 15876
rect 28252 15260 28308 15316
rect 28476 15538 28532 15540
rect 28476 15486 28478 15538
rect 28478 15486 28530 15538
rect 28530 15486 28532 15538
rect 28476 15484 28532 15486
rect 27916 14306 27972 14308
rect 27916 14254 27918 14306
rect 27918 14254 27970 14306
rect 27970 14254 27972 14306
rect 27916 14252 27972 14254
rect 26684 13580 26740 13636
rect 26908 13692 26964 13748
rect 26460 13468 26516 13524
rect 26796 13522 26852 13524
rect 26796 13470 26798 13522
rect 26798 13470 26850 13522
rect 26850 13470 26852 13522
rect 26796 13468 26852 13470
rect 27916 13692 27972 13748
rect 27356 13132 27412 13188
rect 26572 13074 26628 13076
rect 26572 13022 26574 13074
rect 26574 13022 26626 13074
rect 26626 13022 26628 13074
rect 26572 13020 26628 13022
rect 25788 12796 25844 12852
rect 24008 11786 24064 11788
rect 24112 11786 24168 11788
rect 24008 11734 24024 11786
rect 24024 11734 24064 11786
rect 24112 11734 24148 11786
rect 24148 11734 24168 11786
rect 24008 11732 24064 11734
rect 24112 11732 24168 11734
rect 24216 11732 24272 11788
rect 24320 11786 24376 11788
rect 24424 11786 24480 11788
rect 24528 11786 24584 11788
rect 24320 11734 24324 11786
rect 24324 11734 24376 11786
rect 24424 11734 24448 11786
rect 24448 11734 24480 11786
rect 24528 11734 24572 11786
rect 24572 11734 24584 11786
rect 24320 11732 24376 11734
rect 24424 11732 24480 11734
rect 24528 11732 24584 11734
rect 24632 11786 24688 11788
rect 24736 11786 24792 11788
rect 24840 11786 24896 11788
rect 24632 11734 24644 11786
rect 24644 11734 24688 11786
rect 24736 11734 24768 11786
rect 24768 11734 24792 11786
rect 24840 11734 24892 11786
rect 24892 11734 24896 11786
rect 24632 11732 24688 11734
rect 24736 11732 24792 11734
rect 24840 11732 24896 11734
rect 24944 11732 25000 11788
rect 25048 11786 25104 11788
rect 25152 11786 25208 11788
rect 25048 11734 25068 11786
rect 25068 11734 25104 11786
rect 25152 11734 25192 11786
rect 25192 11734 25208 11786
rect 25048 11732 25104 11734
rect 25152 11732 25208 11734
rect 25452 11452 25508 11508
rect 26124 11506 26180 11508
rect 26124 11454 26126 11506
rect 26126 11454 26178 11506
rect 26178 11454 26180 11506
rect 26124 11452 26180 11454
rect 27356 12348 27412 12404
rect 26684 11452 26740 11508
rect 23660 10834 23716 10836
rect 23660 10782 23662 10834
rect 23662 10782 23714 10834
rect 23714 10782 23716 10834
rect 23660 10780 23716 10782
rect 25004 10780 25060 10836
rect 22316 10668 22372 10724
rect 16380 10332 16436 10388
rect 17612 8428 17668 8484
rect 16828 7698 16884 7700
rect 16828 7646 16830 7698
rect 16830 7646 16882 7698
rect 16882 7646 16884 7698
rect 16828 7644 16884 7646
rect 13580 7420 13636 7476
rect 14588 7474 14644 7476
rect 14588 7422 14590 7474
rect 14590 7422 14642 7474
rect 14642 7422 14644 7474
rect 14588 7420 14644 7422
rect 15148 7474 15204 7476
rect 15148 7422 15150 7474
rect 15150 7422 15202 7474
rect 15202 7422 15204 7474
rect 15148 7420 15204 7422
rect 14252 6748 14308 6804
rect 15036 6802 15092 6804
rect 15036 6750 15038 6802
rect 15038 6750 15090 6802
rect 15090 6750 15092 6802
rect 15036 6748 15092 6750
rect 13244 6636 13300 6692
rect 10108 5628 10164 5684
rect 8316 3666 8372 3668
rect 8316 3614 8318 3666
rect 8318 3614 8370 3666
rect 8370 3614 8372 3666
rect 8316 3612 8372 3614
rect 9660 4338 9716 4340
rect 9660 4286 9662 4338
rect 9662 4286 9714 4338
rect 9714 4286 9716 4338
rect 9660 4284 9716 4286
rect 11340 5234 11396 5236
rect 11340 5182 11342 5234
rect 11342 5182 11394 5234
rect 11394 5182 11396 5234
rect 11340 5180 11396 5182
rect 13020 6578 13076 6580
rect 13020 6526 13022 6578
rect 13022 6526 13074 6578
rect 13074 6526 13076 6578
rect 13020 6524 13076 6526
rect 16716 6636 16772 6692
rect 13916 6578 13972 6580
rect 13916 6526 13918 6578
rect 13918 6526 13970 6578
rect 13970 6526 13972 6578
rect 13916 6524 13972 6526
rect 16828 6578 16884 6580
rect 16828 6526 16830 6578
rect 16830 6526 16882 6578
rect 16882 6526 16884 6578
rect 16828 6524 16884 6526
rect 16492 6466 16548 6468
rect 16492 6414 16494 6466
rect 16494 6414 16546 6466
rect 16546 6414 16548 6466
rect 16492 6412 16548 6414
rect 14008 6298 14064 6300
rect 14112 6298 14168 6300
rect 14008 6246 14024 6298
rect 14024 6246 14064 6298
rect 14112 6246 14148 6298
rect 14148 6246 14168 6298
rect 14008 6244 14064 6246
rect 14112 6244 14168 6246
rect 14216 6244 14272 6300
rect 14320 6298 14376 6300
rect 14424 6298 14480 6300
rect 14528 6298 14584 6300
rect 14320 6246 14324 6298
rect 14324 6246 14376 6298
rect 14424 6246 14448 6298
rect 14448 6246 14480 6298
rect 14528 6246 14572 6298
rect 14572 6246 14584 6298
rect 14320 6244 14376 6246
rect 14424 6244 14480 6246
rect 14528 6244 14584 6246
rect 14632 6298 14688 6300
rect 14736 6298 14792 6300
rect 14840 6298 14896 6300
rect 14632 6246 14644 6298
rect 14644 6246 14688 6298
rect 14736 6246 14768 6298
rect 14768 6246 14792 6298
rect 14840 6246 14892 6298
rect 14892 6246 14896 6298
rect 14632 6244 14688 6246
rect 14736 6244 14792 6246
rect 14840 6244 14896 6246
rect 14944 6244 15000 6300
rect 15048 6298 15104 6300
rect 15152 6298 15208 6300
rect 15048 6246 15068 6298
rect 15068 6246 15104 6298
rect 15152 6246 15192 6298
rect 15192 6246 15208 6298
rect 15048 6244 15104 6246
rect 15152 6244 15208 6246
rect 13132 5682 13188 5684
rect 13132 5630 13134 5682
rect 13134 5630 13186 5682
rect 13186 5630 13188 5682
rect 13132 5628 13188 5630
rect 11900 5180 11956 5236
rect 13580 5234 13636 5236
rect 13580 5182 13582 5234
rect 13582 5182 13634 5234
rect 13634 5182 13636 5234
rect 13580 5180 13636 5182
rect 10332 5122 10388 5124
rect 10332 5070 10334 5122
rect 10334 5070 10386 5122
rect 10386 5070 10388 5122
rect 10332 5068 10388 5070
rect 10892 5122 10948 5124
rect 10892 5070 10894 5122
rect 10894 5070 10946 5122
rect 10946 5070 10948 5122
rect 10892 5068 10948 5070
rect 13244 4956 13300 5012
rect 12572 4562 12628 4564
rect 12572 4510 12574 4562
rect 12574 4510 12626 4562
rect 12626 4510 12628 4562
rect 12572 4508 12628 4510
rect 16380 5906 16436 5908
rect 16380 5854 16382 5906
rect 16382 5854 16434 5906
rect 16434 5854 16436 5906
rect 16380 5852 16436 5854
rect 17500 6412 17556 6468
rect 19404 8482 19460 8484
rect 19404 8430 19406 8482
rect 19406 8430 19458 8482
rect 19458 8430 19460 8482
rect 19404 8428 19460 8430
rect 18956 8316 19012 8372
rect 18620 8204 18676 8260
rect 18060 8146 18116 8148
rect 18060 8094 18062 8146
rect 18062 8094 18114 8146
rect 18114 8094 18116 8146
rect 18060 8092 18116 8094
rect 17276 5906 17332 5908
rect 17276 5854 17278 5906
rect 17278 5854 17330 5906
rect 17330 5854 17332 5906
rect 17276 5852 17332 5854
rect 18732 8146 18788 8148
rect 18732 8094 18734 8146
rect 18734 8094 18786 8146
rect 18786 8094 18788 8146
rect 18732 8092 18788 8094
rect 18060 6524 18116 6580
rect 18620 6130 18676 6132
rect 18620 6078 18622 6130
rect 18622 6078 18674 6130
rect 18674 6078 18676 6130
rect 18620 6076 18676 6078
rect 14028 5234 14084 5236
rect 14028 5182 14030 5234
rect 14030 5182 14082 5234
rect 14082 5182 14084 5234
rect 14028 5180 14084 5182
rect 15372 5010 15428 5012
rect 15372 4958 15374 5010
rect 15374 4958 15426 5010
rect 15426 4958 15428 5010
rect 15372 4956 15428 4958
rect 16828 4956 16884 5012
rect 13804 4844 13860 4900
rect 14008 4730 14064 4732
rect 14112 4730 14168 4732
rect 14008 4678 14024 4730
rect 14024 4678 14064 4730
rect 14112 4678 14148 4730
rect 14148 4678 14168 4730
rect 14008 4676 14064 4678
rect 14112 4676 14168 4678
rect 14216 4676 14272 4732
rect 14320 4730 14376 4732
rect 14424 4730 14480 4732
rect 14528 4730 14584 4732
rect 14320 4678 14324 4730
rect 14324 4678 14376 4730
rect 14424 4678 14448 4730
rect 14448 4678 14480 4730
rect 14528 4678 14572 4730
rect 14572 4678 14584 4730
rect 14320 4676 14376 4678
rect 14424 4676 14480 4678
rect 14528 4676 14584 4678
rect 14632 4730 14688 4732
rect 14736 4730 14792 4732
rect 14840 4730 14896 4732
rect 14632 4678 14644 4730
rect 14644 4678 14688 4730
rect 14736 4678 14768 4730
rect 14768 4678 14792 4730
rect 14840 4678 14892 4730
rect 14892 4678 14896 4730
rect 14632 4676 14688 4678
rect 14736 4676 14792 4678
rect 14840 4676 14896 4678
rect 14944 4676 15000 4732
rect 15048 4730 15104 4732
rect 15152 4730 15208 4732
rect 15048 4678 15068 4730
rect 15068 4678 15104 4730
rect 15152 4678 15192 4730
rect 15192 4678 15208 4730
rect 15048 4676 15104 4678
rect 15152 4676 15208 4678
rect 13804 4508 13860 4564
rect 16380 4562 16436 4564
rect 16380 4510 16382 4562
rect 16382 4510 16434 4562
rect 16434 4510 16436 4562
rect 16380 4508 16436 4510
rect 18060 4450 18116 4452
rect 18060 4398 18062 4450
rect 18062 4398 18114 4450
rect 18114 4398 18116 4450
rect 18060 4396 18116 4398
rect 13244 4338 13300 4340
rect 13244 4286 13246 4338
rect 13246 4286 13298 4338
rect 13298 4286 13300 4338
rect 13244 4284 13300 4286
rect 13132 4114 13188 4116
rect 13132 4062 13134 4114
rect 13134 4062 13186 4114
rect 13186 4062 13188 4114
rect 13132 4060 13188 4062
rect 9324 3612 9380 3668
rect 16940 3948 16996 4004
rect 17276 3724 17332 3780
rect 17948 4060 18004 4116
rect 13916 3612 13972 3668
rect 16940 3666 16996 3668
rect 16940 3614 16942 3666
rect 16942 3614 16994 3666
rect 16994 3614 16996 3666
rect 16940 3612 16996 3614
rect 9884 3388 9940 3444
rect 13244 3442 13300 3444
rect 13244 3390 13246 3442
rect 13246 3390 13298 3442
rect 13298 3390 13300 3442
rect 13244 3388 13300 3390
rect 13692 3442 13748 3444
rect 13692 3390 13694 3442
rect 13694 3390 13746 3442
rect 13746 3390 13748 3442
rect 13692 3388 13748 3390
rect 16156 3442 16212 3444
rect 16156 3390 16158 3442
rect 16158 3390 16210 3442
rect 16210 3390 16212 3442
rect 16156 3388 16212 3390
rect 19516 8204 19572 8260
rect 19740 8316 19796 8372
rect 19516 8034 19572 8036
rect 19516 7982 19518 8034
rect 19518 7982 19570 8034
rect 19570 7982 19572 8034
rect 19516 7980 19572 7982
rect 21196 8204 21252 8260
rect 19964 8146 20020 8148
rect 19964 8094 19966 8146
rect 19966 8094 20018 8146
rect 20018 8094 20020 8146
rect 19964 8092 20020 8094
rect 19292 7644 19348 7700
rect 19740 7644 19796 7700
rect 20076 7532 20132 7588
rect 18172 3948 18228 4004
rect 19068 4396 19124 4452
rect 18732 3442 18788 3444
rect 18732 3390 18734 3442
rect 18734 3390 18786 3442
rect 18786 3390 18788 3442
rect 18732 3388 18788 3390
rect 20300 7980 20356 8036
rect 23996 10722 24052 10724
rect 23996 10670 23998 10722
rect 23998 10670 24050 10722
rect 24050 10670 24052 10722
rect 23996 10668 24052 10670
rect 26572 10668 26628 10724
rect 24008 10218 24064 10220
rect 24112 10218 24168 10220
rect 24008 10166 24024 10218
rect 24024 10166 24064 10218
rect 24112 10166 24148 10218
rect 24148 10166 24168 10218
rect 24008 10164 24064 10166
rect 24112 10164 24168 10166
rect 24216 10164 24272 10220
rect 24320 10218 24376 10220
rect 24424 10218 24480 10220
rect 24528 10218 24584 10220
rect 24320 10166 24324 10218
rect 24324 10166 24376 10218
rect 24424 10166 24448 10218
rect 24448 10166 24480 10218
rect 24528 10166 24572 10218
rect 24572 10166 24584 10218
rect 24320 10164 24376 10166
rect 24424 10164 24480 10166
rect 24528 10164 24584 10166
rect 24632 10218 24688 10220
rect 24736 10218 24792 10220
rect 24840 10218 24896 10220
rect 24632 10166 24644 10218
rect 24644 10166 24688 10218
rect 24736 10166 24768 10218
rect 24768 10166 24792 10218
rect 24840 10166 24892 10218
rect 24892 10166 24896 10218
rect 24632 10164 24688 10166
rect 24736 10164 24792 10166
rect 24840 10164 24896 10166
rect 24944 10164 25000 10220
rect 25048 10218 25104 10220
rect 25152 10218 25208 10220
rect 25048 10166 25068 10218
rect 25068 10166 25104 10218
rect 25152 10166 25192 10218
rect 25192 10166 25208 10218
rect 25048 10164 25104 10166
rect 25152 10164 25208 10166
rect 25788 9884 25844 9940
rect 25340 9042 25396 9044
rect 25340 8990 25342 9042
rect 25342 8990 25394 9042
rect 25394 8990 25396 9042
rect 25340 8988 25396 8990
rect 25900 9660 25956 9716
rect 24008 8650 24064 8652
rect 24112 8650 24168 8652
rect 24008 8598 24024 8650
rect 24024 8598 24064 8650
rect 24112 8598 24148 8650
rect 24148 8598 24168 8650
rect 24008 8596 24064 8598
rect 24112 8596 24168 8598
rect 24216 8596 24272 8652
rect 24320 8650 24376 8652
rect 24424 8650 24480 8652
rect 24528 8650 24584 8652
rect 24320 8598 24324 8650
rect 24324 8598 24376 8650
rect 24424 8598 24448 8650
rect 24448 8598 24480 8650
rect 24528 8598 24572 8650
rect 24572 8598 24584 8650
rect 24320 8596 24376 8598
rect 24424 8596 24480 8598
rect 24528 8596 24584 8598
rect 24632 8650 24688 8652
rect 24736 8650 24792 8652
rect 24840 8650 24896 8652
rect 24632 8598 24644 8650
rect 24644 8598 24688 8650
rect 24736 8598 24768 8650
rect 24768 8598 24792 8650
rect 24840 8598 24892 8650
rect 24892 8598 24896 8650
rect 24632 8596 24688 8598
rect 24736 8596 24792 8598
rect 24840 8596 24896 8598
rect 24944 8596 25000 8652
rect 25048 8650 25104 8652
rect 25152 8650 25208 8652
rect 25048 8598 25068 8650
rect 25068 8598 25104 8650
rect 25152 8598 25192 8650
rect 25192 8598 25208 8650
rect 25048 8596 25104 8598
rect 25152 8596 25208 8598
rect 27020 9938 27076 9940
rect 27020 9886 27022 9938
rect 27022 9886 27074 9938
rect 27074 9886 27076 9938
rect 27020 9884 27076 9886
rect 28252 12402 28308 12404
rect 28252 12350 28254 12402
rect 28254 12350 28306 12402
rect 28306 12350 28308 12402
rect 28252 12348 28308 12350
rect 28028 9714 28084 9716
rect 28028 9662 28030 9714
rect 28030 9662 28082 9714
rect 28082 9662 28084 9714
rect 28028 9660 28084 9662
rect 28252 9100 28308 9156
rect 25340 7756 25396 7812
rect 20636 7532 20692 7588
rect 21420 7698 21476 7700
rect 21420 7646 21422 7698
rect 21422 7646 21474 7698
rect 21474 7646 21476 7698
rect 21420 7644 21476 7646
rect 20300 6860 20356 6916
rect 21308 6914 21364 6916
rect 21308 6862 21310 6914
rect 21310 6862 21362 6914
rect 21362 6862 21364 6914
rect 21308 6860 21364 6862
rect 21084 6636 21140 6692
rect 20188 6076 20244 6132
rect 20748 6076 20804 6132
rect 20412 5122 20468 5124
rect 20412 5070 20414 5122
rect 20414 5070 20466 5122
rect 20466 5070 20468 5122
rect 20412 5068 20468 5070
rect 20076 4508 20132 4564
rect 24668 7196 24724 7252
rect 24008 7082 24064 7084
rect 24112 7082 24168 7084
rect 24008 7030 24024 7082
rect 24024 7030 24064 7082
rect 24112 7030 24148 7082
rect 24148 7030 24168 7082
rect 24008 7028 24064 7030
rect 24112 7028 24168 7030
rect 24216 7028 24272 7084
rect 24320 7082 24376 7084
rect 24424 7082 24480 7084
rect 24528 7082 24584 7084
rect 24320 7030 24324 7082
rect 24324 7030 24376 7082
rect 24424 7030 24448 7082
rect 24448 7030 24480 7082
rect 24528 7030 24572 7082
rect 24572 7030 24584 7082
rect 24320 7028 24376 7030
rect 24424 7028 24480 7030
rect 24528 7028 24584 7030
rect 24632 7082 24688 7084
rect 24736 7082 24792 7084
rect 24840 7082 24896 7084
rect 24632 7030 24644 7082
rect 24644 7030 24688 7082
rect 24736 7030 24768 7082
rect 24768 7030 24792 7082
rect 24840 7030 24892 7082
rect 24892 7030 24896 7082
rect 24632 7028 24688 7030
rect 24736 7028 24792 7030
rect 24840 7028 24896 7030
rect 24944 7028 25000 7084
rect 25048 7082 25104 7084
rect 25152 7082 25208 7084
rect 25048 7030 25068 7082
rect 25068 7030 25104 7082
rect 25152 7030 25192 7082
rect 25192 7030 25208 7082
rect 25048 7028 25104 7030
rect 25152 7028 25208 7030
rect 26348 7756 26404 7812
rect 26012 7586 26068 7588
rect 26012 7534 26014 7586
rect 26014 7534 26066 7586
rect 26066 7534 26068 7586
rect 26012 7532 26068 7534
rect 26908 7756 26964 7812
rect 25676 7196 25732 7252
rect 22092 6690 22148 6692
rect 22092 6638 22094 6690
rect 22094 6638 22146 6690
rect 22146 6638 22148 6690
rect 22092 6636 22148 6638
rect 21532 6076 21588 6132
rect 25340 6636 25396 6692
rect 24332 5906 24388 5908
rect 24332 5854 24334 5906
rect 24334 5854 24386 5906
rect 24386 5854 24388 5906
rect 24332 5852 24388 5854
rect 25564 6578 25620 6580
rect 25564 6526 25566 6578
rect 25566 6526 25618 6578
rect 25618 6526 25620 6578
rect 25564 6524 25620 6526
rect 24008 5514 24064 5516
rect 24112 5514 24168 5516
rect 24008 5462 24024 5514
rect 24024 5462 24064 5514
rect 24112 5462 24148 5514
rect 24148 5462 24168 5514
rect 24008 5460 24064 5462
rect 24112 5460 24168 5462
rect 24216 5460 24272 5516
rect 24320 5514 24376 5516
rect 24424 5514 24480 5516
rect 24528 5514 24584 5516
rect 24320 5462 24324 5514
rect 24324 5462 24376 5514
rect 24424 5462 24448 5514
rect 24448 5462 24480 5514
rect 24528 5462 24572 5514
rect 24572 5462 24584 5514
rect 24320 5460 24376 5462
rect 24424 5460 24480 5462
rect 24528 5460 24584 5462
rect 24632 5514 24688 5516
rect 24736 5514 24792 5516
rect 24840 5514 24896 5516
rect 24632 5462 24644 5514
rect 24644 5462 24688 5514
rect 24736 5462 24768 5514
rect 24768 5462 24792 5514
rect 24840 5462 24892 5514
rect 24892 5462 24896 5514
rect 24632 5460 24688 5462
rect 24736 5460 24792 5462
rect 24840 5460 24896 5462
rect 24944 5460 25000 5516
rect 25048 5514 25104 5516
rect 25152 5514 25208 5516
rect 25048 5462 25068 5514
rect 25068 5462 25104 5514
rect 25152 5462 25192 5514
rect 25192 5462 25208 5514
rect 25048 5460 25104 5462
rect 25152 5460 25208 5462
rect 22316 5068 22372 5124
rect 23996 4450 24052 4452
rect 23996 4398 23998 4450
rect 23998 4398 24050 4450
rect 24050 4398 24052 4450
rect 23996 4396 24052 4398
rect 24780 4450 24836 4452
rect 24780 4398 24782 4450
rect 24782 4398 24834 4450
rect 24834 4398 24836 4450
rect 24780 4396 24836 4398
rect 19852 3948 19908 4004
rect 20860 3724 20916 3780
rect 26012 6466 26068 6468
rect 26012 6414 26014 6466
rect 26014 6414 26066 6466
rect 26066 6414 26068 6466
rect 26012 6412 26068 6414
rect 26012 5852 26068 5908
rect 30604 18620 30660 18676
rect 30940 19906 30996 19908
rect 30940 19854 30942 19906
rect 30942 19854 30994 19906
rect 30994 19854 30996 19906
rect 30940 19852 30996 19854
rect 31612 23436 31668 23492
rect 33628 22652 33684 22708
rect 34008 28250 34064 28252
rect 34112 28250 34168 28252
rect 34008 28198 34024 28250
rect 34024 28198 34064 28250
rect 34112 28198 34148 28250
rect 34148 28198 34168 28250
rect 34008 28196 34064 28198
rect 34112 28196 34168 28198
rect 34216 28196 34272 28252
rect 34320 28250 34376 28252
rect 34424 28250 34480 28252
rect 34528 28250 34584 28252
rect 34320 28198 34324 28250
rect 34324 28198 34376 28250
rect 34424 28198 34448 28250
rect 34448 28198 34480 28250
rect 34528 28198 34572 28250
rect 34572 28198 34584 28250
rect 34320 28196 34376 28198
rect 34424 28196 34480 28198
rect 34528 28196 34584 28198
rect 34632 28250 34688 28252
rect 34736 28250 34792 28252
rect 34840 28250 34896 28252
rect 34632 28198 34644 28250
rect 34644 28198 34688 28250
rect 34736 28198 34768 28250
rect 34768 28198 34792 28250
rect 34840 28198 34892 28250
rect 34892 28198 34896 28250
rect 34632 28196 34688 28198
rect 34736 28196 34792 28198
rect 34840 28196 34896 28198
rect 34944 28196 35000 28252
rect 35048 28250 35104 28252
rect 35152 28250 35208 28252
rect 35048 28198 35068 28250
rect 35068 28198 35104 28250
rect 35152 28198 35192 28250
rect 35192 28198 35208 28250
rect 35048 28196 35104 28198
rect 35152 28196 35208 28198
rect 33964 28028 34020 28084
rect 34008 26682 34064 26684
rect 34112 26682 34168 26684
rect 34008 26630 34024 26682
rect 34024 26630 34064 26682
rect 34112 26630 34148 26682
rect 34148 26630 34168 26682
rect 34008 26628 34064 26630
rect 34112 26628 34168 26630
rect 34216 26628 34272 26684
rect 34320 26682 34376 26684
rect 34424 26682 34480 26684
rect 34528 26682 34584 26684
rect 34320 26630 34324 26682
rect 34324 26630 34376 26682
rect 34424 26630 34448 26682
rect 34448 26630 34480 26682
rect 34528 26630 34572 26682
rect 34572 26630 34584 26682
rect 34320 26628 34376 26630
rect 34424 26628 34480 26630
rect 34528 26628 34584 26630
rect 34632 26682 34688 26684
rect 34736 26682 34792 26684
rect 34840 26682 34896 26684
rect 34632 26630 34644 26682
rect 34644 26630 34688 26682
rect 34736 26630 34768 26682
rect 34768 26630 34792 26682
rect 34840 26630 34892 26682
rect 34892 26630 34896 26682
rect 34632 26628 34688 26630
rect 34736 26628 34792 26630
rect 34840 26628 34896 26630
rect 34944 26628 35000 26684
rect 35048 26682 35104 26684
rect 35152 26682 35208 26684
rect 35048 26630 35068 26682
rect 35068 26630 35104 26682
rect 35152 26630 35192 26682
rect 35192 26630 35208 26682
rect 35048 26628 35104 26630
rect 35152 26628 35208 26630
rect 34188 25730 34244 25732
rect 34188 25678 34190 25730
rect 34190 25678 34242 25730
rect 34242 25678 34244 25730
rect 34188 25676 34244 25678
rect 34008 25114 34064 25116
rect 34112 25114 34168 25116
rect 34008 25062 34024 25114
rect 34024 25062 34064 25114
rect 34112 25062 34148 25114
rect 34148 25062 34168 25114
rect 34008 25060 34064 25062
rect 34112 25060 34168 25062
rect 34216 25060 34272 25116
rect 34320 25114 34376 25116
rect 34424 25114 34480 25116
rect 34528 25114 34584 25116
rect 34320 25062 34324 25114
rect 34324 25062 34376 25114
rect 34424 25062 34448 25114
rect 34448 25062 34480 25114
rect 34528 25062 34572 25114
rect 34572 25062 34584 25114
rect 34320 25060 34376 25062
rect 34424 25060 34480 25062
rect 34528 25060 34584 25062
rect 34632 25114 34688 25116
rect 34736 25114 34792 25116
rect 34840 25114 34896 25116
rect 34632 25062 34644 25114
rect 34644 25062 34688 25114
rect 34736 25062 34768 25114
rect 34768 25062 34792 25114
rect 34840 25062 34892 25114
rect 34892 25062 34896 25114
rect 34632 25060 34688 25062
rect 34736 25060 34792 25062
rect 34840 25060 34896 25062
rect 34944 25060 35000 25116
rect 35048 25114 35104 25116
rect 35152 25114 35208 25116
rect 35048 25062 35068 25114
rect 35068 25062 35104 25114
rect 35152 25062 35192 25114
rect 35192 25062 35208 25114
rect 35048 25060 35104 25062
rect 35152 25060 35208 25062
rect 34008 23546 34064 23548
rect 34112 23546 34168 23548
rect 34008 23494 34024 23546
rect 34024 23494 34064 23546
rect 34112 23494 34148 23546
rect 34148 23494 34168 23546
rect 34008 23492 34064 23494
rect 34112 23492 34168 23494
rect 34216 23492 34272 23548
rect 34320 23546 34376 23548
rect 34424 23546 34480 23548
rect 34528 23546 34584 23548
rect 34320 23494 34324 23546
rect 34324 23494 34376 23546
rect 34424 23494 34448 23546
rect 34448 23494 34480 23546
rect 34528 23494 34572 23546
rect 34572 23494 34584 23546
rect 34320 23492 34376 23494
rect 34424 23492 34480 23494
rect 34528 23492 34584 23494
rect 34632 23546 34688 23548
rect 34736 23546 34792 23548
rect 34840 23546 34896 23548
rect 34632 23494 34644 23546
rect 34644 23494 34688 23546
rect 34736 23494 34768 23546
rect 34768 23494 34792 23546
rect 34840 23494 34892 23546
rect 34892 23494 34896 23546
rect 34632 23492 34688 23494
rect 34736 23492 34792 23494
rect 34840 23492 34896 23494
rect 34944 23492 35000 23548
rect 35048 23546 35104 23548
rect 35152 23546 35208 23548
rect 35048 23494 35068 23546
rect 35068 23494 35104 23546
rect 35152 23494 35192 23546
rect 35192 23494 35208 23546
rect 35048 23492 35104 23494
rect 35152 23492 35208 23494
rect 33852 22540 33908 22596
rect 34008 21978 34064 21980
rect 34112 21978 34168 21980
rect 34008 21926 34024 21978
rect 34024 21926 34064 21978
rect 34112 21926 34148 21978
rect 34148 21926 34168 21978
rect 34008 21924 34064 21926
rect 34112 21924 34168 21926
rect 34216 21924 34272 21980
rect 34320 21978 34376 21980
rect 34424 21978 34480 21980
rect 34528 21978 34584 21980
rect 34320 21926 34324 21978
rect 34324 21926 34376 21978
rect 34424 21926 34448 21978
rect 34448 21926 34480 21978
rect 34528 21926 34572 21978
rect 34572 21926 34584 21978
rect 34320 21924 34376 21926
rect 34424 21924 34480 21926
rect 34528 21924 34584 21926
rect 34632 21978 34688 21980
rect 34736 21978 34792 21980
rect 34840 21978 34896 21980
rect 34632 21926 34644 21978
rect 34644 21926 34688 21978
rect 34736 21926 34768 21978
rect 34768 21926 34792 21978
rect 34840 21926 34892 21978
rect 34892 21926 34896 21978
rect 34632 21924 34688 21926
rect 34736 21924 34792 21926
rect 34840 21924 34896 21926
rect 34944 21924 35000 21980
rect 35048 21978 35104 21980
rect 35152 21978 35208 21980
rect 35048 21926 35068 21978
rect 35068 21926 35104 21978
rect 35152 21926 35192 21978
rect 35192 21926 35208 21978
rect 35048 21924 35104 21926
rect 35152 21924 35208 21926
rect 31836 20636 31892 20692
rect 32732 20690 32788 20692
rect 32732 20638 32734 20690
rect 32734 20638 32786 20690
rect 32786 20638 32788 20690
rect 32732 20636 32788 20638
rect 31948 20130 32004 20132
rect 31948 20078 31950 20130
rect 31950 20078 32002 20130
rect 32002 20078 32004 20130
rect 31948 20076 32004 20078
rect 34008 20410 34064 20412
rect 34112 20410 34168 20412
rect 34008 20358 34024 20410
rect 34024 20358 34064 20410
rect 34112 20358 34148 20410
rect 34148 20358 34168 20410
rect 34008 20356 34064 20358
rect 34112 20356 34168 20358
rect 34216 20356 34272 20412
rect 34320 20410 34376 20412
rect 34424 20410 34480 20412
rect 34528 20410 34584 20412
rect 34320 20358 34324 20410
rect 34324 20358 34376 20410
rect 34424 20358 34448 20410
rect 34448 20358 34480 20410
rect 34528 20358 34572 20410
rect 34572 20358 34584 20410
rect 34320 20356 34376 20358
rect 34424 20356 34480 20358
rect 34528 20356 34584 20358
rect 34632 20410 34688 20412
rect 34736 20410 34792 20412
rect 34840 20410 34896 20412
rect 34632 20358 34644 20410
rect 34644 20358 34688 20410
rect 34736 20358 34768 20410
rect 34768 20358 34792 20410
rect 34840 20358 34892 20410
rect 34892 20358 34896 20410
rect 34632 20356 34688 20358
rect 34736 20356 34792 20358
rect 34840 20356 34896 20358
rect 34944 20356 35000 20412
rect 35048 20410 35104 20412
rect 35152 20410 35208 20412
rect 35048 20358 35068 20410
rect 35068 20358 35104 20410
rect 35152 20358 35192 20410
rect 35192 20358 35208 20410
rect 35048 20356 35104 20358
rect 35152 20356 35208 20358
rect 33628 20076 33684 20132
rect 31500 19628 31556 19684
rect 32284 19740 32340 19796
rect 32732 19234 32788 19236
rect 32732 19182 32734 19234
rect 32734 19182 32786 19234
rect 32786 19182 32788 19234
rect 32732 19180 32788 19182
rect 34008 18842 34064 18844
rect 34112 18842 34168 18844
rect 34008 18790 34024 18842
rect 34024 18790 34064 18842
rect 34112 18790 34148 18842
rect 34148 18790 34168 18842
rect 34008 18788 34064 18790
rect 34112 18788 34168 18790
rect 34216 18788 34272 18844
rect 34320 18842 34376 18844
rect 34424 18842 34480 18844
rect 34528 18842 34584 18844
rect 34320 18790 34324 18842
rect 34324 18790 34376 18842
rect 34424 18790 34448 18842
rect 34448 18790 34480 18842
rect 34528 18790 34572 18842
rect 34572 18790 34584 18842
rect 34320 18788 34376 18790
rect 34424 18788 34480 18790
rect 34528 18788 34584 18790
rect 34632 18842 34688 18844
rect 34736 18842 34792 18844
rect 34840 18842 34896 18844
rect 34632 18790 34644 18842
rect 34644 18790 34688 18842
rect 34736 18790 34768 18842
rect 34768 18790 34792 18842
rect 34840 18790 34892 18842
rect 34892 18790 34896 18842
rect 34632 18788 34688 18790
rect 34736 18788 34792 18790
rect 34840 18788 34896 18790
rect 34944 18788 35000 18844
rect 35048 18842 35104 18844
rect 35152 18842 35208 18844
rect 35048 18790 35068 18842
rect 35068 18790 35104 18842
rect 35152 18790 35192 18842
rect 35192 18790 35208 18842
rect 35048 18788 35104 18790
rect 35152 18788 35208 18790
rect 30828 18508 30884 18564
rect 30156 18338 30212 18340
rect 30156 18286 30158 18338
rect 30158 18286 30210 18338
rect 30210 18286 30212 18338
rect 30156 18284 30212 18286
rect 29708 17388 29764 17444
rect 29372 16268 29428 16324
rect 34008 17274 34064 17276
rect 34112 17274 34168 17276
rect 34008 17222 34024 17274
rect 34024 17222 34064 17274
rect 34112 17222 34148 17274
rect 34148 17222 34168 17274
rect 34008 17220 34064 17222
rect 34112 17220 34168 17222
rect 34216 17220 34272 17276
rect 34320 17274 34376 17276
rect 34424 17274 34480 17276
rect 34528 17274 34584 17276
rect 34320 17222 34324 17274
rect 34324 17222 34376 17274
rect 34424 17222 34448 17274
rect 34448 17222 34480 17274
rect 34528 17222 34572 17274
rect 34572 17222 34584 17274
rect 34320 17220 34376 17222
rect 34424 17220 34480 17222
rect 34528 17220 34584 17222
rect 34632 17274 34688 17276
rect 34736 17274 34792 17276
rect 34840 17274 34896 17276
rect 34632 17222 34644 17274
rect 34644 17222 34688 17274
rect 34736 17222 34768 17274
rect 34768 17222 34792 17274
rect 34840 17222 34892 17274
rect 34892 17222 34896 17274
rect 34632 17220 34688 17222
rect 34736 17220 34792 17222
rect 34840 17220 34896 17222
rect 34944 17220 35000 17276
rect 35048 17274 35104 17276
rect 35152 17274 35208 17276
rect 35048 17222 35068 17274
rect 35068 17222 35104 17274
rect 35152 17222 35192 17274
rect 35192 17222 35208 17274
rect 35048 17220 35104 17222
rect 35152 17220 35208 17222
rect 30380 16322 30436 16324
rect 30380 16270 30382 16322
rect 30382 16270 30434 16322
rect 30434 16270 30436 16322
rect 30380 16268 30436 16270
rect 34008 15706 34064 15708
rect 34112 15706 34168 15708
rect 34008 15654 34024 15706
rect 34024 15654 34064 15706
rect 34112 15654 34148 15706
rect 34148 15654 34168 15706
rect 34008 15652 34064 15654
rect 34112 15652 34168 15654
rect 34216 15652 34272 15708
rect 34320 15706 34376 15708
rect 34424 15706 34480 15708
rect 34528 15706 34584 15708
rect 34320 15654 34324 15706
rect 34324 15654 34376 15706
rect 34424 15654 34448 15706
rect 34448 15654 34480 15706
rect 34528 15654 34572 15706
rect 34572 15654 34584 15706
rect 34320 15652 34376 15654
rect 34424 15652 34480 15654
rect 34528 15652 34584 15654
rect 34632 15706 34688 15708
rect 34736 15706 34792 15708
rect 34840 15706 34896 15708
rect 34632 15654 34644 15706
rect 34644 15654 34688 15706
rect 34736 15654 34768 15706
rect 34768 15654 34792 15706
rect 34840 15654 34892 15706
rect 34892 15654 34896 15706
rect 34632 15652 34688 15654
rect 34736 15652 34792 15654
rect 34840 15652 34896 15654
rect 34944 15652 35000 15708
rect 35048 15706 35104 15708
rect 35152 15706 35208 15708
rect 35048 15654 35068 15706
rect 35068 15654 35104 15706
rect 35152 15654 35192 15706
rect 35192 15654 35208 15706
rect 35048 15652 35104 15654
rect 35152 15652 35208 15654
rect 29260 15484 29316 15540
rect 29932 15260 29988 15316
rect 28476 14252 28532 14308
rect 34008 14138 34064 14140
rect 34112 14138 34168 14140
rect 34008 14086 34024 14138
rect 34024 14086 34064 14138
rect 34112 14086 34148 14138
rect 34148 14086 34168 14138
rect 34008 14084 34064 14086
rect 34112 14084 34168 14086
rect 34216 14084 34272 14140
rect 34320 14138 34376 14140
rect 34424 14138 34480 14140
rect 34528 14138 34584 14140
rect 34320 14086 34324 14138
rect 34324 14086 34376 14138
rect 34424 14086 34448 14138
rect 34448 14086 34480 14138
rect 34528 14086 34572 14138
rect 34572 14086 34584 14138
rect 34320 14084 34376 14086
rect 34424 14084 34480 14086
rect 34528 14084 34584 14086
rect 34632 14138 34688 14140
rect 34736 14138 34792 14140
rect 34840 14138 34896 14140
rect 34632 14086 34644 14138
rect 34644 14086 34688 14138
rect 34736 14086 34768 14138
rect 34768 14086 34792 14138
rect 34840 14086 34892 14138
rect 34892 14086 34896 14138
rect 34632 14084 34688 14086
rect 34736 14084 34792 14086
rect 34840 14084 34896 14086
rect 34944 14084 35000 14140
rect 35048 14138 35104 14140
rect 35152 14138 35208 14140
rect 35048 14086 35068 14138
rect 35068 14086 35104 14138
rect 35152 14086 35192 14138
rect 35192 14086 35208 14138
rect 35048 14084 35104 14086
rect 35152 14084 35208 14086
rect 34008 12570 34064 12572
rect 34112 12570 34168 12572
rect 34008 12518 34024 12570
rect 34024 12518 34064 12570
rect 34112 12518 34148 12570
rect 34148 12518 34168 12570
rect 34008 12516 34064 12518
rect 34112 12516 34168 12518
rect 34216 12516 34272 12572
rect 34320 12570 34376 12572
rect 34424 12570 34480 12572
rect 34528 12570 34584 12572
rect 34320 12518 34324 12570
rect 34324 12518 34376 12570
rect 34424 12518 34448 12570
rect 34448 12518 34480 12570
rect 34528 12518 34572 12570
rect 34572 12518 34584 12570
rect 34320 12516 34376 12518
rect 34424 12516 34480 12518
rect 34528 12516 34584 12518
rect 34632 12570 34688 12572
rect 34736 12570 34792 12572
rect 34840 12570 34896 12572
rect 34632 12518 34644 12570
rect 34644 12518 34688 12570
rect 34736 12518 34768 12570
rect 34768 12518 34792 12570
rect 34840 12518 34892 12570
rect 34892 12518 34896 12570
rect 34632 12516 34688 12518
rect 34736 12516 34792 12518
rect 34840 12516 34896 12518
rect 34944 12516 35000 12572
rect 35048 12570 35104 12572
rect 35152 12570 35208 12572
rect 35048 12518 35068 12570
rect 35068 12518 35104 12570
rect 35152 12518 35192 12570
rect 35192 12518 35208 12570
rect 35048 12516 35104 12518
rect 35152 12516 35208 12518
rect 34008 11002 34064 11004
rect 34112 11002 34168 11004
rect 34008 10950 34024 11002
rect 34024 10950 34064 11002
rect 34112 10950 34148 11002
rect 34148 10950 34168 11002
rect 34008 10948 34064 10950
rect 34112 10948 34168 10950
rect 34216 10948 34272 11004
rect 34320 11002 34376 11004
rect 34424 11002 34480 11004
rect 34528 11002 34584 11004
rect 34320 10950 34324 11002
rect 34324 10950 34376 11002
rect 34424 10950 34448 11002
rect 34448 10950 34480 11002
rect 34528 10950 34572 11002
rect 34572 10950 34584 11002
rect 34320 10948 34376 10950
rect 34424 10948 34480 10950
rect 34528 10948 34584 10950
rect 34632 11002 34688 11004
rect 34736 11002 34792 11004
rect 34840 11002 34896 11004
rect 34632 10950 34644 11002
rect 34644 10950 34688 11002
rect 34736 10950 34768 11002
rect 34768 10950 34792 11002
rect 34840 10950 34892 11002
rect 34892 10950 34896 11002
rect 34632 10948 34688 10950
rect 34736 10948 34792 10950
rect 34840 10948 34896 10950
rect 34944 10948 35000 11004
rect 35048 11002 35104 11004
rect 35152 11002 35208 11004
rect 35048 10950 35068 11002
rect 35068 10950 35104 11002
rect 35152 10950 35192 11002
rect 35192 10950 35208 11002
rect 35048 10948 35104 10950
rect 35152 10948 35208 10950
rect 34008 9434 34064 9436
rect 34112 9434 34168 9436
rect 34008 9382 34024 9434
rect 34024 9382 34064 9434
rect 34112 9382 34148 9434
rect 34148 9382 34168 9434
rect 34008 9380 34064 9382
rect 34112 9380 34168 9382
rect 34216 9380 34272 9436
rect 34320 9434 34376 9436
rect 34424 9434 34480 9436
rect 34528 9434 34584 9436
rect 34320 9382 34324 9434
rect 34324 9382 34376 9434
rect 34424 9382 34448 9434
rect 34448 9382 34480 9434
rect 34528 9382 34572 9434
rect 34572 9382 34584 9434
rect 34320 9380 34376 9382
rect 34424 9380 34480 9382
rect 34528 9380 34584 9382
rect 34632 9434 34688 9436
rect 34736 9434 34792 9436
rect 34840 9434 34896 9436
rect 34632 9382 34644 9434
rect 34644 9382 34688 9434
rect 34736 9382 34768 9434
rect 34768 9382 34792 9434
rect 34840 9382 34892 9434
rect 34892 9382 34896 9434
rect 34632 9380 34688 9382
rect 34736 9380 34792 9382
rect 34840 9380 34896 9382
rect 34944 9380 35000 9436
rect 35048 9434 35104 9436
rect 35152 9434 35208 9436
rect 35048 9382 35068 9434
rect 35068 9382 35104 9434
rect 35152 9382 35192 9434
rect 35192 9382 35208 9434
rect 35048 9380 35104 9382
rect 35152 9380 35208 9382
rect 29036 9154 29092 9156
rect 29036 9102 29038 9154
rect 29038 9102 29090 9154
rect 29090 9102 29092 9154
rect 29036 9100 29092 9102
rect 28364 8988 28420 9044
rect 29596 9042 29652 9044
rect 29596 8990 29598 9042
rect 29598 8990 29650 9042
rect 29650 8990 29652 9042
rect 29596 8988 29652 8990
rect 34008 7866 34064 7868
rect 34112 7866 34168 7868
rect 27580 7756 27636 7812
rect 28140 7756 28196 7812
rect 34008 7814 34024 7866
rect 34024 7814 34064 7866
rect 34112 7814 34148 7866
rect 34148 7814 34168 7866
rect 34008 7812 34064 7814
rect 34112 7812 34168 7814
rect 34216 7812 34272 7868
rect 34320 7866 34376 7868
rect 34424 7866 34480 7868
rect 34528 7866 34584 7868
rect 34320 7814 34324 7866
rect 34324 7814 34376 7866
rect 34424 7814 34448 7866
rect 34448 7814 34480 7866
rect 34528 7814 34572 7866
rect 34572 7814 34584 7866
rect 34320 7812 34376 7814
rect 34424 7812 34480 7814
rect 34528 7812 34584 7814
rect 34632 7866 34688 7868
rect 34736 7866 34792 7868
rect 34840 7866 34896 7868
rect 34632 7814 34644 7866
rect 34644 7814 34688 7866
rect 34736 7814 34768 7866
rect 34768 7814 34792 7866
rect 34840 7814 34892 7866
rect 34892 7814 34896 7866
rect 34632 7812 34688 7814
rect 34736 7812 34792 7814
rect 34840 7812 34896 7814
rect 34944 7812 35000 7868
rect 35048 7866 35104 7868
rect 35152 7866 35208 7868
rect 35048 7814 35068 7866
rect 35068 7814 35104 7866
rect 35152 7814 35192 7866
rect 35192 7814 35208 7866
rect 35048 7812 35104 7814
rect 35152 7812 35208 7814
rect 27804 6578 27860 6580
rect 27804 6526 27806 6578
rect 27806 6526 27858 6578
rect 27858 6526 27860 6578
rect 27804 6524 27860 6526
rect 27020 6076 27076 6132
rect 29820 6412 29876 6468
rect 28812 6130 28868 6132
rect 28812 6078 28814 6130
rect 28814 6078 28866 6130
rect 28866 6078 28868 6130
rect 28812 6076 28868 6078
rect 25900 4450 25956 4452
rect 25900 4398 25902 4450
rect 25902 4398 25954 4450
rect 25954 4398 25956 4450
rect 25900 4396 25956 4398
rect 25452 4060 25508 4116
rect 24008 3946 24064 3948
rect 24112 3946 24168 3948
rect 24008 3894 24024 3946
rect 24024 3894 24064 3946
rect 24112 3894 24148 3946
rect 24148 3894 24168 3946
rect 24008 3892 24064 3894
rect 24112 3892 24168 3894
rect 24216 3892 24272 3948
rect 24320 3946 24376 3948
rect 24424 3946 24480 3948
rect 24528 3946 24584 3948
rect 24320 3894 24324 3946
rect 24324 3894 24376 3946
rect 24424 3894 24448 3946
rect 24448 3894 24480 3946
rect 24528 3894 24572 3946
rect 24572 3894 24584 3946
rect 24320 3892 24376 3894
rect 24424 3892 24480 3894
rect 24528 3892 24584 3894
rect 24632 3946 24688 3948
rect 24736 3946 24792 3948
rect 24840 3946 24896 3948
rect 24632 3894 24644 3946
rect 24644 3894 24688 3946
rect 24736 3894 24768 3946
rect 24768 3894 24792 3946
rect 24840 3894 24892 3946
rect 24892 3894 24896 3946
rect 24632 3892 24688 3894
rect 24736 3892 24792 3894
rect 24840 3892 24896 3894
rect 24944 3892 25000 3948
rect 25048 3946 25104 3948
rect 25152 3946 25208 3948
rect 25048 3894 25068 3946
rect 25068 3894 25104 3946
rect 25152 3894 25192 3946
rect 25192 3894 25208 3946
rect 25048 3892 25104 3894
rect 25152 3892 25208 3894
rect 26572 4114 26628 4116
rect 26572 4062 26574 4114
rect 26574 4062 26626 4114
rect 26626 4062 26628 4114
rect 26572 4060 26628 4062
rect 25452 3500 25508 3556
rect 14008 3162 14064 3164
rect 14112 3162 14168 3164
rect 14008 3110 14024 3162
rect 14024 3110 14064 3162
rect 14112 3110 14148 3162
rect 14148 3110 14168 3162
rect 14008 3108 14064 3110
rect 14112 3108 14168 3110
rect 14216 3108 14272 3164
rect 14320 3162 14376 3164
rect 14424 3162 14480 3164
rect 14528 3162 14584 3164
rect 14320 3110 14324 3162
rect 14324 3110 14376 3162
rect 14424 3110 14448 3162
rect 14448 3110 14480 3162
rect 14528 3110 14572 3162
rect 14572 3110 14584 3162
rect 14320 3108 14376 3110
rect 14424 3108 14480 3110
rect 14528 3108 14584 3110
rect 14632 3162 14688 3164
rect 14736 3162 14792 3164
rect 14840 3162 14896 3164
rect 14632 3110 14644 3162
rect 14644 3110 14688 3162
rect 14736 3110 14768 3162
rect 14768 3110 14792 3162
rect 14840 3110 14892 3162
rect 14892 3110 14896 3162
rect 14632 3108 14688 3110
rect 14736 3108 14792 3110
rect 14840 3108 14896 3110
rect 14944 3108 15000 3164
rect 15048 3162 15104 3164
rect 15152 3162 15208 3164
rect 15048 3110 15068 3162
rect 15068 3110 15104 3162
rect 15152 3110 15192 3162
rect 15192 3110 15208 3162
rect 15048 3108 15104 3110
rect 15152 3108 15208 3110
rect 34008 6298 34064 6300
rect 34112 6298 34168 6300
rect 34008 6246 34024 6298
rect 34024 6246 34064 6298
rect 34112 6246 34148 6298
rect 34148 6246 34168 6298
rect 34008 6244 34064 6246
rect 34112 6244 34168 6246
rect 34216 6244 34272 6300
rect 34320 6298 34376 6300
rect 34424 6298 34480 6300
rect 34528 6298 34584 6300
rect 34320 6246 34324 6298
rect 34324 6246 34376 6298
rect 34424 6246 34448 6298
rect 34448 6246 34480 6298
rect 34528 6246 34572 6298
rect 34572 6246 34584 6298
rect 34320 6244 34376 6246
rect 34424 6244 34480 6246
rect 34528 6244 34584 6246
rect 34632 6298 34688 6300
rect 34736 6298 34792 6300
rect 34840 6298 34896 6300
rect 34632 6246 34644 6298
rect 34644 6246 34688 6298
rect 34736 6246 34768 6298
rect 34768 6246 34792 6298
rect 34840 6246 34892 6298
rect 34892 6246 34896 6298
rect 34632 6244 34688 6246
rect 34736 6244 34792 6246
rect 34840 6244 34896 6246
rect 34944 6244 35000 6300
rect 35048 6298 35104 6300
rect 35152 6298 35208 6300
rect 35048 6246 35068 6298
rect 35068 6246 35104 6298
rect 35152 6246 35192 6298
rect 35192 6246 35208 6298
rect 35048 6244 35104 6246
rect 35152 6244 35208 6246
rect 34008 4730 34064 4732
rect 34112 4730 34168 4732
rect 34008 4678 34024 4730
rect 34024 4678 34064 4730
rect 34112 4678 34148 4730
rect 34148 4678 34168 4730
rect 34008 4676 34064 4678
rect 34112 4676 34168 4678
rect 34216 4676 34272 4732
rect 34320 4730 34376 4732
rect 34424 4730 34480 4732
rect 34528 4730 34584 4732
rect 34320 4678 34324 4730
rect 34324 4678 34376 4730
rect 34424 4678 34448 4730
rect 34448 4678 34480 4730
rect 34528 4678 34572 4730
rect 34572 4678 34584 4730
rect 34320 4676 34376 4678
rect 34424 4676 34480 4678
rect 34528 4676 34584 4678
rect 34632 4730 34688 4732
rect 34736 4730 34792 4732
rect 34840 4730 34896 4732
rect 34632 4678 34644 4730
rect 34644 4678 34688 4730
rect 34736 4678 34768 4730
rect 34768 4678 34792 4730
rect 34840 4678 34892 4730
rect 34892 4678 34896 4730
rect 34632 4676 34688 4678
rect 34736 4676 34792 4678
rect 34840 4676 34896 4678
rect 34944 4676 35000 4732
rect 35048 4730 35104 4732
rect 35152 4730 35208 4732
rect 35048 4678 35068 4730
rect 35068 4678 35104 4730
rect 35152 4678 35192 4730
rect 35192 4678 35208 4730
rect 35048 4676 35104 4678
rect 35152 4676 35208 4678
rect 34008 3162 34064 3164
rect 34112 3162 34168 3164
rect 34008 3110 34024 3162
rect 34024 3110 34064 3162
rect 34112 3110 34148 3162
rect 34148 3110 34168 3162
rect 34008 3108 34064 3110
rect 34112 3108 34168 3110
rect 34216 3108 34272 3164
rect 34320 3162 34376 3164
rect 34424 3162 34480 3164
rect 34528 3162 34584 3164
rect 34320 3110 34324 3162
rect 34324 3110 34376 3162
rect 34424 3110 34448 3162
rect 34448 3110 34480 3162
rect 34528 3110 34572 3162
rect 34572 3110 34584 3162
rect 34320 3108 34376 3110
rect 34424 3108 34480 3110
rect 34528 3108 34584 3110
rect 34632 3162 34688 3164
rect 34736 3162 34792 3164
rect 34840 3162 34896 3164
rect 34632 3110 34644 3162
rect 34644 3110 34688 3162
rect 34736 3110 34768 3162
rect 34768 3110 34792 3162
rect 34840 3110 34892 3162
rect 34892 3110 34896 3162
rect 34632 3108 34688 3110
rect 34736 3108 34792 3110
rect 34840 3108 34896 3110
rect 34944 3108 35000 3164
rect 35048 3162 35104 3164
rect 35152 3162 35208 3164
rect 35048 3110 35068 3162
rect 35068 3110 35104 3162
rect 35152 3110 35192 3162
rect 35192 3110 35208 3162
rect 35048 3108 35104 3110
rect 35152 3108 35208 3110
<< metal3 >>
rect 3998 96404 4008 96460
rect 4064 96404 4112 96460
rect 4168 96404 4216 96460
rect 4272 96404 4320 96460
rect 4376 96404 4424 96460
rect 4480 96404 4528 96460
rect 4584 96404 4632 96460
rect 4688 96404 4736 96460
rect 4792 96404 4840 96460
rect 4896 96404 4944 96460
rect 5000 96404 5048 96460
rect 5104 96404 5152 96460
rect 5208 96404 5218 96460
rect 23998 96404 24008 96460
rect 24064 96404 24112 96460
rect 24168 96404 24216 96460
rect 24272 96404 24320 96460
rect 24376 96404 24424 96460
rect 24480 96404 24528 96460
rect 24584 96404 24632 96460
rect 24688 96404 24736 96460
rect 24792 96404 24840 96460
rect 24896 96404 24944 96460
rect 25000 96404 25048 96460
rect 25104 96404 25152 96460
rect 25208 96404 25218 96460
rect 13998 95620 14008 95676
rect 14064 95620 14112 95676
rect 14168 95620 14216 95676
rect 14272 95620 14320 95676
rect 14376 95620 14424 95676
rect 14480 95620 14528 95676
rect 14584 95620 14632 95676
rect 14688 95620 14736 95676
rect 14792 95620 14840 95676
rect 14896 95620 14944 95676
rect 15000 95620 15048 95676
rect 15104 95620 15152 95676
rect 15208 95620 15218 95676
rect 33998 95620 34008 95676
rect 34064 95620 34112 95676
rect 34168 95620 34216 95676
rect 34272 95620 34320 95676
rect 34376 95620 34424 95676
rect 34480 95620 34528 95676
rect 34584 95620 34632 95676
rect 34688 95620 34736 95676
rect 34792 95620 34840 95676
rect 34896 95620 34944 95676
rect 35000 95620 35048 95676
rect 35104 95620 35152 95676
rect 35208 95620 35218 95676
rect 0 95284 800 95312
rect 0 95228 1708 95284
rect 1764 95228 1774 95284
rect 0 95200 800 95228
rect 3998 94836 4008 94892
rect 4064 94836 4112 94892
rect 4168 94836 4216 94892
rect 4272 94836 4320 94892
rect 4376 94836 4424 94892
rect 4480 94836 4528 94892
rect 4584 94836 4632 94892
rect 4688 94836 4736 94892
rect 4792 94836 4840 94892
rect 4896 94836 4944 94892
rect 5000 94836 5048 94892
rect 5104 94836 5152 94892
rect 5208 94836 5218 94892
rect 23998 94836 24008 94892
rect 24064 94836 24112 94892
rect 24168 94836 24216 94892
rect 24272 94836 24320 94892
rect 24376 94836 24424 94892
rect 24480 94836 24528 94892
rect 24584 94836 24632 94892
rect 24688 94836 24736 94892
rect 24792 94836 24840 94892
rect 24896 94836 24944 94892
rect 25000 94836 25048 94892
rect 25104 94836 25152 94892
rect 25208 94836 25218 94892
rect 1698 94220 1708 94276
rect 1764 94220 1774 94276
rect 0 94164 800 94192
rect 1708 94164 1764 94220
rect 0 94108 1764 94164
rect 9874 94108 9884 94164
rect 9940 94108 12908 94164
rect 12964 94108 12974 94164
rect 0 94080 800 94108
rect 13998 94052 14008 94108
rect 14064 94052 14112 94108
rect 14168 94052 14216 94108
rect 14272 94052 14320 94108
rect 14376 94052 14424 94108
rect 14480 94052 14528 94108
rect 14584 94052 14632 94108
rect 14688 94052 14736 94108
rect 14792 94052 14840 94108
rect 14896 94052 14944 94108
rect 15000 94052 15048 94108
rect 15104 94052 15152 94108
rect 15208 94052 15218 94108
rect 33998 94052 34008 94108
rect 34064 94052 34112 94108
rect 34168 94052 34216 94108
rect 34272 94052 34320 94108
rect 34376 94052 34424 94108
rect 34480 94052 34528 94108
rect 34584 94052 34632 94108
rect 34688 94052 34736 94108
rect 34792 94052 34840 94108
rect 34896 94052 34944 94108
rect 35000 94052 35048 94108
rect 35104 94052 35152 94108
rect 35208 94052 35218 94108
rect 3998 93268 4008 93324
rect 4064 93268 4112 93324
rect 4168 93268 4216 93324
rect 4272 93268 4320 93324
rect 4376 93268 4424 93324
rect 4480 93268 4528 93324
rect 4584 93268 4632 93324
rect 4688 93268 4736 93324
rect 4792 93268 4840 93324
rect 4896 93268 4944 93324
rect 5000 93268 5048 93324
rect 5104 93268 5152 93324
rect 5208 93268 5218 93324
rect 23998 93268 24008 93324
rect 24064 93268 24112 93324
rect 24168 93268 24216 93324
rect 24272 93268 24320 93324
rect 24376 93268 24424 93324
rect 24480 93268 24528 93324
rect 24584 93268 24632 93324
rect 24688 93268 24736 93324
rect 24792 93268 24840 93324
rect 24896 93268 24944 93324
rect 25000 93268 25048 93324
rect 25104 93268 25152 93324
rect 25208 93268 25218 93324
rect 0 93044 800 93072
rect 0 92988 1708 93044
rect 1764 92988 1774 93044
rect 0 92960 800 92988
rect 13998 92484 14008 92540
rect 14064 92484 14112 92540
rect 14168 92484 14216 92540
rect 14272 92484 14320 92540
rect 14376 92484 14424 92540
rect 14480 92484 14528 92540
rect 14584 92484 14632 92540
rect 14688 92484 14736 92540
rect 14792 92484 14840 92540
rect 14896 92484 14944 92540
rect 15000 92484 15048 92540
rect 15104 92484 15152 92540
rect 15208 92484 15218 92540
rect 33998 92484 34008 92540
rect 34064 92484 34112 92540
rect 34168 92484 34216 92540
rect 34272 92484 34320 92540
rect 34376 92484 34424 92540
rect 34480 92484 34528 92540
rect 34584 92484 34632 92540
rect 34688 92484 34736 92540
rect 34792 92484 34840 92540
rect 34896 92484 34944 92540
rect 35000 92484 35048 92540
rect 35104 92484 35152 92540
rect 35208 92484 35218 92540
rect 0 91924 800 91952
rect 0 91868 1708 91924
rect 1764 91868 1774 91924
rect 0 91840 800 91868
rect 3998 91700 4008 91756
rect 4064 91700 4112 91756
rect 4168 91700 4216 91756
rect 4272 91700 4320 91756
rect 4376 91700 4424 91756
rect 4480 91700 4528 91756
rect 4584 91700 4632 91756
rect 4688 91700 4736 91756
rect 4792 91700 4840 91756
rect 4896 91700 4944 91756
rect 5000 91700 5048 91756
rect 5104 91700 5152 91756
rect 5208 91700 5218 91756
rect 23998 91700 24008 91756
rect 24064 91700 24112 91756
rect 24168 91700 24216 91756
rect 24272 91700 24320 91756
rect 24376 91700 24424 91756
rect 24480 91700 24528 91756
rect 24584 91700 24632 91756
rect 24688 91700 24736 91756
rect 24792 91700 24840 91756
rect 24896 91700 24944 91756
rect 25000 91700 25048 91756
rect 25104 91700 25152 91756
rect 25208 91700 25218 91756
rect 13998 90916 14008 90972
rect 14064 90916 14112 90972
rect 14168 90916 14216 90972
rect 14272 90916 14320 90972
rect 14376 90916 14424 90972
rect 14480 90916 14528 90972
rect 14584 90916 14632 90972
rect 14688 90916 14736 90972
rect 14792 90916 14840 90972
rect 14896 90916 14944 90972
rect 15000 90916 15048 90972
rect 15104 90916 15152 90972
rect 15208 90916 15218 90972
rect 33998 90916 34008 90972
rect 34064 90916 34112 90972
rect 34168 90916 34216 90972
rect 34272 90916 34320 90972
rect 34376 90916 34424 90972
rect 34480 90916 34528 90972
rect 34584 90916 34632 90972
rect 34688 90916 34736 90972
rect 34792 90916 34840 90972
rect 34896 90916 34944 90972
rect 35000 90916 35048 90972
rect 35104 90916 35152 90972
rect 35208 90916 35218 90972
rect 0 90804 800 90832
rect 0 90748 1708 90804
rect 1764 90748 1774 90804
rect 0 90720 800 90748
rect 3998 90132 4008 90188
rect 4064 90132 4112 90188
rect 4168 90132 4216 90188
rect 4272 90132 4320 90188
rect 4376 90132 4424 90188
rect 4480 90132 4528 90188
rect 4584 90132 4632 90188
rect 4688 90132 4736 90188
rect 4792 90132 4840 90188
rect 4896 90132 4944 90188
rect 5000 90132 5048 90188
rect 5104 90132 5152 90188
rect 5208 90132 5218 90188
rect 23998 90132 24008 90188
rect 24064 90132 24112 90188
rect 24168 90132 24216 90188
rect 24272 90132 24320 90188
rect 24376 90132 24424 90188
rect 24480 90132 24528 90188
rect 24584 90132 24632 90188
rect 24688 90132 24736 90188
rect 24792 90132 24840 90188
rect 24896 90132 24944 90188
rect 25000 90132 25048 90188
rect 25104 90132 25152 90188
rect 25208 90132 25218 90188
rect 0 89684 800 89712
rect 0 89628 1708 89684
rect 1764 89628 1774 89684
rect 0 89600 800 89628
rect 13998 89348 14008 89404
rect 14064 89348 14112 89404
rect 14168 89348 14216 89404
rect 14272 89348 14320 89404
rect 14376 89348 14424 89404
rect 14480 89348 14528 89404
rect 14584 89348 14632 89404
rect 14688 89348 14736 89404
rect 14792 89348 14840 89404
rect 14896 89348 14944 89404
rect 15000 89348 15048 89404
rect 15104 89348 15152 89404
rect 15208 89348 15218 89404
rect 33998 89348 34008 89404
rect 34064 89348 34112 89404
rect 34168 89348 34216 89404
rect 34272 89348 34320 89404
rect 34376 89348 34424 89404
rect 34480 89348 34528 89404
rect 34584 89348 34632 89404
rect 34688 89348 34736 89404
rect 34792 89348 34840 89404
rect 34896 89348 34944 89404
rect 35000 89348 35048 89404
rect 35104 89348 35152 89404
rect 35208 89348 35218 89404
rect 12338 88844 12348 88900
rect 12404 88844 13916 88900
rect 13972 88844 14252 88900
rect 14308 88844 14318 88900
rect 0 88564 800 88592
rect 3998 88564 4008 88620
rect 4064 88564 4112 88620
rect 4168 88564 4216 88620
rect 4272 88564 4320 88620
rect 4376 88564 4424 88620
rect 4480 88564 4528 88620
rect 4584 88564 4632 88620
rect 4688 88564 4736 88620
rect 4792 88564 4840 88620
rect 4896 88564 4944 88620
rect 5000 88564 5048 88620
rect 5104 88564 5152 88620
rect 5208 88564 5218 88620
rect 23998 88564 24008 88620
rect 24064 88564 24112 88620
rect 24168 88564 24216 88620
rect 24272 88564 24320 88620
rect 24376 88564 24424 88620
rect 24480 88564 24528 88620
rect 24584 88564 24632 88620
rect 24688 88564 24736 88620
rect 24792 88564 24840 88620
rect 24896 88564 24944 88620
rect 25000 88564 25048 88620
rect 25104 88564 25152 88620
rect 25208 88564 25218 88620
rect 0 88508 1708 88564
rect 1764 88508 1774 88564
rect 0 88480 800 88508
rect 9762 88172 9772 88228
rect 9828 88172 10332 88228
rect 10388 88172 10398 88228
rect 13234 88172 13244 88228
rect 13300 88172 13916 88228
rect 13972 88172 13982 88228
rect 14690 88060 14700 88116
rect 14756 88060 15596 88116
rect 15652 88060 15662 88116
rect 8418 87948 8428 88004
rect 8484 87948 10444 88004
rect 10500 87948 12012 88004
rect 12068 87948 12078 88004
rect 12562 87948 12572 88004
rect 12628 87948 13580 88004
rect 13636 87948 13646 88004
rect 14242 87948 14252 88004
rect 14308 87948 17276 88004
rect 17332 87948 17342 88004
rect 13998 87780 14008 87836
rect 14064 87780 14112 87836
rect 14168 87780 14216 87836
rect 14272 87780 14320 87836
rect 14376 87780 14424 87836
rect 14480 87780 14528 87836
rect 14584 87780 14632 87836
rect 14688 87780 14736 87836
rect 14792 87780 14840 87836
rect 14896 87780 14944 87836
rect 15000 87780 15048 87836
rect 15104 87780 15152 87836
rect 15208 87780 15218 87836
rect 33998 87780 34008 87836
rect 34064 87780 34112 87836
rect 34168 87780 34216 87836
rect 34272 87780 34320 87836
rect 34376 87780 34424 87836
rect 34480 87780 34528 87836
rect 34584 87780 34632 87836
rect 34688 87780 34736 87836
rect 34792 87780 34840 87836
rect 34896 87780 34944 87836
rect 35000 87780 35048 87836
rect 35104 87780 35152 87836
rect 35208 87780 35218 87836
rect 15362 87724 15372 87780
rect 15428 87724 16436 87780
rect 16380 87668 16436 87724
rect 9874 87612 9884 87668
rect 9940 87612 11452 87668
rect 11508 87612 15876 87668
rect 16370 87612 16380 87668
rect 16436 87612 16716 87668
rect 16772 87612 20412 87668
rect 20468 87612 20478 87668
rect 15820 87556 15876 87612
rect 15820 87500 20524 87556
rect 20580 87500 20590 87556
rect 0 87444 800 87472
rect 0 87388 1708 87444
rect 1764 87388 1774 87444
rect 5618 87388 5628 87444
rect 5684 87388 6524 87444
rect 6580 87388 8876 87444
rect 8932 87388 8942 87444
rect 19394 87388 19404 87444
rect 19460 87388 20972 87444
rect 21028 87388 21038 87444
rect 0 87360 800 87388
rect 16930 87276 16940 87332
rect 16996 87276 17388 87332
rect 17444 87276 17454 87332
rect 20402 87276 20412 87332
rect 20468 87276 21308 87332
rect 21364 87276 21374 87332
rect 10658 87164 10668 87220
rect 10724 87164 12796 87220
rect 12852 87164 12862 87220
rect 3998 86996 4008 87052
rect 4064 86996 4112 87052
rect 4168 86996 4216 87052
rect 4272 86996 4320 87052
rect 4376 86996 4424 87052
rect 4480 86996 4528 87052
rect 4584 86996 4632 87052
rect 4688 86996 4736 87052
rect 4792 86996 4840 87052
rect 4896 86996 4944 87052
rect 5000 86996 5048 87052
rect 5104 86996 5152 87052
rect 5208 86996 5218 87052
rect 23998 86996 24008 87052
rect 24064 86996 24112 87052
rect 24168 86996 24216 87052
rect 24272 86996 24320 87052
rect 24376 86996 24424 87052
rect 24480 86996 24528 87052
rect 24584 86996 24632 87052
rect 24688 86996 24736 87052
rect 24792 86996 24840 87052
rect 24896 86996 24944 87052
rect 25000 86996 25048 87052
rect 25104 86996 25152 87052
rect 25208 86996 25218 87052
rect 6066 86828 6076 86884
rect 6132 86828 7644 86884
rect 7700 86828 7710 86884
rect 8754 86604 8764 86660
rect 8820 86604 9324 86660
rect 9380 86604 9884 86660
rect 9940 86604 10892 86660
rect 10948 86604 12460 86660
rect 12516 86604 12526 86660
rect 12898 86604 12908 86660
rect 12964 86604 13580 86660
rect 13636 86604 13646 86660
rect 13794 86604 13804 86660
rect 13860 86604 14364 86660
rect 14420 86604 16044 86660
rect 16100 86604 16110 86660
rect 7298 86492 7308 86548
rect 7364 86492 8540 86548
rect 8596 86492 8606 86548
rect 10210 86492 10220 86548
rect 10276 86492 11004 86548
rect 11060 86492 11900 86548
rect 11956 86492 11966 86548
rect 1698 86380 1708 86436
rect 1764 86380 1774 86436
rect 7970 86380 7980 86436
rect 8036 86380 9100 86436
rect 9156 86380 11116 86436
rect 11172 86380 11182 86436
rect 0 86324 800 86352
rect 1708 86324 1764 86380
rect 0 86268 1764 86324
rect 0 86240 800 86268
rect 13998 86212 14008 86268
rect 14064 86212 14112 86268
rect 14168 86212 14216 86268
rect 14272 86212 14320 86268
rect 14376 86212 14424 86268
rect 14480 86212 14528 86268
rect 14584 86212 14632 86268
rect 14688 86212 14736 86268
rect 14792 86212 14840 86268
rect 14896 86212 14944 86268
rect 15000 86212 15048 86268
rect 15104 86212 15152 86268
rect 15208 86212 15218 86268
rect 33998 86212 34008 86268
rect 34064 86212 34112 86268
rect 34168 86212 34216 86268
rect 34272 86212 34320 86268
rect 34376 86212 34424 86268
rect 34480 86212 34528 86268
rect 34584 86212 34632 86268
rect 34688 86212 34736 86268
rect 34792 86212 34840 86268
rect 34896 86212 34944 86268
rect 35000 86212 35048 86268
rect 35104 86212 35152 86268
rect 35208 86212 35218 86268
rect 8530 86156 8540 86212
rect 8596 86156 13580 86212
rect 13636 86156 13646 86212
rect 9650 86044 9660 86100
rect 9716 86044 10220 86100
rect 10276 86044 18284 86100
rect 18340 86044 18350 86100
rect 21298 86044 21308 86100
rect 21364 86044 21374 86100
rect 21308 85988 21364 86044
rect 16594 85932 16604 85988
rect 16660 85932 18060 85988
rect 18116 85932 18126 85988
rect 21308 85932 23100 85988
rect 23156 85932 23996 85988
rect 24052 85932 24062 85988
rect 12338 85820 12348 85876
rect 12404 85820 13468 85876
rect 13524 85820 13804 85876
rect 13860 85820 14140 85876
rect 14196 85820 14206 85876
rect 14466 85820 14476 85876
rect 14532 85820 15036 85876
rect 15092 85820 15102 85876
rect 20066 85820 20076 85876
rect 20132 85820 23884 85876
rect 23940 85820 24556 85876
rect 24612 85820 24622 85876
rect 13570 85708 13580 85764
rect 13636 85708 14252 85764
rect 14308 85708 14318 85764
rect 14802 85708 14812 85764
rect 14868 85708 15372 85764
rect 15428 85708 16156 85764
rect 16212 85708 16828 85764
rect 16884 85708 18620 85764
rect 18676 85708 18956 85764
rect 19012 85708 20188 85764
rect 22530 85708 22540 85764
rect 22596 85708 23660 85764
rect 23716 85708 23726 85764
rect 23986 85708 23996 85764
rect 24052 85708 25340 85764
rect 25396 85708 25406 85764
rect 20132 85540 20188 85708
rect 13682 85484 13692 85540
rect 13748 85484 14812 85540
rect 14868 85484 14878 85540
rect 20132 85484 20748 85540
rect 20804 85484 20814 85540
rect 3998 85428 4008 85484
rect 4064 85428 4112 85484
rect 4168 85428 4216 85484
rect 4272 85428 4320 85484
rect 4376 85428 4424 85484
rect 4480 85428 4528 85484
rect 4584 85428 4632 85484
rect 4688 85428 4736 85484
rect 4792 85428 4840 85484
rect 4896 85428 4944 85484
rect 5000 85428 5048 85484
rect 5104 85428 5152 85484
rect 5208 85428 5218 85484
rect 23998 85428 24008 85484
rect 24064 85428 24112 85484
rect 24168 85428 24216 85484
rect 24272 85428 24320 85484
rect 24376 85428 24424 85484
rect 24480 85428 24528 85484
rect 24584 85428 24632 85484
rect 24688 85428 24736 85484
rect 24792 85428 24840 85484
rect 24896 85428 24944 85484
rect 25000 85428 25048 85484
rect 25104 85428 25152 85484
rect 25208 85428 25218 85484
rect 0 85204 800 85232
rect 0 85148 1708 85204
rect 1764 85148 1774 85204
rect 4834 85148 4844 85204
rect 4900 85148 5404 85204
rect 5460 85148 13692 85204
rect 13748 85148 13758 85204
rect 14242 85148 14252 85204
rect 14308 85148 15372 85204
rect 15428 85148 15438 85204
rect 0 85120 800 85148
rect 3826 85036 3836 85092
rect 3892 85036 6524 85092
rect 6580 85036 7196 85092
rect 7252 85036 7262 85092
rect 6738 84924 6748 84980
rect 6804 84924 9212 84980
rect 9268 84924 10444 84980
rect 10500 84924 10510 84980
rect 13682 84924 13692 84980
rect 13748 84924 13916 84980
rect 13972 84924 13982 84980
rect 20738 84924 20748 84980
rect 20804 84924 21980 84980
rect 22036 84924 22046 84980
rect 13010 84812 13020 84868
rect 13076 84812 14476 84868
rect 14532 84812 18172 84868
rect 18228 84812 19292 84868
rect 19348 84812 20300 84868
rect 20356 84812 20366 84868
rect 13998 84644 14008 84700
rect 14064 84644 14112 84700
rect 14168 84644 14216 84700
rect 14272 84644 14320 84700
rect 14376 84644 14424 84700
rect 14480 84644 14528 84700
rect 14584 84644 14632 84700
rect 14688 84644 14736 84700
rect 14792 84644 14840 84700
rect 14896 84644 14944 84700
rect 15000 84644 15048 84700
rect 15104 84644 15152 84700
rect 15208 84644 15218 84700
rect 33998 84644 34008 84700
rect 34064 84644 34112 84700
rect 34168 84644 34216 84700
rect 34272 84644 34320 84700
rect 34376 84644 34424 84700
rect 34480 84644 34528 84700
rect 34584 84644 34632 84700
rect 34688 84644 34736 84700
rect 34792 84644 34840 84700
rect 34896 84644 34944 84700
rect 35000 84644 35048 84700
rect 35104 84644 35152 84700
rect 35208 84644 35218 84700
rect 6962 84476 6972 84532
rect 7028 84476 8316 84532
rect 8372 84476 8382 84532
rect 14578 84476 14588 84532
rect 14644 84476 15596 84532
rect 15652 84476 15662 84532
rect 14466 84364 14476 84420
rect 14532 84364 15036 84420
rect 15092 84364 15102 84420
rect 11778 84252 11788 84308
rect 11844 84252 12572 84308
rect 12628 84252 13020 84308
rect 13076 84252 13692 84308
rect 13748 84252 13758 84308
rect 20290 84252 20300 84308
rect 20356 84252 20972 84308
rect 21028 84252 21038 84308
rect 16482 84140 16492 84196
rect 16548 84140 16716 84196
rect 16772 84140 17500 84196
rect 17556 84140 17566 84196
rect 20626 84140 20636 84196
rect 20692 84140 21756 84196
rect 21812 84140 21822 84196
rect 0 84084 800 84112
rect 0 84028 1708 84084
rect 1764 84028 1774 84084
rect 5842 84028 5852 84084
rect 5908 84028 6860 84084
rect 6916 84028 13580 84084
rect 13636 84028 13646 84084
rect 18274 84028 18284 84084
rect 18340 84028 19068 84084
rect 19124 84028 19292 84084
rect 19348 84028 19358 84084
rect 0 84000 800 84028
rect 3998 83860 4008 83916
rect 4064 83860 4112 83916
rect 4168 83860 4216 83916
rect 4272 83860 4320 83916
rect 4376 83860 4424 83916
rect 4480 83860 4528 83916
rect 4584 83860 4632 83916
rect 4688 83860 4736 83916
rect 4792 83860 4840 83916
rect 4896 83860 4944 83916
rect 5000 83860 5048 83916
rect 5104 83860 5152 83916
rect 5208 83860 5218 83916
rect 23998 83860 24008 83916
rect 24064 83860 24112 83916
rect 24168 83860 24216 83916
rect 24272 83860 24320 83916
rect 24376 83860 24424 83916
rect 24480 83860 24528 83916
rect 24584 83860 24632 83916
rect 24688 83860 24736 83916
rect 24792 83860 24840 83916
rect 24896 83860 24944 83916
rect 25000 83860 25048 83916
rect 25104 83860 25152 83916
rect 25208 83860 25218 83916
rect 3826 83692 3836 83748
rect 3892 83692 5964 83748
rect 6020 83692 6030 83748
rect 6290 83692 6300 83748
rect 6356 83692 7308 83748
rect 7364 83692 10220 83748
rect 10276 83692 10892 83748
rect 10948 83692 10958 83748
rect 18722 83692 18732 83748
rect 18788 83692 19628 83748
rect 19684 83692 19694 83748
rect 5618 83580 5628 83636
rect 5684 83580 22316 83636
rect 22372 83580 22382 83636
rect 4274 83468 4284 83524
rect 4340 83468 5404 83524
rect 5460 83468 5470 83524
rect 13458 83468 13468 83524
rect 13524 83468 15932 83524
rect 15988 83468 15998 83524
rect 18274 83468 18284 83524
rect 18340 83468 18956 83524
rect 19012 83468 19022 83524
rect 4498 83356 4508 83412
rect 4564 83356 5292 83412
rect 5348 83356 5358 83412
rect 8194 83356 8204 83412
rect 8260 83356 8764 83412
rect 8820 83356 8830 83412
rect 14466 83356 14476 83412
rect 14532 83356 15260 83412
rect 15316 83356 15326 83412
rect 18386 83356 18396 83412
rect 18452 83356 19068 83412
rect 19124 83356 19134 83412
rect 2258 83244 2268 83300
rect 2324 83244 3388 83300
rect 3444 83244 3454 83300
rect 7074 83244 7084 83300
rect 7140 83244 7644 83300
rect 7700 83244 8428 83300
rect 8484 83244 9212 83300
rect 9268 83244 9278 83300
rect 13794 83244 13804 83300
rect 13860 83244 14028 83300
rect 14084 83244 14094 83300
rect 16258 83244 16268 83300
rect 16324 83244 17052 83300
rect 17108 83244 17118 83300
rect 22530 83244 22540 83300
rect 22596 83244 22876 83300
rect 22932 83244 22942 83300
rect 13654 83132 13692 83188
rect 13748 83132 13758 83188
rect 13998 83076 14008 83132
rect 14064 83076 14112 83132
rect 14168 83076 14216 83132
rect 14272 83076 14320 83132
rect 14376 83076 14424 83132
rect 14480 83076 14528 83132
rect 14584 83076 14632 83132
rect 14688 83076 14736 83132
rect 14792 83076 14840 83132
rect 14896 83076 14944 83132
rect 15000 83076 15048 83132
rect 15104 83076 15152 83132
rect 15208 83076 15218 83132
rect 33998 83076 34008 83132
rect 34064 83076 34112 83132
rect 34168 83076 34216 83132
rect 34272 83076 34320 83132
rect 34376 83076 34424 83132
rect 34480 83076 34528 83132
rect 34584 83076 34632 83132
rect 34688 83076 34736 83132
rect 34792 83076 34840 83132
rect 34896 83076 34944 83132
rect 35000 83076 35048 83132
rect 35104 83076 35152 83132
rect 35208 83076 35218 83132
rect 0 82964 800 82992
rect 0 82908 1708 82964
rect 1764 82908 1774 82964
rect 12562 82908 12572 82964
rect 12628 82908 15148 82964
rect 15204 82908 15214 82964
rect 0 82880 800 82908
rect 4722 82796 4732 82852
rect 4788 82796 5068 82852
rect 5124 82796 8204 82852
rect 8260 82796 8270 82852
rect 13010 82796 13020 82852
rect 13076 82796 15260 82852
rect 15316 82796 15708 82852
rect 15764 82796 16268 82852
rect 16324 82796 16334 82852
rect 10658 82684 10668 82740
rect 10724 82684 12796 82740
rect 12852 82684 12862 82740
rect 13794 82684 13804 82740
rect 13860 82684 14140 82740
rect 14196 82684 14206 82740
rect 14466 82684 14476 82740
rect 14532 82684 15372 82740
rect 15428 82684 15438 82740
rect 16818 82684 16828 82740
rect 16884 82684 17612 82740
rect 17668 82684 17678 82740
rect 23874 82684 23884 82740
rect 23940 82684 24556 82740
rect 24612 82684 25788 82740
rect 25844 82684 25854 82740
rect 6290 82572 6300 82628
rect 6356 82572 6636 82628
rect 6692 82572 11788 82628
rect 11844 82572 12572 82628
rect 12628 82572 13356 82628
rect 13412 82572 13422 82628
rect 6402 82460 6412 82516
rect 6468 82460 8764 82516
rect 8820 82460 10220 82516
rect 10276 82460 10286 82516
rect 15586 82460 15596 82516
rect 15652 82460 17836 82516
rect 17892 82460 18732 82516
rect 18788 82460 20636 82516
rect 20692 82460 20702 82516
rect 21074 82460 21084 82516
rect 21140 82460 22092 82516
rect 22148 82460 22158 82516
rect 22418 82460 22428 82516
rect 22484 82460 24108 82516
rect 24164 82460 24174 82516
rect 21084 82404 21140 82460
rect 5292 82348 6188 82404
rect 6244 82348 6254 82404
rect 6748 82348 7644 82404
rect 7700 82348 9436 82404
rect 9492 82348 10332 82404
rect 10388 82348 10398 82404
rect 15922 82348 15932 82404
rect 15988 82348 16716 82404
rect 16772 82348 16782 82404
rect 18060 82348 21140 82404
rect 3998 82292 4008 82348
rect 4064 82292 4112 82348
rect 4168 82292 4216 82348
rect 4272 82292 4320 82348
rect 4376 82292 4424 82348
rect 4480 82292 4528 82348
rect 4584 82292 4632 82348
rect 4688 82292 4736 82348
rect 4792 82292 4840 82348
rect 4896 82292 4944 82348
rect 5000 82292 5048 82348
rect 5104 82292 5152 82348
rect 5208 82292 5218 82348
rect 5292 82180 5348 82348
rect 6748 82292 6804 82348
rect 11218 82292 11228 82348
rect 11284 82292 11294 82348
rect 18060 82292 18116 82348
rect 23998 82292 24008 82348
rect 24064 82292 24112 82348
rect 24168 82292 24216 82348
rect 24272 82292 24320 82348
rect 24376 82292 24424 82348
rect 24480 82292 24528 82348
rect 24584 82292 24632 82348
rect 24688 82292 24736 82348
rect 24792 82292 24840 82348
rect 24896 82292 24944 82348
rect 25000 82292 25048 82348
rect 25104 82292 25152 82348
rect 25208 82292 25218 82348
rect 5842 82236 5852 82292
rect 5908 82236 6300 82292
rect 6356 82236 6804 82292
rect 11228 82180 11284 82292
rect 15138 82236 15148 82292
rect 15204 82236 16492 82292
rect 16548 82236 18060 82292
rect 18116 82236 18126 82292
rect 4834 82124 4844 82180
rect 4900 82124 5348 82180
rect 10966 82124 11004 82180
rect 11060 82124 11070 82180
rect 11228 82124 11900 82180
rect 11956 82124 11966 82180
rect 15148 82124 15372 82180
rect 15428 82124 15438 82180
rect 20066 82124 20076 82180
rect 20132 82124 21420 82180
rect 21476 82124 21868 82180
rect 21924 82124 25340 82180
rect 25396 82124 25406 82180
rect 3602 82012 3612 82068
rect 3668 82012 4508 82068
rect 4564 82012 4574 82068
rect 10434 82012 10444 82068
rect 10500 82012 12348 82068
rect 12404 82012 12414 82068
rect 13804 82012 14476 82068
rect 14532 82012 14542 82068
rect 13804 81956 13860 82012
rect 15148 81956 15204 82124
rect 13794 81900 13804 81956
rect 13860 81900 13870 81956
rect 14354 81900 14364 81956
rect 14420 81900 15204 81956
rect 16258 81900 16268 81956
rect 16324 81900 16716 81956
rect 16772 81900 18956 81956
rect 19012 81900 19022 81956
rect 0 81844 800 81872
rect 0 81788 1708 81844
rect 1764 81788 1774 81844
rect 11442 81788 11452 81844
rect 11508 81788 13468 81844
rect 13524 81788 13692 81844
rect 13748 81788 13758 81844
rect 14018 81788 14028 81844
rect 14084 81788 14812 81844
rect 14868 81788 15484 81844
rect 15540 81788 16156 81844
rect 16212 81788 17052 81844
rect 17108 81788 17118 81844
rect 0 81760 800 81788
rect 4386 81676 4396 81732
rect 4452 81676 5180 81732
rect 5236 81676 6636 81732
rect 6692 81676 6702 81732
rect 13804 81676 14700 81732
rect 14756 81676 14766 81732
rect 15250 81676 15260 81732
rect 15316 81676 15764 81732
rect 16482 81676 16492 81732
rect 16548 81676 18844 81732
rect 18900 81676 18910 81732
rect 21970 81676 21980 81732
rect 22036 81676 22540 81732
rect 22596 81676 22606 81732
rect 10182 81452 10220 81508
rect 10276 81452 10286 81508
rect 13804 81284 13860 81676
rect 13998 81508 14008 81564
rect 14064 81508 14112 81564
rect 14168 81508 14216 81564
rect 14272 81508 14320 81564
rect 14376 81508 14424 81564
rect 14480 81508 14528 81564
rect 14584 81508 14632 81564
rect 14688 81508 14736 81564
rect 14792 81508 14840 81564
rect 14896 81508 14944 81564
rect 15000 81508 15048 81564
rect 15104 81508 15152 81564
rect 15208 81508 15218 81564
rect 14690 81340 14700 81396
rect 14756 81340 15484 81396
rect 15540 81340 15550 81396
rect 15708 81284 15764 81676
rect 33998 81508 34008 81564
rect 34064 81508 34112 81564
rect 34168 81508 34216 81564
rect 34272 81508 34320 81564
rect 34376 81508 34424 81564
rect 34480 81508 34528 81564
rect 34584 81508 34632 81564
rect 34688 81508 34736 81564
rect 34792 81508 34840 81564
rect 34896 81508 34944 81564
rect 35000 81508 35048 81564
rect 35104 81508 35152 81564
rect 35208 81508 35218 81564
rect 16482 81452 16492 81508
rect 16548 81452 17724 81508
rect 17780 81452 17790 81508
rect 16034 81340 16044 81396
rect 16100 81340 16716 81396
rect 16772 81340 16782 81396
rect 13804 81228 15036 81284
rect 15092 81228 15102 81284
rect 15250 81228 15260 81284
rect 15316 81228 15764 81284
rect 17042 81228 17052 81284
rect 17108 81228 18284 81284
rect 18340 81228 18350 81284
rect 9762 81116 9772 81172
rect 9828 81116 11676 81172
rect 11732 81116 11742 81172
rect 14130 81116 14140 81172
rect 14196 81116 16492 81172
rect 16548 81116 16558 81172
rect 16706 81116 16716 81172
rect 16772 81116 17388 81172
rect 17444 81116 17454 81172
rect 4610 81004 4620 81060
rect 4676 81004 9884 81060
rect 9940 81004 9950 81060
rect 10658 81004 10668 81060
rect 10724 81004 12124 81060
rect 12180 81004 12190 81060
rect 13794 81004 13804 81060
rect 13860 81004 13916 81060
rect 13972 81004 13982 81060
rect 14578 81004 14588 81060
rect 14644 81004 16380 81060
rect 16436 81004 18060 81060
rect 18116 81004 18126 81060
rect 19170 81004 19180 81060
rect 19236 81004 20076 81060
rect 20132 81004 22316 81060
rect 22372 81004 23660 81060
rect 23716 81004 23726 81060
rect 5506 80892 5516 80948
rect 5572 80892 5964 80948
rect 6020 80892 6030 80948
rect 9884 80836 9940 81004
rect 12786 80892 12796 80948
rect 12852 80892 16716 80948
rect 16772 80892 16782 80948
rect 18834 80892 18844 80948
rect 18900 80892 19292 80948
rect 19348 80892 20524 80948
rect 20580 80892 21980 80948
rect 22036 80892 22046 80948
rect 9884 80780 11004 80836
rect 11060 80780 11070 80836
rect 0 80724 800 80752
rect 3998 80724 4008 80780
rect 4064 80724 4112 80780
rect 4168 80724 4216 80780
rect 4272 80724 4320 80780
rect 4376 80724 4424 80780
rect 4480 80724 4528 80780
rect 4584 80724 4632 80780
rect 4688 80724 4736 80780
rect 4792 80724 4840 80780
rect 4896 80724 4944 80780
rect 5000 80724 5048 80780
rect 5104 80724 5152 80780
rect 5208 80724 5218 80780
rect 23998 80724 24008 80780
rect 24064 80724 24112 80780
rect 24168 80724 24216 80780
rect 24272 80724 24320 80780
rect 24376 80724 24424 80780
rect 24480 80724 24528 80780
rect 24584 80724 24632 80780
rect 24688 80724 24736 80780
rect 24792 80724 24840 80780
rect 24896 80724 24944 80780
rect 25000 80724 25048 80780
rect 25104 80724 25152 80780
rect 25208 80724 25218 80780
rect 0 80668 1708 80724
rect 1764 80668 1774 80724
rect 10322 80668 10332 80724
rect 10388 80668 10780 80724
rect 10836 80668 10846 80724
rect 0 80640 800 80668
rect 1810 80556 1820 80612
rect 1876 80556 5628 80612
rect 5684 80556 5694 80612
rect 14466 80556 14476 80612
rect 14532 80556 15484 80612
rect 15540 80556 15550 80612
rect 18274 80556 18284 80612
rect 18340 80556 19404 80612
rect 19460 80556 19470 80612
rect 10098 80444 10108 80500
rect 10164 80444 11004 80500
rect 11060 80444 11070 80500
rect 13906 80444 13916 80500
rect 13972 80444 14700 80500
rect 14756 80444 17500 80500
rect 17556 80444 19180 80500
rect 19236 80444 19246 80500
rect 6066 80332 6076 80388
rect 6132 80332 7308 80388
rect 7364 80332 7374 80388
rect 10546 80332 10556 80388
rect 10612 80332 11900 80388
rect 11956 80332 11966 80388
rect 14354 80332 14364 80388
rect 14420 80332 15372 80388
rect 15428 80332 15820 80388
rect 15876 80332 15886 80388
rect 6738 80220 6748 80276
rect 6804 80220 8204 80276
rect 8260 80220 9212 80276
rect 9268 80220 18844 80276
rect 18900 80220 19964 80276
rect 20020 80220 20030 80276
rect 7410 80108 7420 80164
rect 7476 80108 8092 80164
rect 8148 80108 9100 80164
rect 9156 80108 9660 80164
rect 9716 80108 9726 80164
rect 10546 80108 10556 80164
rect 10612 80108 11676 80164
rect 11732 80108 11742 80164
rect 12898 80108 12908 80164
rect 12964 80108 13468 80164
rect 13524 80108 13916 80164
rect 13972 80108 14812 80164
rect 14868 80108 14878 80164
rect 13998 79940 14008 79996
rect 14064 79940 14112 79996
rect 14168 79940 14216 79996
rect 14272 79940 14320 79996
rect 14376 79940 14424 79996
rect 14480 79940 14528 79996
rect 14584 79940 14632 79996
rect 14688 79940 14736 79996
rect 14792 79940 14840 79996
rect 14896 79940 14944 79996
rect 15000 79940 15048 79996
rect 15104 79940 15152 79996
rect 15208 79940 15218 79996
rect 33998 79940 34008 79996
rect 34064 79940 34112 79996
rect 34168 79940 34216 79996
rect 34272 79940 34320 79996
rect 34376 79940 34424 79996
rect 34480 79940 34528 79996
rect 34584 79940 34632 79996
rect 34688 79940 34736 79996
rect 34792 79940 34840 79996
rect 34896 79940 34944 79996
rect 35000 79940 35048 79996
rect 35104 79940 35152 79996
rect 35208 79940 35218 79996
rect 4722 79772 4732 79828
rect 4788 79772 5292 79828
rect 5348 79772 6748 79828
rect 6804 79772 6814 79828
rect 11890 79772 11900 79828
rect 11956 79772 15260 79828
rect 15316 79772 15596 79828
rect 15652 79772 15662 79828
rect 0 79604 800 79632
rect 0 79548 1708 79604
rect 1764 79548 1774 79604
rect 10994 79548 11004 79604
rect 11060 79548 14252 79604
rect 14308 79548 14318 79604
rect 0 79520 800 79548
rect 8754 79436 8764 79492
rect 8820 79436 10556 79492
rect 10612 79436 13804 79492
rect 13860 79436 13870 79492
rect 15138 79436 15148 79492
rect 15204 79436 16380 79492
rect 16436 79436 16446 79492
rect 5394 79324 5404 79380
rect 5460 79324 6076 79380
rect 6132 79324 6142 79380
rect 6514 79324 6524 79380
rect 6580 79324 7980 79380
rect 8036 79324 8046 79380
rect 10770 79212 10780 79268
rect 10836 79212 11228 79268
rect 11284 79212 11294 79268
rect 3998 79156 4008 79212
rect 4064 79156 4112 79212
rect 4168 79156 4216 79212
rect 4272 79156 4320 79212
rect 4376 79156 4424 79212
rect 4480 79156 4528 79212
rect 4584 79156 4632 79212
rect 4688 79156 4736 79212
rect 4792 79156 4840 79212
rect 4896 79156 4944 79212
rect 5000 79156 5048 79212
rect 5104 79156 5152 79212
rect 5208 79156 5218 79212
rect 23998 79156 24008 79212
rect 24064 79156 24112 79212
rect 24168 79156 24216 79212
rect 24272 79156 24320 79212
rect 24376 79156 24424 79212
rect 24480 79156 24528 79212
rect 24584 79156 24632 79212
rect 24688 79156 24736 79212
rect 24792 79156 24840 79212
rect 24896 79156 24944 79212
rect 25000 79156 25048 79212
rect 25104 79156 25152 79212
rect 25208 79156 25218 79212
rect 9650 79100 9660 79156
rect 9716 79100 10892 79156
rect 10948 79100 13356 79156
rect 13412 79100 13422 79156
rect 6290 78988 6300 79044
rect 6356 78988 6748 79044
rect 6804 78988 7532 79044
rect 7588 78988 7598 79044
rect 13682 78988 13692 79044
rect 13748 78988 15372 79044
rect 15428 78988 15438 79044
rect 7532 78932 7588 78988
rect 3378 78876 3388 78932
rect 3444 78876 4508 78932
rect 4564 78876 4574 78932
rect 5394 78876 5404 78932
rect 5460 78876 6244 78932
rect 7532 78876 9772 78932
rect 9828 78876 12012 78932
rect 12068 78876 12078 78932
rect 13234 78876 13244 78932
rect 13300 78876 13692 78932
rect 13748 78876 13758 78932
rect 4610 78764 4620 78820
rect 4676 78764 5852 78820
rect 5908 78764 5918 78820
rect 6188 78596 6244 78876
rect 8194 78764 8204 78820
rect 8260 78764 9884 78820
rect 9940 78764 9950 78820
rect 13906 78652 13916 78708
rect 13972 78652 15484 78708
rect 15540 78652 15550 78708
rect 20738 78652 20748 78708
rect 20804 78652 22988 78708
rect 23044 78652 23054 78708
rect 1698 78540 1708 78596
rect 1764 78540 1774 78596
rect 4162 78540 4172 78596
rect 4228 78540 5964 78596
rect 6020 78540 6030 78596
rect 6178 78540 6188 78596
rect 6244 78540 7084 78596
rect 7140 78540 7150 78596
rect 9986 78540 9996 78596
rect 10052 78540 11004 78596
rect 11060 78540 11452 78596
rect 11508 78540 11518 78596
rect 13570 78540 13580 78596
rect 13636 78540 15820 78596
rect 15876 78540 15886 78596
rect 0 78484 800 78512
rect 1708 78484 1764 78540
rect 0 78428 1764 78484
rect 20178 78428 20188 78484
rect 20244 78428 20972 78484
rect 21028 78428 21980 78484
rect 22036 78428 24332 78484
rect 24388 78428 25228 78484
rect 25284 78428 25294 78484
rect 0 78400 800 78428
rect 13998 78372 14008 78428
rect 14064 78372 14112 78428
rect 14168 78372 14216 78428
rect 14272 78372 14320 78428
rect 14376 78372 14424 78428
rect 14480 78372 14528 78428
rect 14584 78372 14632 78428
rect 14688 78372 14736 78428
rect 14792 78372 14840 78428
rect 14896 78372 14944 78428
rect 15000 78372 15048 78428
rect 15104 78372 15152 78428
rect 15208 78372 15218 78428
rect 33998 78372 34008 78428
rect 34064 78372 34112 78428
rect 34168 78372 34216 78428
rect 34272 78372 34320 78428
rect 34376 78372 34424 78428
rect 34480 78372 34528 78428
rect 34584 78372 34632 78428
rect 34688 78372 34736 78428
rect 34792 78372 34840 78428
rect 34896 78372 34944 78428
rect 35000 78372 35048 78428
rect 35104 78372 35152 78428
rect 35208 78372 35218 78428
rect 4498 78316 4508 78372
rect 4564 78316 5292 78372
rect 5348 78316 5358 78372
rect 4722 78204 4732 78260
rect 4788 78204 5292 78260
rect 5348 78204 5404 78260
rect 5460 78204 5470 78260
rect 12898 78204 12908 78260
rect 12964 78204 14700 78260
rect 14756 78204 14766 78260
rect 20290 78204 20300 78260
rect 20356 78204 22204 78260
rect 22260 78204 22270 78260
rect 23874 78204 23884 78260
rect 23940 78204 25340 78260
rect 25396 78204 25406 78260
rect 9202 78092 9212 78148
rect 9268 78092 9278 78148
rect 13570 78092 13580 78148
rect 13636 78092 13692 78148
rect 13748 78092 13758 78148
rect 9212 78036 9268 78092
rect 5842 77980 5852 78036
rect 5908 77980 7756 78036
rect 7812 77980 7822 78036
rect 8642 77980 8652 78036
rect 8708 77980 10108 78036
rect 10164 77980 10556 78036
rect 10612 77980 10622 78036
rect 15362 77980 15372 78036
rect 15428 77980 15484 78036
rect 15540 77980 15550 78036
rect 4834 77868 4844 77924
rect 4900 77868 5908 77924
rect 6066 77868 6076 77924
rect 6132 77868 6748 77924
rect 6804 77868 9660 77924
rect 9716 77868 9726 77924
rect 10658 77868 10668 77924
rect 10724 77868 11340 77924
rect 11396 77868 11406 77924
rect 12450 77868 12460 77924
rect 12516 77868 16380 77924
rect 16436 77868 16446 77924
rect 5852 77812 5908 77868
rect 3602 77756 3612 77812
rect 3668 77756 5628 77812
rect 5684 77756 5694 77812
rect 5852 77756 6132 77812
rect 6514 77756 6524 77812
rect 6580 77756 7308 77812
rect 7364 77756 7374 77812
rect 6076 77700 6132 77756
rect 6066 77644 6076 77700
rect 6132 77644 6142 77700
rect 8306 77644 8316 77700
rect 8372 77644 10108 77700
rect 10164 77644 10174 77700
rect 3998 77588 4008 77644
rect 4064 77588 4112 77644
rect 4168 77588 4216 77644
rect 4272 77588 4320 77644
rect 4376 77588 4424 77644
rect 4480 77588 4528 77644
rect 4584 77588 4632 77644
rect 4688 77588 4736 77644
rect 4792 77588 4840 77644
rect 4896 77588 4944 77644
rect 5000 77588 5048 77644
rect 5104 77588 5152 77644
rect 5208 77588 5218 77644
rect 23998 77588 24008 77644
rect 24064 77588 24112 77644
rect 24168 77588 24216 77644
rect 24272 77588 24320 77644
rect 24376 77588 24424 77644
rect 24480 77588 24528 77644
rect 24584 77588 24632 77644
rect 24688 77588 24736 77644
rect 24792 77588 24840 77644
rect 24896 77588 24944 77644
rect 25000 77588 25048 77644
rect 25104 77588 25152 77644
rect 25208 77588 25218 77644
rect 4274 77420 4284 77476
rect 4340 77420 5292 77476
rect 5348 77420 5358 77476
rect 0 77364 800 77392
rect 0 77308 1708 77364
rect 1764 77308 1774 77364
rect 5954 77308 5964 77364
rect 6020 77308 7420 77364
rect 7476 77308 8876 77364
rect 8932 77308 10052 77364
rect 13010 77308 13020 77364
rect 13076 77308 13804 77364
rect 13860 77308 14588 77364
rect 14644 77308 14654 77364
rect 24770 77308 24780 77364
rect 24836 77308 25676 77364
rect 25732 77308 25742 77364
rect 0 77280 800 77308
rect 9996 77252 10052 77308
rect 5058 77196 5068 77252
rect 5124 77196 6524 77252
rect 6580 77196 6860 77252
rect 6916 77196 6926 77252
rect 9996 77196 12572 77252
rect 12628 77196 12638 77252
rect 13346 77196 13356 77252
rect 13412 77196 13804 77252
rect 13860 77196 13870 77252
rect 14018 77196 14028 77252
rect 14084 77196 17276 77252
rect 17332 77196 17342 77252
rect 19954 77196 19964 77252
rect 20020 77196 21196 77252
rect 21252 77196 21868 77252
rect 21924 77196 21934 77252
rect 22306 77196 22316 77252
rect 22372 77196 24220 77252
rect 24276 77196 24286 77252
rect 6290 77084 6300 77140
rect 6356 77084 6636 77140
rect 6692 77084 6702 77140
rect 15362 77084 15372 77140
rect 15428 77084 16044 77140
rect 16100 77084 16110 77140
rect 11666 76972 11676 77028
rect 11732 76972 12012 77028
rect 12068 76972 12078 77028
rect 15138 76972 15148 77028
rect 15204 76972 15428 77028
rect 15372 76916 15428 76972
rect 15362 76860 15372 76916
rect 15428 76860 15438 76916
rect 16818 76860 16828 76916
rect 16884 76860 17388 76916
rect 17444 76860 20356 76916
rect 13998 76804 14008 76860
rect 14064 76804 14112 76860
rect 14168 76804 14216 76860
rect 14272 76804 14320 76860
rect 14376 76804 14424 76860
rect 14480 76804 14528 76860
rect 14584 76804 14632 76860
rect 14688 76804 14736 76860
rect 14792 76804 14840 76860
rect 14896 76804 14944 76860
rect 15000 76804 15048 76860
rect 15104 76804 15152 76860
rect 15208 76804 15218 76860
rect 15586 76748 15596 76804
rect 15652 76748 16380 76804
rect 16436 76748 17780 76804
rect 17724 76692 17780 76748
rect 20300 76692 20356 76860
rect 33998 76804 34008 76860
rect 34064 76804 34112 76860
rect 34168 76804 34216 76860
rect 34272 76804 34320 76860
rect 34376 76804 34424 76860
rect 34480 76804 34528 76860
rect 34584 76804 34632 76860
rect 34688 76804 34736 76860
rect 34792 76804 34840 76860
rect 34896 76804 34944 76860
rect 35000 76804 35048 76860
rect 35104 76804 35152 76860
rect 35208 76804 35218 76860
rect 3798 76636 3836 76692
rect 3892 76636 4732 76692
rect 4788 76636 4798 76692
rect 8530 76636 8540 76692
rect 8596 76636 9324 76692
rect 9380 76636 9772 76692
rect 9828 76636 12460 76692
rect 12516 76636 12526 76692
rect 14588 76636 15708 76692
rect 15764 76636 15774 76692
rect 17714 76636 17724 76692
rect 17780 76636 18732 76692
rect 18788 76636 18798 76692
rect 20290 76636 20300 76692
rect 20356 76636 21756 76692
rect 21812 76636 21822 76692
rect 14588 76580 14644 76636
rect 12002 76524 12012 76580
rect 12068 76524 14588 76580
rect 14644 76524 14654 76580
rect 15810 76524 15820 76580
rect 15876 76524 23436 76580
rect 23492 76524 23502 76580
rect 11106 76412 11116 76468
rect 11172 76412 13580 76468
rect 13636 76412 15372 76468
rect 15428 76412 16380 76468
rect 16436 76412 16446 76468
rect 18834 76412 18844 76468
rect 18900 76412 20188 76468
rect 20244 76412 20254 76468
rect 5730 76300 5740 76356
rect 5796 76300 6524 76356
rect 6580 76300 6748 76356
rect 6804 76300 6814 76356
rect 10658 76300 10668 76356
rect 10724 76300 12460 76356
rect 12516 76300 12526 76356
rect 16034 76300 16044 76356
rect 16100 76300 18284 76356
rect 18340 76300 18350 76356
rect 19282 76300 19292 76356
rect 19348 76300 20748 76356
rect 20804 76300 21308 76356
rect 21364 76300 21374 76356
rect 0 76244 800 76272
rect 0 76188 1708 76244
rect 1764 76188 1774 76244
rect 0 76160 800 76188
rect 3998 76020 4008 76076
rect 4064 76020 4112 76076
rect 4168 76020 4216 76076
rect 4272 76020 4320 76076
rect 4376 76020 4424 76076
rect 4480 76020 4528 76076
rect 4584 76020 4632 76076
rect 4688 76020 4736 76076
rect 4792 76020 4840 76076
rect 4896 76020 4944 76076
rect 5000 76020 5048 76076
rect 5104 76020 5152 76076
rect 5208 76020 5218 76076
rect 23998 76020 24008 76076
rect 24064 76020 24112 76076
rect 24168 76020 24216 76076
rect 24272 76020 24320 76076
rect 24376 76020 24424 76076
rect 24480 76020 24528 76076
rect 24584 76020 24632 76076
rect 24688 76020 24736 76076
rect 24792 76020 24840 76076
rect 24896 76020 24944 76076
rect 25000 76020 25048 76076
rect 25104 76020 25152 76076
rect 25208 76020 25218 76076
rect 4386 75740 4396 75796
rect 4452 75740 5852 75796
rect 5908 75740 5918 75796
rect 12338 75740 12348 75796
rect 12404 75740 12796 75796
rect 12852 75740 13356 75796
rect 13412 75740 14924 75796
rect 14980 75740 15764 75796
rect 15708 75684 15764 75740
rect 8866 75628 8876 75684
rect 8932 75628 10892 75684
rect 10948 75628 10958 75684
rect 15698 75628 15708 75684
rect 15764 75628 16156 75684
rect 16212 75628 16828 75684
rect 16884 75628 16894 75684
rect 13682 75516 13692 75572
rect 13748 75516 14476 75572
rect 14532 75516 14542 75572
rect 13794 75404 13804 75460
rect 13860 75404 14700 75460
rect 14756 75404 14766 75460
rect 19394 75404 19404 75460
rect 19460 75404 20524 75460
rect 20580 75404 20590 75460
rect 6066 75292 6076 75348
rect 6132 75292 6636 75348
rect 6692 75292 10780 75348
rect 10836 75292 10846 75348
rect 13998 75236 14008 75292
rect 14064 75236 14112 75292
rect 14168 75236 14216 75292
rect 14272 75236 14320 75292
rect 14376 75236 14424 75292
rect 14480 75236 14528 75292
rect 14584 75236 14632 75292
rect 14688 75236 14736 75292
rect 14792 75236 14840 75292
rect 14896 75236 14944 75292
rect 15000 75236 15048 75292
rect 15104 75236 15152 75292
rect 15208 75236 15218 75292
rect 33998 75236 34008 75292
rect 34064 75236 34112 75292
rect 34168 75236 34216 75292
rect 34272 75236 34320 75292
rect 34376 75236 34424 75292
rect 34480 75236 34528 75292
rect 34584 75236 34632 75292
rect 34688 75236 34736 75292
rect 34792 75236 34840 75292
rect 34896 75236 34944 75292
rect 35000 75236 35048 75292
rect 35104 75236 35152 75292
rect 35208 75236 35218 75292
rect 0 75124 800 75152
rect 0 75068 1708 75124
rect 1764 75068 1774 75124
rect 12674 75068 12684 75124
rect 12740 75068 13804 75124
rect 13860 75068 14252 75124
rect 14308 75068 14318 75124
rect 15362 75068 15372 75124
rect 15428 75068 15708 75124
rect 15764 75068 16492 75124
rect 16548 75068 16558 75124
rect 0 75040 800 75068
rect 15372 75012 15428 75068
rect 9986 74956 9996 75012
rect 10052 74956 10892 75012
rect 10948 74956 10958 75012
rect 13122 74956 13132 75012
rect 13188 74956 15428 75012
rect 7970 74844 7980 74900
rect 8036 74844 8652 74900
rect 8708 74844 8988 74900
rect 9044 74844 9054 74900
rect 12226 74844 12236 74900
rect 12292 74844 12572 74900
rect 12628 74844 12638 74900
rect 17938 74732 17948 74788
rect 18004 74732 18508 74788
rect 18564 74732 18574 74788
rect 6178 74620 6188 74676
rect 6244 74620 7420 74676
rect 7476 74620 7486 74676
rect 8082 74620 8092 74676
rect 8148 74620 8876 74676
rect 8932 74620 8942 74676
rect 3998 74452 4008 74508
rect 4064 74452 4112 74508
rect 4168 74452 4216 74508
rect 4272 74452 4320 74508
rect 4376 74452 4424 74508
rect 4480 74452 4528 74508
rect 4584 74452 4632 74508
rect 4688 74452 4736 74508
rect 4792 74452 4840 74508
rect 4896 74452 4944 74508
rect 5000 74452 5048 74508
rect 5104 74452 5152 74508
rect 5208 74452 5218 74508
rect 23998 74452 24008 74508
rect 24064 74452 24112 74508
rect 24168 74452 24216 74508
rect 24272 74452 24320 74508
rect 24376 74452 24424 74508
rect 24480 74452 24528 74508
rect 24584 74452 24632 74508
rect 24688 74452 24736 74508
rect 24792 74452 24840 74508
rect 24896 74452 24944 74508
rect 25000 74452 25048 74508
rect 25104 74452 25152 74508
rect 25208 74452 25218 74508
rect 4050 74284 4060 74340
rect 4116 74284 6636 74340
rect 6692 74284 6702 74340
rect 18386 74284 18396 74340
rect 18452 74284 19516 74340
rect 19572 74284 19582 74340
rect 1810 74172 1820 74228
rect 1876 74172 3164 74228
rect 3220 74172 5740 74228
rect 5796 74172 6972 74228
rect 7028 74172 7038 74228
rect 9426 74172 9436 74228
rect 9492 74172 11228 74228
rect 11284 74172 11294 74228
rect 3826 74060 3836 74116
rect 3892 74060 4060 74116
rect 4116 74060 4126 74116
rect 5964 74060 6188 74116
rect 6244 74060 6254 74116
rect 0 74004 800 74032
rect 0 73948 2156 74004
rect 2212 73948 2222 74004
rect 2482 73948 2492 74004
rect 2548 73948 3500 74004
rect 3556 73948 3566 74004
rect 4610 73948 4620 74004
rect 4676 73948 5292 74004
rect 5348 73948 5358 74004
rect 0 73920 800 73948
rect 5964 73892 6020 74060
rect 13570 73948 13580 74004
rect 13636 73948 17948 74004
rect 18004 73948 18014 74004
rect 4722 73836 4732 73892
rect 4788 73836 6020 73892
rect 11330 73836 11340 73892
rect 11396 73836 13692 73892
rect 13748 73836 13758 73892
rect 14354 73836 14364 73892
rect 14420 73836 15372 73892
rect 15428 73836 15438 73892
rect 13010 73724 13020 73780
rect 13076 73724 13580 73780
rect 13636 73724 13646 73780
rect 13998 73668 14008 73724
rect 14064 73668 14112 73724
rect 14168 73668 14216 73724
rect 14272 73668 14320 73724
rect 14376 73668 14424 73724
rect 14480 73668 14528 73724
rect 14584 73668 14632 73724
rect 14688 73668 14736 73724
rect 14792 73668 14840 73724
rect 14896 73668 14944 73724
rect 15000 73668 15048 73724
rect 15104 73668 15152 73724
rect 15208 73668 15218 73724
rect 33998 73668 34008 73724
rect 34064 73668 34112 73724
rect 34168 73668 34216 73724
rect 34272 73668 34320 73724
rect 34376 73668 34424 73724
rect 34480 73668 34528 73724
rect 34584 73668 34632 73724
rect 34688 73668 34736 73724
rect 34792 73668 34840 73724
rect 34896 73668 34944 73724
rect 35000 73668 35048 73724
rect 35104 73668 35152 73724
rect 35208 73668 35218 73724
rect 7858 73500 7868 73556
rect 7924 73500 9660 73556
rect 9716 73500 9726 73556
rect 13682 73500 13692 73556
rect 13748 73500 14364 73556
rect 14420 73500 15932 73556
rect 15988 73500 18284 73556
rect 18340 73500 18732 73556
rect 18788 73500 19404 73556
rect 19460 73500 21532 73556
rect 21588 73500 21598 73556
rect 20626 73388 20636 73444
rect 20692 73388 23884 73444
rect 23940 73388 23950 73444
rect 6066 73276 6076 73332
rect 6132 73276 7756 73332
rect 7812 73276 7822 73332
rect 10098 73276 10108 73332
rect 10164 73276 11004 73332
rect 11060 73276 11340 73332
rect 11396 73276 11406 73332
rect 21746 73276 21756 73332
rect 21812 73276 22876 73332
rect 22932 73276 22942 73332
rect 8530 73164 8540 73220
rect 8596 73164 9548 73220
rect 9604 73164 9884 73220
rect 9940 73164 10556 73220
rect 10612 73164 11676 73220
rect 11732 73164 11742 73220
rect 23426 73164 23436 73220
rect 23492 73164 24332 73220
rect 24388 73164 24398 73220
rect 0 72884 800 72912
rect 3998 72884 4008 72940
rect 4064 72884 4112 72940
rect 4168 72884 4216 72940
rect 4272 72884 4320 72940
rect 4376 72884 4424 72940
rect 4480 72884 4528 72940
rect 4584 72884 4632 72940
rect 4688 72884 4736 72940
rect 4792 72884 4840 72940
rect 4896 72884 4944 72940
rect 5000 72884 5048 72940
rect 5104 72884 5152 72940
rect 5208 72884 5218 72940
rect 23998 72884 24008 72940
rect 24064 72884 24112 72940
rect 24168 72884 24216 72940
rect 24272 72884 24320 72940
rect 24376 72884 24424 72940
rect 24480 72884 24528 72940
rect 24584 72884 24632 72940
rect 24688 72884 24736 72940
rect 24792 72884 24840 72940
rect 24896 72884 24944 72940
rect 25000 72884 25048 72940
rect 25104 72884 25152 72940
rect 25208 72884 25218 72940
rect 0 72828 1708 72884
rect 1764 72828 1774 72884
rect 0 72800 800 72828
rect 4946 72716 4956 72772
rect 5012 72716 6636 72772
rect 6692 72716 6702 72772
rect 3154 72492 3164 72548
rect 3220 72492 4172 72548
rect 4228 72492 5964 72548
rect 6020 72492 6030 72548
rect 6290 72492 6300 72548
rect 6356 72492 7868 72548
rect 7924 72492 9772 72548
rect 9828 72492 9838 72548
rect 4722 72380 4732 72436
rect 4788 72380 5292 72436
rect 5348 72380 6412 72436
rect 6468 72380 6478 72436
rect 8306 72380 8316 72436
rect 8372 72380 9884 72436
rect 9940 72380 9950 72436
rect 7634 72268 7644 72324
rect 7700 72268 8652 72324
rect 8708 72268 8718 72324
rect 23538 72268 23548 72324
rect 23604 72268 24332 72324
rect 24388 72268 24398 72324
rect 13998 72100 14008 72156
rect 14064 72100 14112 72156
rect 14168 72100 14216 72156
rect 14272 72100 14320 72156
rect 14376 72100 14424 72156
rect 14480 72100 14528 72156
rect 14584 72100 14632 72156
rect 14688 72100 14736 72156
rect 14792 72100 14840 72156
rect 14896 72100 14944 72156
rect 15000 72100 15048 72156
rect 15104 72100 15152 72156
rect 15208 72100 15218 72156
rect 33998 72100 34008 72156
rect 34064 72100 34112 72156
rect 34168 72100 34216 72156
rect 34272 72100 34320 72156
rect 34376 72100 34424 72156
rect 34480 72100 34528 72156
rect 34584 72100 34632 72156
rect 34688 72100 34736 72156
rect 34792 72100 34840 72156
rect 34896 72100 34944 72156
rect 35000 72100 35048 72156
rect 35104 72100 35152 72156
rect 35208 72100 35218 72156
rect 19842 71820 19852 71876
rect 19908 71820 22652 71876
rect 22708 71820 22718 71876
rect 0 71764 800 71792
rect 0 71708 1708 71764
rect 1764 71708 1774 71764
rect 0 71680 800 71708
rect 21186 71596 21196 71652
rect 21252 71596 23436 71652
rect 23492 71596 23502 71652
rect 34962 71484 34972 71540
rect 35028 71484 35308 71540
rect 35364 71484 35374 71540
rect 3998 71316 4008 71372
rect 4064 71316 4112 71372
rect 4168 71316 4216 71372
rect 4272 71316 4320 71372
rect 4376 71316 4424 71372
rect 4480 71316 4528 71372
rect 4584 71316 4632 71372
rect 4688 71316 4736 71372
rect 4792 71316 4840 71372
rect 4896 71316 4944 71372
rect 5000 71316 5048 71372
rect 5104 71316 5152 71372
rect 5208 71316 5218 71372
rect 23998 71316 24008 71372
rect 24064 71316 24112 71372
rect 24168 71316 24216 71372
rect 24272 71316 24320 71372
rect 24376 71316 24424 71372
rect 24480 71316 24528 71372
rect 24584 71316 24632 71372
rect 24688 71316 24736 71372
rect 24792 71316 24840 71372
rect 24896 71316 24944 71372
rect 25000 71316 25048 71372
rect 25104 71316 25152 71372
rect 25208 71316 25218 71372
rect 15250 71036 15260 71092
rect 15316 71036 15932 71092
rect 15988 71036 15998 71092
rect 13468 70924 13580 70980
rect 13636 70924 19292 70980
rect 19348 70924 21420 70980
rect 21476 70924 21486 70980
rect 24210 70924 24220 70980
rect 24276 70924 25116 70980
rect 25172 70924 27356 70980
rect 27412 70924 27422 70980
rect 30146 70924 30156 70980
rect 30212 70924 33068 70980
rect 33124 70924 33852 70980
rect 33908 70924 33918 70980
rect 1698 70700 1708 70756
rect 1764 70700 1774 70756
rect 6962 70700 6972 70756
rect 7028 70700 11116 70756
rect 11172 70700 11182 70756
rect 0 70644 800 70672
rect 1708 70644 1764 70700
rect 13468 70644 13524 70924
rect 15250 70812 15260 70868
rect 15316 70812 15428 70868
rect 0 70588 1764 70644
rect 13458 70588 13468 70644
rect 13524 70588 13534 70644
rect 0 70560 800 70588
rect 13998 70532 14008 70588
rect 14064 70532 14112 70588
rect 14168 70532 14216 70588
rect 14272 70532 14320 70588
rect 14376 70532 14424 70588
rect 14480 70532 14528 70588
rect 14584 70532 14632 70588
rect 14688 70532 14736 70588
rect 14792 70532 14840 70588
rect 14896 70532 14944 70588
rect 15000 70532 15048 70588
rect 15104 70532 15152 70588
rect 15208 70532 15218 70588
rect 15372 70420 15428 70812
rect 23538 70700 23548 70756
rect 23604 70700 23614 70756
rect 31826 70700 31836 70756
rect 31892 70700 35756 70756
rect 35812 70700 35822 70756
rect 23548 70532 23604 70700
rect 33998 70532 34008 70588
rect 34064 70532 34112 70588
rect 34168 70532 34216 70588
rect 34272 70532 34320 70588
rect 34376 70532 34424 70588
rect 34480 70532 34528 70588
rect 34584 70532 34632 70588
rect 34688 70532 34736 70588
rect 34792 70532 34840 70588
rect 34896 70532 34944 70588
rect 35000 70532 35048 70588
rect 35104 70532 35152 70588
rect 35208 70532 35218 70588
rect 22194 70476 22204 70532
rect 22260 70476 23604 70532
rect 23874 70476 23884 70532
rect 23940 70476 25676 70532
rect 25732 70476 25742 70532
rect 32386 70476 32396 70532
rect 32452 70476 33404 70532
rect 33460 70476 33470 70532
rect 35298 70476 35308 70532
rect 35364 70476 35644 70532
rect 35700 70476 35710 70532
rect 13570 70364 13580 70420
rect 13636 70364 15036 70420
rect 15092 70364 15428 70420
rect 23548 70420 23604 70476
rect 23548 70364 27020 70420
rect 27076 70364 27086 70420
rect 33170 70364 33180 70420
rect 33236 70364 33740 70420
rect 33796 70364 33806 70420
rect 34402 70364 34412 70420
rect 34468 70364 35308 70420
rect 35364 70364 35374 70420
rect 9650 70252 9660 70308
rect 9716 70252 10556 70308
rect 10612 70252 16044 70308
rect 16100 70252 16548 70308
rect 16492 70196 16548 70252
rect 32620 70252 33292 70308
rect 33348 70252 36652 70308
rect 36708 70252 36718 70308
rect 8418 70140 8428 70196
rect 8484 70140 9436 70196
rect 9492 70140 9502 70196
rect 16482 70140 16492 70196
rect 16548 70140 16558 70196
rect 16706 70140 16716 70196
rect 16772 70140 18508 70196
rect 18564 70140 18574 70196
rect 25554 70140 25564 70196
rect 25620 70140 26236 70196
rect 26292 70140 26302 70196
rect 27122 70140 27132 70196
rect 27188 70140 27916 70196
rect 27972 70140 28700 70196
rect 28756 70140 31836 70196
rect 31892 70140 31902 70196
rect 32620 70084 32676 70252
rect 36306 70140 36316 70196
rect 36372 70140 38108 70196
rect 38164 70140 38174 70196
rect 6178 70028 6188 70084
rect 6244 70028 7420 70084
rect 7476 70028 8988 70084
rect 9044 70028 9772 70084
rect 9828 70028 10332 70084
rect 10388 70028 10398 70084
rect 17826 70028 17836 70084
rect 17892 70028 19404 70084
rect 19460 70028 19470 70084
rect 23762 70028 23772 70084
rect 23828 70028 24668 70084
rect 24724 70028 25116 70084
rect 25172 70028 25182 70084
rect 26450 70028 26460 70084
rect 26516 70028 27580 70084
rect 27636 70028 27646 70084
rect 29810 70028 29820 70084
rect 29876 70028 32508 70084
rect 32564 70028 32676 70084
rect 35186 70028 35196 70084
rect 35252 70028 37772 70084
rect 37828 70028 37838 70084
rect 36082 69916 36092 69972
rect 36148 69916 37436 69972
rect 37492 69916 37884 69972
rect 37940 69916 37950 69972
rect 33394 69804 33404 69860
rect 33460 69804 34972 69860
rect 35028 69804 35532 69860
rect 35588 69804 35598 69860
rect 3998 69748 4008 69804
rect 4064 69748 4112 69804
rect 4168 69748 4216 69804
rect 4272 69748 4320 69804
rect 4376 69748 4424 69804
rect 4480 69748 4528 69804
rect 4584 69748 4632 69804
rect 4688 69748 4736 69804
rect 4792 69748 4840 69804
rect 4896 69748 4944 69804
rect 5000 69748 5048 69804
rect 5104 69748 5152 69804
rect 5208 69748 5218 69804
rect 23998 69748 24008 69804
rect 24064 69748 24112 69804
rect 24168 69748 24216 69804
rect 24272 69748 24320 69804
rect 24376 69748 24424 69804
rect 24480 69748 24528 69804
rect 24584 69748 24632 69804
rect 24688 69748 24736 69804
rect 24792 69748 24840 69804
rect 24896 69748 24944 69804
rect 25000 69748 25048 69804
rect 25104 69748 25152 69804
rect 25208 69748 25218 69804
rect 13682 69692 13692 69748
rect 13748 69692 13804 69748
rect 13860 69692 13870 69748
rect 12002 69580 12012 69636
rect 12068 69580 14252 69636
rect 14308 69580 14812 69636
rect 14868 69580 15708 69636
rect 15764 69580 15774 69636
rect 24546 69580 24556 69636
rect 24612 69580 25340 69636
rect 25396 69580 25406 69636
rect 33506 69580 33516 69636
rect 33572 69580 34636 69636
rect 34692 69580 34702 69636
rect 0 69524 800 69552
rect 0 69468 1708 69524
rect 1764 69468 1774 69524
rect 14914 69468 14924 69524
rect 14980 69468 15372 69524
rect 15428 69468 15438 69524
rect 15586 69468 15596 69524
rect 15652 69468 15764 69524
rect 16146 69468 16156 69524
rect 16212 69468 18956 69524
rect 19012 69468 19022 69524
rect 25890 69468 25900 69524
rect 25956 69468 29260 69524
rect 29316 69468 29326 69524
rect 0 69440 800 69468
rect 15708 69412 15764 69468
rect 15474 69356 15484 69412
rect 15540 69356 15550 69412
rect 15708 69356 16492 69412
rect 16548 69356 17388 69412
rect 17444 69356 17454 69412
rect 17938 69356 17948 69412
rect 18004 69356 18396 69412
rect 18452 69356 18462 69412
rect 11890 69244 11900 69300
rect 11956 69244 14028 69300
rect 14084 69244 14094 69300
rect 15484 69188 15540 69356
rect 17826 69244 17836 69300
rect 17892 69244 18508 69300
rect 18564 69244 18574 69300
rect 27010 69244 27020 69300
rect 27076 69244 27580 69300
rect 27636 69244 28364 69300
rect 28420 69244 29148 69300
rect 29204 69244 29214 69300
rect 35522 69244 35532 69300
rect 35588 69244 35756 69300
rect 35812 69244 35980 69300
rect 36036 69244 37548 69300
rect 37604 69244 37614 69300
rect 17836 69188 17892 69244
rect 10434 69132 10444 69188
rect 10500 69132 11228 69188
rect 11284 69132 12236 69188
rect 12292 69132 12302 69188
rect 12898 69132 12908 69188
rect 12964 69132 13580 69188
rect 13636 69132 13646 69188
rect 13906 69132 13916 69188
rect 13972 69132 15036 69188
rect 15092 69132 15820 69188
rect 15876 69132 17892 69188
rect 19366 69132 19404 69188
rect 19460 69132 19470 69188
rect 33852 69132 33964 69188
rect 34020 69132 34030 69188
rect 12236 69076 12292 69132
rect 12236 69020 13356 69076
rect 13412 69020 13422 69076
rect 16594 69020 16604 69076
rect 16660 69020 18732 69076
rect 18788 69020 18798 69076
rect 13998 68964 14008 69020
rect 14064 68964 14112 69020
rect 14168 68964 14216 69020
rect 14272 68964 14320 69020
rect 14376 68964 14424 69020
rect 14480 68964 14528 69020
rect 14584 68964 14632 69020
rect 14688 68964 14736 69020
rect 14792 68964 14840 69020
rect 14896 68964 14944 69020
rect 15000 68964 15048 69020
rect 15104 68964 15152 69020
rect 15208 68964 15218 69020
rect 15698 68908 15708 68964
rect 15764 68908 17724 68964
rect 17780 68908 17790 68964
rect 18162 68908 18172 68964
rect 18228 68908 25620 68964
rect 13542 68796 13580 68852
rect 13636 68796 13646 68852
rect 16034 68796 16044 68852
rect 16100 68796 17052 68852
rect 17108 68796 17118 68852
rect 19058 68796 19068 68852
rect 19124 68796 19740 68852
rect 19796 68796 19806 68852
rect 25564 68740 25620 68908
rect 33852 68852 33908 69132
rect 33998 68964 34008 69020
rect 34064 68964 34112 69020
rect 34168 68964 34216 69020
rect 34272 68964 34320 69020
rect 34376 68964 34424 69020
rect 34480 68964 34528 69020
rect 34584 68964 34632 69020
rect 34688 68964 34736 69020
rect 34792 68964 34840 69020
rect 34896 68964 34944 69020
rect 35000 68964 35048 69020
rect 35104 68964 35152 69020
rect 35208 68964 35218 69020
rect 27906 68796 27916 68852
rect 27972 68796 28812 68852
rect 28868 68796 28878 68852
rect 30594 68796 30604 68852
rect 30660 68796 34972 68852
rect 35028 68796 36204 68852
rect 36260 68796 36270 68852
rect 15250 68684 15260 68740
rect 15316 68684 15820 68740
rect 15876 68684 16492 68740
rect 16548 68684 16558 68740
rect 25554 68684 25564 68740
rect 25620 68684 25630 68740
rect 16258 68572 16268 68628
rect 16324 68572 16940 68628
rect 16996 68572 17500 68628
rect 17556 68572 17566 68628
rect 18162 68572 18172 68628
rect 18228 68572 19516 68628
rect 19572 68572 19582 68628
rect 24210 68572 24220 68628
rect 24276 68572 25676 68628
rect 25732 68572 25742 68628
rect 26674 68572 26684 68628
rect 26740 68572 29596 68628
rect 29652 68572 29662 68628
rect 10882 68460 10892 68516
rect 10948 68460 11900 68516
rect 11956 68460 11966 68516
rect 16706 68460 16716 68516
rect 16772 68460 17948 68516
rect 18004 68460 18014 68516
rect 24658 68460 24668 68516
rect 24724 68460 26348 68516
rect 26404 68460 26414 68516
rect 0 68404 800 68432
rect 0 68348 1708 68404
rect 1764 68348 1774 68404
rect 24434 68348 24444 68404
rect 24500 68348 26460 68404
rect 26516 68348 26526 68404
rect 29026 68348 29036 68404
rect 29092 68348 30156 68404
rect 30212 68348 30222 68404
rect 0 68320 800 68348
rect 3998 68180 4008 68236
rect 4064 68180 4112 68236
rect 4168 68180 4216 68236
rect 4272 68180 4320 68236
rect 4376 68180 4424 68236
rect 4480 68180 4528 68236
rect 4584 68180 4632 68236
rect 4688 68180 4736 68236
rect 4792 68180 4840 68236
rect 4896 68180 4944 68236
rect 5000 68180 5048 68236
rect 5104 68180 5152 68236
rect 5208 68180 5218 68236
rect 23998 68180 24008 68236
rect 24064 68180 24112 68236
rect 24168 68180 24216 68236
rect 24272 68180 24320 68236
rect 24376 68180 24424 68236
rect 24480 68180 24528 68236
rect 24584 68180 24632 68236
rect 24688 68180 24736 68236
rect 24792 68180 24840 68236
rect 24896 68180 24944 68236
rect 25000 68180 25048 68236
rect 25104 68180 25152 68236
rect 25208 68180 25218 68236
rect 19170 68124 19180 68180
rect 19236 68124 21420 68180
rect 21476 68124 21486 68180
rect 5842 68012 5852 68068
rect 5908 68012 6860 68068
rect 6916 68012 16268 68068
rect 16324 68012 16334 68068
rect 20738 68012 20748 68068
rect 20804 68012 24444 68068
rect 24500 68012 24510 68068
rect 3042 67788 3052 67844
rect 3108 67788 4172 67844
rect 4228 67788 4238 67844
rect 14466 67788 14476 67844
rect 14532 67788 15372 67844
rect 15428 67788 15438 67844
rect 26450 67788 26460 67844
rect 26516 67788 27804 67844
rect 27860 67788 27870 67844
rect 35858 67788 35868 67844
rect 35924 67788 37100 67844
rect 37156 67788 37166 67844
rect 13458 67676 13468 67732
rect 13524 67676 14028 67732
rect 14084 67676 14588 67732
rect 14644 67676 14654 67732
rect 15586 67676 15596 67732
rect 15652 67676 16492 67732
rect 16548 67676 16716 67732
rect 16772 67676 16782 67732
rect 29362 67676 29372 67732
rect 29428 67676 30716 67732
rect 30772 67676 30782 67732
rect 5282 67564 5292 67620
rect 5348 67564 5628 67620
rect 5684 67564 5694 67620
rect 6402 67564 6412 67620
rect 6468 67564 6972 67620
rect 7028 67564 7038 67620
rect 11218 67564 11228 67620
rect 11284 67564 12572 67620
rect 12628 67564 12638 67620
rect 13234 67564 13244 67620
rect 13300 67564 14252 67620
rect 14308 67564 14318 67620
rect 14802 67564 14812 67620
rect 14868 67564 16156 67620
rect 16212 67564 17388 67620
rect 17444 67564 17454 67620
rect 20066 67564 20076 67620
rect 20132 67564 21532 67620
rect 21588 67564 21598 67620
rect 32050 67564 32060 67620
rect 32116 67564 32956 67620
rect 33012 67564 33022 67620
rect 6066 67452 6076 67508
rect 6132 67452 7420 67508
rect 7476 67452 9884 67508
rect 9940 67452 9950 67508
rect 6486 67340 6524 67396
rect 6580 67340 6590 67396
rect 0 67284 800 67312
rect 13804 67284 13860 67564
rect 13998 67396 14008 67452
rect 14064 67396 14112 67452
rect 14168 67396 14216 67452
rect 14272 67396 14320 67452
rect 14376 67396 14424 67452
rect 14480 67396 14528 67452
rect 14584 67396 14632 67452
rect 14688 67396 14736 67452
rect 14792 67396 14840 67452
rect 14896 67396 14944 67452
rect 15000 67396 15048 67452
rect 15104 67396 15152 67452
rect 15208 67396 15218 67452
rect 33998 67396 34008 67452
rect 34064 67396 34112 67452
rect 34168 67396 34216 67452
rect 34272 67396 34320 67452
rect 34376 67396 34424 67452
rect 34480 67396 34528 67452
rect 34584 67396 34632 67452
rect 34688 67396 34736 67452
rect 34792 67396 34840 67452
rect 34896 67396 34944 67452
rect 35000 67396 35048 67452
rect 35104 67396 35152 67452
rect 35208 67396 35218 67452
rect 0 67228 1708 67284
rect 1764 67228 1774 67284
rect 4946 67228 4956 67284
rect 5012 67228 6580 67284
rect 9090 67228 9100 67284
rect 9156 67228 9660 67284
rect 9716 67228 11452 67284
rect 11508 67228 12236 67284
rect 12292 67228 13468 67284
rect 13524 67228 13534 67284
rect 13804 67228 14924 67284
rect 14980 67228 14990 67284
rect 20962 67228 20972 67284
rect 21028 67228 21038 67284
rect 25330 67228 25340 67284
rect 25396 67228 29036 67284
rect 29092 67228 29102 67284
rect 34514 67228 34524 67284
rect 34580 67228 35308 67284
rect 35364 67228 35374 67284
rect 0 67200 800 67228
rect 6524 67172 6580 67228
rect 20972 67172 21028 67228
rect 4498 67116 4508 67172
rect 4564 67116 5404 67172
rect 5460 67116 6300 67172
rect 6356 67116 6366 67172
rect 6514 67116 6524 67172
rect 6580 67116 6590 67172
rect 12562 67116 12572 67172
rect 12628 67116 13244 67172
rect 13300 67116 13916 67172
rect 13972 67116 13982 67172
rect 15922 67116 15932 67172
rect 15988 67116 17612 67172
rect 17668 67116 17678 67172
rect 19394 67116 19404 67172
rect 19460 67116 19470 67172
rect 20972 67116 21532 67172
rect 21588 67116 21598 67172
rect 31266 67116 31276 67172
rect 31332 67116 32172 67172
rect 32228 67116 33292 67172
rect 33348 67116 33358 67172
rect 19404 67060 19460 67116
rect 11666 67004 11676 67060
rect 11732 67004 13580 67060
rect 13636 67004 13646 67060
rect 16706 67004 16716 67060
rect 16772 67004 17164 67060
rect 17220 67004 17948 67060
rect 18004 67004 18014 67060
rect 19170 67004 19180 67060
rect 19236 67004 19460 67060
rect 3490 66892 3500 66948
rect 3556 66892 4732 66948
rect 4788 66892 5404 66948
rect 5460 66892 6860 66948
rect 6916 66892 8092 66948
rect 8148 66892 8158 66948
rect 15092 66892 18732 66948
rect 18788 66892 18798 66948
rect 15092 66836 15148 66892
rect 2258 66780 2268 66836
rect 2324 66780 3388 66836
rect 3444 66780 3454 66836
rect 7298 66780 7308 66836
rect 7364 66780 8764 66836
rect 8820 66780 10780 66836
rect 10836 66780 15148 66836
rect 17826 66780 17836 66836
rect 17892 66780 19180 66836
rect 19236 66780 19246 66836
rect 20972 66724 21028 67116
rect 23762 66892 23772 66948
rect 23828 66892 25228 66948
rect 25284 66892 25340 66948
rect 25396 66892 26236 66948
rect 26292 66892 26684 66948
rect 26740 66892 26750 66948
rect 31378 66892 31388 66948
rect 31444 66892 33180 66948
rect 33236 66892 33246 66948
rect 22530 66780 22540 66836
rect 22596 66780 24444 66836
rect 24500 66780 24510 66836
rect 31154 66780 31164 66836
rect 31220 66780 31612 66836
rect 31668 66780 32396 66836
rect 32452 66780 32462 66836
rect 6962 66668 6972 66724
rect 7028 66668 21028 66724
rect 3998 66612 4008 66668
rect 4064 66612 4112 66668
rect 4168 66612 4216 66668
rect 4272 66612 4320 66668
rect 4376 66612 4424 66668
rect 4480 66612 4528 66668
rect 4584 66612 4632 66668
rect 4688 66612 4736 66668
rect 4792 66612 4840 66668
rect 4896 66612 4944 66668
rect 5000 66612 5048 66668
rect 5104 66612 5152 66668
rect 5208 66612 5218 66668
rect 23998 66612 24008 66668
rect 24064 66612 24112 66668
rect 24168 66612 24216 66668
rect 24272 66612 24320 66668
rect 24376 66612 24424 66668
rect 24480 66612 24528 66668
rect 24584 66612 24632 66668
rect 24688 66612 24736 66668
rect 24792 66612 24840 66668
rect 24896 66612 24944 66668
rect 25000 66612 25048 66668
rect 25104 66612 25152 66668
rect 25208 66612 25218 66668
rect 7634 66556 7644 66612
rect 7700 66556 8428 66612
rect 8484 66556 8494 66612
rect 10994 66444 11004 66500
rect 11060 66444 13132 66500
rect 13188 66444 13198 66500
rect 18162 66444 18172 66500
rect 18228 66444 19292 66500
rect 19348 66444 19358 66500
rect 10210 66332 10220 66388
rect 10276 66332 11676 66388
rect 11732 66332 11742 66388
rect 35634 66332 35644 66388
rect 35700 66332 36988 66388
rect 37044 66332 37054 66388
rect 6402 66220 6412 66276
rect 6468 66220 6972 66276
rect 7028 66220 7038 66276
rect 8194 66220 8204 66276
rect 8260 66220 17164 66276
rect 17220 66220 18172 66276
rect 18228 66220 18732 66276
rect 18788 66220 19180 66276
rect 19236 66220 19246 66276
rect 20178 66220 20188 66276
rect 20244 66220 20636 66276
rect 20692 66220 25452 66276
rect 25508 66220 25518 66276
rect 29362 66220 29372 66276
rect 29428 66220 31836 66276
rect 31892 66220 31902 66276
rect 0 66164 800 66192
rect 0 66108 2156 66164
rect 2212 66108 2222 66164
rect 3602 66108 3612 66164
rect 3668 66108 4508 66164
rect 4564 66108 4574 66164
rect 9874 66108 9884 66164
rect 9940 66108 11228 66164
rect 11284 66108 11294 66164
rect 18498 66108 18508 66164
rect 18564 66108 19964 66164
rect 20020 66108 20748 66164
rect 20804 66108 20814 66164
rect 21298 66108 21308 66164
rect 21364 66108 22540 66164
rect 22596 66108 22606 66164
rect 28588 66108 31948 66164
rect 32004 66108 33740 66164
rect 33796 66108 36876 66164
rect 36932 66108 36942 66164
rect 0 66080 800 66108
rect 28588 66052 28644 66108
rect 4386 65996 4396 66052
rect 4452 65996 5740 66052
rect 5796 65996 6076 66052
rect 6132 65996 6142 66052
rect 17154 65996 17164 66052
rect 17220 65996 17612 66052
rect 17668 65996 19516 66052
rect 19572 65996 19582 66052
rect 23874 65996 23884 66052
rect 23940 65996 24556 66052
rect 24612 65996 28588 66052
rect 28644 65996 28654 66052
rect 31826 65996 31836 66052
rect 31892 65996 32732 66052
rect 32788 65996 32798 66052
rect 13998 65828 14008 65884
rect 14064 65828 14112 65884
rect 14168 65828 14216 65884
rect 14272 65828 14320 65884
rect 14376 65828 14424 65884
rect 14480 65828 14528 65884
rect 14584 65828 14632 65884
rect 14688 65828 14736 65884
rect 14792 65828 14840 65884
rect 14896 65828 14944 65884
rect 15000 65828 15048 65884
rect 15104 65828 15152 65884
rect 15208 65828 15218 65884
rect 33998 65828 34008 65884
rect 34064 65828 34112 65884
rect 34168 65828 34216 65884
rect 34272 65828 34320 65884
rect 34376 65828 34424 65884
rect 34480 65828 34528 65884
rect 34584 65828 34632 65884
rect 34688 65828 34736 65884
rect 34792 65828 34840 65884
rect 34896 65828 34944 65884
rect 35000 65828 35048 65884
rect 35104 65828 35152 65884
rect 35208 65828 35218 65884
rect 4722 65660 4732 65716
rect 4788 65660 6188 65716
rect 6244 65660 9996 65716
rect 10052 65660 10062 65716
rect 20402 65660 20412 65716
rect 20468 65660 21532 65716
rect 21588 65660 21598 65716
rect 28354 65660 28364 65716
rect 28420 65660 29372 65716
rect 29428 65660 29438 65716
rect 4050 65548 4060 65604
rect 4116 65548 5292 65604
rect 5348 65548 5358 65604
rect 17612 65548 20580 65604
rect 17612 65492 17668 65548
rect 20524 65492 20580 65548
rect 3332 65436 5628 65492
rect 5684 65436 6300 65492
rect 6356 65436 7196 65492
rect 7252 65436 8540 65492
rect 8596 65436 8606 65492
rect 9314 65436 9324 65492
rect 9380 65436 9996 65492
rect 10052 65436 10062 65492
rect 10210 65436 10220 65492
rect 10276 65436 10668 65492
rect 10724 65436 11116 65492
rect 11172 65436 17668 65492
rect 19170 65436 19180 65492
rect 19236 65436 20300 65492
rect 20356 65436 20366 65492
rect 20524 65436 21196 65492
rect 21252 65436 21262 65492
rect 26002 65436 26012 65492
rect 26068 65436 30828 65492
rect 30884 65436 30894 65492
rect 36306 65436 36316 65492
rect 36372 65436 37660 65492
rect 37716 65436 37726 65492
rect 1922 65212 1932 65268
rect 1988 65212 3276 65268
rect 3332 65212 3388 65436
rect 9324 65380 9380 65436
rect 7746 65324 7756 65380
rect 7812 65324 9380 65380
rect 13542 65324 13580 65380
rect 13636 65324 13646 65380
rect 14018 65324 14028 65380
rect 14084 65324 15820 65380
rect 15876 65324 15886 65380
rect 18946 65324 18956 65380
rect 19012 65324 19740 65380
rect 19796 65324 20076 65380
rect 20132 65324 20860 65380
rect 20916 65324 20926 65380
rect 24994 65324 25004 65380
rect 25060 65324 25340 65380
rect 25396 65324 25406 65380
rect 8978 65212 8988 65268
rect 9044 65212 12796 65268
rect 12852 65212 13916 65268
rect 13972 65212 17164 65268
rect 17220 65212 18172 65268
rect 18228 65212 18238 65268
rect 19058 65212 19068 65268
rect 19124 65212 19134 65268
rect 20290 65212 20300 65268
rect 20356 65212 21084 65268
rect 21140 65212 21150 65268
rect 19068 65156 19124 65212
rect 5730 65100 5740 65156
rect 5796 65100 13020 65156
rect 13076 65100 13086 65156
rect 13766 65100 13804 65156
rect 13860 65100 13870 65156
rect 14130 65100 14140 65156
rect 14196 65100 15484 65156
rect 15540 65100 15550 65156
rect 18050 65100 18060 65156
rect 18116 65100 19516 65156
rect 19572 65100 20524 65156
rect 20580 65100 20590 65156
rect 0 65044 800 65072
rect 3998 65044 4008 65100
rect 4064 65044 4112 65100
rect 4168 65044 4216 65100
rect 4272 65044 4320 65100
rect 4376 65044 4424 65100
rect 4480 65044 4528 65100
rect 4584 65044 4632 65100
rect 4688 65044 4736 65100
rect 4792 65044 4840 65100
rect 4896 65044 4944 65100
rect 5000 65044 5048 65100
rect 5104 65044 5152 65100
rect 5208 65044 5218 65100
rect 23998 65044 24008 65100
rect 24064 65044 24112 65100
rect 24168 65044 24216 65100
rect 24272 65044 24320 65100
rect 24376 65044 24424 65100
rect 24480 65044 24528 65100
rect 24584 65044 24632 65100
rect 24688 65044 24736 65100
rect 24792 65044 24840 65100
rect 24896 65044 24944 65100
rect 25000 65044 25048 65100
rect 25104 65044 25152 65100
rect 25208 65044 25218 65100
rect 0 64988 1708 65044
rect 1764 64988 1774 65044
rect 9202 64988 9212 65044
rect 9268 64988 10108 65044
rect 10164 64988 19964 65044
rect 20020 64988 20030 65044
rect 36082 64988 36092 65044
rect 36148 64988 37324 65044
rect 37380 64988 37390 65044
rect 0 64960 800 64988
rect 11330 64876 11340 64932
rect 11396 64876 11788 64932
rect 11844 64876 11854 64932
rect 12226 64876 12236 64932
rect 12292 64876 13244 64932
rect 13300 64876 13916 64932
rect 13972 64876 13982 64932
rect 14802 64876 14812 64932
rect 14868 64876 15428 64932
rect 16146 64876 16156 64932
rect 16212 64876 26796 64932
rect 26852 64876 26862 64932
rect 34626 64876 34636 64932
rect 34692 64876 35532 64932
rect 35588 64876 35598 64932
rect 35858 64876 35868 64932
rect 35924 64876 36988 64932
rect 37044 64876 37054 64932
rect 15372 64820 15428 64876
rect 10434 64764 10444 64820
rect 10500 64764 15148 64820
rect 15362 64764 15372 64820
rect 15428 64764 15438 64820
rect 15092 64708 15148 64764
rect 13122 64652 13132 64708
rect 13188 64652 14588 64708
rect 14644 64652 14654 64708
rect 15092 64652 17276 64708
rect 17332 64652 17342 64708
rect 18274 64652 18284 64708
rect 18340 64652 20188 64708
rect 20244 64652 20254 64708
rect 3154 64540 3164 64596
rect 3220 64540 3724 64596
rect 3780 64540 3790 64596
rect 13458 64540 13468 64596
rect 13524 64540 14700 64596
rect 14756 64540 15372 64596
rect 15428 64540 30268 64596
rect 30324 64540 30334 64596
rect 12002 64428 12012 64484
rect 12068 64428 12572 64484
rect 12628 64428 14476 64484
rect 14532 64428 15428 64484
rect 16706 64428 16716 64484
rect 16772 64428 18284 64484
rect 18340 64428 18350 64484
rect 18498 64428 18508 64484
rect 18564 64428 19180 64484
rect 19236 64428 19292 64484
rect 19348 64428 19358 64484
rect 8418 64316 8428 64372
rect 8484 64316 12236 64372
rect 12292 64316 12302 64372
rect 13998 64260 14008 64316
rect 14064 64260 14112 64316
rect 14168 64260 14216 64316
rect 14272 64260 14320 64316
rect 14376 64260 14424 64316
rect 14480 64260 14528 64316
rect 14584 64260 14632 64316
rect 14688 64260 14736 64316
rect 14792 64260 14840 64316
rect 14896 64260 14944 64316
rect 15000 64260 15048 64316
rect 15104 64260 15152 64316
rect 15208 64260 15218 64316
rect 15372 64260 15428 64428
rect 33998 64260 34008 64316
rect 34064 64260 34112 64316
rect 34168 64260 34216 64316
rect 34272 64260 34320 64316
rect 34376 64260 34424 64316
rect 34480 64260 34528 64316
rect 34584 64260 34632 64316
rect 34688 64260 34736 64316
rect 34792 64260 34840 64316
rect 34896 64260 34944 64316
rect 35000 64260 35048 64316
rect 35104 64260 35152 64316
rect 35208 64260 35218 64316
rect 15362 64204 15372 64260
rect 15428 64204 15438 64260
rect 5282 64092 5292 64148
rect 5348 64092 6188 64148
rect 6244 64092 6254 64148
rect 8530 64092 8540 64148
rect 8596 64092 8988 64148
rect 9044 64092 9054 64148
rect 13682 64092 13692 64148
rect 13748 64092 14700 64148
rect 14756 64092 14766 64148
rect 15250 64092 15260 64148
rect 15316 64092 15372 64148
rect 15428 64092 15438 64148
rect 4834 63980 4844 64036
rect 4900 63980 5404 64036
rect 5460 63980 5852 64036
rect 5908 63980 5918 64036
rect 12908 63980 16156 64036
rect 16212 63980 16222 64036
rect 19926 63980 19964 64036
rect 20020 63980 20030 64036
rect 0 63924 800 63952
rect 12908 63924 12964 63980
rect 0 63868 1708 63924
rect 1764 63868 1774 63924
rect 5394 63868 5404 63924
rect 5460 63868 12964 63924
rect 13122 63868 13132 63924
rect 13188 63868 13916 63924
rect 13972 63868 15596 63924
rect 15652 63868 15662 63924
rect 17602 63868 17612 63924
rect 17668 63868 18284 63924
rect 18340 63868 18956 63924
rect 19012 63868 20412 63924
rect 20468 63868 20478 63924
rect 27010 63868 27020 63924
rect 27076 63868 28812 63924
rect 28868 63868 29260 63924
rect 29316 63868 29326 63924
rect 34850 63868 34860 63924
rect 34916 63868 37324 63924
rect 37380 63868 37390 63924
rect 0 63840 800 63868
rect 5618 63756 5628 63812
rect 5684 63756 5694 63812
rect 8306 63756 8316 63812
rect 8372 63756 10444 63812
rect 10500 63756 10510 63812
rect 3998 63476 4008 63532
rect 4064 63476 4112 63532
rect 4168 63476 4216 63532
rect 4272 63476 4320 63532
rect 4376 63476 4424 63532
rect 4480 63476 4528 63532
rect 4584 63476 4632 63532
rect 4688 63476 4736 63532
rect 4792 63476 4840 63532
rect 4896 63476 4944 63532
rect 5000 63476 5048 63532
rect 5104 63476 5152 63532
rect 5208 63476 5218 63532
rect 5628 63364 5684 63756
rect 12908 63700 12964 63868
rect 13794 63756 13804 63812
rect 13860 63756 14924 63812
rect 14980 63756 14990 63812
rect 29922 63756 29932 63812
rect 29988 63756 31836 63812
rect 31892 63756 31902 63812
rect 12908 63644 13692 63700
rect 13748 63644 13804 63700
rect 13860 63644 13870 63700
rect 14242 63644 14252 63700
rect 14308 63644 15820 63700
rect 15876 63644 15886 63700
rect 13682 63532 13692 63588
rect 13748 63532 13804 63588
rect 13860 63532 13870 63588
rect 23998 63476 24008 63532
rect 24064 63476 24112 63532
rect 24168 63476 24216 63532
rect 24272 63476 24320 63532
rect 24376 63476 24424 63532
rect 24480 63476 24528 63532
rect 24584 63476 24632 63532
rect 24688 63476 24736 63532
rect 24792 63476 24840 63532
rect 24896 63476 24944 63532
rect 25000 63476 25048 63532
rect 25104 63476 25152 63532
rect 25208 63476 25218 63532
rect 13570 63420 13580 63476
rect 13636 63420 13646 63476
rect 13580 63364 13636 63420
rect 2370 63308 2380 63364
rect 2436 63308 3836 63364
rect 3892 63308 3902 63364
rect 4722 63308 4732 63364
rect 4788 63308 5684 63364
rect 7522 63308 7532 63364
rect 7588 63308 9212 63364
rect 9268 63308 9278 63364
rect 10434 63308 10444 63364
rect 10500 63308 11004 63364
rect 11060 63308 11070 63364
rect 13580 63308 13692 63364
rect 13748 63308 15148 63364
rect 15092 63252 15148 63308
rect 4162 63196 4172 63252
rect 4228 63196 5404 63252
rect 5460 63196 5470 63252
rect 6850 63196 6860 63252
rect 6916 63196 8764 63252
rect 8820 63196 8830 63252
rect 10098 63196 10108 63252
rect 10164 63196 13580 63252
rect 13636 63196 13646 63252
rect 15092 63196 17276 63252
rect 17332 63196 17342 63252
rect 24770 63196 24780 63252
rect 24836 63196 25676 63252
rect 25732 63196 25742 63252
rect 33842 63196 33852 63252
rect 33908 63196 34748 63252
rect 34804 63196 34814 63252
rect 13580 63140 13636 63196
rect 4946 63084 4956 63140
rect 5012 63084 6188 63140
rect 6244 63084 9548 63140
rect 9604 63084 9884 63140
rect 9940 63084 9950 63140
rect 13580 63084 23436 63140
rect 23492 63084 23502 63140
rect 23762 63084 23772 63140
rect 23828 63084 24892 63140
rect 24948 63084 24958 63140
rect 30482 63084 30492 63140
rect 30548 63084 31052 63140
rect 31108 63084 31118 63140
rect 3490 62972 3500 63028
rect 3556 62972 4732 63028
rect 4788 62972 4798 63028
rect 12450 62972 12460 63028
rect 12516 62972 13580 63028
rect 13636 62972 14476 63028
rect 14532 62972 14542 63028
rect 15250 62972 15260 63028
rect 15316 62972 15484 63028
rect 15540 62972 15550 63028
rect 16370 62972 16380 63028
rect 16436 62972 16828 63028
rect 16884 62972 16894 63028
rect 19394 62972 19404 63028
rect 19460 62972 20636 63028
rect 20692 62972 20702 63028
rect 24098 62972 24108 63028
rect 24164 62972 24668 63028
rect 24724 62972 25340 63028
rect 25396 62972 26572 63028
rect 26628 62972 27132 63028
rect 27188 62972 27198 63028
rect 35074 62972 35084 63028
rect 35140 62972 35868 63028
rect 35924 62972 35934 63028
rect 1698 62860 1708 62916
rect 1764 62860 1774 62916
rect 10882 62860 10892 62916
rect 10948 62860 12348 62916
rect 12404 62860 14028 62916
rect 14084 62860 16604 62916
rect 16660 62860 16670 62916
rect 19954 62860 19964 62916
rect 20020 62860 20076 62916
rect 20132 62860 20142 62916
rect 25218 62860 25228 62916
rect 25284 62860 26796 62916
rect 26852 62860 26862 62916
rect 31042 62860 31052 62916
rect 31108 62860 31500 62916
rect 31556 62860 35532 62916
rect 35588 62860 35598 62916
rect 35746 62860 35756 62916
rect 35812 62860 37548 62916
rect 37604 62860 37614 62916
rect 0 62804 800 62832
rect 1708 62804 1764 62860
rect 0 62748 1764 62804
rect 20290 62748 20300 62804
rect 20356 62748 20748 62804
rect 20804 62748 28588 62804
rect 28644 62748 30716 62804
rect 30772 62748 31276 62804
rect 31332 62748 31342 62804
rect 0 62720 800 62748
rect 13998 62692 14008 62748
rect 14064 62692 14112 62748
rect 14168 62692 14216 62748
rect 14272 62692 14320 62748
rect 14376 62692 14424 62748
rect 14480 62692 14528 62748
rect 14584 62692 14632 62748
rect 14688 62692 14736 62748
rect 14792 62692 14840 62748
rect 14896 62692 14944 62748
rect 15000 62692 15048 62748
rect 15104 62692 15152 62748
rect 15208 62692 15218 62748
rect 33998 62692 34008 62748
rect 34064 62692 34112 62748
rect 34168 62692 34216 62748
rect 34272 62692 34320 62748
rect 34376 62692 34424 62748
rect 34480 62692 34528 62748
rect 34584 62692 34632 62748
rect 34688 62692 34736 62748
rect 34792 62692 34840 62748
rect 34896 62692 34944 62748
rect 35000 62692 35048 62748
rect 35104 62692 35152 62748
rect 35208 62692 35218 62748
rect 13766 62636 13804 62692
rect 13860 62636 13870 62692
rect 17154 62636 17164 62692
rect 17220 62636 18172 62692
rect 18228 62636 19628 62692
rect 19684 62636 19852 62692
rect 19908 62636 19918 62692
rect 12898 62524 12908 62580
rect 12964 62524 14364 62580
rect 14420 62524 15932 62580
rect 15988 62524 15998 62580
rect 19366 62524 19404 62580
rect 19460 62524 19470 62580
rect 24098 62524 24108 62580
rect 24164 62524 25732 62580
rect 25676 62468 25732 62524
rect 26852 62524 28252 62580
rect 28308 62524 29596 62580
rect 29652 62524 29662 62580
rect 33618 62524 33628 62580
rect 33684 62524 36764 62580
rect 36820 62524 36830 62580
rect 26852 62468 26908 62524
rect 4834 62412 4844 62468
rect 4900 62412 5516 62468
rect 5572 62412 5582 62468
rect 7074 62412 7084 62468
rect 7140 62412 8876 62468
rect 8932 62412 8942 62468
rect 12786 62412 12796 62468
rect 12852 62412 13356 62468
rect 13412 62412 13580 62468
rect 13636 62412 14588 62468
rect 14644 62412 14654 62468
rect 14924 62412 15708 62468
rect 15764 62412 16380 62468
rect 16436 62412 16446 62468
rect 19058 62412 19068 62468
rect 19124 62412 19292 62468
rect 19348 62412 20300 62468
rect 20356 62412 20366 62468
rect 20514 62412 20524 62468
rect 20580 62412 22316 62468
rect 22372 62412 24668 62468
rect 24724 62412 24734 62468
rect 25666 62412 25676 62468
rect 25732 62412 26908 62468
rect 33842 62412 33852 62468
rect 33908 62412 34412 62468
rect 34468 62412 34478 62468
rect 5516 62356 5572 62412
rect 14924 62356 14980 62412
rect 4386 62300 4396 62356
rect 4452 62300 5292 62356
rect 5348 62300 5358 62356
rect 5516 62300 7420 62356
rect 7476 62300 7486 62356
rect 9762 62300 9772 62356
rect 9828 62300 10892 62356
rect 10948 62300 10958 62356
rect 13234 62300 13244 62356
rect 13300 62300 14924 62356
rect 14980 62300 14990 62356
rect 15362 62300 15372 62356
rect 15428 62300 16044 62356
rect 16100 62300 17052 62356
rect 17108 62300 17118 62356
rect 19506 62300 19516 62356
rect 19572 62300 20188 62356
rect 20244 62300 20254 62356
rect 25330 62300 25340 62356
rect 25396 62300 29148 62356
rect 29204 62300 30044 62356
rect 30100 62300 33404 62356
rect 33460 62300 33740 62356
rect 33796 62300 33806 62356
rect 4834 62188 4844 62244
rect 4900 62188 7196 62244
rect 7252 62188 7262 62244
rect 8306 62188 8316 62244
rect 8372 62188 9996 62244
rect 10052 62188 10062 62244
rect 13906 62188 13916 62244
rect 13972 62188 14588 62244
rect 14644 62188 14654 62244
rect 15026 62188 15036 62244
rect 15092 62188 16940 62244
rect 16996 62188 17006 62244
rect 26012 62188 28812 62244
rect 28868 62188 30492 62244
rect 30548 62188 30558 62244
rect 26012 62132 26068 62188
rect 4946 62076 4956 62132
rect 5012 62076 5292 62132
rect 5348 62076 5358 62132
rect 10210 62076 10220 62132
rect 10276 62076 12796 62132
rect 12852 62076 12862 62132
rect 13570 62076 13580 62132
rect 13636 62076 16828 62132
rect 16884 62076 16894 62132
rect 26002 62076 26012 62132
rect 26068 62076 26078 62132
rect 36754 62076 36764 62132
rect 36820 62076 37772 62132
rect 37828 62076 37838 62132
rect 14578 61964 14588 62020
rect 14644 61964 15372 62020
rect 15428 61964 15438 62020
rect 3998 61908 4008 61964
rect 4064 61908 4112 61964
rect 4168 61908 4216 61964
rect 4272 61908 4320 61964
rect 4376 61908 4424 61964
rect 4480 61908 4528 61964
rect 4584 61908 4632 61964
rect 4688 61908 4736 61964
rect 4792 61908 4840 61964
rect 4896 61908 4944 61964
rect 5000 61908 5048 61964
rect 5104 61908 5152 61964
rect 5208 61908 5218 61964
rect 23998 61908 24008 61964
rect 24064 61908 24112 61964
rect 24168 61908 24216 61964
rect 24272 61908 24320 61964
rect 24376 61908 24424 61964
rect 24480 61908 24528 61964
rect 24584 61908 24632 61964
rect 24688 61908 24736 61964
rect 24792 61908 24840 61964
rect 24896 61908 24944 61964
rect 25000 61908 25048 61964
rect 25104 61908 25152 61964
rect 25208 61908 25218 61964
rect 11218 61852 11228 61908
rect 11284 61852 12124 61908
rect 12180 61852 12190 61908
rect 13122 61852 13132 61908
rect 13188 61852 15596 61908
rect 15652 61852 15662 61908
rect 25778 61852 25788 61908
rect 25844 61852 26124 61908
rect 26180 61852 26190 61908
rect 7420 61740 24220 61796
rect 24276 61740 25228 61796
rect 25284 61740 25294 61796
rect 0 61684 800 61712
rect 7420 61684 7476 61740
rect 0 61628 1708 61684
rect 1764 61628 1774 61684
rect 5954 61628 5964 61684
rect 6020 61628 7476 61684
rect 13766 61628 13804 61684
rect 13860 61628 13870 61684
rect 14914 61628 14924 61684
rect 14980 61628 15484 61684
rect 15540 61628 15550 61684
rect 16930 61628 16940 61684
rect 16996 61628 17724 61684
rect 17780 61628 17790 61684
rect 0 61600 800 61628
rect 4050 61516 4060 61572
rect 4116 61516 5628 61572
rect 5684 61516 5694 61572
rect 10322 61516 10332 61572
rect 10388 61516 11004 61572
rect 11060 61516 19292 61572
rect 19348 61516 19358 61572
rect 36194 61516 36204 61572
rect 36260 61516 37324 61572
rect 37380 61516 37390 61572
rect 3826 61404 3836 61460
rect 3892 61404 4620 61460
rect 4676 61404 5292 61460
rect 5348 61404 13972 61460
rect 24546 61404 24556 61460
rect 24612 61404 25340 61460
rect 25396 61404 25788 61460
rect 25844 61404 26908 61460
rect 26964 61404 26974 61460
rect 28466 61404 28476 61460
rect 28532 61404 30604 61460
rect 30660 61404 30670 61460
rect 13916 61348 13972 61404
rect 2258 61292 2268 61348
rect 2324 61292 3724 61348
rect 3780 61292 3790 61348
rect 4722 61292 4732 61348
rect 4788 61292 5404 61348
rect 5460 61292 5740 61348
rect 5796 61292 8316 61348
rect 8372 61292 8382 61348
rect 9874 61292 9884 61348
rect 9940 61292 10780 61348
rect 10836 61292 11116 61348
rect 11172 61292 12348 61348
rect 12404 61292 12414 61348
rect 13654 61292 13692 61348
rect 13748 61292 13758 61348
rect 13916 61292 21420 61348
rect 21476 61292 21980 61348
rect 22036 61292 22046 61348
rect 28578 61292 28588 61348
rect 28644 61292 29596 61348
rect 29652 61292 29662 61348
rect 32498 61292 32508 61348
rect 32564 61292 33628 61348
rect 33684 61292 33852 61348
rect 33908 61292 34412 61348
rect 34468 61292 34478 61348
rect 6626 61180 6636 61236
rect 6692 61180 7084 61236
rect 7140 61180 7150 61236
rect 10994 61180 11004 61236
rect 11060 61180 11340 61236
rect 11396 61180 11406 61236
rect 13998 61124 14008 61180
rect 14064 61124 14112 61180
rect 14168 61124 14216 61180
rect 14272 61124 14320 61180
rect 14376 61124 14424 61180
rect 14480 61124 14528 61180
rect 14584 61124 14632 61180
rect 14688 61124 14736 61180
rect 14792 61124 14840 61180
rect 14896 61124 14944 61180
rect 15000 61124 15048 61180
rect 15104 61124 15152 61180
rect 15208 61124 15218 61180
rect 33998 61124 34008 61180
rect 34064 61124 34112 61180
rect 34168 61124 34216 61180
rect 34272 61124 34320 61180
rect 34376 61124 34424 61180
rect 34480 61124 34528 61180
rect 34584 61124 34632 61180
rect 34688 61124 34736 61180
rect 34792 61124 34840 61180
rect 34896 61124 34944 61180
rect 35000 61124 35048 61180
rect 35104 61124 35152 61180
rect 35208 61124 35218 61180
rect 30146 61068 30156 61124
rect 30212 61068 30828 61124
rect 30884 61068 30894 61124
rect 15922 60956 15932 61012
rect 15988 60956 16268 61012
rect 16324 60956 16334 61012
rect 26674 60956 26684 61012
rect 26740 60956 26908 61012
rect 28578 60956 28588 61012
rect 28644 60956 29932 61012
rect 29988 60956 33180 61012
rect 33236 60956 33246 61012
rect 5842 60844 5852 60900
rect 5908 60844 7532 60900
rect 7588 60844 7598 60900
rect 26852 60788 26908 60956
rect 30594 60844 30604 60900
rect 30660 60844 31724 60900
rect 31780 60844 33068 60900
rect 33124 60844 33134 60900
rect 7410 60732 7420 60788
rect 7476 60732 8540 60788
rect 8596 60732 16492 60788
rect 16548 60732 16558 60788
rect 26852 60732 27020 60788
rect 27076 60732 27086 60788
rect 31490 60732 31500 60788
rect 31556 60732 33292 60788
rect 33348 60732 33358 60788
rect 8194 60620 8204 60676
rect 8260 60620 8988 60676
rect 9044 60620 9054 60676
rect 10098 60620 10108 60676
rect 10164 60620 12684 60676
rect 12740 60620 12750 60676
rect 25330 60620 25340 60676
rect 25396 60620 26012 60676
rect 26068 60620 26078 60676
rect 31042 60620 31052 60676
rect 31108 60620 32060 60676
rect 32116 60620 33404 60676
rect 33460 60620 33740 60676
rect 33796 60620 33806 60676
rect 0 60564 800 60592
rect 0 60508 1708 60564
rect 1764 60508 1774 60564
rect 9090 60508 9100 60564
rect 9156 60508 13580 60564
rect 13636 60508 13646 60564
rect 16146 60508 16156 60564
rect 16212 60508 16604 60564
rect 16660 60508 16670 60564
rect 29586 60508 29596 60564
rect 29652 60508 33180 60564
rect 33236 60508 33246 60564
rect 0 60480 800 60508
rect 28690 60396 28700 60452
rect 28756 60396 29372 60452
rect 29428 60396 30268 60452
rect 30324 60396 30334 60452
rect 3998 60340 4008 60396
rect 4064 60340 4112 60396
rect 4168 60340 4216 60396
rect 4272 60340 4320 60396
rect 4376 60340 4424 60396
rect 4480 60340 4528 60396
rect 4584 60340 4632 60396
rect 4688 60340 4736 60396
rect 4792 60340 4840 60396
rect 4896 60340 4944 60396
rect 5000 60340 5048 60396
rect 5104 60340 5152 60396
rect 5208 60340 5218 60396
rect 23998 60340 24008 60396
rect 24064 60340 24112 60396
rect 24168 60340 24216 60396
rect 24272 60340 24320 60396
rect 24376 60340 24424 60396
rect 24480 60340 24528 60396
rect 24584 60340 24632 60396
rect 24688 60340 24736 60396
rect 24792 60340 24840 60396
rect 24896 60340 24944 60396
rect 25000 60340 25048 60396
rect 25104 60340 25152 60396
rect 25208 60340 25218 60396
rect 32386 60172 32396 60228
rect 32452 60172 33964 60228
rect 34020 60172 34030 60228
rect 36194 60172 36204 60228
rect 36260 60172 37548 60228
rect 37604 60172 38332 60228
rect 38388 60172 38398 60228
rect 5730 60060 5740 60116
rect 5796 60060 6636 60116
rect 6692 60060 9660 60116
rect 9716 60060 11676 60116
rect 11732 60060 11742 60116
rect 15092 60060 20524 60116
rect 20580 60060 20590 60116
rect 30034 60060 30044 60116
rect 30100 60060 32284 60116
rect 32340 60060 32350 60116
rect 15092 60004 15148 60060
rect 7074 59948 7084 60004
rect 7140 59948 15148 60004
rect 30930 59948 30940 60004
rect 30996 59948 31724 60004
rect 31780 59948 31790 60004
rect 36418 59948 36428 60004
rect 36484 59948 37324 60004
rect 37380 59948 37390 60004
rect 30034 59836 30044 59892
rect 30100 59836 30716 59892
rect 30772 59836 31668 59892
rect 31612 59780 31668 59836
rect 6178 59724 6188 59780
rect 6244 59724 6524 59780
rect 6580 59724 6590 59780
rect 23426 59724 23436 59780
rect 23492 59724 23772 59780
rect 23828 59724 26684 59780
rect 26740 59724 26750 59780
rect 28354 59724 28364 59780
rect 28420 59724 31052 59780
rect 31108 59724 31118 59780
rect 31602 59724 31612 59780
rect 31668 59724 31678 59780
rect 33170 59724 33180 59780
rect 33236 59724 34300 59780
rect 34356 59724 34366 59780
rect 13998 59556 14008 59612
rect 14064 59556 14112 59612
rect 14168 59556 14216 59612
rect 14272 59556 14320 59612
rect 14376 59556 14424 59612
rect 14480 59556 14528 59612
rect 14584 59556 14632 59612
rect 14688 59556 14736 59612
rect 14792 59556 14840 59612
rect 14896 59556 14944 59612
rect 15000 59556 15048 59612
rect 15104 59556 15152 59612
rect 15208 59556 15218 59612
rect 33998 59556 34008 59612
rect 34064 59556 34112 59612
rect 34168 59556 34216 59612
rect 34272 59556 34320 59612
rect 34376 59556 34424 59612
rect 34480 59556 34528 59612
rect 34584 59556 34632 59612
rect 34688 59556 34736 59612
rect 34792 59556 34840 59612
rect 34896 59556 34944 59612
rect 35000 59556 35048 59612
rect 35104 59556 35152 59612
rect 35208 59556 35218 59612
rect 19030 59500 19068 59556
rect 19124 59500 19740 59556
rect 19796 59500 20188 59556
rect 20244 59500 20254 59556
rect 0 59444 800 59472
rect 0 59388 1708 59444
rect 1764 59388 1774 59444
rect 13570 59388 13580 59444
rect 13636 59388 13916 59444
rect 13972 59388 13982 59444
rect 14914 59388 14924 59444
rect 14980 59388 15372 59444
rect 15428 59388 15438 59444
rect 17266 59388 17276 59444
rect 17332 59388 18396 59444
rect 18452 59388 18462 59444
rect 19842 59388 19852 59444
rect 19908 59388 22092 59444
rect 22148 59388 22158 59444
rect 23874 59388 23884 59444
rect 23940 59388 25340 59444
rect 25396 59388 28812 59444
rect 28868 59388 29932 59444
rect 29988 59388 30492 59444
rect 30548 59388 32508 59444
rect 32564 59388 33180 59444
rect 33236 59388 33246 59444
rect 0 59360 800 59388
rect 9314 59276 9324 59332
rect 9380 59276 13020 59332
rect 13076 59276 13086 59332
rect 30146 59276 30156 59332
rect 30212 59276 31276 59332
rect 31332 59276 33068 59332
rect 33124 59276 33134 59332
rect 12562 59164 12572 59220
rect 12628 59164 15372 59220
rect 15428 59164 15438 59220
rect 18722 59164 18732 59220
rect 18788 59164 20524 59220
rect 20580 59164 20590 59220
rect 21522 59164 21532 59220
rect 21588 59164 21598 59220
rect 19506 59052 19516 59108
rect 19572 59052 20636 59108
rect 20692 59052 20702 59108
rect 21532 58996 21588 59164
rect 21746 59052 21756 59108
rect 21812 59052 22204 59108
rect 22260 59052 27244 59108
rect 27300 59052 27310 59108
rect 13794 58940 13804 58996
rect 13860 58940 14700 58996
rect 14756 58940 14766 58996
rect 20178 58940 20188 58996
rect 20244 58940 20748 58996
rect 20804 58940 21588 58996
rect 14018 58828 14028 58884
rect 14084 58828 18956 58884
rect 19012 58828 19022 58884
rect 19254 58828 19292 58884
rect 19348 58828 20860 58884
rect 20916 58828 20926 58884
rect 27794 58828 27804 58884
rect 27860 58828 29708 58884
rect 29764 58828 30380 58884
rect 30436 58828 31052 58884
rect 31108 58828 33292 58884
rect 33348 58828 33358 58884
rect 3998 58772 4008 58828
rect 4064 58772 4112 58828
rect 4168 58772 4216 58828
rect 4272 58772 4320 58828
rect 4376 58772 4424 58828
rect 4480 58772 4528 58828
rect 4584 58772 4632 58828
rect 4688 58772 4736 58828
rect 4792 58772 4840 58828
rect 4896 58772 4944 58828
rect 5000 58772 5048 58828
rect 5104 58772 5152 58828
rect 5208 58772 5218 58828
rect 23998 58772 24008 58828
rect 24064 58772 24112 58828
rect 24168 58772 24216 58828
rect 24272 58772 24320 58828
rect 24376 58772 24424 58828
rect 24480 58772 24528 58828
rect 24584 58772 24632 58828
rect 24688 58772 24736 58828
rect 24792 58772 24840 58828
rect 24896 58772 24944 58828
rect 25000 58772 25048 58828
rect 25104 58772 25152 58828
rect 25208 58772 25218 58828
rect 6514 58716 6524 58772
rect 6580 58716 13468 58772
rect 13524 58716 13534 58772
rect 19058 58716 19068 58772
rect 19124 58716 19460 58772
rect 19702 58716 19740 58772
rect 19796 58716 19806 58772
rect 7382 58604 7420 58660
rect 7476 58604 7486 58660
rect 18498 58604 18508 58660
rect 18564 58604 18844 58660
rect 18900 58604 18910 58660
rect 19404 58548 19460 58716
rect 19590 58604 19628 58660
rect 19684 58604 19694 58660
rect 3714 58492 3724 58548
rect 3780 58492 3948 58548
rect 4004 58492 10220 58548
rect 10276 58492 10286 58548
rect 12450 58492 12460 58548
rect 12516 58492 13580 58548
rect 13636 58492 13646 58548
rect 19394 58492 19404 58548
rect 19460 58492 19470 58548
rect 31602 58492 31612 58548
rect 31668 58492 32284 58548
rect 32340 58492 32350 58548
rect 13906 58380 13916 58436
rect 13972 58380 14812 58436
rect 14868 58380 17164 58436
rect 17220 58380 17230 58436
rect 18498 58380 18508 58436
rect 18564 58380 19852 58436
rect 19908 58380 19918 58436
rect 20290 58380 20300 58436
rect 20356 58380 21644 58436
rect 21700 58380 21710 58436
rect 26002 58380 26012 58436
rect 26068 58380 26572 58436
rect 26628 58380 27356 58436
rect 27412 58380 28140 58436
rect 28196 58380 28206 58436
rect 28466 58380 28476 58436
rect 28532 58380 29932 58436
rect 29988 58380 29998 58436
rect 33394 58380 33404 58436
rect 33460 58380 35196 58436
rect 35252 58380 35262 58436
rect 0 58324 800 58352
rect 0 58268 2492 58324
rect 2548 58268 2940 58324
rect 2996 58268 3006 58324
rect 13692 58268 15036 58324
rect 15092 58268 15708 58324
rect 15764 58268 15774 58324
rect 16146 58268 16156 58324
rect 16212 58268 16380 58324
rect 16436 58268 16604 58324
rect 16660 58268 18172 58324
rect 18228 58268 18396 58324
rect 18452 58268 18462 58324
rect 25666 58268 25676 58324
rect 25732 58268 26684 58324
rect 26740 58268 26750 58324
rect 34402 58268 34412 58324
rect 34468 58268 35084 58324
rect 35140 58268 35150 58324
rect 35522 58268 35532 58324
rect 35588 58268 36876 58324
rect 36932 58268 36942 58324
rect 0 58240 800 58268
rect 7522 58156 7532 58212
rect 7588 58156 8204 58212
rect 8260 58156 8270 58212
rect 8754 58156 8764 58212
rect 8820 58156 9436 58212
rect 9492 58156 9502 58212
rect 13692 57988 13748 58268
rect 17724 58212 17780 58268
rect 14914 58156 14924 58212
rect 14980 58156 15372 58212
rect 15428 58156 15438 58212
rect 17714 58156 17724 58212
rect 17780 58156 17790 58212
rect 18834 58156 18844 58212
rect 18900 58156 23660 58212
rect 23716 58156 23726 58212
rect 30370 58156 30380 58212
rect 30436 58156 30940 58212
rect 30996 58156 31388 58212
rect 31444 58156 32732 58212
rect 32788 58156 32798 58212
rect 33852 58156 34972 58212
rect 35028 58156 35038 58212
rect 36418 58156 36428 58212
rect 36484 58156 37100 58212
rect 37156 58156 37166 58212
rect 18386 58044 18396 58100
rect 18452 58044 19068 58100
rect 19124 58044 19134 58100
rect 13998 57988 14008 58044
rect 14064 57988 14112 58044
rect 14168 57988 14216 58044
rect 14272 57988 14320 58044
rect 14376 57988 14424 58044
rect 14480 57988 14528 58044
rect 14584 57988 14632 58044
rect 14688 57988 14736 58044
rect 14792 57988 14840 58044
rect 14896 57988 14944 58044
rect 15000 57988 15048 58044
rect 15104 57988 15152 58044
rect 15208 57988 15218 58044
rect 13682 57932 13692 57988
rect 13748 57932 13758 57988
rect 16604 57932 25452 57988
rect 25508 57932 26236 57988
rect 26292 57932 26302 57988
rect 15026 57820 15036 57876
rect 15092 57820 16044 57876
rect 16100 57820 16110 57876
rect 16604 57764 16660 57932
rect 33852 57876 33908 58156
rect 33998 57988 34008 58044
rect 34064 57988 34112 58044
rect 34168 57988 34216 58044
rect 34272 57988 34320 58044
rect 34376 57988 34424 58044
rect 34480 57988 34528 58044
rect 34584 57988 34632 58044
rect 34688 57988 34736 58044
rect 34792 57988 34840 58044
rect 34896 57988 34944 58044
rect 35000 57988 35048 58044
rect 35104 57988 35152 58044
rect 35208 57988 35218 58044
rect 26786 57820 26796 57876
rect 26852 57820 28140 57876
rect 28196 57820 28206 57876
rect 28578 57820 28588 57876
rect 28644 57820 30828 57876
rect 30884 57820 30894 57876
rect 33852 57820 34300 57876
rect 34356 57820 34366 57876
rect 9426 57708 9436 57764
rect 9492 57708 10556 57764
rect 10612 57708 16660 57764
rect 19954 57708 19964 57764
rect 20020 57708 24780 57764
rect 24836 57708 24846 57764
rect 11330 57596 11340 57652
rect 11396 57596 11788 57652
rect 11844 57596 12348 57652
rect 12404 57596 12414 57652
rect 12786 57596 12796 57652
rect 12852 57596 14364 57652
rect 14420 57596 14430 57652
rect 17602 57596 17612 57652
rect 17668 57596 18620 57652
rect 18676 57596 18686 57652
rect 19394 57596 19404 57652
rect 19460 57596 20748 57652
rect 20804 57596 21532 57652
rect 21588 57596 21598 57652
rect 23650 57596 23660 57652
rect 23716 57596 25676 57652
rect 25732 57596 25742 57652
rect 33394 57596 33404 57652
rect 33460 57596 34076 57652
rect 34132 57596 34142 57652
rect 6066 57484 6076 57540
rect 6132 57484 6972 57540
rect 7028 57484 7038 57540
rect 9090 57484 9100 57540
rect 9156 57484 10780 57540
rect 10836 57484 10846 57540
rect 13804 57428 13860 57596
rect 16818 57484 16828 57540
rect 16884 57484 18172 57540
rect 18228 57484 19180 57540
rect 19236 57484 20524 57540
rect 20580 57484 20590 57540
rect 11732 57372 12460 57428
rect 12516 57372 12796 57428
rect 12852 57372 12862 57428
rect 13794 57372 13804 57428
rect 13860 57372 13870 57428
rect 14242 57372 14252 57428
rect 14308 57372 18620 57428
rect 18676 57372 19292 57428
rect 19348 57372 19358 57428
rect 19702 57372 19740 57428
rect 19796 57372 19806 57428
rect 6850 57260 6860 57316
rect 6916 57260 6926 57316
rect 0 57204 800 57232
rect 3998 57204 4008 57260
rect 4064 57204 4112 57260
rect 4168 57204 4216 57260
rect 4272 57204 4320 57260
rect 4376 57204 4424 57260
rect 4480 57204 4528 57260
rect 4584 57204 4632 57260
rect 4688 57204 4736 57260
rect 4792 57204 4840 57260
rect 4896 57204 4944 57260
rect 5000 57204 5048 57260
rect 5104 57204 5152 57260
rect 5208 57204 5218 57260
rect 0 57148 2604 57204
rect 2660 57148 2670 57204
rect 0 57120 800 57148
rect 6860 57092 6916 57260
rect 11732 57204 11788 57372
rect 25330 57260 25340 57316
rect 25396 57260 25900 57316
rect 25956 57260 25966 57316
rect 34850 57260 34860 57316
rect 34916 57260 35532 57316
rect 35588 57260 35598 57316
rect 23998 57204 24008 57260
rect 24064 57204 24112 57260
rect 24168 57204 24216 57260
rect 24272 57204 24320 57260
rect 24376 57204 24424 57260
rect 24480 57204 24528 57260
rect 24584 57204 24632 57260
rect 24688 57204 24736 57260
rect 24792 57204 24840 57260
rect 24896 57204 24944 57260
rect 25000 57204 25048 57260
rect 25104 57204 25152 57260
rect 25208 57204 25218 57260
rect 7074 57148 7084 57204
rect 7140 57148 7868 57204
rect 7924 57148 7934 57204
rect 8194 57148 8204 57204
rect 8260 57148 9660 57204
rect 9716 57148 9726 57204
rect 10770 57148 10780 57204
rect 10836 57148 11116 57204
rect 11172 57148 11564 57204
rect 11620 57148 11788 57204
rect 17714 57148 17724 57204
rect 17780 57148 20300 57204
rect 20356 57148 20366 57204
rect 6860 57036 7980 57092
rect 8036 57036 8046 57092
rect 11890 57036 11900 57092
rect 11956 57036 13580 57092
rect 13636 57036 15372 57092
rect 15428 57036 15820 57092
rect 15876 57036 15886 57092
rect 36194 57036 36204 57092
rect 36260 57036 36988 57092
rect 37044 57036 37054 57092
rect 9650 56924 9660 56980
rect 9716 56924 11676 56980
rect 11732 56924 11742 56980
rect 12114 56924 12124 56980
rect 12180 56924 12460 56980
rect 12516 56924 12526 56980
rect 34738 56924 34748 56980
rect 34804 56924 36764 56980
rect 36820 56924 36830 56980
rect 9986 56812 9996 56868
rect 10052 56812 11340 56868
rect 11396 56812 13132 56868
rect 13188 56812 13198 56868
rect 13794 56812 13804 56868
rect 13860 56812 14252 56868
rect 14308 56812 16828 56868
rect 16884 56812 16894 56868
rect 21522 56812 21532 56868
rect 21588 56812 25116 56868
rect 25172 56812 25182 56868
rect 4386 56700 4396 56756
rect 4452 56700 5292 56756
rect 5348 56700 6636 56756
rect 6692 56700 6702 56756
rect 13458 56700 13468 56756
rect 13524 56700 14364 56756
rect 14420 56700 14430 56756
rect 18050 56700 18060 56756
rect 18116 56700 19740 56756
rect 19796 56700 19806 56756
rect 23090 56700 23100 56756
rect 23156 56700 23548 56756
rect 36978 56700 36988 56756
rect 37044 56700 37436 56756
rect 37492 56700 37502 56756
rect 23492 56644 23548 56700
rect 2258 56588 2268 56644
rect 2324 56588 3276 56644
rect 3332 56588 3342 56644
rect 4274 56588 4284 56644
rect 4340 56588 4956 56644
rect 5012 56588 5292 56644
rect 5348 56588 5358 56644
rect 6514 56588 6524 56644
rect 6580 56588 7532 56644
rect 7588 56588 7598 56644
rect 10434 56588 10444 56644
rect 10500 56588 11340 56644
rect 11396 56588 11406 56644
rect 12572 56588 16828 56644
rect 16884 56588 17388 56644
rect 17444 56588 17454 56644
rect 23492 56588 23996 56644
rect 24052 56588 26124 56644
rect 26180 56588 26190 56644
rect 31154 56588 31164 56644
rect 31220 56588 33852 56644
rect 33908 56588 34300 56644
rect 34356 56588 35084 56644
rect 35140 56588 35980 56644
rect 36036 56588 36428 56644
rect 36484 56588 36494 56644
rect 9650 56476 9660 56532
rect 9716 56476 10556 56532
rect 10612 56476 12236 56532
rect 12292 56476 12302 56532
rect 12572 56420 12628 56588
rect 13998 56420 14008 56476
rect 14064 56420 14112 56476
rect 14168 56420 14216 56476
rect 14272 56420 14320 56476
rect 14376 56420 14424 56476
rect 14480 56420 14528 56476
rect 14584 56420 14632 56476
rect 14688 56420 14736 56476
rect 14792 56420 14840 56476
rect 14896 56420 14944 56476
rect 15000 56420 15048 56476
rect 15104 56420 15152 56476
rect 15208 56420 15218 56476
rect 33998 56420 34008 56476
rect 34064 56420 34112 56476
rect 34168 56420 34216 56476
rect 34272 56420 34320 56476
rect 34376 56420 34424 56476
rect 34480 56420 34528 56476
rect 34584 56420 34632 56476
rect 34688 56420 34736 56476
rect 34792 56420 34840 56476
rect 34896 56420 34944 56476
rect 35000 56420 35048 56476
rect 35104 56420 35152 56476
rect 35208 56420 35218 56476
rect 12562 56364 12572 56420
rect 12628 56364 12638 56420
rect 16370 56364 16380 56420
rect 16436 56364 19852 56420
rect 19908 56364 19918 56420
rect 4162 56252 4172 56308
rect 4228 56252 5740 56308
rect 5796 56252 5806 56308
rect 10098 56252 10108 56308
rect 10164 56252 12460 56308
rect 12516 56252 12526 56308
rect 12674 56252 12684 56308
rect 12740 56252 14028 56308
rect 14084 56252 14094 56308
rect 18470 56252 18508 56308
rect 18564 56252 18574 56308
rect 18946 56252 18956 56308
rect 19012 56252 20076 56308
rect 20132 56252 20142 56308
rect 22754 56252 22764 56308
rect 22820 56252 26348 56308
rect 26404 56252 26414 56308
rect 11778 56140 11788 56196
rect 11844 56140 13580 56196
rect 13636 56140 13916 56196
rect 13972 56140 13982 56196
rect 15026 56140 15036 56196
rect 15092 56140 20748 56196
rect 20804 56140 22204 56196
rect 22260 56140 22270 56196
rect 22418 56140 22428 56196
rect 22484 56140 22988 56196
rect 23044 56140 24668 56196
rect 24724 56140 24734 56196
rect 26450 56140 26460 56196
rect 26516 56140 27692 56196
rect 27748 56140 28140 56196
rect 28196 56140 30268 56196
rect 30324 56140 32060 56196
rect 32116 56140 33684 56196
rect 0 56084 800 56112
rect 33628 56084 33684 56140
rect 35252 56084 35308 56308
rect 35364 56252 36204 56308
rect 36260 56252 37660 56308
rect 37716 56252 37726 56308
rect 0 56028 2380 56084
rect 2436 56028 2828 56084
rect 2884 56028 2894 56084
rect 7746 56028 7756 56084
rect 7812 56028 8428 56084
rect 8484 56028 8764 56084
rect 8820 56028 8830 56084
rect 11666 56028 11676 56084
rect 11732 56028 12908 56084
rect 12964 56028 13468 56084
rect 13524 56028 13534 56084
rect 17042 56028 17052 56084
rect 17108 56028 17388 56084
rect 17444 56028 17454 56084
rect 20290 56028 20300 56084
rect 20356 56028 21420 56084
rect 21476 56028 22316 56084
rect 22372 56028 22382 56084
rect 31154 56028 31164 56084
rect 31220 56028 32508 56084
rect 32564 56028 33292 56084
rect 33348 56028 33358 56084
rect 33618 56028 33628 56084
rect 33684 56028 35308 56084
rect 0 56000 800 56028
rect 33292 55972 33348 56028
rect 3266 55916 3276 55972
rect 3332 55916 10444 55972
rect 10500 55916 10510 55972
rect 10658 55916 10668 55972
rect 10724 55916 14252 55972
rect 14308 55916 14588 55972
rect 14644 55916 14654 55972
rect 15092 55916 20860 55972
rect 20916 55916 21644 55972
rect 21700 55916 22092 55972
rect 22148 55916 22158 55972
rect 33292 55916 33852 55972
rect 33908 55916 33918 55972
rect 35746 55916 35756 55972
rect 35812 55916 37100 55972
rect 37156 55916 37166 55972
rect 15092 55860 15148 55916
rect 12450 55804 12460 55860
rect 12516 55804 15148 55860
rect 16818 55804 16828 55860
rect 16884 55804 18060 55860
rect 18116 55804 18126 55860
rect 13010 55692 13020 55748
rect 13076 55692 13692 55748
rect 13748 55692 13804 55748
rect 13860 55692 14588 55748
rect 14644 55692 14654 55748
rect 15474 55692 15484 55748
rect 15540 55692 17836 55748
rect 17892 55692 17902 55748
rect 3998 55636 4008 55692
rect 4064 55636 4112 55692
rect 4168 55636 4216 55692
rect 4272 55636 4320 55692
rect 4376 55636 4424 55692
rect 4480 55636 4528 55692
rect 4584 55636 4632 55692
rect 4688 55636 4736 55692
rect 4792 55636 4840 55692
rect 4896 55636 4944 55692
rect 5000 55636 5048 55692
rect 5104 55636 5152 55692
rect 5208 55636 5218 55692
rect 23998 55636 24008 55692
rect 24064 55636 24112 55692
rect 24168 55636 24216 55692
rect 24272 55636 24320 55692
rect 24376 55636 24424 55692
rect 24480 55636 24528 55692
rect 24584 55636 24632 55692
rect 24688 55636 24736 55692
rect 24792 55636 24840 55692
rect 24896 55636 24944 55692
rect 25000 55636 25048 55692
rect 25104 55636 25152 55692
rect 25208 55636 25218 55692
rect 7186 55468 7196 55524
rect 7252 55468 7868 55524
rect 7924 55468 7934 55524
rect 8754 55468 8764 55524
rect 8820 55468 8830 55524
rect 10070 55468 10108 55524
rect 10164 55468 10174 55524
rect 11666 55468 11676 55524
rect 11732 55468 12572 55524
rect 12628 55468 12638 55524
rect 8764 55412 8820 55468
rect 1810 55356 1820 55412
rect 1876 55356 3724 55412
rect 3780 55356 3790 55412
rect 8194 55356 8204 55412
rect 8260 55356 12348 55412
rect 12404 55356 12414 55412
rect 13458 55356 13468 55412
rect 13524 55356 14252 55412
rect 14308 55356 14318 55412
rect 15092 55356 19068 55412
rect 19124 55356 19134 55412
rect 15092 55300 15148 55356
rect 3266 55244 3276 55300
rect 0 54964 800 54992
rect 3332 54964 3388 55300
rect 3602 55244 3612 55300
rect 3668 55244 4844 55300
rect 4900 55244 6188 55300
rect 6244 55244 15148 55300
rect 16370 55244 16380 55300
rect 16436 55244 18844 55300
rect 18900 55244 19516 55300
rect 19572 55244 21756 55300
rect 21812 55244 21822 55300
rect 36418 55244 36428 55300
rect 36484 55244 37100 55300
rect 37156 55244 37166 55300
rect 4946 55132 4956 55188
rect 5012 55132 7084 55188
rect 7140 55132 7150 55188
rect 10210 55132 10220 55188
rect 10276 55132 10668 55188
rect 10724 55132 10734 55188
rect 12450 55132 12460 55188
rect 12516 55132 13804 55188
rect 13860 55132 14028 55188
rect 14084 55132 14094 55188
rect 15092 55132 15932 55188
rect 15988 55132 15998 55188
rect 18386 55132 18396 55188
rect 18452 55132 18732 55188
rect 18788 55132 19628 55188
rect 19684 55132 20300 55188
rect 20356 55132 20366 55188
rect 21074 55132 21084 55188
rect 21140 55132 22540 55188
rect 22596 55132 22606 55188
rect 5730 55020 5740 55076
rect 5796 55020 6636 55076
rect 6692 55020 6860 55076
rect 6916 55020 6926 55076
rect 10108 55020 11004 55076
rect 11060 55020 11070 55076
rect 11442 55020 11452 55076
rect 11508 55020 12012 55076
rect 12068 55020 15036 55076
rect 15092 55020 15148 55132
rect 15474 55020 15484 55076
rect 15540 55020 16044 55076
rect 16100 55020 16110 55076
rect 10108 54964 10164 55020
rect 0 54908 2604 54964
rect 2660 54908 2670 54964
rect 3332 54908 10108 54964
rect 10164 54908 10174 54964
rect 0 54880 800 54908
rect 13998 54852 14008 54908
rect 14064 54852 14112 54908
rect 14168 54852 14216 54908
rect 14272 54852 14320 54908
rect 14376 54852 14424 54908
rect 14480 54852 14528 54908
rect 14584 54852 14632 54908
rect 14688 54852 14736 54908
rect 14792 54852 14840 54908
rect 14896 54852 14944 54908
rect 15000 54852 15048 54908
rect 15104 54852 15152 54908
rect 15208 54852 15218 54908
rect 33998 54852 34008 54908
rect 34064 54852 34112 54908
rect 34168 54852 34216 54908
rect 34272 54852 34320 54908
rect 34376 54852 34424 54908
rect 34480 54852 34528 54908
rect 34584 54852 34632 54908
rect 34688 54852 34736 54908
rect 34792 54852 34840 54908
rect 34896 54852 34944 54908
rect 35000 54852 35048 54908
rect 35104 54852 35152 54908
rect 35208 54852 35218 54908
rect 3714 54684 3724 54740
rect 3780 54684 5628 54740
rect 5684 54684 6748 54740
rect 6804 54684 7868 54740
rect 7924 54684 7934 54740
rect 9986 54684 9996 54740
rect 10052 54684 11564 54740
rect 11620 54684 13692 54740
rect 13748 54684 14364 54740
rect 14420 54684 14430 54740
rect 21186 54684 21196 54740
rect 21252 54684 22092 54740
rect 22148 54684 22876 54740
rect 22932 54684 22942 54740
rect 6262 54572 6300 54628
rect 6356 54572 6366 54628
rect 7186 54572 7196 54628
rect 7252 54572 8092 54628
rect 8148 54572 8158 54628
rect 8978 54572 8988 54628
rect 9044 54572 9212 54628
rect 9268 54572 10780 54628
rect 10836 54572 10846 54628
rect 11330 54572 11340 54628
rect 11396 54572 23548 54628
rect 23604 54572 23614 54628
rect 6178 54460 6188 54516
rect 6244 54460 7644 54516
rect 7700 54460 8876 54516
rect 8932 54460 8942 54516
rect 9436 54460 15036 54516
rect 15092 54460 15102 54516
rect 27346 54460 27356 54516
rect 27412 54460 30380 54516
rect 30436 54460 30446 54516
rect 9436 54404 9492 54460
rect 6514 54348 6524 54404
rect 6580 54348 7196 54404
rect 7252 54348 7262 54404
rect 7410 54348 7420 54404
rect 7476 54348 9492 54404
rect 10210 54348 10220 54404
rect 10276 54348 11452 54404
rect 11508 54348 11518 54404
rect 13916 54348 15372 54404
rect 15428 54348 15438 54404
rect 4722 54236 4732 54292
rect 4788 54236 5740 54292
rect 5796 54236 6300 54292
rect 6356 54236 6366 54292
rect 13468 54236 13692 54292
rect 13748 54236 13758 54292
rect 13468 54180 13524 54236
rect 13458 54124 13468 54180
rect 13524 54124 13534 54180
rect 3998 54068 4008 54124
rect 4064 54068 4112 54124
rect 4168 54068 4216 54124
rect 4272 54068 4320 54124
rect 4376 54068 4424 54124
rect 4480 54068 4528 54124
rect 4584 54068 4632 54124
rect 4688 54068 4736 54124
rect 4792 54068 4840 54124
rect 4896 54068 4944 54124
rect 5000 54068 5048 54124
rect 5104 54068 5152 54124
rect 5208 54068 5218 54124
rect 13916 54068 13972 54348
rect 15026 54124 15036 54180
rect 15092 54124 18172 54180
rect 18228 54124 18238 54180
rect 23998 54068 24008 54124
rect 24064 54068 24112 54124
rect 24168 54068 24216 54124
rect 24272 54068 24320 54124
rect 24376 54068 24424 54124
rect 24480 54068 24528 54124
rect 24584 54068 24632 54124
rect 24688 54068 24736 54124
rect 24792 54068 24840 54124
rect 24896 54068 24944 54124
rect 25000 54068 25048 54124
rect 25104 54068 25152 54124
rect 25208 54068 25218 54124
rect 8530 54012 8540 54068
rect 8596 54012 9660 54068
rect 9716 54012 9726 54068
rect 13906 54012 13916 54068
rect 13972 54012 13982 54068
rect 18274 54012 18284 54068
rect 18340 54012 19964 54068
rect 20020 54012 20030 54068
rect 13794 53900 13804 53956
rect 13860 53900 14476 53956
rect 14532 53900 14542 53956
rect 15026 53900 15036 53956
rect 15092 53900 15372 53956
rect 15428 53900 15438 53956
rect 19618 53900 19628 53956
rect 19684 53900 20076 53956
rect 20132 53900 20142 53956
rect 24668 53900 26460 53956
rect 26516 53900 26526 53956
rect 26786 53900 26796 53956
rect 26852 53900 27692 53956
rect 27748 53900 27758 53956
rect 0 53844 800 53872
rect 24668 53844 24724 53900
rect 0 53788 2492 53844
rect 2548 53788 2558 53844
rect 3266 53788 3276 53844
rect 3332 53788 10332 53844
rect 10388 53788 10398 53844
rect 16818 53788 16828 53844
rect 16884 53788 20188 53844
rect 20244 53788 20254 53844
rect 23538 53788 23548 53844
rect 23604 53788 24668 53844
rect 24724 53788 24734 53844
rect 26562 53788 26572 53844
rect 26628 53788 27356 53844
rect 27412 53788 27422 53844
rect 0 53760 800 53788
rect 4050 53676 4060 53732
rect 4116 53676 5628 53732
rect 5684 53676 5694 53732
rect 7858 53676 7868 53732
rect 7924 53676 9772 53732
rect 9828 53676 9838 53732
rect 11442 53676 11452 53732
rect 11508 53676 12236 53732
rect 12292 53676 12302 53732
rect 21634 53676 21644 53732
rect 21700 53676 22876 53732
rect 22932 53676 23660 53732
rect 23716 53676 23726 53732
rect 30930 53676 30940 53732
rect 30996 53676 31276 53732
rect 31332 53676 31342 53732
rect 5730 53564 5740 53620
rect 5796 53564 6188 53620
rect 6244 53564 6254 53620
rect 10658 53564 10668 53620
rect 10724 53564 11900 53620
rect 11956 53564 11966 53620
rect 15026 53564 15036 53620
rect 15092 53508 15148 53620
rect 18946 53564 18956 53620
rect 19012 53564 19404 53620
rect 19460 53564 21532 53620
rect 21588 53564 21598 53620
rect 25666 53564 25676 53620
rect 25732 53564 26908 53620
rect 28466 53564 28476 53620
rect 28532 53564 30268 53620
rect 30324 53564 30334 53620
rect 30818 53564 30828 53620
rect 30884 53564 31388 53620
rect 31444 53564 31948 53620
rect 32004 53564 32014 53620
rect 26852 53508 26908 53564
rect 10882 53452 10892 53508
rect 10948 53452 12348 53508
rect 12404 53452 12414 53508
rect 15092 53452 15372 53508
rect 15428 53452 15438 53508
rect 25106 53452 25116 53508
rect 25172 53452 25900 53508
rect 25956 53452 25966 53508
rect 26852 53452 29372 53508
rect 29428 53452 29438 53508
rect 13998 53284 14008 53340
rect 14064 53284 14112 53340
rect 14168 53284 14216 53340
rect 14272 53284 14320 53340
rect 14376 53284 14424 53340
rect 14480 53284 14528 53340
rect 14584 53284 14632 53340
rect 14688 53284 14736 53340
rect 14792 53284 14840 53340
rect 14896 53284 14944 53340
rect 15000 53284 15048 53340
rect 15104 53284 15152 53340
rect 15208 53284 15218 53340
rect 33998 53284 34008 53340
rect 34064 53284 34112 53340
rect 34168 53284 34216 53340
rect 34272 53284 34320 53340
rect 34376 53284 34424 53340
rect 34480 53284 34528 53340
rect 34584 53284 34632 53340
rect 34688 53284 34736 53340
rect 34792 53284 34840 53340
rect 34896 53284 34944 53340
rect 35000 53284 35048 53340
rect 35104 53284 35152 53340
rect 35208 53284 35218 53340
rect 3266 53228 3276 53284
rect 3332 53228 11228 53284
rect 11284 53228 11564 53284
rect 11620 53228 11630 53284
rect 22194 53228 22204 53284
rect 22260 53228 22652 53284
rect 22708 53228 23772 53284
rect 23828 53228 24220 53284
rect 24276 53228 24286 53284
rect 3462 53116 3500 53172
rect 3556 53116 3566 53172
rect 5170 53116 5180 53172
rect 5236 53116 5852 53172
rect 5908 53116 6524 53172
rect 6580 53116 7308 53172
rect 7364 53116 7420 53172
rect 7476 53116 7486 53172
rect 10098 53116 10108 53172
rect 10164 53116 25340 53172
rect 25396 53116 26460 53172
rect 26516 53116 26526 53172
rect 28466 53116 28476 53172
rect 28532 53116 31276 53172
rect 31332 53116 31342 53172
rect 6066 53004 6076 53060
rect 6132 53004 6300 53060
rect 6356 53004 6366 53060
rect 12562 53004 12572 53060
rect 12628 53004 13580 53060
rect 13636 53004 13646 53060
rect 18274 53004 18284 53060
rect 18340 53004 23660 53060
rect 23716 53004 23726 53060
rect 2482 52892 2492 52948
rect 2548 52892 3500 52948
rect 3556 52892 3566 52948
rect 9426 52892 9436 52948
rect 9492 52892 10780 52948
rect 10836 52892 13916 52948
rect 13972 52892 13982 52948
rect 14130 52892 14140 52948
rect 14196 52892 22316 52948
rect 22372 52892 22382 52948
rect 30258 52892 30268 52948
rect 30324 52892 30828 52948
rect 30884 52892 30894 52948
rect 4722 52780 4732 52836
rect 4788 52780 5292 52836
rect 5348 52780 5358 52836
rect 10994 52780 11004 52836
rect 11060 52780 18956 52836
rect 19012 52780 19022 52836
rect 0 52724 800 52752
rect 0 52668 2044 52724
rect 2100 52668 2828 52724
rect 2884 52668 2894 52724
rect 3164 52668 10556 52724
rect 10612 52668 11788 52724
rect 11844 52668 14140 52724
rect 14196 52668 14206 52724
rect 0 52640 800 52668
rect 3164 52612 3220 52668
rect 3154 52556 3164 52612
rect 3220 52556 3230 52612
rect 6178 52556 6188 52612
rect 6244 52556 19852 52612
rect 19908 52556 20412 52612
rect 20468 52556 21644 52612
rect 21700 52556 21710 52612
rect 3998 52500 4008 52556
rect 4064 52500 4112 52556
rect 4168 52500 4216 52556
rect 4272 52500 4320 52556
rect 4376 52500 4424 52556
rect 4480 52500 4528 52556
rect 4584 52500 4632 52556
rect 4688 52500 4736 52556
rect 4792 52500 4840 52556
rect 4896 52500 4944 52556
rect 5000 52500 5048 52556
rect 5104 52500 5152 52556
rect 5208 52500 5218 52556
rect 23998 52500 24008 52556
rect 24064 52500 24112 52556
rect 24168 52500 24216 52556
rect 24272 52500 24320 52556
rect 24376 52500 24424 52556
rect 24480 52500 24528 52556
rect 24584 52500 24632 52556
rect 24688 52500 24736 52556
rect 24792 52500 24840 52556
rect 24896 52500 24944 52556
rect 25000 52500 25048 52556
rect 25104 52500 25152 52556
rect 25208 52500 25218 52556
rect 11218 52444 11228 52500
rect 11284 52444 13468 52500
rect 13524 52444 13534 52500
rect 22530 52444 22540 52500
rect 22596 52444 22606 52500
rect 10098 52220 10108 52276
rect 10164 52220 11004 52276
rect 11060 52220 11070 52276
rect 11442 52220 11452 52276
rect 11508 52220 11788 52276
rect 11844 52220 11854 52276
rect 22540 52164 22596 52444
rect 23874 52220 23884 52276
rect 23940 52220 25452 52276
rect 25508 52220 25518 52276
rect 30034 52220 30044 52276
rect 30100 52220 31052 52276
rect 31108 52220 31118 52276
rect 10892 52108 11900 52164
rect 11956 52108 12124 52164
rect 12180 52108 12572 52164
rect 12628 52108 12638 52164
rect 19954 52108 19964 52164
rect 20020 52108 21868 52164
rect 21924 52108 23772 52164
rect 23828 52108 24220 52164
rect 24276 52108 25676 52164
rect 25732 52108 25742 52164
rect 30258 52108 30268 52164
rect 30324 52108 31612 52164
rect 31668 52108 31678 52164
rect 10892 52052 10948 52108
rect 4946 51996 4956 52052
rect 5012 51996 5852 52052
rect 5908 51996 5918 52052
rect 10882 51996 10892 52052
rect 10948 51996 10958 52052
rect 11676 51940 11732 52108
rect 13458 51996 13468 52052
rect 13524 51996 14028 52052
rect 14084 51996 14364 52052
rect 14420 51996 14430 52052
rect 15362 51996 15372 52052
rect 15428 51996 16268 52052
rect 16324 51996 16334 52052
rect 19394 51996 19404 52052
rect 19460 51996 20188 52052
rect 20244 51996 21532 52052
rect 21588 51996 21598 52052
rect 23314 51996 23324 52052
rect 23380 51996 25788 52052
rect 25844 51996 27580 52052
rect 27636 51996 27646 52052
rect 30706 51996 30716 52052
rect 30772 51996 31724 52052
rect 31780 51996 31790 52052
rect 3378 51884 3388 51940
rect 3444 51884 3454 51940
rect 6178 51884 6188 51940
rect 6244 51884 8540 51940
rect 8596 51884 9660 51940
rect 9716 51884 9726 51940
rect 11666 51884 11676 51940
rect 11732 51884 11742 51940
rect 15474 51884 15484 51940
rect 15540 51884 21420 51940
rect 21476 51884 21980 51940
rect 22036 51884 23436 51940
rect 23492 51884 23502 51940
rect 30818 51884 30828 51940
rect 30884 51884 32172 51940
rect 32228 51884 32238 51940
rect 33170 51884 33180 51940
rect 33236 51884 34860 51940
rect 34916 51884 34926 51940
rect 3388 51828 3444 51884
rect 3388 51772 3612 51828
rect 3668 51772 3678 51828
rect 13998 51716 14008 51772
rect 14064 51716 14112 51772
rect 14168 51716 14216 51772
rect 14272 51716 14320 51772
rect 14376 51716 14424 51772
rect 14480 51716 14528 51772
rect 14584 51716 14632 51772
rect 14688 51716 14736 51772
rect 14792 51716 14840 51772
rect 14896 51716 14944 51772
rect 15000 51716 15048 51772
rect 15104 51716 15152 51772
rect 15208 51716 15218 51772
rect 33998 51716 34008 51772
rect 34064 51716 34112 51772
rect 34168 51716 34216 51772
rect 34272 51716 34320 51772
rect 34376 51716 34424 51772
rect 34480 51716 34528 51772
rect 34584 51716 34632 51772
rect 34688 51716 34736 51772
rect 34792 51716 34840 51772
rect 34896 51716 34944 51772
rect 35000 51716 35048 51772
rect 35104 51716 35152 51772
rect 35208 51716 35218 51772
rect 3378 51660 3388 51716
rect 3444 51660 3500 51716
rect 3556 51660 3566 51716
rect 4050 51660 4060 51716
rect 4116 51660 5292 51716
rect 5348 51660 6300 51716
rect 6356 51660 6366 51716
rect 9202 51660 9212 51716
rect 9268 51660 13804 51716
rect 13860 51660 13870 51716
rect 0 51604 800 51632
rect 0 51548 1932 51604
rect 1988 51548 1998 51604
rect 4722 51548 4732 51604
rect 4788 51548 6188 51604
rect 6244 51548 6254 51604
rect 13570 51548 13580 51604
rect 13636 51548 14252 51604
rect 14308 51548 14318 51604
rect 22866 51548 22876 51604
rect 22932 51548 23772 51604
rect 23828 51548 24892 51604
rect 24948 51548 25788 51604
rect 25844 51548 26236 51604
rect 26292 51548 26302 51604
rect 30930 51548 30940 51604
rect 30996 51548 33852 51604
rect 33908 51548 33918 51604
rect 0 51520 800 51548
rect 26898 51436 26908 51492
rect 26964 51436 27580 51492
rect 27636 51436 27646 51492
rect 2370 51324 2380 51380
rect 2436 51324 3276 51380
rect 3332 51324 3342 51380
rect 6066 51324 6076 51380
rect 6132 51324 6636 51380
rect 6692 51324 8540 51380
rect 8596 51324 8606 51380
rect 29362 51324 29372 51380
rect 29428 51324 31948 51380
rect 32004 51324 32620 51380
rect 32676 51324 33180 51380
rect 33236 51324 33246 51380
rect 17602 51212 17612 51268
rect 17668 51212 18172 51268
rect 18228 51212 18238 51268
rect 15474 51100 15484 51156
rect 15540 51100 15550 51156
rect 3998 50932 4008 50988
rect 4064 50932 4112 50988
rect 4168 50932 4216 50988
rect 4272 50932 4320 50988
rect 4376 50932 4424 50988
rect 4480 50932 4528 50988
rect 4584 50932 4632 50988
rect 4688 50932 4736 50988
rect 4792 50932 4840 50988
rect 4896 50932 4944 50988
rect 5000 50932 5048 50988
rect 5104 50932 5152 50988
rect 5208 50932 5218 50988
rect 15484 50820 15540 51100
rect 23998 50932 24008 50988
rect 24064 50932 24112 50988
rect 24168 50932 24216 50988
rect 24272 50932 24320 50988
rect 24376 50932 24424 50988
rect 24480 50932 24528 50988
rect 24584 50932 24632 50988
rect 24688 50932 24736 50988
rect 24792 50932 24840 50988
rect 24896 50932 24944 50988
rect 25000 50932 25048 50988
rect 25104 50932 25152 50988
rect 25208 50932 25218 50988
rect 15138 50764 15148 50820
rect 15204 50764 15540 50820
rect 18610 50652 18620 50708
rect 18676 50652 19628 50708
rect 19684 50652 19852 50708
rect 19908 50652 19918 50708
rect 22418 50652 22428 50708
rect 22484 50652 23100 50708
rect 23156 50652 24332 50708
rect 24388 50652 24892 50708
rect 24948 50652 25564 50708
rect 25620 50652 25630 50708
rect 30146 50652 30156 50708
rect 30212 50652 30716 50708
rect 30772 50652 30782 50708
rect 6738 50540 6748 50596
rect 6804 50540 7980 50596
rect 8036 50540 8046 50596
rect 13794 50540 13804 50596
rect 13860 50540 15484 50596
rect 15540 50540 15550 50596
rect 17378 50540 17388 50596
rect 17444 50540 18844 50596
rect 18900 50540 18910 50596
rect 0 50484 800 50512
rect 0 50428 2156 50484
rect 2212 50428 2222 50484
rect 4946 50428 4956 50484
rect 5012 50428 6636 50484
rect 6692 50428 6972 50484
rect 7028 50428 7038 50484
rect 7298 50428 7308 50484
rect 7364 50428 8316 50484
rect 8372 50428 8382 50484
rect 14802 50428 14812 50484
rect 14868 50428 17276 50484
rect 17332 50428 17342 50484
rect 19282 50428 19292 50484
rect 19348 50428 23996 50484
rect 24052 50428 24062 50484
rect 33814 50428 33852 50484
rect 33908 50428 34524 50484
rect 34580 50428 34590 50484
rect 0 50400 800 50428
rect 15922 50372 15932 50428
rect 15988 50372 15998 50428
rect 13570 50316 13580 50372
rect 13636 50316 13916 50372
rect 13972 50316 13982 50372
rect 14354 50316 14364 50372
rect 14420 50316 15708 50372
rect 15764 50316 15774 50372
rect 27122 50316 27132 50372
rect 27188 50316 28028 50372
rect 28084 50316 28094 50372
rect 13998 50148 14008 50204
rect 14064 50148 14112 50204
rect 14168 50148 14216 50204
rect 14272 50148 14320 50204
rect 14376 50148 14424 50204
rect 14480 50148 14528 50204
rect 14584 50148 14632 50204
rect 14688 50148 14736 50204
rect 14792 50148 14840 50204
rect 14896 50148 14944 50204
rect 15000 50148 15048 50204
rect 15104 50148 15152 50204
rect 15208 50148 15218 50204
rect 33998 50148 34008 50204
rect 34064 50148 34112 50204
rect 34168 50148 34216 50204
rect 34272 50148 34320 50204
rect 34376 50148 34424 50204
rect 34480 50148 34528 50204
rect 34584 50148 34632 50204
rect 34688 50148 34736 50204
rect 34792 50148 34840 50204
rect 34896 50148 34944 50204
rect 35000 50148 35048 50204
rect 35104 50148 35152 50204
rect 35208 50148 35218 50204
rect 4498 49980 4508 50036
rect 4564 49980 5516 50036
rect 5572 49980 5582 50036
rect 8642 49980 8652 50036
rect 8708 49980 9660 50036
rect 9716 49980 10220 50036
rect 10276 49980 10286 50036
rect 3602 49868 3612 49924
rect 3668 49868 26460 49924
rect 26516 49868 27692 49924
rect 27748 49868 27758 49924
rect 11218 49756 11228 49812
rect 11284 49756 11676 49812
rect 11732 49756 11742 49812
rect 16482 49756 16492 49812
rect 16548 49756 18956 49812
rect 19012 49756 19022 49812
rect 9762 49644 9772 49700
rect 9828 49644 10332 49700
rect 10388 49644 13468 49700
rect 13524 49644 13534 49700
rect 14242 49644 14252 49700
rect 14308 49644 15708 49700
rect 15764 49644 15774 49700
rect 15922 49644 15932 49700
rect 15988 49644 17500 49700
rect 17556 49644 17566 49700
rect 31154 49644 31164 49700
rect 31220 49644 33180 49700
rect 33236 49644 33740 49700
rect 33796 49644 33806 49700
rect 7634 49532 7644 49588
rect 7700 49532 8540 49588
rect 8596 49532 8606 49588
rect 0 49364 800 49392
rect 3998 49364 4008 49420
rect 4064 49364 4112 49420
rect 4168 49364 4216 49420
rect 4272 49364 4320 49420
rect 4376 49364 4424 49420
rect 4480 49364 4528 49420
rect 4584 49364 4632 49420
rect 4688 49364 4736 49420
rect 4792 49364 4840 49420
rect 4896 49364 4944 49420
rect 5000 49364 5048 49420
rect 5104 49364 5152 49420
rect 5208 49364 5218 49420
rect 23998 49364 24008 49420
rect 24064 49364 24112 49420
rect 24168 49364 24216 49420
rect 24272 49364 24320 49420
rect 24376 49364 24424 49420
rect 24480 49364 24528 49420
rect 24584 49364 24632 49420
rect 24688 49364 24736 49420
rect 24792 49364 24840 49420
rect 24896 49364 24944 49420
rect 25000 49364 25048 49420
rect 25104 49364 25152 49420
rect 25208 49364 25218 49420
rect 0 49308 2492 49364
rect 2548 49308 2558 49364
rect 11218 49308 11228 49364
rect 11284 49308 11564 49364
rect 11620 49308 11788 49364
rect 11844 49308 11854 49364
rect 0 49280 800 49308
rect 11732 49252 11788 49308
rect 11732 49196 12908 49252
rect 12964 49196 20188 49252
rect 20244 49196 20254 49252
rect 25442 49196 25452 49252
rect 25508 49196 26236 49252
rect 26292 49196 26302 49252
rect 26852 49196 29596 49252
rect 29652 49196 29662 49252
rect 31714 49196 31724 49252
rect 31780 49196 33516 49252
rect 33572 49196 33582 49252
rect 18834 49084 18844 49140
rect 18900 49084 20076 49140
rect 20132 49084 20142 49140
rect 26852 49028 26908 49196
rect 31042 49084 31052 49140
rect 31108 49084 32172 49140
rect 32228 49084 32238 49140
rect 13794 48972 13804 49028
rect 13860 48972 13916 49028
rect 13972 48972 13982 49028
rect 15362 48972 15372 49028
rect 15428 48972 15820 49028
rect 15876 48972 16156 49028
rect 16212 48972 17052 49028
rect 17108 48972 17118 49028
rect 24322 48972 24332 49028
rect 24388 48972 25676 49028
rect 25732 48972 26684 49028
rect 26740 48972 26908 49028
rect 27010 48972 27020 49028
rect 27076 48972 27086 49028
rect 33058 48972 33068 49028
rect 33124 48972 33628 49028
rect 33684 48972 33694 49028
rect 27020 48916 27076 48972
rect 3826 48860 3836 48916
rect 3892 48860 5628 48916
rect 5684 48860 5694 48916
rect 12786 48860 12796 48916
rect 12852 48860 14252 48916
rect 14308 48860 14318 48916
rect 14690 48860 14700 48916
rect 14756 48860 15652 48916
rect 17938 48860 17948 48916
rect 18004 48860 18620 48916
rect 18676 48860 18686 48916
rect 25330 48860 25340 48916
rect 25396 48860 26236 48916
rect 26292 48860 27076 48916
rect 31602 48860 31612 48916
rect 31668 48860 32284 48916
rect 32340 48860 32350 48916
rect 15596 48804 15652 48860
rect 5730 48748 5740 48804
rect 5796 48748 11788 48804
rect 11844 48748 13524 48804
rect 13682 48748 13692 48804
rect 13748 48748 15372 48804
rect 15428 48748 15438 48804
rect 15586 48748 15596 48804
rect 15652 48748 16716 48804
rect 16772 48748 16782 48804
rect 17714 48748 17724 48804
rect 17780 48748 19628 48804
rect 19684 48748 26908 48804
rect 26964 48748 28588 48804
rect 28644 48748 31836 48804
rect 31892 48748 31902 48804
rect 33842 48748 33852 48804
rect 33908 48748 34300 48804
rect 34356 48748 35364 48804
rect 13468 48692 13524 48748
rect 35308 48692 35364 48748
rect 13468 48636 13580 48692
rect 13636 48636 13646 48692
rect 22306 48636 22316 48692
rect 22372 48636 23324 48692
rect 23380 48636 23390 48692
rect 35308 48636 36428 48692
rect 36484 48636 36494 48692
rect 13998 48580 14008 48636
rect 14064 48580 14112 48636
rect 14168 48580 14216 48636
rect 14272 48580 14320 48636
rect 14376 48580 14424 48636
rect 14480 48580 14528 48636
rect 14584 48580 14632 48636
rect 14688 48580 14736 48636
rect 14792 48580 14840 48636
rect 14896 48580 14944 48636
rect 15000 48580 15048 48636
rect 15104 48580 15152 48636
rect 15208 48580 15218 48636
rect 33998 48580 34008 48636
rect 34064 48580 34112 48636
rect 34168 48580 34216 48636
rect 34272 48580 34320 48636
rect 34376 48580 34424 48636
rect 34480 48580 34528 48636
rect 34584 48580 34632 48636
rect 34688 48580 34736 48636
rect 34792 48580 34840 48636
rect 34896 48580 34944 48636
rect 35000 48580 35048 48636
rect 35104 48580 35152 48636
rect 35208 48580 35218 48636
rect 3266 48524 3276 48580
rect 3332 48524 9436 48580
rect 9492 48524 9502 48580
rect 30370 48524 30380 48580
rect 30436 48524 31276 48580
rect 31332 48524 31342 48580
rect 6850 48412 6860 48468
rect 6916 48412 11004 48468
rect 11060 48412 11070 48468
rect 22866 48412 22876 48468
rect 22932 48412 23884 48468
rect 23940 48412 24444 48468
rect 24500 48412 24510 48468
rect 28690 48412 28700 48468
rect 28756 48412 30828 48468
rect 30884 48412 30894 48468
rect 23650 48300 23660 48356
rect 23716 48300 25340 48356
rect 25396 48300 27020 48356
rect 27076 48300 27086 48356
rect 30482 48300 30492 48356
rect 30548 48300 31276 48356
rect 31332 48300 31342 48356
rect 0 48244 800 48272
rect 0 48188 2492 48244
rect 2548 48188 2940 48244
rect 2996 48188 3006 48244
rect 8530 48188 8540 48244
rect 8596 48188 9996 48244
rect 10052 48188 10062 48244
rect 11666 48188 11676 48244
rect 11732 48188 15932 48244
rect 15988 48188 15998 48244
rect 20962 48188 20972 48244
rect 21028 48188 23772 48244
rect 23828 48188 23838 48244
rect 27346 48188 27356 48244
rect 27412 48188 31164 48244
rect 31220 48188 31230 48244
rect 31826 48188 31836 48244
rect 31892 48188 32060 48244
rect 32116 48188 32126 48244
rect 32498 48188 32508 48244
rect 32564 48188 34076 48244
rect 34132 48188 34142 48244
rect 0 48160 800 48188
rect 4610 48076 4620 48132
rect 4676 48076 5292 48132
rect 5348 48076 5358 48132
rect 8978 48076 8988 48132
rect 9044 48076 9884 48132
rect 9940 48076 9950 48132
rect 13346 48076 13356 48132
rect 13412 48076 14588 48132
rect 14644 48076 15372 48132
rect 15428 48076 15438 48132
rect 3998 47796 4008 47852
rect 4064 47796 4112 47852
rect 4168 47796 4216 47852
rect 4272 47796 4320 47852
rect 4376 47796 4424 47852
rect 4480 47796 4528 47852
rect 4584 47796 4632 47852
rect 4688 47796 4736 47852
rect 4792 47796 4840 47852
rect 4896 47796 4944 47852
rect 5000 47796 5048 47852
rect 5104 47796 5152 47852
rect 5208 47796 5218 47852
rect 23998 47796 24008 47852
rect 24064 47796 24112 47852
rect 24168 47796 24216 47852
rect 24272 47796 24320 47852
rect 24376 47796 24424 47852
rect 24480 47796 24528 47852
rect 24584 47796 24632 47852
rect 24688 47796 24736 47852
rect 24792 47796 24840 47852
rect 24896 47796 24944 47852
rect 25000 47796 25048 47852
rect 25104 47796 25152 47852
rect 25208 47796 25218 47852
rect 8754 47628 8764 47684
rect 8820 47628 9884 47684
rect 9940 47628 9950 47684
rect 3378 47516 3388 47572
rect 3444 47516 3482 47572
rect 12114 47516 12124 47572
rect 12180 47516 13580 47572
rect 13636 47516 13646 47572
rect 21410 47516 21420 47572
rect 21476 47516 22092 47572
rect 22148 47516 22158 47572
rect 23762 47516 23772 47572
rect 23828 47516 24444 47572
rect 24500 47516 25788 47572
rect 25844 47516 29260 47572
rect 29316 47516 29326 47572
rect 3266 47404 3276 47460
rect 3332 47404 10108 47460
rect 10164 47404 10668 47460
rect 10724 47404 10734 47460
rect 13794 47404 13804 47460
rect 13860 47404 13916 47460
rect 13972 47404 13982 47460
rect 15092 47404 17612 47460
rect 17668 47404 17678 47460
rect 22530 47404 22540 47460
rect 22596 47404 23660 47460
rect 23716 47404 23726 47460
rect 30706 47404 30716 47460
rect 30772 47404 31500 47460
rect 31556 47404 32172 47460
rect 32228 47404 32238 47460
rect 2594 47292 2604 47348
rect 2660 47292 3388 47348
rect 3444 47292 3724 47348
rect 3780 47292 3790 47348
rect 9090 47292 9100 47348
rect 9156 47292 11228 47348
rect 11284 47292 13580 47348
rect 13636 47292 13646 47348
rect 15092 47236 15148 47404
rect 29474 47292 29484 47348
rect 29540 47292 30380 47348
rect 30436 47292 30446 47348
rect 7074 47180 7084 47236
rect 7140 47180 8092 47236
rect 8148 47180 8158 47236
rect 13468 47180 14700 47236
rect 14756 47180 15148 47236
rect 19842 47180 19852 47236
rect 19908 47180 21644 47236
rect 21700 47180 21980 47236
rect 22036 47180 23996 47236
rect 24052 47180 25340 47236
rect 25396 47180 25406 47236
rect 31266 47180 31276 47236
rect 31332 47180 32172 47236
rect 32228 47180 32238 47236
rect 0 47124 800 47152
rect 0 47068 2156 47124
rect 2212 47068 2828 47124
rect 2884 47068 2894 47124
rect 4946 47068 4956 47124
rect 5012 47068 5292 47124
rect 5348 47068 9436 47124
rect 9492 47068 9502 47124
rect 0 47040 800 47068
rect 13468 47012 13524 47180
rect 27122 47068 27132 47124
rect 27188 47068 27198 47124
rect 13998 47012 14008 47068
rect 14064 47012 14112 47068
rect 14168 47012 14216 47068
rect 14272 47012 14320 47068
rect 14376 47012 14424 47068
rect 14480 47012 14528 47068
rect 14584 47012 14632 47068
rect 14688 47012 14736 47068
rect 14792 47012 14840 47068
rect 14896 47012 14944 47068
rect 15000 47012 15048 47068
rect 15104 47012 15152 47068
rect 15208 47012 15218 47068
rect 18610 47012 18620 47068
rect 18676 47012 18686 47068
rect 27132 47012 27188 47068
rect 33998 47012 34008 47068
rect 34064 47012 34112 47068
rect 34168 47012 34216 47068
rect 34272 47012 34320 47068
rect 34376 47012 34424 47068
rect 34480 47012 34528 47068
rect 34584 47012 34632 47068
rect 34688 47012 34736 47068
rect 34792 47012 34840 47068
rect 34896 47012 34944 47068
rect 35000 47012 35048 47068
rect 35104 47012 35152 47068
rect 35208 47012 35218 47068
rect 4834 46956 4844 47012
rect 4900 46956 5628 47012
rect 5684 46956 13244 47012
rect 13300 46956 13524 47012
rect 15362 46956 15372 47012
rect 15428 46956 17276 47012
rect 17332 46956 17342 47012
rect 18386 46956 18396 47012
rect 18452 46956 18676 47012
rect 27132 46956 28364 47012
rect 28420 46956 28430 47012
rect 28690 46956 28700 47012
rect 28756 46956 29596 47012
rect 29652 46956 32732 47012
rect 32788 46956 32798 47012
rect 5506 46844 5516 46900
rect 5572 46844 7420 46900
rect 7476 46844 7486 46900
rect 13906 46844 13916 46900
rect 13972 46844 18956 46900
rect 19012 46844 19022 46900
rect 22754 46844 22764 46900
rect 22820 46844 23772 46900
rect 23828 46844 23838 46900
rect 26450 46844 26460 46900
rect 26516 46844 27916 46900
rect 27972 46844 27982 46900
rect 31602 46844 31612 46900
rect 31668 46844 32172 46900
rect 32228 46844 36316 46900
rect 36372 46844 36382 46900
rect 5730 46732 5740 46788
rect 5796 46732 6412 46788
rect 6468 46732 6860 46788
rect 6916 46732 6926 46788
rect 18274 46732 18284 46788
rect 18340 46732 22876 46788
rect 22932 46732 22942 46788
rect 26562 46732 26572 46788
rect 26628 46732 27468 46788
rect 27524 46732 27534 46788
rect 32386 46732 32396 46788
rect 32452 46732 34524 46788
rect 34580 46732 34590 46788
rect 2482 46620 2492 46676
rect 2548 46620 3836 46676
rect 3892 46620 3902 46676
rect 9426 46620 9436 46676
rect 9492 46620 9996 46676
rect 10052 46620 11004 46676
rect 11060 46620 11788 46676
rect 11844 46620 11854 46676
rect 32610 46620 32620 46676
rect 32676 46620 34188 46676
rect 34244 46620 36204 46676
rect 36260 46620 37100 46676
rect 37156 46620 37884 46676
rect 37940 46620 37950 46676
rect 9090 46508 9100 46564
rect 9156 46508 11452 46564
rect 11508 46508 11518 46564
rect 17574 46508 17612 46564
rect 17668 46508 17678 46564
rect 26002 46508 26012 46564
rect 26068 46508 26572 46564
rect 26628 46508 26638 46564
rect 31938 46508 31948 46564
rect 32004 46508 33180 46564
rect 33236 46508 35756 46564
rect 35812 46508 35822 46564
rect 33618 46396 33628 46452
rect 33684 46396 35308 46452
rect 35364 46396 35644 46452
rect 35700 46396 35980 46452
rect 36036 46396 37548 46452
rect 37604 46396 37614 46452
rect 32274 46284 32284 46340
rect 32340 46284 34636 46340
rect 34692 46284 35532 46340
rect 35588 46284 36316 46340
rect 36372 46284 37996 46340
rect 38052 46284 38062 46340
rect 3998 46228 4008 46284
rect 4064 46228 4112 46284
rect 4168 46228 4216 46284
rect 4272 46228 4320 46284
rect 4376 46228 4424 46284
rect 4480 46228 4528 46284
rect 4584 46228 4632 46284
rect 4688 46228 4736 46284
rect 4792 46228 4840 46284
rect 4896 46228 4944 46284
rect 5000 46228 5048 46284
rect 5104 46228 5152 46284
rect 5208 46228 5218 46284
rect 23998 46228 24008 46284
rect 24064 46228 24112 46284
rect 24168 46228 24216 46284
rect 24272 46228 24320 46284
rect 24376 46228 24424 46284
rect 24480 46228 24528 46284
rect 24584 46228 24632 46284
rect 24688 46228 24736 46284
rect 24792 46228 24840 46284
rect 24896 46228 24944 46284
rect 25000 46228 25048 46284
rect 25104 46228 25152 46284
rect 25208 46228 25218 46284
rect 30146 46060 30156 46116
rect 30212 46060 30940 46116
rect 30996 46060 31006 46116
rect 0 46004 800 46032
rect 0 45948 2492 46004
rect 2548 45948 2558 46004
rect 3266 45948 3276 46004
rect 3332 45948 9324 46004
rect 9380 45948 9390 46004
rect 25750 45948 25788 46004
rect 25844 45948 25854 46004
rect 0 45920 800 45948
rect 11778 45836 11788 45892
rect 11844 45836 13132 45892
rect 13188 45836 13804 45892
rect 13860 45836 13870 45892
rect 16370 45836 16380 45892
rect 16436 45836 17500 45892
rect 17556 45836 17566 45892
rect 21298 45836 21308 45892
rect 21364 45836 22204 45892
rect 22260 45836 22270 45892
rect 24770 45836 24780 45892
rect 24836 45836 26236 45892
rect 26292 45836 26302 45892
rect 35746 45836 35756 45892
rect 35812 45836 37100 45892
rect 37156 45836 37166 45892
rect 4946 45724 4956 45780
rect 5012 45724 5516 45780
rect 5572 45724 5582 45780
rect 16594 45724 16604 45780
rect 16660 45724 17612 45780
rect 17668 45724 17678 45780
rect 24098 45724 24108 45780
rect 24164 45724 26012 45780
rect 26068 45724 26078 45780
rect 27794 45724 27804 45780
rect 27860 45724 28700 45780
rect 28756 45724 30044 45780
rect 30100 45724 30110 45780
rect 35410 45724 35420 45780
rect 35476 45724 36988 45780
rect 37044 45724 37054 45780
rect 18722 45612 18732 45668
rect 18788 45612 18798 45668
rect 19618 45612 19628 45668
rect 19684 45612 21532 45668
rect 21588 45612 21868 45668
rect 21924 45612 24332 45668
rect 24388 45612 24398 45668
rect 28130 45612 28140 45668
rect 28196 45612 29260 45668
rect 29316 45612 29820 45668
rect 29876 45612 33180 45668
rect 33236 45612 33246 45668
rect 13998 45444 14008 45500
rect 14064 45444 14112 45500
rect 14168 45444 14216 45500
rect 14272 45444 14320 45500
rect 14376 45444 14424 45500
rect 14480 45444 14528 45500
rect 14584 45444 14632 45500
rect 14688 45444 14736 45500
rect 14792 45444 14840 45500
rect 14896 45444 14944 45500
rect 15000 45444 15048 45500
rect 15104 45444 15152 45500
rect 15208 45444 15218 45500
rect 5842 45388 5852 45444
rect 5908 45388 7196 45444
rect 7252 45388 8204 45444
rect 8260 45388 10892 45444
rect 10948 45388 11788 45444
rect 11844 45388 11854 45444
rect 18732 45332 18788 45612
rect 19282 45500 19292 45556
rect 19348 45500 29372 45556
rect 29428 45500 29438 45556
rect 33998 45444 34008 45500
rect 34064 45444 34112 45500
rect 34168 45444 34216 45500
rect 34272 45444 34320 45500
rect 34376 45444 34424 45500
rect 34480 45444 34528 45500
rect 34584 45444 34632 45500
rect 34688 45444 34736 45500
rect 34792 45444 34840 45500
rect 34896 45444 34944 45500
rect 35000 45444 35048 45500
rect 35104 45444 35152 45500
rect 35208 45444 35218 45500
rect 26852 45388 33628 45444
rect 33684 45388 33908 45444
rect 26852 45332 26908 45388
rect 7298 45276 7308 45332
rect 7364 45276 11340 45332
rect 11396 45276 11406 45332
rect 13654 45276 13692 45332
rect 13748 45276 14140 45332
rect 14196 45276 14206 45332
rect 15922 45276 15932 45332
rect 15988 45276 16380 45332
rect 16436 45276 16446 45332
rect 16594 45276 16604 45332
rect 16660 45276 17724 45332
rect 17780 45276 17790 45332
rect 18274 45276 18284 45332
rect 18340 45276 19180 45332
rect 19236 45276 19246 45332
rect 22306 45276 22316 45332
rect 22372 45276 23548 45332
rect 23604 45276 23614 45332
rect 24322 45276 24332 45332
rect 24388 45276 26908 45332
rect 33852 45332 33908 45388
rect 33852 45276 34300 45332
rect 34356 45276 34366 45332
rect 16380 45220 16436 45276
rect 3266 45164 3276 45220
rect 3332 44996 3388 45220
rect 4162 45164 4172 45220
rect 4228 45164 5628 45220
rect 5684 45164 5694 45220
rect 9986 45164 9996 45220
rect 10052 45164 11788 45220
rect 11844 45164 15820 45220
rect 15876 45164 15886 45220
rect 16380 45164 17388 45220
rect 17444 45164 17454 45220
rect 18284 45108 18340 45276
rect 24332 45220 24388 45276
rect 23426 45164 23436 45220
rect 23492 45164 24388 45220
rect 34850 45164 34860 45220
rect 34916 45164 35980 45220
rect 36036 45164 36046 45220
rect 7634 45052 7644 45108
rect 7700 45052 7980 45108
rect 8036 45052 8046 45108
rect 9650 45052 9660 45108
rect 9716 45052 10556 45108
rect 10612 45052 10780 45108
rect 10836 45052 10846 45108
rect 13122 45052 13132 45108
rect 13188 45052 13804 45108
rect 13860 45052 13870 45108
rect 14130 45052 14140 45108
rect 14196 45052 14206 45108
rect 14354 45052 14364 45108
rect 14420 45052 15148 45108
rect 15204 45052 15214 45108
rect 15362 45052 15372 45108
rect 15428 45052 18340 45108
rect 21746 45052 21756 45108
rect 21812 45052 25788 45108
rect 25844 45052 25854 45108
rect 26338 45052 26348 45108
rect 26404 45052 27692 45108
rect 27748 45052 27758 45108
rect 14140 44996 14196 45052
rect 3332 44940 6076 44996
rect 6132 44940 8036 44996
rect 14140 44940 15484 44996
rect 15540 44940 16828 44996
rect 16884 44940 16894 44996
rect 22306 44940 22316 44996
rect 22372 44940 25452 44996
rect 25508 44940 26124 44996
rect 26180 44940 27244 44996
rect 27300 44940 27580 44996
rect 27636 44940 27646 44996
rect 32498 44940 32508 44996
rect 32564 44940 33852 44996
rect 33908 44940 33918 44996
rect 0 44884 800 44912
rect 0 44828 2492 44884
rect 2548 44828 2558 44884
rect 3836 44828 4396 44884
rect 4452 44828 4462 44884
rect 5282 44828 5292 44884
rect 5348 44828 5964 44884
rect 6020 44828 6030 44884
rect 0 44800 800 44828
rect 3836 44548 3892 44828
rect 7298 44716 7308 44772
rect 7364 44716 7644 44772
rect 7700 44716 7710 44772
rect 3998 44660 4008 44716
rect 4064 44660 4112 44716
rect 4168 44660 4216 44716
rect 4272 44660 4320 44716
rect 4376 44660 4424 44716
rect 4480 44660 4528 44716
rect 4584 44660 4632 44716
rect 4688 44660 4736 44716
rect 4792 44660 4840 44716
rect 4896 44660 4944 44716
rect 5000 44660 5048 44716
rect 5104 44660 5152 44716
rect 5208 44660 5218 44716
rect 3798 44492 3836 44548
rect 3892 44492 4396 44548
rect 4452 44492 4462 44548
rect 6738 44380 6748 44436
rect 6804 44380 7308 44436
rect 7364 44380 7374 44436
rect 7644 44324 7700 44716
rect 7980 44660 8036 44940
rect 13682 44828 13692 44884
rect 13748 44828 15932 44884
rect 15988 44828 15998 44884
rect 17378 44828 17388 44884
rect 17444 44828 18620 44884
rect 18676 44828 19852 44884
rect 19908 44828 19918 44884
rect 25106 44828 25116 44884
rect 25172 44828 26236 44884
rect 26292 44828 26302 44884
rect 34738 44828 34748 44884
rect 34804 44828 35980 44884
rect 36036 44828 36046 44884
rect 13794 44716 13804 44772
rect 13860 44716 14364 44772
rect 14420 44716 14430 44772
rect 15092 44716 15372 44772
rect 15428 44716 15438 44772
rect 15092 44660 15148 44716
rect 23998 44660 24008 44716
rect 24064 44660 24112 44716
rect 24168 44660 24216 44716
rect 24272 44660 24320 44716
rect 24376 44660 24424 44716
rect 24480 44660 24528 44716
rect 24584 44660 24632 44716
rect 24688 44660 24736 44716
rect 24792 44660 24840 44716
rect 24896 44660 24944 44716
rect 25000 44660 25048 44716
rect 25104 44660 25152 44716
rect 25208 44660 25218 44716
rect 7980 44604 15148 44660
rect 17602 44492 17612 44548
rect 17668 44492 18956 44548
rect 19012 44492 19022 44548
rect 10994 44380 11004 44436
rect 11060 44380 11676 44436
rect 11732 44380 12908 44436
rect 12964 44380 13468 44436
rect 13524 44380 13534 44436
rect 17714 44380 17724 44436
rect 17780 44380 18508 44436
rect 18564 44380 18574 44436
rect 23762 44380 23772 44436
rect 23828 44380 23884 44436
rect 23940 44380 23950 44436
rect 7644 44268 8092 44324
rect 8148 44268 8158 44324
rect 8306 44268 8316 44324
rect 8372 44268 9660 44324
rect 9716 44268 9726 44324
rect 10098 44268 10108 44324
rect 10164 44268 10174 44324
rect 21970 44268 21980 44324
rect 22036 44268 26012 44324
rect 26068 44268 26078 44324
rect 33506 44268 33516 44324
rect 33572 44268 33740 44324
rect 33796 44268 34524 44324
rect 34580 44268 34590 44324
rect 35858 44268 35868 44324
rect 35924 44268 37548 44324
rect 37604 44268 37614 44324
rect 4946 44156 4956 44212
rect 5012 44156 5292 44212
rect 5348 44156 6412 44212
rect 6468 44156 6478 44212
rect 10108 44100 10164 44268
rect 21980 44212 22036 44268
rect 10546 44156 10556 44212
rect 10612 44156 11452 44212
rect 11508 44156 11518 44212
rect 17602 44156 17612 44212
rect 17668 44156 18172 44212
rect 18228 44156 19068 44212
rect 19124 44156 19134 44212
rect 19954 44156 19964 44212
rect 20020 44156 20412 44212
rect 20468 44156 22036 44212
rect 33628 44156 34636 44212
rect 34692 44156 34702 44212
rect 33628 44100 33684 44156
rect 2258 44044 2268 44100
rect 2324 44044 3836 44100
rect 3892 44044 3902 44100
rect 6514 44044 6524 44100
rect 6580 44044 11004 44100
rect 11060 44044 11340 44100
rect 11396 44044 12572 44100
rect 12628 44044 12638 44100
rect 22978 44044 22988 44100
rect 23044 44044 23660 44100
rect 23716 44044 23726 44100
rect 33618 44044 33628 44100
rect 33684 44044 33694 44100
rect 33842 44044 33852 44100
rect 33908 44044 35308 44100
rect 35364 44044 35374 44100
rect 3378 43932 3388 43988
rect 3444 43932 10388 43988
rect 18610 43932 18620 43988
rect 18676 43932 18900 43988
rect 1596 43820 3388 43876
rect 3444 43820 3454 43876
rect 4722 43820 4732 43876
rect 4788 43820 6076 43876
rect 6132 43820 6142 43876
rect 0 43764 800 43792
rect 1596 43764 1652 43820
rect 10332 43764 10388 43932
rect 13998 43876 14008 43932
rect 14064 43876 14112 43932
rect 14168 43876 14216 43932
rect 14272 43876 14320 43932
rect 14376 43876 14424 43932
rect 14480 43876 14528 43932
rect 14584 43876 14632 43932
rect 14688 43876 14736 43932
rect 14792 43876 14840 43932
rect 14896 43876 14944 43932
rect 15000 43876 15048 43932
rect 15104 43876 15152 43932
rect 15208 43876 15218 43932
rect 18844 43876 18900 43932
rect 33998 43876 34008 43932
rect 34064 43876 34112 43932
rect 34168 43876 34216 43932
rect 34272 43876 34320 43932
rect 34376 43876 34424 43932
rect 34480 43876 34528 43932
rect 34584 43876 34632 43932
rect 34688 43876 34736 43932
rect 34792 43876 34840 43932
rect 34896 43876 34944 43932
rect 35000 43876 35048 43932
rect 35104 43876 35152 43932
rect 35208 43876 35218 43932
rect 18834 43820 18844 43876
rect 18900 43820 19516 43876
rect 19572 43820 19582 43876
rect 0 43708 1652 43764
rect 1810 43708 1820 43764
rect 1876 43708 5628 43764
rect 5684 43708 6972 43764
rect 7028 43708 7038 43764
rect 8082 43708 8092 43764
rect 8148 43708 10108 43764
rect 10164 43708 10174 43764
rect 10332 43708 20972 43764
rect 21028 43708 21532 43764
rect 21588 43708 21598 43764
rect 0 43680 800 43708
rect 3378 43596 3388 43652
rect 3444 43596 3482 43652
rect 11106 43596 11116 43652
rect 11172 43596 13916 43652
rect 13972 43596 14252 43652
rect 14308 43596 14318 43652
rect 15474 43596 15484 43652
rect 15540 43596 17388 43652
rect 17444 43596 17454 43652
rect 18050 43596 18060 43652
rect 18116 43596 19740 43652
rect 19796 43596 19806 43652
rect 29138 43596 29148 43652
rect 29204 43596 30492 43652
rect 30548 43596 30558 43652
rect 36418 43596 36428 43652
rect 36484 43596 37660 43652
rect 37716 43596 37884 43652
rect 37940 43596 37950 43652
rect 10658 43484 10668 43540
rect 10724 43484 12348 43540
rect 12404 43484 12414 43540
rect 14466 43484 14476 43540
rect 14532 43484 19292 43540
rect 19348 43484 19358 43540
rect 19516 43484 20188 43540
rect 20244 43484 20254 43540
rect 29474 43484 29484 43540
rect 29540 43484 30156 43540
rect 30212 43484 30222 43540
rect 19516 43428 19572 43484
rect 4162 43372 4172 43428
rect 4228 43372 5740 43428
rect 5796 43372 5806 43428
rect 8194 43372 8204 43428
rect 8260 43372 8540 43428
rect 8596 43372 11452 43428
rect 11508 43372 12796 43428
rect 12852 43372 12862 43428
rect 13346 43372 13356 43428
rect 13412 43372 14140 43428
rect 14196 43372 14206 43428
rect 16594 43372 16604 43428
rect 16660 43372 18956 43428
rect 19012 43372 19572 43428
rect 19842 43372 19852 43428
rect 19908 43372 21756 43428
rect 21812 43372 21822 43428
rect 29362 43372 29372 43428
rect 29428 43372 30940 43428
rect 30996 43372 32508 43428
rect 32564 43372 32574 43428
rect 33506 43372 33516 43428
rect 33572 43372 34636 43428
rect 34692 43372 34702 43428
rect 16146 43260 16156 43316
rect 16212 43260 18396 43316
rect 18452 43260 21420 43316
rect 21476 43260 26012 43316
rect 26068 43260 26796 43316
rect 26852 43260 26862 43316
rect 16706 43148 16716 43204
rect 16772 43148 17500 43204
rect 17556 43148 17566 43204
rect 3998 43092 4008 43148
rect 4064 43092 4112 43148
rect 4168 43092 4216 43148
rect 4272 43092 4320 43148
rect 4376 43092 4424 43148
rect 4480 43092 4528 43148
rect 4584 43092 4632 43148
rect 4688 43092 4736 43148
rect 4792 43092 4840 43148
rect 4896 43092 4944 43148
rect 5000 43092 5048 43148
rect 5104 43092 5152 43148
rect 5208 43092 5218 43148
rect 23998 43092 24008 43148
rect 24064 43092 24112 43148
rect 24168 43092 24216 43148
rect 24272 43092 24320 43148
rect 24376 43092 24424 43148
rect 24480 43092 24528 43148
rect 24584 43092 24632 43148
rect 24688 43092 24736 43148
rect 24792 43092 24840 43148
rect 24896 43092 24944 43148
rect 25000 43092 25048 43148
rect 25104 43092 25152 43148
rect 25208 43092 25218 43148
rect 9986 43036 9996 43092
rect 10052 43036 10062 43092
rect 33394 43036 33404 43092
rect 33460 43036 33852 43092
rect 33908 43036 33918 43092
rect 9996 42980 10052 43036
rect 9202 42924 9212 42980
rect 9268 42924 11676 42980
rect 11732 42924 13580 42980
rect 13636 42924 13646 42980
rect 5058 42812 5068 42868
rect 5124 42812 6076 42868
rect 6132 42812 6142 42868
rect 6290 42812 6300 42868
rect 6356 42812 7420 42868
rect 7476 42812 7486 42868
rect 8530 42812 8540 42868
rect 8596 42812 8876 42868
rect 8932 42812 8942 42868
rect 9650 42812 9660 42868
rect 9716 42812 9996 42868
rect 10052 42812 10062 42868
rect 22530 42812 22540 42868
rect 22596 42812 23324 42868
rect 23380 42812 23390 42868
rect 23538 42812 23548 42868
rect 23604 42812 23884 42868
rect 23940 42812 25004 42868
rect 25060 42812 25070 42868
rect 26114 42812 26124 42868
rect 26180 42812 26572 42868
rect 26628 42812 28140 42868
rect 28196 42812 29596 42868
rect 29652 42812 30268 42868
rect 30324 42812 30334 42868
rect 33618 42812 33628 42868
rect 33684 42812 34300 42868
rect 34356 42812 34972 42868
rect 35028 42812 35038 42868
rect 3154 42700 3164 42756
rect 3220 42700 19292 42756
rect 19348 42700 19358 42756
rect 20738 42700 20748 42756
rect 20804 42700 22316 42756
rect 22372 42700 22382 42756
rect 27010 42700 27020 42756
rect 27076 42700 27580 42756
rect 27636 42700 30492 42756
rect 30548 42700 33740 42756
rect 33796 42700 33806 42756
rect 33954 42700 33964 42756
rect 34020 42700 34412 42756
rect 34468 42700 34478 42756
rect 36306 42700 36316 42756
rect 36372 42700 36988 42756
rect 37044 42700 37660 42756
rect 37716 42700 37726 42756
rect 0 42644 800 42672
rect 0 42588 3500 42644
rect 3556 42588 3566 42644
rect 6738 42588 6748 42644
rect 6804 42588 7196 42644
rect 7252 42588 8204 42644
rect 8260 42588 8270 42644
rect 12786 42588 12796 42644
rect 12852 42588 13580 42644
rect 13636 42588 13804 42644
rect 13860 42588 13870 42644
rect 14130 42588 14140 42644
rect 14196 42588 19124 42644
rect 23650 42588 23660 42644
rect 23716 42588 24556 42644
rect 24612 42588 24622 42644
rect 33618 42588 33628 42644
rect 33684 42588 35084 42644
rect 35140 42588 35150 42644
rect 36418 42588 36428 42644
rect 36484 42588 37100 42644
rect 37156 42588 37166 42644
rect 0 42560 800 42588
rect 8642 42476 8652 42532
rect 8708 42476 9660 42532
rect 9716 42476 9726 42532
rect 13998 42308 14008 42364
rect 14064 42308 14112 42364
rect 14168 42308 14216 42364
rect 14272 42308 14320 42364
rect 14376 42308 14424 42364
rect 14480 42308 14528 42364
rect 14584 42308 14632 42364
rect 14688 42308 14736 42364
rect 14792 42308 14840 42364
rect 14896 42308 14944 42364
rect 15000 42308 15048 42364
rect 15104 42308 15152 42364
rect 15208 42308 15218 42364
rect 19068 42196 19124 42588
rect 20178 42476 20188 42532
rect 20244 42476 20972 42532
rect 21028 42476 21038 42532
rect 30146 42476 30156 42532
rect 30212 42476 31276 42532
rect 31332 42476 31724 42532
rect 31780 42476 31790 42532
rect 33506 42476 33516 42532
rect 33572 42476 35364 42532
rect 36082 42476 36092 42532
rect 36148 42476 37660 42532
rect 37716 42476 37726 42532
rect 37874 42476 37884 42532
rect 37940 42476 38220 42532
rect 38276 42476 38286 42532
rect 35308 42420 35364 42476
rect 35308 42364 37772 42420
rect 37828 42364 37838 42420
rect 33998 42308 34008 42364
rect 34064 42308 34112 42364
rect 34168 42308 34216 42364
rect 34272 42308 34320 42364
rect 34376 42308 34424 42364
rect 34480 42308 34528 42364
rect 34584 42308 34632 42364
rect 34688 42308 34736 42364
rect 34792 42308 34840 42364
rect 34896 42308 34944 42364
rect 35000 42308 35048 42364
rect 35104 42308 35152 42364
rect 35208 42308 35218 42364
rect 9202 42140 9212 42196
rect 9268 42140 10108 42196
rect 10164 42140 10174 42196
rect 17826 42140 17836 42196
rect 17892 42140 18060 42196
rect 18116 42140 18126 42196
rect 19058 42140 19068 42196
rect 19124 42140 19964 42196
rect 20020 42140 20748 42196
rect 20804 42140 20814 42196
rect 30818 42140 30828 42196
rect 30884 42140 32172 42196
rect 32228 42140 33180 42196
rect 33236 42140 35532 42196
rect 35588 42140 35598 42196
rect 9986 42028 9996 42084
rect 10052 42028 10892 42084
rect 10948 42028 10958 42084
rect 17714 42028 17724 42084
rect 17780 42028 18396 42084
rect 18452 42028 18462 42084
rect 35186 42028 35196 42084
rect 35252 42028 37548 42084
rect 37604 42028 37614 42084
rect 18396 41972 18452 42028
rect 8418 41916 8428 41972
rect 8484 41916 9212 41972
rect 9268 41916 11564 41972
rect 11620 41916 11630 41972
rect 18396 41916 18732 41972
rect 18788 41916 18798 41972
rect 22530 41916 22540 41972
rect 22596 41916 24444 41972
rect 24500 41916 25340 41972
rect 25396 41916 25406 41972
rect 26226 41916 26236 41972
rect 26292 41916 27020 41972
rect 27076 41916 27086 41972
rect 29250 41916 29260 41972
rect 29316 41916 29932 41972
rect 29988 41916 29998 41972
rect 30258 41916 30268 41972
rect 30324 41916 31052 41972
rect 31108 41916 31118 41972
rect 33954 41916 33964 41972
rect 34020 41916 35084 41972
rect 35140 41916 35150 41972
rect 35298 41916 35308 41972
rect 35364 41916 36988 41972
rect 37044 41916 37054 41972
rect 37202 41916 37212 41972
rect 37268 41916 37278 41972
rect 37212 41860 37268 41916
rect 8306 41804 8316 41860
rect 8372 41804 9772 41860
rect 9828 41804 10668 41860
rect 10724 41804 10734 41860
rect 35746 41804 35756 41860
rect 35812 41804 37884 41860
rect 37940 41804 37950 41860
rect 25442 41692 25452 41748
rect 25508 41692 27132 41748
rect 27188 41692 27198 41748
rect 31714 41580 31724 41636
rect 31780 41580 33180 41636
rect 33236 41580 33246 41636
rect 33740 41580 33852 41636
rect 33908 41580 33918 41636
rect 0 41524 800 41552
rect 3998 41524 4008 41580
rect 4064 41524 4112 41580
rect 4168 41524 4216 41580
rect 4272 41524 4320 41580
rect 4376 41524 4424 41580
rect 4480 41524 4528 41580
rect 4584 41524 4632 41580
rect 4688 41524 4736 41580
rect 4792 41524 4840 41580
rect 4896 41524 4944 41580
rect 5000 41524 5048 41580
rect 5104 41524 5152 41580
rect 5208 41524 5218 41580
rect 23998 41524 24008 41580
rect 24064 41524 24112 41580
rect 24168 41524 24216 41580
rect 24272 41524 24320 41580
rect 24376 41524 24424 41580
rect 24480 41524 24528 41580
rect 24584 41524 24632 41580
rect 24688 41524 24736 41580
rect 24792 41524 24840 41580
rect 24896 41524 24944 41580
rect 25000 41524 25048 41580
rect 25104 41524 25152 41580
rect 25208 41524 25218 41580
rect 33740 41524 33796 41580
rect 0 41468 2604 41524
rect 2660 41468 2670 41524
rect 33730 41468 33740 41524
rect 33796 41468 33806 41524
rect 0 41440 800 41468
rect 11106 41356 11116 41412
rect 11172 41356 12348 41412
rect 12404 41356 12414 41412
rect 16482 41356 16492 41412
rect 16548 41356 17500 41412
rect 17556 41356 17566 41412
rect 25442 41356 25452 41412
rect 25508 41356 25788 41412
rect 25844 41356 25854 41412
rect 27346 41356 27356 41412
rect 27412 41356 29764 41412
rect 30818 41356 30828 41412
rect 30884 41356 32172 41412
rect 32228 41356 32238 41412
rect 33282 41356 33292 41412
rect 33348 41356 37100 41412
rect 37156 41356 37166 41412
rect 29708 41300 29764 41356
rect 10210 41244 10220 41300
rect 10276 41244 21532 41300
rect 21588 41244 22652 41300
rect 22708 41244 22718 41300
rect 24658 41244 24668 41300
rect 24724 41244 26012 41300
rect 26068 41244 27804 41300
rect 27860 41244 27870 41300
rect 29698 41244 29708 41300
rect 29764 41244 30268 41300
rect 30324 41244 30334 41300
rect 30594 41244 30604 41300
rect 30660 41244 32396 41300
rect 32452 41244 37660 41300
rect 37716 41244 37726 41300
rect 7522 41132 7532 41188
rect 7588 41132 7980 41188
rect 8036 41132 8046 41188
rect 10658 41132 10668 41188
rect 10724 41132 12012 41188
rect 12068 41132 12078 41188
rect 20738 41132 20748 41188
rect 20804 41132 21868 41188
rect 21924 41132 21934 41188
rect 22082 41132 22092 41188
rect 22148 41132 24780 41188
rect 24836 41132 25452 41188
rect 25508 41132 25518 41188
rect 25778 41132 25788 41188
rect 25844 41132 26908 41188
rect 26964 41132 28476 41188
rect 28532 41132 28542 41188
rect 30706 41132 30716 41188
rect 30772 41132 32060 41188
rect 32116 41132 32126 41188
rect 32274 41132 32284 41188
rect 32340 41132 35308 41188
rect 35364 41132 35374 41188
rect 8194 41020 8204 41076
rect 8260 41020 10556 41076
rect 10612 41020 10622 41076
rect 24546 41020 24556 41076
rect 24612 41020 25228 41076
rect 25284 41020 25294 41076
rect 33842 41020 33852 41076
rect 33908 41020 34748 41076
rect 34804 41020 37212 41076
rect 37268 41020 37278 41076
rect 5282 40908 5292 40964
rect 5348 40908 7980 40964
rect 8036 40908 8046 40964
rect 23874 40908 23884 40964
rect 23940 40908 24444 40964
rect 24500 40908 27916 40964
rect 27972 40908 29148 40964
rect 29204 40908 29214 40964
rect 33170 40908 33180 40964
rect 33236 40908 35868 40964
rect 35924 40908 37996 40964
rect 38052 40908 38062 40964
rect 13998 40740 14008 40796
rect 14064 40740 14112 40796
rect 14168 40740 14216 40796
rect 14272 40740 14320 40796
rect 14376 40740 14424 40796
rect 14480 40740 14528 40796
rect 14584 40740 14632 40796
rect 14688 40740 14736 40796
rect 14792 40740 14840 40796
rect 14896 40740 14944 40796
rect 15000 40740 15048 40796
rect 15104 40740 15152 40796
rect 15208 40740 15218 40796
rect 33998 40740 34008 40796
rect 34064 40740 34112 40796
rect 34168 40740 34216 40796
rect 34272 40740 34320 40796
rect 34376 40740 34424 40796
rect 34480 40740 34528 40796
rect 34584 40740 34632 40796
rect 34688 40740 34736 40796
rect 34792 40740 34840 40796
rect 34896 40740 34944 40796
rect 35000 40740 35048 40796
rect 35104 40740 35152 40796
rect 35208 40740 35218 40796
rect 4722 40684 4732 40740
rect 4788 40684 5740 40740
rect 5796 40684 7196 40740
rect 7252 40684 7262 40740
rect 23622 40684 23660 40740
rect 23716 40684 23726 40740
rect 29026 40684 29036 40740
rect 29092 40684 29932 40740
rect 29988 40684 30604 40740
rect 30660 40684 30670 40740
rect 6738 40572 6748 40628
rect 6804 40572 7420 40628
rect 7476 40572 7486 40628
rect 7644 40572 7980 40628
rect 8036 40572 8764 40628
rect 8820 40572 8830 40628
rect 9314 40572 9324 40628
rect 9380 40572 11788 40628
rect 11844 40572 11854 40628
rect 13458 40572 13468 40628
rect 13524 40572 13804 40628
rect 13860 40572 14140 40628
rect 14196 40572 14206 40628
rect 15138 40572 15148 40628
rect 15204 40572 17612 40628
rect 17668 40572 17678 40628
rect 21970 40572 21980 40628
rect 22036 40572 22204 40628
rect 22260 40572 23100 40628
rect 23156 40572 23166 40628
rect 25442 40572 25452 40628
rect 25508 40572 26796 40628
rect 7644 40516 7700 40572
rect 3938 40460 3948 40516
rect 4004 40460 5740 40516
rect 5796 40460 5806 40516
rect 6626 40460 6636 40516
rect 6692 40460 7700 40516
rect 7858 40460 7868 40516
rect 7924 40460 8316 40516
rect 8372 40460 9996 40516
rect 10052 40460 10062 40516
rect 0 40404 800 40432
rect 14140 40404 14196 40572
rect 26852 40516 26908 40628
rect 30258 40572 30268 40628
rect 30324 40572 31612 40628
rect 31668 40572 32844 40628
rect 32900 40572 32910 40628
rect 33618 40572 33628 40628
rect 33684 40572 33740 40628
rect 33796 40572 33964 40628
rect 34020 40572 37772 40628
rect 37828 40572 38220 40628
rect 38276 40572 38286 40628
rect 26852 40460 30156 40516
rect 30212 40460 32228 40516
rect 33282 40460 33292 40516
rect 33348 40460 34076 40516
rect 34132 40460 34142 40516
rect 32172 40404 32228 40460
rect 0 40348 2604 40404
rect 2660 40348 2670 40404
rect 14140 40348 14924 40404
rect 14980 40348 15932 40404
rect 15988 40348 21532 40404
rect 21588 40348 25788 40404
rect 25844 40348 25854 40404
rect 27010 40348 27020 40404
rect 27076 40348 27804 40404
rect 27860 40348 29932 40404
rect 29988 40348 30940 40404
rect 30996 40348 31006 40404
rect 32162 40348 32172 40404
rect 32228 40348 33068 40404
rect 33124 40348 35644 40404
rect 35700 40348 35710 40404
rect 0 40320 800 40348
rect 7522 40236 7532 40292
rect 7588 40236 8036 40292
rect 13570 40236 13580 40292
rect 13636 40236 15036 40292
rect 15092 40236 15102 40292
rect 23650 40236 23660 40292
rect 23716 40236 24332 40292
rect 24388 40236 25452 40292
rect 25508 40236 25518 40292
rect 31490 40236 31500 40292
rect 31556 40236 33292 40292
rect 33348 40236 33358 40292
rect 7980 40068 8036 40236
rect 32386 40124 32396 40180
rect 32452 40124 33404 40180
rect 33460 40124 33470 40180
rect 7970 40012 7980 40068
rect 8036 40012 8046 40068
rect 3998 39956 4008 40012
rect 4064 39956 4112 40012
rect 4168 39956 4216 40012
rect 4272 39956 4320 40012
rect 4376 39956 4424 40012
rect 4480 39956 4528 40012
rect 4584 39956 4632 40012
rect 4688 39956 4736 40012
rect 4792 39956 4840 40012
rect 4896 39956 4944 40012
rect 5000 39956 5048 40012
rect 5104 39956 5152 40012
rect 5208 39956 5218 40012
rect 23998 39956 24008 40012
rect 24064 39956 24112 40012
rect 24168 39956 24216 40012
rect 24272 39956 24320 40012
rect 24376 39956 24424 40012
rect 24480 39956 24528 40012
rect 24584 39956 24632 40012
rect 24688 39956 24736 40012
rect 24792 39956 24840 40012
rect 24896 39956 24944 40012
rect 25000 39956 25048 40012
rect 25104 39956 25152 40012
rect 25208 39956 25218 40012
rect 2258 39788 2268 39844
rect 2324 39788 3724 39844
rect 3780 39788 3790 39844
rect 23538 39788 23548 39844
rect 23604 39788 24108 39844
rect 24164 39788 24174 39844
rect 33506 39788 33516 39844
rect 33572 39788 33964 39844
rect 34020 39788 34030 39844
rect 36306 39788 36316 39844
rect 36372 39788 38108 39844
rect 38164 39788 38174 39844
rect 9986 39676 9996 39732
rect 10052 39676 10780 39732
rect 10836 39676 11228 39732
rect 11284 39676 11294 39732
rect 19170 39676 19180 39732
rect 19236 39676 20972 39732
rect 21028 39676 21756 39732
rect 21812 39676 23548 39732
rect 23604 39676 26124 39732
rect 26180 39676 26190 39732
rect 29474 39676 29484 39732
rect 29540 39676 30156 39732
rect 30212 39676 30492 39732
rect 30548 39676 30558 39732
rect 33618 39676 33628 39732
rect 33684 39676 34636 39732
rect 34692 39676 34702 39732
rect 3826 39564 3836 39620
rect 3892 39564 4284 39620
rect 4340 39564 6188 39620
rect 6244 39564 6254 39620
rect 6514 39564 6524 39620
rect 6580 39564 7308 39620
rect 7364 39564 7374 39620
rect 8754 39564 8764 39620
rect 8820 39564 9660 39620
rect 9716 39564 9726 39620
rect 23090 39564 23100 39620
rect 23156 39564 23660 39620
rect 23716 39564 24556 39620
rect 24612 39564 25676 39620
rect 25732 39564 28252 39620
rect 28308 39564 28318 39620
rect 3154 39452 3164 39508
rect 3220 39452 5964 39508
rect 6020 39452 15148 39508
rect 15092 39396 15148 39452
rect 6178 39340 6188 39396
rect 6244 39340 6972 39396
rect 7028 39340 7038 39396
rect 8978 39340 8988 39396
rect 9044 39340 9548 39396
rect 9604 39340 9614 39396
rect 15092 39340 19516 39396
rect 19572 39340 19582 39396
rect 0 39284 800 39312
rect 0 39228 2492 39284
rect 2548 39228 2558 39284
rect 0 39200 800 39228
rect 13998 39172 14008 39228
rect 14064 39172 14112 39228
rect 14168 39172 14216 39228
rect 14272 39172 14320 39228
rect 14376 39172 14424 39228
rect 14480 39172 14528 39228
rect 14584 39172 14632 39228
rect 14688 39172 14736 39228
rect 14792 39172 14840 39228
rect 14896 39172 14944 39228
rect 15000 39172 15048 39228
rect 15104 39172 15152 39228
rect 15208 39172 15218 39228
rect 33998 39172 34008 39228
rect 34064 39172 34112 39228
rect 34168 39172 34216 39228
rect 34272 39172 34320 39228
rect 34376 39172 34424 39228
rect 34480 39172 34528 39228
rect 34584 39172 34632 39228
rect 34688 39172 34736 39228
rect 34792 39172 34840 39228
rect 34896 39172 34944 39228
rect 35000 39172 35048 39228
rect 35104 39172 35152 39228
rect 35208 39172 35218 39228
rect 7522 39116 7532 39172
rect 7588 39116 8652 39172
rect 8708 39116 8718 39172
rect 36418 39116 36428 39172
rect 36484 39116 37100 39172
rect 37156 39116 37166 39172
rect 3154 39004 3164 39060
rect 3220 39004 6076 39060
rect 6132 39004 6524 39060
rect 6580 39004 6590 39060
rect 6962 39004 6972 39060
rect 7028 39004 8092 39060
rect 8148 39004 9436 39060
rect 9492 39004 9502 39060
rect 11218 39004 11228 39060
rect 11284 39004 14924 39060
rect 14980 39004 14990 39060
rect 32274 39004 32284 39060
rect 32340 39004 33740 39060
rect 33796 39004 33852 39060
rect 33908 39004 33918 39060
rect 34290 39004 34300 39060
rect 34356 39004 37212 39060
rect 37268 39004 37278 39060
rect 3266 38892 3276 38948
rect 3332 38892 5404 38948
rect 5460 38892 16156 38948
rect 16212 38892 16716 38948
rect 16772 38892 16782 38948
rect 32386 38892 32396 38948
rect 32452 38892 34188 38948
rect 34244 38892 34254 38948
rect 34962 38892 34972 38948
rect 35028 38892 38108 38948
rect 38164 38892 38174 38948
rect 4610 38780 4620 38836
rect 4676 38780 5740 38836
rect 5796 38780 8316 38836
rect 8372 38780 8382 38836
rect 11330 38780 11340 38836
rect 11396 38780 11564 38836
rect 11620 38780 15484 38836
rect 15540 38780 15550 38836
rect 16818 38780 16828 38836
rect 16884 38780 17388 38836
rect 17444 38780 17454 38836
rect 32610 38780 32620 38836
rect 32676 38780 34748 38836
rect 34804 38780 34814 38836
rect 8316 38668 8988 38724
rect 9044 38668 9054 38724
rect 13346 38668 13356 38724
rect 13412 38668 16492 38724
rect 16548 38668 17948 38724
rect 18004 38668 19852 38724
rect 19908 38668 19918 38724
rect 31826 38668 31836 38724
rect 31892 38668 33516 38724
rect 33572 38668 33582 38724
rect 35186 38668 35196 38724
rect 35252 38668 35868 38724
rect 35924 38668 35934 38724
rect 8316 38612 8372 38668
rect 8082 38556 8092 38612
rect 8148 38556 8372 38612
rect 15250 38556 15260 38612
rect 15316 38556 16380 38612
rect 16436 38556 18620 38612
rect 18676 38556 19068 38612
rect 19124 38556 19134 38612
rect 17574 38444 17612 38500
rect 17668 38444 17678 38500
rect 33506 38444 33516 38500
rect 33572 38444 33852 38500
rect 33908 38444 33918 38500
rect 3998 38388 4008 38444
rect 4064 38388 4112 38444
rect 4168 38388 4216 38444
rect 4272 38388 4320 38444
rect 4376 38388 4424 38444
rect 4480 38388 4528 38444
rect 4584 38388 4632 38444
rect 4688 38388 4736 38444
rect 4792 38388 4840 38444
rect 4896 38388 4944 38444
rect 5000 38388 5048 38444
rect 5104 38388 5152 38444
rect 5208 38388 5218 38444
rect 23998 38388 24008 38444
rect 24064 38388 24112 38444
rect 24168 38388 24216 38444
rect 24272 38388 24320 38444
rect 24376 38388 24424 38444
rect 24480 38388 24528 38444
rect 24584 38388 24632 38444
rect 24688 38388 24736 38444
rect 24792 38388 24840 38444
rect 24896 38388 24944 38444
rect 25000 38388 25048 38444
rect 25104 38388 25152 38444
rect 25208 38388 25218 38444
rect 37314 38332 37324 38388
rect 37380 38332 37884 38388
rect 37940 38332 37950 38388
rect 8642 38220 8652 38276
rect 8708 38220 9884 38276
rect 9940 38220 9950 38276
rect 18274 38220 18284 38276
rect 18340 38220 18732 38276
rect 18788 38220 18798 38276
rect 32050 38220 32060 38276
rect 32116 38220 35644 38276
rect 35700 38220 35710 38276
rect 0 38164 800 38192
rect 0 38108 2492 38164
rect 2548 38108 2558 38164
rect 24882 38108 24892 38164
rect 24948 38108 25564 38164
rect 25620 38108 25630 38164
rect 31938 38108 31948 38164
rect 32004 38108 33740 38164
rect 33796 38108 34076 38164
rect 34132 38108 34142 38164
rect 36082 38108 36092 38164
rect 36148 38108 37660 38164
rect 37716 38108 37996 38164
rect 38052 38108 38062 38164
rect 0 38080 800 38108
rect 19618 37996 19628 38052
rect 19684 37996 22092 38052
rect 22148 37996 22158 38052
rect 31714 37996 31724 38052
rect 31780 37996 32620 38052
rect 32676 37996 32686 38052
rect 7298 37772 7308 37828
rect 7364 37772 8876 37828
rect 8932 37772 8942 37828
rect 16034 37772 16044 37828
rect 16100 37772 17948 37828
rect 18004 37772 18956 37828
rect 19012 37772 19022 37828
rect 27570 37772 27580 37828
rect 27636 37772 30492 37828
rect 30548 37772 31052 37828
rect 31108 37772 31118 37828
rect 15372 37660 22204 37716
rect 22260 37660 22270 37716
rect 33394 37660 33404 37716
rect 33460 37660 33852 37716
rect 33908 37660 33918 37716
rect 13998 37604 14008 37660
rect 14064 37604 14112 37660
rect 14168 37604 14216 37660
rect 14272 37604 14320 37660
rect 14376 37604 14424 37660
rect 14480 37604 14528 37660
rect 14584 37604 14632 37660
rect 14688 37604 14736 37660
rect 14792 37604 14840 37660
rect 14896 37604 14944 37660
rect 15000 37604 15048 37660
rect 15104 37604 15152 37660
rect 15208 37604 15218 37660
rect 15372 37492 15428 37660
rect 33998 37604 34008 37660
rect 34064 37604 34112 37660
rect 34168 37604 34216 37660
rect 34272 37604 34320 37660
rect 34376 37604 34424 37660
rect 34480 37604 34528 37660
rect 34584 37604 34632 37660
rect 34688 37604 34736 37660
rect 34792 37604 34840 37660
rect 34896 37604 34944 37660
rect 35000 37604 35048 37660
rect 35104 37604 35152 37660
rect 35208 37604 35218 37660
rect 26450 37548 26460 37604
rect 26516 37548 28028 37604
rect 28084 37548 31948 37604
rect 32004 37548 32014 37604
rect 14802 37436 14812 37492
rect 14868 37436 15428 37492
rect 15698 37436 15708 37492
rect 15764 37436 17836 37492
rect 17892 37436 17902 37492
rect 21858 37436 21868 37492
rect 21924 37436 24668 37492
rect 24724 37436 25900 37492
rect 25956 37436 26684 37492
rect 26740 37436 26750 37492
rect 28242 37436 28252 37492
rect 28308 37436 30604 37492
rect 30660 37436 31164 37492
rect 31220 37436 31230 37492
rect 34514 37436 34524 37492
rect 34580 37436 37324 37492
rect 37380 37436 37390 37492
rect 3154 37324 3164 37380
rect 3220 37324 7420 37380
rect 7476 37324 7486 37380
rect 12562 37324 12572 37380
rect 12628 37324 14028 37380
rect 14084 37324 14094 37380
rect 16818 37324 16828 37380
rect 16884 37324 18732 37380
rect 18788 37324 18798 37380
rect 21074 37324 21084 37380
rect 21140 37324 21532 37380
rect 21588 37324 22428 37380
rect 22484 37324 22494 37380
rect 23650 37324 23660 37380
rect 23716 37324 23772 37380
rect 23828 37324 23838 37380
rect 12226 37212 12236 37268
rect 12292 37212 13244 37268
rect 13300 37212 13310 37268
rect 14242 37212 14252 37268
rect 14308 37212 16492 37268
rect 16548 37212 18060 37268
rect 18116 37212 19628 37268
rect 19684 37212 19694 37268
rect 26460 37156 26516 37436
rect 26982 37324 27020 37380
rect 27076 37324 27580 37380
rect 27636 37324 27646 37380
rect 33506 37324 33516 37380
rect 33572 37324 36204 37380
rect 36260 37324 37436 37380
rect 37492 37324 37996 37380
rect 38052 37324 38062 37380
rect 26674 37212 26684 37268
rect 26740 37212 26908 37268
rect 26964 37212 27916 37268
rect 27972 37212 28252 37268
rect 28308 37212 28318 37268
rect 30482 37212 30492 37268
rect 30548 37212 31724 37268
rect 31780 37212 31790 37268
rect 32498 37212 32508 37268
rect 32564 37212 35196 37268
rect 35252 37212 35262 37268
rect 10434 37100 10444 37156
rect 10500 37100 11452 37156
rect 11508 37100 12796 37156
rect 12852 37100 12862 37156
rect 16818 37100 16828 37156
rect 16884 37100 17500 37156
rect 17556 37100 17566 37156
rect 26460 37100 28028 37156
rect 28084 37100 28094 37156
rect 31154 37100 31164 37156
rect 31220 37100 33628 37156
rect 33684 37100 33694 37156
rect 36306 37100 36316 37156
rect 36372 37100 36988 37156
rect 37044 37100 37054 37156
rect 0 37044 800 37072
rect 0 36988 2492 37044
rect 2548 36988 2558 37044
rect 26450 36988 26460 37044
rect 26516 36988 27356 37044
rect 27412 36988 27422 37044
rect 27794 36988 27804 37044
rect 27860 36988 29484 37044
rect 29540 36988 29820 37044
rect 29876 36988 29886 37044
rect 0 36960 800 36988
rect 13682 36876 13692 36932
rect 13748 36876 15036 36932
rect 15092 36876 15102 36932
rect 32386 36876 32396 36932
rect 32452 36876 33068 36932
rect 33124 36876 33134 36932
rect 33730 36876 33740 36932
rect 33796 36876 34188 36932
rect 34244 36876 34254 36932
rect 3998 36820 4008 36876
rect 4064 36820 4112 36876
rect 4168 36820 4216 36876
rect 4272 36820 4320 36876
rect 4376 36820 4424 36876
rect 4480 36820 4528 36876
rect 4584 36820 4632 36876
rect 4688 36820 4736 36876
rect 4792 36820 4840 36876
rect 4896 36820 4944 36876
rect 5000 36820 5048 36876
rect 5104 36820 5152 36876
rect 5208 36820 5218 36876
rect 23998 36820 24008 36876
rect 24064 36820 24112 36876
rect 24168 36820 24216 36876
rect 24272 36820 24320 36876
rect 24376 36820 24424 36876
rect 24480 36820 24528 36876
rect 24584 36820 24632 36876
rect 24688 36820 24736 36876
rect 24792 36820 24840 36876
rect 24896 36820 24944 36876
rect 25000 36820 25048 36876
rect 25104 36820 25152 36876
rect 25208 36820 25218 36876
rect 27682 36652 27692 36708
rect 27748 36652 29036 36708
rect 29092 36652 29102 36708
rect 6962 36540 6972 36596
rect 7028 36540 7532 36596
rect 7588 36540 7598 36596
rect 8418 36540 8428 36596
rect 8484 36540 10892 36596
rect 10948 36540 10958 36596
rect 15092 36540 16044 36596
rect 16100 36540 16110 36596
rect 32162 36540 32172 36596
rect 32228 36540 33292 36596
rect 33348 36540 33358 36596
rect 7074 36428 7084 36484
rect 7140 36428 8316 36484
rect 8372 36428 8382 36484
rect 8978 36428 8988 36484
rect 9044 36428 10332 36484
rect 10388 36428 10398 36484
rect 12562 36428 12572 36484
rect 12628 36428 13580 36484
rect 13636 36428 13646 36484
rect 15092 36372 15148 36540
rect 26852 36428 27020 36484
rect 27076 36428 27692 36484
rect 27748 36428 27758 36484
rect 26852 36372 26908 36428
rect 5170 36316 5180 36372
rect 5236 36316 5852 36372
rect 5908 36316 5918 36372
rect 7858 36316 7868 36372
rect 7924 36316 8764 36372
rect 8820 36316 9548 36372
rect 9604 36316 9614 36372
rect 11330 36316 11340 36372
rect 11396 36316 12124 36372
rect 12180 36316 14812 36372
rect 14868 36316 15148 36372
rect 23426 36316 23436 36372
rect 23492 36316 26908 36372
rect 31714 36316 31724 36372
rect 31780 36316 37324 36372
rect 37380 36316 37390 36372
rect 4050 36204 4060 36260
rect 4116 36204 4956 36260
rect 5012 36204 5022 36260
rect 6178 36204 6188 36260
rect 6244 36204 7532 36260
rect 7588 36204 7598 36260
rect 12898 36204 12908 36260
rect 12964 36204 13692 36260
rect 13748 36204 13758 36260
rect 18834 36204 18844 36260
rect 18900 36204 20188 36260
rect 20244 36204 20254 36260
rect 23062 36204 23100 36260
rect 23156 36204 23166 36260
rect 33068 36204 34188 36260
rect 34244 36204 34254 36260
rect 36418 36204 36428 36260
rect 36484 36204 38108 36260
rect 38164 36204 38174 36260
rect 33068 36148 33124 36204
rect 31714 36092 31724 36148
rect 31780 36092 32172 36148
rect 32228 36092 33068 36148
rect 33124 36092 33134 36148
rect 36978 36092 36988 36148
rect 37044 36092 37054 36148
rect 13998 36036 14008 36092
rect 14064 36036 14112 36092
rect 14168 36036 14216 36092
rect 14272 36036 14320 36092
rect 14376 36036 14424 36092
rect 14480 36036 14528 36092
rect 14584 36036 14632 36092
rect 14688 36036 14736 36092
rect 14792 36036 14840 36092
rect 14896 36036 14944 36092
rect 15000 36036 15048 36092
rect 15104 36036 15152 36092
rect 15208 36036 15218 36092
rect 33998 36036 34008 36092
rect 34064 36036 34112 36092
rect 34168 36036 34216 36092
rect 34272 36036 34320 36092
rect 34376 36036 34424 36092
rect 34480 36036 34528 36092
rect 34584 36036 34632 36092
rect 34688 36036 34736 36092
rect 34792 36036 34840 36092
rect 34896 36036 34944 36092
rect 35000 36036 35048 36092
rect 35104 36036 35152 36092
rect 35208 36036 35218 36092
rect 4834 35980 4844 36036
rect 4900 35980 7084 36036
rect 7140 35980 7150 36036
rect 0 35924 800 35952
rect 36988 35924 37044 36092
rect 0 35868 2492 35924
rect 2548 35868 2558 35924
rect 4946 35868 4956 35924
rect 5012 35868 5292 35924
rect 5348 35868 6300 35924
rect 6356 35868 9100 35924
rect 9156 35868 9166 35924
rect 20290 35868 20300 35924
rect 20356 35868 22876 35924
rect 22932 35868 23548 35924
rect 23604 35868 23614 35924
rect 31836 35868 32396 35924
rect 32452 35868 32462 35924
rect 33730 35868 33740 35924
rect 33796 35868 34300 35924
rect 34356 35868 34366 35924
rect 35186 35868 35196 35924
rect 35252 35868 37044 35924
rect 0 35840 800 35868
rect 31836 35812 31892 35868
rect 8642 35756 8652 35812
rect 8708 35756 9660 35812
rect 9716 35756 9726 35812
rect 13570 35756 13580 35812
rect 13636 35756 14924 35812
rect 14980 35756 14990 35812
rect 16370 35756 16380 35812
rect 16436 35756 25340 35812
rect 25396 35756 25900 35812
rect 25956 35756 27356 35812
rect 27412 35756 27804 35812
rect 27860 35756 27870 35812
rect 28466 35756 28476 35812
rect 28532 35756 31836 35812
rect 31892 35756 31902 35812
rect 33058 35756 33068 35812
rect 33124 35756 34636 35812
rect 34692 35756 34702 35812
rect 8418 35644 8428 35700
rect 8484 35644 9716 35700
rect 12786 35644 12796 35700
rect 12852 35644 14028 35700
rect 14084 35644 14094 35700
rect 14578 35644 14588 35700
rect 14644 35644 15148 35700
rect 15204 35644 15214 35700
rect 21522 35644 21532 35700
rect 21588 35644 23996 35700
rect 24052 35644 24062 35700
rect 31378 35644 31388 35700
rect 31444 35644 33628 35700
rect 33684 35644 35420 35700
rect 35476 35644 35486 35700
rect 36306 35644 36316 35700
rect 36372 35644 37212 35700
rect 37268 35644 37278 35700
rect 9660 35588 9716 35644
rect 7410 35532 7420 35588
rect 7476 35532 8652 35588
rect 8708 35532 8718 35588
rect 9660 35532 15148 35588
rect 18610 35532 18620 35588
rect 18676 35532 19404 35588
rect 19460 35532 23436 35588
rect 23492 35532 24444 35588
rect 24500 35532 24510 35588
rect 33730 35532 33740 35588
rect 33796 35532 36204 35588
rect 36260 35532 36540 35588
rect 36596 35532 38108 35588
rect 38164 35532 38174 35588
rect 3154 35420 3164 35476
rect 3220 35420 5404 35476
rect 5460 35420 5470 35476
rect 9538 35420 9548 35476
rect 9604 35420 10332 35476
rect 10388 35420 10892 35476
rect 10948 35420 12460 35476
rect 12516 35420 12526 35476
rect 15092 35364 15148 35532
rect 23538 35420 23548 35476
rect 23604 35420 25340 35476
rect 25396 35420 25406 35476
rect 26674 35420 26684 35476
rect 26740 35420 27244 35476
rect 27300 35420 27310 35476
rect 31154 35420 31164 35476
rect 31220 35420 31724 35476
rect 31780 35420 31948 35476
rect 32004 35420 32014 35476
rect 32162 35420 32172 35476
rect 32228 35420 32844 35476
rect 32900 35420 34300 35476
rect 34356 35420 34366 35476
rect 8754 35308 8764 35364
rect 8820 35308 9996 35364
rect 10052 35308 10062 35364
rect 10220 35308 12012 35364
rect 12068 35308 12078 35364
rect 15092 35308 17052 35364
rect 17108 35308 17118 35364
rect 30818 35308 30828 35364
rect 30884 35308 31612 35364
rect 31668 35308 31678 35364
rect 32498 35308 32508 35364
rect 32564 35308 36988 35364
rect 37044 35308 37054 35364
rect 3998 35252 4008 35308
rect 4064 35252 4112 35308
rect 4168 35252 4216 35308
rect 4272 35252 4320 35308
rect 4376 35252 4424 35308
rect 4480 35252 4528 35308
rect 4584 35252 4632 35308
rect 4688 35252 4736 35308
rect 4792 35252 4840 35308
rect 4896 35252 4944 35308
rect 5000 35252 5048 35308
rect 5104 35252 5152 35308
rect 5208 35252 5218 35308
rect 8764 35252 8820 35308
rect 10220 35252 10276 35308
rect 23998 35252 24008 35308
rect 24064 35252 24112 35308
rect 24168 35252 24216 35308
rect 24272 35252 24320 35308
rect 24376 35252 24424 35308
rect 24480 35252 24528 35308
rect 24584 35252 24632 35308
rect 24688 35252 24736 35308
rect 24792 35252 24840 35308
rect 24896 35252 24944 35308
rect 25000 35252 25048 35308
rect 25104 35252 25152 35308
rect 25208 35252 25218 35308
rect 6626 35196 6636 35252
rect 6692 35196 8820 35252
rect 9426 35196 9436 35252
rect 9492 35196 10276 35252
rect 14690 35196 14700 35252
rect 14756 35196 15036 35252
rect 15092 35196 17500 35252
rect 17556 35196 18620 35252
rect 18676 35196 18686 35252
rect 19516 35196 23660 35252
rect 23716 35196 23726 35252
rect 37762 35196 37772 35252
rect 37828 35196 38108 35252
rect 38164 35196 38174 35252
rect 19516 35140 19572 35196
rect 3042 35084 3052 35140
rect 3108 35084 4732 35140
rect 4788 35084 6412 35140
rect 6468 35084 6478 35140
rect 9874 35084 9884 35140
rect 9940 35084 10892 35140
rect 10948 35084 10958 35140
rect 13794 35084 13804 35140
rect 13860 35084 14588 35140
rect 14644 35084 14654 35140
rect 15092 35084 19572 35140
rect 19842 35084 19852 35140
rect 19908 35084 20636 35140
rect 20692 35084 20702 35140
rect 37314 35084 37324 35140
rect 37380 35084 37884 35140
rect 37940 35084 37950 35140
rect 4610 34972 4620 35028
rect 4676 34972 5292 35028
rect 5348 34972 5358 35028
rect 7186 34972 7196 35028
rect 7252 34972 7308 35028
rect 7364 34972 7374 35028
rect 13654 34972 13692 35028
rect 13748 34972 13758 35028
rect 15092 34916 15148 35084
rect 33506 34972 33516 35028
rect 33572 34972 35868 35028
rect 35924 34972 35934 35028
rect 4162 34860 4172 34916
rect 4228 34860 5628 34916
rect 5684 34860 5694 34916
rect 7298 34860 7308 34916
rect 7364 34860 7374 34916
rect 9762 34860 9772 34916
rect 9828 34860 11116 34916
rect 11172 34860 11182 34916
rect 11778 34860 11788 34916
rect 11844 34860 15148 34916
rect 23090 34860 23100 34916
rect 23156 34860 26012 34916
rect 26068 34860 26908 34916
rect 26964 34860 28252 34916
rect 28308 34860 28318 34916
rect 33618 34860 33628 34916
rect 33684 34860 34524 34916
rect 34580 34860 34590 34916
rect 36418 34860 36428 34916
rect 36484 34860 36876 34916
rect 36932 34860 37548 34916
rect 37604 34860 37996 34916
rect 38052 34860 38062 34916
rect 0 34804 800 34832
rect 7308 34804 7364 34860
rect 0 34748 2604 34804
rect 2660 34748 2670 34804
rect 4946 34748 4956 34804
rect 5012 34748 5292 34804
rect 5348 34748 6076 34804
rect 6132 34748 6142 34804
rect 7074 34748 7084 34804
rect 7140 34748 7364 34804
rect 8978 34748 8988 34804
rect 9044 34748 10556 34804
rect 10612 34748 10622 34804
rect 11218 34748 11228 34804
rect 11284 34748 11676 34804
rect 11732 34748 12068 34804
rect 12450 34748 12460 34804
rect 12516 34748 16772 34804
rect 16930 34748 16940 34804
rect 16996 34748 17612 34804
rect 17668 34748 17678 34804
rect 19058 34748 19068 34804
rect 19124 34748 19516 34804
rect 19572 34748 21644 34804
rect 21700 34748 21710 34804
rect 23202 34748 23212 34804
rect 23268 34748 25788 34804
rect 25844 34748 27804 34804
rect 27860 34748 27870 34804
rect 32386 34748 32396 34804
rect 32452 34748 35084 34804
rect 35140 34748 37212 34804
rect 37268 34748 37278 34804
rect 0 34720 800 34748
rect 12012 34692 12068 34748
rect 16716 34692 16772 34748
rect 2258 34636 2268 34692
rect 2324 34636 3836 34692
rect 3892 34636 3902 34692
rect 5730 34636 5740 34692
rect 5796 34636 6188 34692
rect 6244 34636 6254 34692
rect 6402 34636 6412 34692
rect 6468 34636 7644 34692
rect 7700 34636 7710 34692
rect 12012 34636 16212 34692
rect 16706 34636 16716 34692
rect 16772 34636 17836 34692
rect 17892 34636 27132 34692
rect 27188 34636 27198 34692
rect 33058 34636 33068 34692
rect 33124 34636 33852 34692
rect 33908 34636 33918 34692
rect 34850 34636 34860 34692
rect 34916 34636 37548 34692
rect 37604 34636 37614 34692
rect 16156 34580 16212 34636
rect 13010 34524 13020 34580
rect 13076 34524 13580 34580
rect 13636 34524 13804 34580
rect 13860 34524 13870 34580
rect 16156 34524 25452 34580
rect 25508 34524 25518 34580
rect 13998 34468 14008 34524
rect 14064 34468 14112 34524
rect 14168 34468 14216 34524
rect 14272 34468 14320 34524
rect 14376 34468 14424 34524
rect 14480 34468 14528 34524
rect 14584 34468 14632 34524
rect 14688 34468 14736 34524
rect 14792 34468 14840 34524
rect 14896 34468 14944 34524
rect 15000 34468 15048 34524
rect 15104 34468 15152 34524
rect 15208 34468 15218 34524
rect 6188 34412 6524 34468
rect 6580 34412 6590 34468
rect 7298 34412 7308 34468
rect 7364 34412 7644 34468
rect 7700 34412 7710 34468
rect 6188 34356 6244 34412
rect 33852 34356 33908 34636
rect 35858 34524 35868 34580
rect 35924 34524 36988 34580
rect 37044 34524 37054 34580
rect 33998 34468 34008 34524
rect 34064 34468 34112 34524
rect 34168 34468 34216 34524
rect 34272 34468 34320 34524
rect 34376 34468 34424 34524
rect 34480 34468 34528 34524
rect 34584 34468 34632 34524
rect 34688 34468 34736 34524
rect 34792 34468 34840 34524
rect 34896 34468 34944 34524
rect 35000 34468 35048 34524
rect 35104 34468 35152 34524
rect 35208 34468 35218 34524
rect 6178 34300 6188 34356
rect 6244 34300 6254 34356
rect 8418 34300 8428 34356
rect 8484 34300 9884 34356
rect 9940 34300 9950 34356
rect 10658 34300 10668 34356
rect 10724 34300 12124 34356
rect 12180 34300 12460 34356
rect 12516 34300 12526 34356
rect 15810 34300 15820 34356
rect 15876 34300 16716 34356
rect 16772 34300 16782 34356
rect 17826 34300 17836 34356
rect 17892 34300 18172 34356
rect 18228 34300 18238 34356
rect 28354 34300 28364 34356
rect 28420 34300 29708 34356
rect 29764 34300 30156 34356
rect 30212 34300 30222 34356
rect 33852 34300 37436 34356
rect 37492 34300 37772 34356
rect 37828 34300 37838 34356
rect 3266 34188 3276 34244
rect 3332 34020 3388 34244
rect 6514 34188 6524 34244
rect 6580 34188 6972 34244
rect 7028 34188 7038 34244
rect 7634 34188 7644 34244
rect 7700 34188 8204 34244
rect 8260 34188 8270 34244
rect 16492 34132 16548 34300
rect 32498 34188 32508 34244
rect 32564 34188 33628 34244
rect 33684 34188 34412 34244
rect 34468 34188 34478 34244
rect 6850 34076 6860 34132
rect 6916 34076 7196 34132
rect 7252 34076 7262 34132
rect 7522 34076 7532 34132
rect 7588 34076 9548 34132
rect 9604 34076 9614 34132
rect 16482 34076 16492 34132
rect 16548 34076 16558 34132
rect 3332 33964 5516 34020
rect 5572 33964 6524 34020
rect 6580 33964 6590 34020
rect 7074 33964 7084 34020
rect 7140 33964 7868 34020
rect 7924 33964 7934 34020
rect 10770 33964 10780 34020
rect 10836 33964 11676 34020
rect 11732 33964 11742 34020
rect 20066 33964 20076 34020
rect 20132 33964 21756 34020
rect 21812 33964 21822 34020
rect 34178 33964 34188 34020
rect 34244 33964 37884 34020
rect 37940 33964 37950 34020
rect 8642 33852 8652 33908
rect 8708 33852 12236 33908
rect 12292 33852 12908 33908
rect 12964 33852 13468 33908
rect 13524 33852 13534 33908
rect 16370 33852 16380 33908
rect 16436 33852 17164 33908
rect 17220 33852 17230 33908
rect 33506 33740 33516 33796
rect 33572 33740 35084 33796
rect 35140 33740 36988 33796
rect 37044 33740 37054 33796
rect 0 33684 800 33712
rect 3998 33684 4008 33740
rect 4064 33684 4112 33740
rect 4168 33684 4216 33740
rect 4272 33684 4320 33740
rect 4376 33684 4424 33740
rect 4480 33684 4528 33740
rect 4584 33684 4632 33740
rect 4688 33684 4736 33740
rect 4792 33684 4840 33740
rect 4896 33684 4944 33740
rect 5000 33684 5048 33740
rect 5104 33684 5152 33740
rect 5208 33684 5218 33740
rect 23998 33684 24008 33740
rect 24064 33684 24112 33740
rect 24168 33684 24216 33740
rect 24272 33684 24320 33740
rect 24376 33684 24424 33740
rect 24480 33684 24528 33740
rect 24584 33684 24632 33740
rect 24688 33684 24736 33740
rect 24792 33684 24840 33740
rect 24896 33684 24944 33740
rect 25000 33684 25048 33740
rect 25104 33684 25152 33740
rect 25208 33684 25218 33740
rect 0 33628 3500 33684
rect 3556 33628 3566 33684
rect 18050 33628 18060 33684
rect 18116 33628 18956 33684
rect 19012 33628 21196 33684
rect 21252 33628 21262 33684
rect 23202 33628 23212 33684
rect 23268 33628 23940 33684
rect 28242 33628 28252 33684
rect 28308 33628 30268 33684
rect 30324 33628 30334 33684
rect 33282 33628 33292 33684
rect 33348 33628 34076 33684
rect 34132 33628 37156 33684
rect 0 33600 800 33628
rect 23884 33572 23940 33628
rect 37100 33572 37156 33628
rect 5254 33516 5292 33572
rect 5348 33516 5358 33572
rect 21298 33516 21308 33572
rect 21364 33516 22204 33572
rect 22260 33516 23436 33572
rect 23492 33516 23502 33572
rect 23884 33516 23996 33572
rect 24052 33516 24062 33572
rect 31378 33516 31388 33572
rect 31444 33516 31948 33572
rect 32004 33516 32956 33572
rect 33012 33516 33022 33572
rect 33170 33516 33180 33572
rect 33236 33516 33964 33572
rect 34020 33516 35420 33572
rect 35476 33516 36876 33572
rect 36932 33516 36942 33572
rect 37100 33516 37212 33572
rect 37268 33516 37278 33572
rect 32956 33460 33012 33516
rect 2482 33404 2492 33460
rect 2548 33404 3388 33460
rect 5058 33404 5068 33460
rect 5124 33404 6748 33460
rect 6804 33404 6814 33460
rect 12002 33404 12012 33460
rect 12068 33404 15372 33460
rect 15428 33404 15438 33460
rect 19282 33404 19292 33460
rect 19348 33404 22540 33460
rect 22596 33404 23884 33460
rect 23940 33404 23950 33460
rect 25442 33404 25452 33460
rect 25508 33404 26236 33460
rect 26292 33404 27020 33460
rect 27076 33404 27086 33460
rect 32956 33404 35084 33460
rect 35140 33404 35532 33460
rect 35588 33404 37100 33460
rect 37156 33404 37166 33460
rect 3332 33348 3388 33404
rect 3332 33292 5180 33348
rect 5236 33292 5246 33348
rect 8306 33292 8316 33348
rect 8372 33292 10556 33348
rect 10612 33292 10622 33348
rect 13906 33292 13916 33348
rect 13972 33292 16268 33348
rect 16324 33292 16334 33348
rect 32834 33292 32844 33348
rect 32900 33292 34748 33348
rect 34804 33292 37324 33348
rect 37380 33292 37390 33348
rect 3154 33180 3164 33236
rect 3220 33180 3388 33236
rect 6626 33180 6636 33236
rect 6692 33180 7420 33236
rect 7476 33180 7486 33236
rect 33730 33180 33740 33236
rect 33796 33180 34076 33236
rect 34132 33180 34142 33236
rect 3332 33124 3388 33180
rect 33740 33124 33796 33180
rect 3332 33068 4172 33124
rect 4228 33068 5964 33124
rect 6020 33068 6030 33124
rect 8306 33068 8316 33124
rect 8372 33068 9324 33124
rect 9380 33068 9390 33124
rect 13804 33068 14476 33124
rect 14532 33068 14542 33124
rect 17042 33068 17052 33124
rect 17108 33068 17612 33124
rect 17668 33068 18508 33124
rect 18564 33068 22428 33124
rect 22484 33068 22494 33124
rect 24658 33068 24668 33124
rect 24724 33068 25228 33124
rect 25284 33068 31836 33124
rect 31892 33068 32172 33124
rect 32228 33068 32732 33124
rect 32788 33068 33404 33124
rect 33460 33068 33796 33124
rect 5170 32956 5180 33012
rect 5236 32956 5740 33012
rect 5796 32956 5806 33012
rect 6850 32956 6860 33012
rect 6916 32956 8036 33012
rect 1810 32732 1820 32788
rect 1876 32732 4732 32788
rect 4788 32732 4798 32788
rect 0 32564 800 32592
rect 7980 32564 8036 32956
rect 13804 32788 13860 33068
rect 15922 32956 15932 33012
rect 15988 32956 16380 33012
rect 16436 32956 27020 33012
rect 27076 32956 30940 33012
rect 30996 32956 31612 33012
rect 31668 32956 31678 33012
rect 33702 32956 33740 33012
rect 33796 32956 33806 33012
rect 13998 32900 14008 32956
rect 14064 32900 14112 32956
rect 14168 32900 14216 32956
rect 14272 32900 14320 32956
rect 14376 32900 14424 32956
rect 14480 32900 14528 32956
rect 14584 32900 14632 32956
rect 14688 32900 14736 32956
rect 14792 32900 14840 32956
rect 14896 32900 14944 32956
rect 15000 32900 15048 32956
rect 15104 32900 15152 32956
rect 15208 32900 15218 32956
rect 33998 32900 34008 32956
rect 34064 32900 34112 32956
rect 34168 32900 34216 32956
rect 34272 32900 34320 32956
rect 34376 32900 34424 32956
rect 34480 32900 34528 32956
rect 34584 32900 34632 32956
rect 34688 32900 34736 32956
rect 34792 32900 34840 32956
rect 34896 32900 34944 32956
rect 35000 32900 35048 32956
rect 35104 32900 35152 32956
rect 35208 32900 35218 32956
rect 23986 32844 23996 32900
rect 24052 32844 25340 32900
rect 25396 32844 25406 32900
rect 13804 32732 14476 32788
rect 14532 32732 14542 32788
rect 15362 32732 15372 32788
rect 15428 32732 15484 32788
rect 15540 32732 16268 32788
rect 16324 32732 16334 32788
rect 23426 32732 23436 32788
rect 23492 32732 25788 32788
rect 25844 32732 25854 32788
rect 30146 32732 30156 32788
rect 30212 32732 31164 32788
rect 31220 32732 32396 32788
rect 32452 32732 32462 32788
rect 33506 32732 33516 32788
rect 33572 32732 34076 32788
rect 34132 32732 34142 32788
rect 36082 32732 36092 32788
rect 36148 32732 36988 32788
rect 37044 32732 37054 32788
rect 22978 32620 22988 32676
rect 23044 32620 23660 32676
rect 23716 32620 24444 32676
rect 24500 32620 26236 32676
rect 26292 32620 27244 32676
rect 27300 32620 27310 32676
rect 29922 32620 29932 32676
rect 29988 32620 31388 32676
rect 31444 32620 31454 32676
rect 0 32508 1820 32564
rect 1876 32508 1886 32564
rect 7970 32508 7980 32564
rect 8036 32508 8046 32564
rect 12898 32508 12908 32564
rect 12964 32508 13580 32564
rect 13636 32508 13646 32564
rect 20850 32508 20860 32564
rect 20916 32508 21308 32564
rect 21364 32508 21374 32564
rect 33506 32508 33516 32564
rect 33572 32508 34524 32564
rect 34580 32508 34590 32564
rect 0 32480 800 32508
rect 3826 32396 3836 32452
rect 3892 32396 5516 32452
rect 5572 32396 6188 32452
rect 6244 32396 6636 32452
rect 6692 32396 7532 32452
rect 7588 32396 8316 32452
rect 8372 32396 15820 32452
rect 15876 32396 15886 32452
rect 23874 32284 23884 32340
rect 23940 32284 24780 32340
rect 24836 32284 26236 32340
rect 26292 32284 26302 32340
rect 32386 32284 32396 32340
rect 32452 32284 33404 32340
rect 33460 32284 33470 32340
rect 3998 32116 4008 32172
rect 4064 32116 4112 32172
rect 4168 32116 4216 32172
rect 4272 32116 4320 32172
rect 4376 32116 4424 32172
rect 4480 32116 4528 32172
rect 4584 32116 4632 32172
rect 4688 32116 4736 32172
rect 4792 32116 4840 32172
rect 4896 32116 4944 32172
rect 5000 32116 5048 32172
rect 5104 32116 5152 32172
rect 5208 32116 5218 32172
rect 23998 32116 24008 32172
rect 24064 32116 24112 32172
rect 24168 32116 24216 32172
rect 24272 32116 24320 32172
rect 24376 32116 24424 32172
rect 24480 32116 24528 32172
rect 24584 32116 24632 32172
rect 24688 32116 24736 32172
rect 24792 32116 24840 32172
rect 24896 32116 24944 32172
rect 25000 32116 25048 32172
rect 25104 32116 25152 32172
rect 25208 32116 25218 32172
rect 3602 32060 3612 32116
rect 3668 32060 3836 32116
rect 3892 32060 3902 32116
rect 35298 31948 35308 32004
rect 35364 31948 36092 32004
rect 36148 31948 36158 32004
rect 5394 31836 5404 31892
rect 5460 31836 5852 31892
rect 5908 31836 6524 31892
rect 6580 31836 6590 31892
rect 7522 31836 7532 31892
rect 7588 31836 7980 31892
rect 8036 31836 8876 31892
rect 8932 31836 8942 31892
rect 9986 31836 9996 31892
rect 10052 31836 12684 31892
rect 12740 31836 21532 31892
rect 21588 31836 21598 31892
rect 21746 31836 21756 31892
rect 21812 31836 22988 31892
rect 23044 31836 23054 31892
rect 23884 31836 23996 31892
rect 24052 31836 25452 31892
rect 25508 31836 25518 31892
rect 26338 31836 26348 31892
rect 26404 31836 29820 31892
rect 29876 31836 29886 31892
rect 34738 31836 34748 31892
rect 34804 31836 36204 31892
rect 36260 31836 36270 31892
rect 5058 31724 5068 31780
rect 5124 31724 6076 31780
rect 6132 31724 6142 31780
rect 8876 31668 8932 31836
rect 23884 31780 23940 31836
rect 10210 31724 10220 31780
rect 10276 31724 13020 31780
rect 13076 31724 13086 31780
rect 16594 31724 16604 31780
rect 16660 31724 17052 31780
rect 17108 31724 18172 31780
rect 18228 31724 18238 31780
rect 22530 31724 22540 31780
rect 22596 31724 23940 31780
rect 26852 31724 27692 31780
rect 27748 31724 27758 31780
rect 28466 31724 28476 31780
rect 28532 31724 32620 31780
rect 32676 31724 33516 31780
rect 33572 31724 34188 31780
rect 34244 31724 34254 31780
rect 26852 31668 26908 31724
rect 8876 31612 13692 31668
rect 13748 31612 13758 31668
rect 14130 31612 14140 31668
rect 14196 31612 14924 31668
rect 14980 31612 15372 31668
rect 15428 31612 15438 31668
rect 15586 31612 15596 31668
rect 15652 31612 17276 31668
rect 17332 31612 17342 31668
rect 21410 31612 21420 31668
rect 21476 31612 25564 31668
rect 25620 31612 26908 31668
rect 27122 31612 27132 31668
rect 27188 31612 28028 31668
rect 28084 31612 28094 31668
rect 13692 31556 13748 31612
rect 13692 31500 15820 31556
rect 15876 31500 15886 31556
rect 17378 31500 17388 31556
rect 17444 31500 18732 31556
rect 18788 31500 18798 31556
rect 26534 31500 26572 31556
rect 26628 31500 26638 31556
rect 27346 31500 27356 31556
rect 27412 31500 29596 31556
rect 29652 31500 29662 31556
rect 31602 31500 31612 31556
rect 31668 31500 32396 31556
rect 32452 31500 32462 31556
rect 33852 31500 33964 31556
rect 34020 31500 34030 31556
rect 0 31444 800 31472
rect 33852 31444 33908 31500
rect 0 31388 2156 31444
rect 2212 31388 2828 31444
rect 2884 31388 2894 31444
rect 27794 31388 27804 31444
rect 27860 31388 30380 31444
rect 30436 31388 32284 31444
rect 32340 31388 33292 31444
rect 33348 31388 33908 31444
rect 0 31360 800 31388
rect 13998 31332 14008 31388
rect 14064 31332 14112 31388
rect 14168 31332 14216 31388
rect 14272 31332 14320 31388
rect 14376 31332 14424 31388
rect 14480 31332 14528 31388
rect 14584 31332 14632 31388
rect 14688 31332 14736 31388
rect 14792 31332 14840 31388
rect 14896 31332 14944 31388
rect 15000 31332 15048 31388
rect 15104 31332 15152 31388
rect 15208 31332 15218 31388
rect 33998 31332 34008 31388
rect 34064 31332 34112 31388
rect 34168 31332 34216 31388
rect 34272 31332 34320 31388
rect 34376 31332 34424 31388
rect 34480 31332 34528 31388
rect 34584 31332 34632 31388
rect 34688 31332 34736 31388
rect 34792 31332 34840 31388
rect 34896 31332 34944 31388
rect 35000 31332 35048 31388
rect 35104 31332 35152 31388
rect 35208 31332 35218 31388
rect 16370 31164 16380 31220
rect 16436 31164 17500 31220
rect 17556 31164 17566 31220
rect 3154 31052 3164 31108
rect 3220 31052 13692 31108
rect 13748 31052 13758 31108
rect 27458 31052 27468 31108
rect 27524 31052 29036 31108
rect 29092 31052 30492 31108
rect 30548 31052 30558 31108
rect 32498 31052 32508 31108
rect 32564 31052 34076 31108
rect 34132 31052 34142 31108
rect 4498 30940 4508 30996
rect 4564 30940 5516 30996
rect 5572 30940 7308 30996
rect 7364 30940 7374 30996
rect 8978 30940 8988 30996
rect 9044 30940 9660 30996
rect 9716 30940 9726 30996
rect 32386 30940 32396 30996
rect 32452 30940 35196 30996
rect 35252 30940 35262 30996
rect 7308 30884 7364 30940
rect 7308 30828 13356 30884
rect 13412 30828 13422 30884
rect 28354 30828 28364 30884
rect 28420 30828 29372 30884
rect 29428 30828 29438 30884
rect 31714 30828 31724 30884
rect 31780 30828 32508 30884
rect 32564 30828 32574 30884
rect 3154 30716 3164 30772
rect 3220 30716 14364 30772
rect 14420 30716 14430 30772
rect 15586 30716 15596 30772
rect 15652 30716 17388 30772
rect 17444 30716 17454 30772
rect 3998 30548 4008 30604
rect 4064 30548 4112 30604
rect 4168 30548 4216 30604
rect 4272 30548 4320 30604
rect 4376 30548 4424 30604
rect 4480 30548 4528 30604
rect 4584 30548 4632 30604
rect 4688 30548 4736 30604
rect 4792 30548 4840 30604
rect 4896 30548 4944 30604
rect 5000 30548 5048 30604
rect 5104 30548 5152 30604
rect 5208 30548 5218 30604
rect 23998 30548 24008 30604
rect 24064 30548 24112 30604
rect 24168 30548 24216 30604
rect 24272 30548 24320 30604
rect 24376 30548 24424 30604
rect 24480 30548 24528 30604
rect 24584 30548 24632 30604
rect 24688 30548 24736 30604
rect 24792 30548 24840 30604
rect 24896 30548 24944 30604
rect 25000 30548 25048 30604
rect 25104 30548 25152 30604
rect 25208 30548 25218 30604
rect 2268 30380 2828 30436
rect 2884 30380 2894 30436
rect 0 30324 800 30352
rect 2268 30324 2324 30380
rect 0 30268 2324 30324
rect 5170 30268 5180 30324
rect 5236 30268 6076 30324
rect 6132 30268 7532 30324
rect 7588 30268 7598 30324
rect 7970 30268 7980 30324
rect 8036 30268 10220 30324
rect 10276 30268 10286 30324
rect 14690 30268 14700 30324
rect 14756 30268 15596 30324
rect 15652 30268 16044 30324
rect 16100 30268 16110 30324
rect 17164 30268 23212 30324
rect 23268 30268 26012 30324
rect 26068 30268 26078 30324
rect 26852 30268 28364 30324
rect 28420 30268 28430 30324
rect 29810 30268 29820 30324
rect 29876 30268 30268 30324
rect 30324 30268 31556 30324
rect 0 30240 800 30268
rect 17164 30212 17220 30268
rect 26852 30212 26908 30268
rect 31500 30212 31556 30268
rect 2594 30156 2604 30212
rect 2660 30156 2670 30212
rect 3154 30156 3164 30212
rect 3220 30156 3724 30212
rect 3780 30156 3790 30212
rect 4722 30156 4732 30212
rect 4788 30156 5292 30212
rect 5348 30156 5358 30212
rect 5842 30156 5852 30212
rect 5908 30156 7308 30212
rect 7364 30156 7868 30212
rect 7924 30156 7934 30212
rect 11666 30156 11676 30212
rect 11732 30156 13020 30212
rect 13076 30156 13086 30212
rect 13346 30156 13356 30212
rect 13412 30156 14252 30212
rect 14308 30156 17164 30212
rect 17220 30156 17230 30212
rect 17826 30156 17836 30212
rect 17892 30156 19740 30212
rect 19796 30156 19806 30212
rect 20066 30156 20076 30212
rect 20132 30156 21420 30212
rect 21476 30156 21486 30212
rect 25330 30156 25340 30212
rect 25396 30156 26684 30212
rect 26740 30156 26908 30212
rect 31490 30156 31500 30212
rect 31556 30156 31836 30212
rect 31892 30156 31902 30212
rect 2604 30100 2660 30156
rect 2604 30044 3948 30100
rect 4004 30044 4014 30100
rect 10322 30044 10332 30100
rect 10388 30044 12460 30100
rect 12516 30044 13468 30100
rect 13524 30044 13534 30100
rect 26852 30044 27692 30100
rect 27748 30044 28588 30100
rect 28644 30044 29820 30100
rect 29876 30044 29886 30100
rect 26852 29988 26908 30044
rect 3266 29932 3276 29988
rect 3332 29932 3724 29988
rect 3780 29932 3790 29988
rect 7746 29932 7756 29988
rect 7812 29932 9772 29988
rect 9828 29932 9838 29988
rect 9986 29932 9996 29988
rect 10052 29932 11340 29988
rect 11396 29932 11406 29988
rect 13458 29932 13468 29988
rect 13524 29932 14364 29988
rect 14420 29932 15708 29988
rect 15764 29932 15774 29988
rect 25442 29932 25452 29988
rect 25508 29932 26124 29988
rect 26180 29932 26908 29988
rect 27570 29932 27580 29988
rect 27636 29932 29260 29988
rect 29316 29932 29326 29988
rect 31612 29932 34636 29988
rect 34692 29932 34702 29988
rect 2146 29820 2156 29876
rect 2212 29820 4060 29876
rect 4116 29820 4126 29876
rect 13998 29764 14008 29820
rect 14064 29764 14112 29820
rect 14168 29764 14216 29820
rect 14272 29764 14320 29820
rect 14376 29764 14424 29820
rect 14480 29764 14528 29820
rect 14584 29764 14632 29820
rect 14688 29764 14736 29820
rect 14792 29764 14840 29820
rect 14896 29764 14944 29820
rect 15000 29764 15048 29820
rect 15104 29764 15152 29820
rect 15208 29764 15218 29820
rect 31612 29764 31668 29932
rect 33998 29764 34008 29820
rect 34064 29764 34112 29820
rect 34168 29764 34216 29820
rect 34272 29764 34320 29820
rect 34376 29764 34424 29820
rect 34480 29764 34528 29820
rect 34584 29764 34632 29820
rect 34688 29764 34736 29820
rect 34792 29764 34840 29820
rect 34896 29764 34944 29820
rect 35000 29764 35048 29820
rect 35104 29764 35152 29820
rect 35208 29764 35218 29820
rect 31602 29708 31612 29764
rect 31668 29708 31678 29764
rect 3938 29596 3948 29652
rect 4004 29596 7084 29652
rect 7140 29596 10780 29652
rect 10836 29596 12348 29652
rect 12404 29596 12414 29652
rect 14466 29596 14476 29652
rect 14532 29596 15484 29652
rect 15540 29596 15596 29652
rect 15652 29596 17276 29652
rect 17332 29596 19292 29652
rect 19348 29596 19740 29652
rect 19796 29596 19806 29652
rect 14476 29540 14532 29596
rect 2034 29484 2044 29540
rect 2100 29484 4620 29540
rect 4676 29484 4686 29540
rect 6850 29484 6860 29540
rect 6916 29484 8092 29540
rect 8148 29484 8876 29540
rect 8932 29484 8942 29540
rect 12450 29484 12460 29540
rect 12516 29484 13804 29540
rect 13860 29484 14532 29540
rect 19842 29484 19852 29540
rect 19908 29484 22316 29540
rect 22372 29484 23324 29540
rect 23380 29484 23390 29540
rect 3826 29372 3836 29428
rect 3892 29372 4508 29428
rect 4564 29372 4574 29428
rect 11890 29372 11900 29428
rect 11956 29372 13580 29428
rect 13636 29372 13646 29428
rect 16034 29372 16044 29428
rect 16100 29372 17388 29428
rect 17444 29372 17454 29428
rect 18722 29372 18732 29428
rect 18788 29372 21084 29428
rect 21140 29372 25452 29428
rect 25508 29372 25518 29428
rect 27122 29372 27132 29428
rect 27188 29372 30268 29428
rect 30324 29372 30940 29428
rect 30996 29372 31006 29428
rect 33058 29372 33068 29428
rect 33124 29372 33516 29428
rect 33572 29372 33582 29428
rect 3490 29260 3500 29316
rect 3556 29260 4732 29316
rect 4788 29260 4798 29316
rect 7410 29260 7420 29316
rect 7476 29260 9660 29316
rect 9716 29260 9726 29316
rect 0 29204 800 29232
rect 0 29148 2156 29204
rect 2212 29148 2222 29204
rect 3836 29148 3948 29204
rect 4004 29148 4014 29204
rect 4834 29148 4844 29204
rect 4900 29148 5348 29204
rect 14690 29148 14700 29204
rect 14756 29148 15372 29204
rect 15428 29148 15438 29204
rect 0 29120 800 29148
rect 2482 28924 2492 28980
rect 2548 28924 3220 28980
rect 3164 28868 3220 28924
rect 3836 28868 3892 29148
rect 3998 28980 4008 29036
rect 4064 28980 4112 29036
rect 4168 28980 4216 29036
rect 4272 28980 4320 29036
rect 4376 28980 4424 29036
rect 4480 28980 4528 29036
rect 4584 28980 4632 29036
rect 4688 28980 4736 29036
rect 4792 28980 4840 29036
rect 4896 28980 4944 29036
rect 5000 28980 5048 29036
rect 5104 28980 5152 29036
rect 5208 28980 5218 29036
rect 5292 28868 5348 29148
rect 13906 29036 13916 29092
rect 13972 29036 14924 29092
rect 14980 29036 14990 29092
rect 23998 28980 24008 29036
rect 24064 28980 24112 29036
rect 24168 28980 24216 29036
rect 24272 28980 24320 29036
rect 24376 28980 24424 29036
rect 24480 28980 24528 29036
rect 24584 28980 24632 29036
rect 24688 28980 24736 29036
rect 24792 28980 24840 29036
rect 24896 28980 24944 29036
rect 25000 28980 25048 29036
rect 25104 28980 25152 29036
rect 25208 28980 25218 29036
rect 13458 28924 13468 28980
rect 13524 28924 14420 28980
rect 3154 28812 3164 28868
rect 3220 28812 3230 28868
rect 3602 28812 3612 28868
rect 3668 28812 4172 28868
rect 4228 28812 4238 28868
rect 4722 28812 4732 28868
rect 4788 28812 5348 28868
rect 3332 28700 9884 28756
rect 9940 28700 9950 28756
rect 3332 28644 3388 28700
rect 14364 28644 14420 28924
rect 21634 28812 21644 28868
rect 21700 28812 22988 28868
rect 23044 28812 23054 28868
rect 20066 28700 20076 28756
rect 20132 28700 21980 28756
rect 22036 28700 23436 28756
rect 23492 28700 23502 28756
rect 2818 28588 2828 28644
rect 2884 28588 3388 28644
rect 3798 28588 3836 28644
rect 3892 28588 4508 28644
rect 4564 28588 4574 28644
rect 7074 28588 7084 28644
rect 7140 28588 7868 28644
rect 7924 28588 7934 28644
rect 9538 28588 9548 28644
rect 9604 28588 11564 28644
rect 11620 28588 11630 28644
rect 14354 28588 14364 28644
rect 14420 28588 14430 28644
rect 15474 28588 15484 28644
rect 15540 28588 18284 28644
rect 18340 28588 18350 28644
rect 25442 28588 25452 28644
rect 25508 28588 28140 28644
rect 28196 28588 28206 28644
rect 29698 28588 29708 28644
rect 29764 28588 31612 28644
rect 31668 28588 33068 28644
rect 33124 28588 33134 28644
rect 11564 28532 11620 28588
rect 1586 28476 1596 28532
rect 1652 28476 3948 28532
rect 4004 28476 4844 28532
rect 4900 28476 4910 28532
rect 5170 28476 5180 28532
rect 5236 28476 5852 28532
rect 5908 28476 5918 28532
rect 6066 28476 6076 28532
rect 6132 28476 6170 28532
rect 11564 28476 13692 28532
rect 13748 28476 13758 28532
rect 16370 28476 16380 28532
rect 16436 28476 16828 28532
rect 16884 28476 17612 28532
rect 17668 28476 17678 28532
rect 31378 28476 31388 28532
rect 31444 28476 33292 28532
rect 33348 28476 33358 28532
rect 16380 28420 16436 28476
rect 2930 28364 2940 28420
rect 2996 28364 3612 28420
rect 3668 28364 3678 28420
rect 3826 28364 3836 28420
rect 3892 28364 5516 28420
rect 5572 28364 5582 28420
rect 6178 28364 6188 28420
rect 6244 28364 8316 28420
rect 8372 28364 8382 28420
rect 13122 28364 13132 28420
rect 13188 28364 15260 28420
rect 15316 28364 16436 28420
rect 31714 28364 31724 28420
rect 31780 28364 32060 28420
rect 32116 28364 32126 28420
rect 13430 28252 13468 28308
rect 13524 28252 13534 28308
rect 13998 28196 14008 28252
rect 14064 28196 14112 28252
rect 14168 28196 14216 28252
rect 14272 28196 14320 28252
rect 14376 28196 14424 28252
rect 14480 28196 14528 28252
rect 14584 28196 14632 28252
rect 14688 28196 14736 28252
rect 14792 28196 14840 28252
rect 14896 28196 14944 28252
rect 15000 28196 15048 28252
rect 15104 28196 15152 28252
rect 15208 28196 15218 28252
rect 5506 28140 5516 28196
rect 5572 28140 6748 28196
rect 6804 28140 6814 28196
rect 0 28084 800 28112
rect 33292 28084 33348 28476
rect 33998 28196 34008 28252
rect 34064 28196 34112 28252
rect 34168 28196 34216 28252
rect 34272 28196 34320 28252
rect 34376 28196 34424 28252
rect 34480 28196 34528 28252
rect 34584 28196 34632 28252
rect 34688 28196 34736 28252
rect 34792 28196 34840 28252
rect 34896 28196 34944 28252
rect 35000 28196 35048 28252
rect 35104 28196 35152 28252
rect 35208 28196 35218 28252
rect 0 28028 1876 28084
rect 18386 28028 18396 28084
rect 18452 28028 20076 28084
rect 20132 28028 20142 28084
rect 23650 28028 23660 28084
rect 23716 28028 25340 28084
rect 25396 28028 26012 28084
rect 26068 28028 26078 28084
rect 33292 28028 33964 28084
rect 34020 28028 34030 28084
rect 0 28000 800 28028
rect 1820 27972 1876 28028
rect 1810 27916 1820 27972
rect 1876 27916 1886 27972
rect 8082 27916 8092 27972
rect 8148 27916 8540 27972
rect 8596 27916 9548 27972
rect 9604 27916 9614 27972
rect 13570 27916 13580 27972
rect 13636 27916 14028 27972
rect 14084 27916 14094 27972
rect 14578 27916 14588 27972
rect 14644 27916 15708 27972
rect 15764 27916 15774 27972
rect 30034 27916 30044 27972
rect 30100 27916 32956 27972
rect 33012 27916 33022 27972
rect 5730 27804 5740 27860
rect 5796 27804 6412 27860
rect 6468 27804 6478 27860
rect 11554 27804 11564 27860
rect 11620 27804 12684 27860
rect 12740 27804 13916 27860
rect 13972 27804 13982 27860
rect 15810 27804 15820 27860
rect 15876 27804 17836 27860
rect 17892 27804 17902 27860
rect 19282 27804 19292 27860
rect 19348 27804 20972 27860
rect 21028 27804 21038 27860
rect 23874 27804 23884 27860
rect 23940 27804 25676 27860
rect 25732 27804 25742 27860
rect 5618 27692 5628 27748
rect 5684 27692 6076 27748
rect 6132 27692 6142 27748
rect 9874 27692 9884 27748
rect 9940 27692 12348 27748
rect 12404 27692 12414 27748
rect 13682 27692 13692 27748
rect 13748 27692 15260 27748
rect 15316 27692 15326 27748
rect 23538 27692 23548 27748
rect 23604 27692 24444 27748
rect 24500 27692 24510 27748
rect 3836 27580 4956 27636
rect 5012 27580 5022 27636
rect 5506 27580 5516 27636
rect 5572 27580 6188 27636
rect 6244 27580 6254 27636
rect 6738 27580 6748 27636
rect 6804 27580 9772 27636
rect 9828 27580 9838 27636
rect 30146 27580 30156 27636
rect 30212 27580 30828 27636
rect 30884 27580 30894 27636
rect 3836 27300 3892 27580
rect 8642 27468 8652 27524
rect 8708 27468 12460 27524
rect 12516 27468 12526 27524
rect 3998 27412 4008 27468
rect 4064 27412 4112 27468
rect 4168 27412 4216 27468
rect 4272 27412 4320 27468
rect 4376 27412 4424 27468
rect 4480 27412 4528 27468
rect 4584 27412 4632 27468
rect 4688 27412 4736 27468
rect 4792 27412 4840 27468
rect 4896 27412 4944 27468
rect 5000 27412 5048 27468
rect 5104 27412 5152 27468
rect 5208 27412 5218 27468
rect 23998 27412 24008 27468
rect 24064 27412 24112 27468
rect 24168 27412 24216 27468
rect 24272 27412 24320 27468
rect 24376 27412 24424 27468
rect 24480 27412 24528 27468
rect 24584 27412 24632 27468
rect 24688 27412 24736 27468
rect 24792 27412 24840 27468
rect 24896 27412 24944 27468
rect 25000 27412 25048 27468
rect 25104 27412 25152 27468
rect 25208 27412 25218 27468
rect 5926 27356 5964 27412
rect 6020 27356 6030 27412
rect 3378 27244 3388 27300
rect 3444 27244 4284 27300
rect 4340 27244 4350 27300
rect 4722 27244 4732 27300
rect 4788 27244 5516 27300
rect 5572 27244 5582 27300
rect 6402 27244 6412 27300
rect 6468 27244 6972 27300
rect 7028 27244 9324 27300
rect 9380 27244 9390 27300
rect 20962 27244 20972 27300
rect 21028 27244 22316 27300
rect 22372 27244 25788 27300
rect 25844 27244 25854 27300
rect 5058 27132 5068 27188
rect 5124 27132 6076 27188
rect 6132 27132 6142 27188
rect 8316 27132 11564 27188
rect 11620 27132 11630 27188
rect 14018 27132 14028 27188
rect 14084 27132 15148 27188
rect 15204 27132 15214 27188
rect 25666 27132 25676 27188
rect 25732 27132 26348 27188
rect 26404 27132 26414 27188
rect 8316 27076 8372 27132
rect 2930 27020 2940 27076
rect 2996 27020 3276 27076
rect 3332 27020 3342 27076
rect 4284 27020 4844 27076
rect 4900 27020 5292 27076
rect 5348 27020 5358 27076
rect 5730 27020 5740 27076
rect 5796 27020 5806 27076
rect 6178 27020 6188 27076
rect 6244 27020 6300 27076
rect 6356 27020 6366 27076
rect 7074 27020 7084 27076
rect 7140 27020 8316 27076
rect 8372 27020 8382 27076
rect 8866 27020 8876 27076
rect 8932 27020 13804 27076
rect 13860 27020 15484 27076
rect 15540 27020 15550 27076
rect 29698 27020 29708 27076
rect 29764 27020 30156 27076
rect 30212 27020 30222 27076
rect 0 26964 800 26992
rect 4284 26964 4340 27020
rect 5740 26964 5796 27020
rect 0 26908 3388 26964
rect 3444 26908 3454 26964
rect 3938 26908 3948 26964
rect 4004 26908 4340 26964
rect 4396 26908 4508 26964
rect 4564 26908 5796 26964
rect 7270 26908 7308 26964
rect 7364 26908 7374 26964
rect 12226 26908 12236 26964
rect 12292 26908 14364 26964
rect 14420 26908 14700 26964
rect 14756 26908 16380 26964
rect 16436 26908 16446 26964
rect 0 26880 800 26908
rect 4396 26852 4452 26908
rect 3154 26796 3164 26852
rect 3220 26796 4452 26852
rect 5730 26796 5740 26852
rect 5796 26796 5964 26852
rect 6020 26796 6636 26852
rect 6692 26796 7084 26852
rect 7140 26796 7150 26852
rect 29810 26796 29820 26852
rect 29876 26796 30940 26852
rect 30996 26796 31006 26852
rect 21186 26684 21196 26740
rect 21252 26684 21980 26740
rect 22036 26684 23660 26740
rect 23716 26684 23726 26740
rect 13998 26628 14008 26684
rect 14064 26628 14112 26684
rect 14168 26628 14216 26684
rect 14272 26628 14320 26684
rect 14376 26628 14424 26684
rect 14480 26628 14528 26684
rect 14584 26628 14632 26684
rect 14688 26628 14736 26684
rect 14792 26628 14840 26684
rect 14896 26628 14944 26684
rect 15000 26628 15048 26684
rect 15104 26628 15152 26684
rect 15208 26628 15218 26684
rect 33998 26628 34008 26684
rect 34064 26628 34112 26684
rect 34168 26628 34216 26684
rect 34272 26628 34320 26684
rect 34376 26628 34424 26684
rect 34480 26628 34528 26684
rect 34584 26628 34632 26684
rect 34688 26628 34736 26684
rect 34792 26628 34840 26684
rect 34896 26628 34944 26684
rect 35000 26628 35048 26684
rect 35104 26628 35152 26684
rect 35208 26628 35218 26684
rect 1810 26572 1820 26628
rect 1876 26572 3612 26628
rect 3668 26572 3678 26628
rect 6038 26572 6076 26628
rect 6132 26572 6142 26628
rect 21410 26572 21420 26628
rect 21476 26572 23212 26628
rect 23268 26572 23278 26628
rect 2594 26460 2604 26516
rect 2660 26460 3836 26516
rect 3892 26460 5292 26516
rect 5348 26460 5852 26516
rect 5908 26460 7756 26516
rect 7812 26460 8092 26516
rect 8148 26460 8158 26516
rect 20402 26460 20412 26516
rect 20468 26460 21756 26516
rect 21812 26460 22092 26516
rect 22148 26460 22158 26516
rect 3266 26236 3276 26292
rect 3332 26236 4620 26292
rect 4676 26236 7196 26292
rect 7252 26236 7262 26292
rect 29586 26236 29596 26292
rect 29652 26236 30716 26292
rect 30772 26236 30782 26292
rect 22642 26124 22652 26180
rect 22708 26124 23772 26180
rect 23828 26124 25676 26180
rect 25732 26124 29260 26180
rect 29316 26124 30604 26180
rect 30660 26124 30670 26180
rect 3042 26012 3052 26068
rect 3108 26012 4956 26068
rect 5012 26012 5628 26068
rect 5684 26012 5964 26068
rect 6020 26012 6030 26068
rect 7186 25900 7196 25956
rect 7252 25900 7644 25956
rect 7700 25900 7710 25956
rect 0 25844 800 25872
rect 3998 25844 4008 25900
rect 4064 25844 4112 25900
rect 4168 25844 4216 25900
rect 4272 25844 4320 25900
rect 4376 25844 4424 25900
rect 4480 25844 4528 25900
rect 4584 25844 4632 25900
rect 4688 25844 4736 25900
rect 4792 25844 4840 25900
rect 4896 25844 4944 25900
rect 5000 25844 5048 25900
rect 5104 25844 5152 25900
rect 5208 25844 5218 25900
rect 23998 25844 24008 25900
rect 24064 25844 24112 25900
rect 24168 25844 24216 25900
rect 24272 25844 24320 25900
rect 24376 25844 24424 25900
rect 24480 25844 24528 25900
rect 24584 25844 24632 25900
rect 24688 25844 24736 25900
rect 24792 25844 24840 25900
rect 24896 25844 24944 25900
rect 25000 25844 25048 25900
rect 25104 25844 25152 25900
rect 25208 25844 25218 25900
rect 0 25788 1708 25844
rect 1764 25788 1774 25844
rect 3154 25788 3164 25844
rect 3220 25788 3892 25844
rect 0 25760 800 25788
rect 3836 25732 3892 25788
rect 6188 25788 11788 25844
rect 6188 25732 6244 25788
rect 3462 25676 3500 25732
rect 3556 25676 3566 25732
rect 3836 25676 6244 25732
rect 7634 25676 7644 25732
rect 7700 25676 8876 25732
rect 8932 25676 8942 25732
rect 11732 25620 11788 25788
rect 20290 25676 20300 25732
rect 20356 25676 20748 25732
rect 20804 25676 23772 25732
rect 23828 25676 27356 25732
rect 27412 25676 27422 25732
rect 32946 25676 32956 25732
rect 33012 25676 34188 25732
rect 34244 25676 34254 25732
rect 3826 25564 3836 25620
rect 3892 25564 4172 25620
rect 4228 25564 4238 25620
rect 5394 25564 5404 25620
rect 5460 25564 8092 25620
rect 8148 25564 8158 25620
rect 11732 25564 13692 25620
rect 13748 25564 14028 25620
rect 14084 25564 14476 25620
rect 14532 25564 14542 25620
rect 29362 25564 29372 25620
rect 29428 25564 30156 25620
rect 30212 25564 33740 25620
rect 33796 25564 33806 25620
rect 3154 25452 3164 25508
rect 3220 25452 6076 25508
rect 6132 25452 6300 25508
rect 6356 25452 6366 25508
rect 29698 25452 29708 25508
rect 29764 25452 30268 25508
rect 30324 25452 30716 25508
rect 30772 25452 30782 25508
rect 4722 25340 4732 25396
rect 4788 25340 5292 25396
rect 5348 25340 5358 25396
rect 26852 25340 27580 25396
rect 27636 25340 27916 25396
rect 27972 25340 27982 25396
rect 26852 25284 26908 25340
rect 5282 25228 5292 25284
rect 5348 25228 6860 25284
rect 6916 25228 7196 25284
rect 7252 25228 9212 25284
rect 9268 25228 10220 25284
rect 10276 25228 12572 25284
rect 12628 25228 13580 25284
rect 13636 25228 13646 25284
rect 15026 25228 15036 25284
rect 15092 25228 15484 25284
rect 15540 25228 15550 25284
rect 21410 25228 21420 25284
rect 21476 25228 22316 25284
rect 22372 25228 22382 25284
rect 23426 25228 23436 25284
rect 23492 25228 24556 25284
rect 24612 25228 26908 25284
rect 27458 25228 27468 25284
rect 27524 25228 28252 25284
rect 28308 25228 28318 25284
rect 31378 25228 31388 25284
rect 31444 25228 33404 25284
rect 33460 25228 33470 25284
rect 26562 25116 26572 25172
rect 26628 25116 26796 25172
rect 26852 25116 26862 25172
rect 27010 25116 27020 25172
rect 27076 25116 28812 25172
rect 28868 25116 28878 25172
rect 13998 25060 14008 25116
rect 14064 25060 14112 25116
rect 14168 25060 14216 25116
rect 14272 25060 14320 25116
rect 14376 25060 14424 25116
rect 14480 25060 14528 25116
rect 14584 25060 14632 25116
rect 14688 25060 14736 25116
rect 14792 25060 14840 25116
rect 14896 25060 14944 25116
rect 15000 25060 15048 25116
rect 15104 25060 15152 25116
rect 15208 25060 15218 25116
rect 33998 25060 34008 25116
rect 34064 25060 34112 25116
rect 34168 25060 34216 25116
rect 34272 25060 34320 25116
rect 34376 25060 34424 25116
rect 34480 25060 34528 25116
rect 34584 25060 34632 25116
rect 34688 25060 34736 25116
rect 34792 25060 34840 25116
rect 34896 25060 34944 25116
rect 35000 25060 35048 25116
rect 35104 25060 35152 25116
rect 35208 25060 35218 25116
rect 26674 25004 26684 25060
rect 26740 25004 29932 25060
rect 29988 25004 29998 25060
rect 6178 24892 6188 24948
rect 6244 24892 18732 24948
rect 18788 24892 19516 24948
rect 19572 24892 19582 24948
rect 27122 24892 27132 24948
rect 27188 24892 28476 24948
rect 28532 24892 29148 24948
rect 29204 24892 29214 24948
rect 12562 24780 12572 24836
rect 12628 24780 14028 24836
rect 14084 24780 15148 24836
rect 24658 24780 24668 24836
rect 24724 24780 25452 24836
rect 25508 24780 26012 24836
rect 26068 24780 27244 24836
rect 27300 24780 27310 24836
rect 0 24724 800 24752
rect 0 24668 2940 24724
rect 2996 24668 3006 24724
rect 3154 24668 3164 24724
rect 3220 24668 3258 24724
rect 3826 24668 3836 24724
rect 3892 24668 6636 24724
rect 6692 24668 8988 24724
rect 9044 24668 10556 24724
rect 10612 24668 10622 24724
rect 0 24640 800 24668
rect 2034 24556 2044 24612
rect 2100 24556 2492 24612
rect 2548 24556 2558 24612
rect 15092 24500 15148 24780
rect 27794 24668 27804 24724
rect 27860 24668 28812 24724
rect 28868 24668 28878 24724
rect 29474 24668 29484 24724
rect 29540 24668 30492 24724
rect 30548 24668 30558 24724
rect 18274 24556 18284 24612
rect 18340 24556 19740 24612
rect 19796 24556 20188 24612
rect 20244 24556 20254 24612
rect 25778 24556 25788 24612
rect 25844 24556 27916 24612
rect 27972 24556 27982 24612
rect 28140 24500 28196 24668
rect 29586 24556 29596 24612
rect 29652 24556 30268 24612
rect 30324 24556 30334 24612
rect 8306 24444 8316 24500
rect 8372 24444 9660 24500
rect 9716 24444 9726 24500
rect 15092 24444 15372 24500
rect 15428 24444 15438 24500
rect 23090 24444 23100 24500
rect 23156 24444 25228 24500
rect 25284 24444 25294 24500
rect 26674 24444 26684 24500
rect 26740 24444 28196 24500
rect 10770 24332 10780 24388
rect 10836 24332 11564 24388
rect 11620 24332 16492 24388
rect 16548 24332 16558 24388
rect 3998 24276 4008 24332
rect 4064 24276 4112 24332
rect 4168 24276 4216 24332
rect 4272 24276 4320 24332
rect 4376 24276 4424 24332
rect 4480 24276 4528 24332
rect 4584 24276 4632 24332
rect 4688 24276 4736 24332
rect 4792 24276 4840 24332
rect 4896 24276 4944 24332
rect 5000 24276 5048 24332
rect 5104 24276 5152 24332
rect 5208 24276 5218 24332
rect 23998 24276 24008 24332
rect 24064 24276 24112 24332
rect 24168 24276 24216 24332
rect 24272 24276 24320 24332
rect 24376 24276 24424 24332
rect 24480 24276 24528 24332
rect 24584 24276 24632 24332
rect 24688 24276 24736 24332
rect 24792 24276 24840 24332
rect 24896 24276 24944 24332
rect 25000 24276 25048 24332
rect 25104 24276 25152 24332
rect 25208 24276 25218 24332
rect 26002 24108 26012 24164
rect 26068 24108 30604 24164
rect 30660 24108 30670 24164
rect 22866 23996 22876 24052
rect 22932 23996 24556 24052
rect 24612 23996 24622 24052
rect 27234 23996 27244 24052
rect 27300 23996 27916 24052
rect 27972 23996 29484 24052
rect 29540 23996 31052 24052
rect 31108 23996 31118 24052
rect 24882 23884 24892 23940
rect 24948 23884 27020 23940
rect 27076 23884 27086 23940
rect 28130 23884 28140 23940
rect 28196 23884 29148 23940
rect 29204 23884 29214 23940
rect 28140 23828 28196 23884
rect 2706 23772 2716 23828
rect 2772 23772 4508 23828
rect 4564 23772 4574 23828
rect 11666 23772 11676 23828
rect 11732 23772 12236 23828
rect 12292 23772 12302 23828
rect 13794 23772 13804 23828
rect 13860 23772 14364 23828
rect 14420 23772 14430 23828
rect 16594 23772 16604 23828
rect 16660 23772 18844 23828
rect 18900 23772 19852 23828
rect 19908 23772 19918 23828
rect 20402 23772 20412 23828
rect 20468 23772 21756 23828
rect 21812 23772 22764 23828
rect 22820 23772 22830 23828
rect 26852 23772 28196 23828
rect 3266 23660 3276 23716
rect 3332 23660 3388 23716
rect 3444 23660 3454 23716
rect 11218 23660 11228 23716
rect 11284 23660 11900 23716
rect 11956 23660 11966 23716
rect 13570 23660 13580 23716
rect 13636 23660 13916 23716
rect 13972 23660 13982 23716
rect 16482 23660 16492 23716
rect 16548 23660 17836 23716
rect 17892 23660 20636 23716
rect 20692 23660 20702 23716
rect 23762 23660 23772 23716
rect 23828 23660 24444 23716
rect 24500 23660 24510 23716
rect 24658 23660 24668 23716
rect 24724 23660 26684 23716
rect 26740 23660 26750 23716
rect 0 23604 800 23632
rect 24444 23604 24500 23660
rect 26852 23604 26908 23772
rect 27010 23660 27020 23716
rect 27076 23660 29708 23716
rect 29764 23660 29774 23716
rect 30258 23660 30268 23716
rect 30324 23660 31500 23716
rect 31556 23660 31948 23716
rect 32004 23660 32014 23716
rect 0 23548 2156 23604
rect 2212 23548 2222 23604
rect 4498 23548 4508 23604
rect 4564 23548 6412 23604
rect 6468 23548 6478 23604
rect 15474 23548 15484 23604
rect 15540 23548 16268 23604
rect 16324 23548 18284 23604
rect 18340 23548 18350 23604
rect 24444 23548 26908 23604
rect 27794 23548 27804 23604
rect 27860 23548 29372 23604
rect 29428 23548 29438 23604
rect 0 23520 800 23548
rect 3266 23492 3276 23548
rect 3332 23492 3342 23548
rect 13998 23492 14008 23548
rect 14064 23492 14112 23548
rect 14168 23492 14216 23548
rect 14272 23492 14320 23548
rect 14376 23492 14424 23548
rect 14480 23492 14528 23548
rect 14584 23492 14632 23548
rect 14688 23492 14736 23548
rect 14792 23492 14840 23548
rect 14896 23492 14944 23548
rect 15000 23492 15048 23548
rect 15104 23492 15152 23548
rect 15208 23492 15218 23548
rect 33998 23492 34008 23548
rect 34064 23492 34112 23548
rect 34168 23492 34216 23548
rect 34272 23492 34320 23548
rect 34376 23492 34424 23548
rect 34480 23492 34528 23548
rect 34584 23492 34632 23548
rect 34688 23492 34736 23548
rect 34792 23492 34840 23548
rect 34896 23492 34944 23548
rect 35000 23492 35048 23548
rect 35104 23492 35152 23548
rect 35208 23492 35218 23548
rect 1810 23436 1820 23492
rect 1876 23436 2828 23492
rect 2884 23436 2894 23492
rect 3042 23436 3052 23492
rect 3108 23436 3332 23492
rect 3826 23436 3836 23492
rect 3892 23436 5180 23492
rect 5236 23436 6188 23492
rect 6244 23436 6254 23492
rect 6402 23436 6412 23492
rect 6468 23436 6636 23492
rect 6692 23436 6702 23492
rect 13654 23436 13692 23492
rect 13748 23436 13758 23492
rect 28140 23436 31388 23492
rect 31444 23436 31612 23492
rect 31668 23436 31678 23492
rect 28140 23380 28196 23436
rect 1708 23324 15932 23380
rect 15988 23324 15998 23380
rect 20962 23324 20972 23380
rect 21028 23324 21868 23380
rect 21924 23324 23436 23380
rect 23492 23324 23502 23380
rect 27570 23324 27580 23380
rect 27636 23324 28140 23380
rect 28196 23324 28206 23380
rect 29586 23324 29596 23380
rect 29652 23324 30604 23380
rect 30660 23324 30670 23380
rect 1708 23156 1764 23324
rect 1922 23212 1932 23268
rect 1988 23212 3612 23268
rect 3668 23212 3678 23268
rect 3826 23212 3836 23268
rect 3892 23212 3948 23268
rect 4004 23212 4014 23268
rect 5394 23212 5404 23268
rect 5460 23212 6636 23268
rect 6692 23212 6702 23268
rect 13346 23212 13356 23268
rect 13412 23212 21980 23268
rect 22036 23212 24108 23268
rect 24164 23212 25340 23268
rect 25396 23212 25406 23268
rect 1708 23100 2268 23156
rect 2324 23100 2334 23156
rect 9650 23100 9660 23156
rect 9716 23100 11116 23156
rect 11172 23100 13468 23156
rect 13524 23100 13534 23156
rect 13794 23100 13804 23156
rect 13860 23100 14588 23156
rect 14644 23100 14654 23156
rect 13804 23044 13860 23100
rect 3378 22988 3388 23044
rect 3444 22988 7756 23044
rect 7812 22988 7822 23044
rect 12450 22988 12460 23044
rect 12516 22988 13860 23044
rect 18386 22988 18396 23044
rect 18452 22988 21308 23044
rect 21364 22988 23660 23044
rect 23716 22988 23726 23044
rect 1698 22876 1708 22932
rect 1764 22876 2268 22932
rect 2324 22876 2334 22932
rect 3164 22876 3948 22932
rect 4004 22876 4014 22932
rect 4498 22876 4508 22932
rect 4564 22876 5292 22932
rect 5348 22876 5358 22932
rect 13682 22876 13692 22932
rect 13748 22876 13916 22932
rect 13972 22876 13982 22932
rect 3164 22820 3220 22876
rect 2370 22764 2380 22820
rect 2436 22764 3220 22820
rect 3998 22708 4008 22764
rect 4064 22708 4112 22764
rect 4168 22708 4216 22764
rect 4272 22708 4320 22764
rect 4376 22708 4424 22764
rect 4480 22708 4528 22764
rect 4584 22708 4632 22764
rect 4688 22708 4736 22764
rect 4792 22708 4840 22764
rect 4896 22708 4944 22764
rect 5000 22708 5048 22764
rect 5104 22708 5152 22764
rect 5208 22708 5218 22764
rect 23998 22708 24008 22764
rect 24064 22708 24112 22764
rect 24168 22708 24216 22764
rect 24272 22708 24320 22764
rect 24376 22708 24424 22764
rect 24480 22708 24528 22764
rect 24584 22708 24632 22764
rect 24688 22708 24736 22764
rect 24792 22708 24840 22764
rect 24896 22708 24944 22764
rect 25000 22708 25048 22764
rect 25104 22708 25152 22764
rect 25208 22708 25218 22764
rect 13766 22652 13804 22708
rect 13860 22652 13870 22708
rect 30034 22652 30044 22708
rect 30100 22652 30492 22708
rect 30548 22652 31388 22708
rect 31444 22652 33628 22708
rect 33684 22652 33694 22708
rect 2482 22540 2492 22596
rect 2548 22540 4172 22596
rect 4228 22540 4238 22596
rect 10546 22540 10556 22596
rect 10612 22540 13692 22596
rect 13748 22540 13758 22596
rect 23986 22540 23996 22596
rect 24052 22540 26908 22596
rect 26964 22540 27580 22596
rect 27636 22540 27646 22596
rect 28130 22540 28140 22596
rect 28196 22540 33852 22596
rect 33908 22540 33918 22596
rect 0 22484 800 22512
rect 0 22428 1708 22484
rect 1764 22428 1774 22484
rect 7298 22428 7308 22484
rect 7364 22428 20860 22484
rect 20916 22428 21756 22484
rect 21812 22428 21822 22484
rect 23874 22428 23884 22484
rect 23940 22428 25452 22484
rect 25508 22428 25518 22484
rect 27346 22428 27356 22484
rect 27412 22428 29484 22484
rect 29540 22428 29550 22484
rect 0 22400 800 22428
rect 2482 22316 2492 22372
rect 2548 22316 2828 22372
rect 2884 22316 2894 22372
rect 11778 22316 11788 22372
rect 11844 22316 12460 22372
rect 12516 22316 12526 22372
rect 15362 22316 15372 22372
rect 15428 22316 17500 22372
rect 17556 22316 17566 22372
rect 20402 22316 20412 22372
rect 20468 22316 23100 22372
rect 23156 22316 28924 22372
rect 28980 22316 28990 22372
rect 11554 22204 11564 22260
rect 11620 22204 12124 22260
rect 12180 22204 12190 22260
rect 13682 22204 13692 22260
rect 13748 22204 14140 22260
rect 14196 22204 14206 22260
rect 14690 22204 14700 22260
rect 14756 22204 17052 22260
rect 17108 22204 17118 22260
rect 20178 22204 20188 22260
rect 20244 22204 21980 22260
rect 22036 22204 22046 22260
rect 24882 22204 24892 22260
rect 24948 22204 25228 22260
rect 25284 22204 25340 22260
rect 25396 22204 27356 22260
rect 27412 22204 27422 22260
rect 29698 22204 29708 22260
rect 29764 22204 30044 22260
rect 30100 22204 30110 22260
rect 4834 22092 4844 22148
rect 4900 22092 5404 22148
rect 5460 22092 6076 22148
rect 6132 22092 6142 22148
rect 12226 22092 12236 22148
rect 12292 22092 13692 22148
rect 13748 22092 13758 22148
rect 13998 21924 14008 21980
rect 14064 21924 14112 21980
rect 14168 21924 14216 21980
rect 14272 21924 14320 21980
rect 14376 21924 14424 21980
rect 14480 21924 14528 21980
rect 14584 21924 14632 21980
rect 14688 21924 14736 21980
rect 14792 21924 14840 21980
rect 14896 21924 14944 21980
rect 15000 21924 15048 21980
rect 15104 21924 15152 21980
rect 15208 21924 15218 21980
rect 15372 21812 15428 22204
rect 18498 22092 18508 22148
rect 18564 22092 19404 22148
rect 19460 22092 20972 22148
rect 21028 22092 23324 22148
rect 23380 22092 23996 22148
rect 24052 22092 24062 22148
rect 25442 22092 25452 22148
rect 25508 22092 26348 22148
rect 26404 22092 27020 22148
rect 27076 22092 29260 22148
rect 29316 22092 29326 22148
rect 30146 22092 30156 22148
rect 30212 22092 30492 22148
rect 30548 22092 30558 22148
rect 23426 21980 23436 22036
rect 23492 21980 26460 22036
rect 26516 21980 26526 22036
rect 27570 21980 27580 22036
rect 27636 21980 29708 22036
rect 29764 21980 29774 22036
rect 33998 21924 34008 21980
rect 34064 21924 34112 21980
rect 34168 21924 34216 21980
rect 34272 21924 34320 21980
rect 34376 21924 34424 21980
rect 34480 21924 34528 21980
rect 34584 21924 34632 21980
rect 34688 21924 34736 21980
rect 34792 21924 34840 21980
rect 34896 21924 34944 21980
rect 35000 21924 35048 21980
rect 35104 21924 35152 21980
rect 35208 21924 35218 21980
rect 28578 21868 28588 21924
rect 28644 21868 30044 21924
rect 30100 21868 31052 21924
rect 31108 21868 31118 21924
rect 4834 21756 4844 21812
rect 4900 21756 6188 21812
rect 6244 21756 6254 21812
rect 6738 21756 6748 21812
rect 6804 21756 8428 21812
rect 8484 21756 8876 21812
rect 8932 21756 8942 21812
rect 15250 21756 15260 21812
rect 15316 21756 15428 21812
rect 23538 21756 23548 21812
rect 23604 21756 24668 21812
rect 24724 21756 24734 21812
rect 26786 21756 26796 21812
rect 26852 21756 29148 21812
rect 29204 21756 29214 21812
rect 3826 21644 3836 21700
rect 3892 21644 6188 21700
rect 6244 21644 6254 21700
rect 6962 21644 6972 21700
rect 7028 21644 8764 21700
rect 8820 21644 8830 21700
rect 16706 21644 16716 21700
rect 16772 21644 18620 21700
rect 18676 21644 18686 21700
rect 1698 21532 1708 21588
rect 1764 21532 5628 21588
rect 5684 21532 5694 21588
rect 6402 21532 6412 21588
rect 6468 21532 6860 21588
rect 6916 21532 7532 21588
rect 7588 21532 7598 21588
rect 16594 21532 16604 21588
rect 16660 21532 17500 21588
rect 17556 21532 21532 21588
rect 21588 21532 21598 21588
rect 6412 21476 6468 21532
rect 5394 21420 5404 21476
rect 5460 21420 6468 21476
rect 12562 21420 12572 21476
rect 12628 21420 15148 21476
rect 29698 21420 29708 21476
rect 29764 21420 30156 21476
rect 30212 21420 30222 21476
rect 0 21364 800 21392
rect 0 21308 1820 21364
rect 1876 21308 2604 21364
rect 2660 21308 2670 21364
rect 10322 21308 10332 21364
rect 10388 21308 13132 21364
rect 13188 21308 13198 21364
rect 15092 21308 15148 21420
rect 15204 21308 15596 21364
rect 15652 21308 15662 21364
rect 22978 21308 22988 21364
rect 23044 21308 24780 21364
rect 24836 21308 27692 21364
rect 27748 21308 27758 21364
rect 0 21280 800 21308
rect 13682 21196 13692 21252
rect 13748 21196 16380 21252
rect 16436 21196 16446 21252
rect 3998 21140 4008 21196
rect 4064 21140 4112 21196
rect 4168 21140 4216 21196
rect 4272 21140 4320 21196
rect 4376 21140 4424 21196
rect 4480 21140 4528 21196
rect 4584 21140 4632 21196
rect 4688 21140 4736 21196
rect 4792 21140 4840 21196
rect 4896 21140 4944 21196
rect 5000 21140 5048 21196
rect 5104 21140 5152 21196
rect 5208 21140 5218 21196
rect 23998 21140 24008 21196
rect 24064 21140 24112 21196
rect 24168 21140 24216 21196
rect 24272 21140 24320 21196
rect 24376 21140 24424 21196
rect 24480 21140 24528 21196
rect 24584 21140 24632 21196
rect 24688 21140 24736 21196
rect 24792 21140 24840 21196
rect 24896 21140 24944 21196
rect 25000 21140 25048 21196
rect 25104 21140 25152 21196
rect 25208 21140 25218 21196
rect 4498 20972 4508 21028
rect 4564 20972 5292 21028
rect 5348 20972 5358 21028
rect 13682 20972 13692 21028
rect 13748 20972 14140 21028
rect 14196 20972 14206 21028
rect 21410 20972 21420 21028
rect 21476 20972 22204 21028
rect 22260 20972 22270 21028
rect 24210 20972 24220 21028
rect 24276 20972 25788 21028
rect 25844 20972 25854 21028
rect 13682 20860 13692 20916
rect 13748 20860 15148 20916
rect 15204 20860 16716 20916
rect 16772 20860 16782 20916
rect 20738 20860 20748 20916
rect 20804 20860 24108 20916
rect 24164 20860 24668 20916
rect 24724 20860 24734 20916
rect 25218 20860 25228 20916
rect 25284 20860 25676 20916
rect 25732 20860 26236 20916
rect 26292 20860 26302 20916
rect 26852 20860 28588 20916
rect 28644 20860 28654 20916
rect 26852 20804 26908 20860
rect 4610 20748 4620 20804
rect 4676 20748 5404 20804
rect 5460 20748 6076 20804
rect 6132 20748 6142 20804
rect 8418 20748 8428 20804
rect 8484 20748 9100 20804
rect 9156 20748 9772 20804
rect 9828 20748 12908 20804
rect 12964 20748 12974 20804
rect 21522 20748 21532 20804
rect 21588 20748 22428 20804
rect 22484 20748 22494 20804
rect 23202 20748 23212 20804
rect 23268 20748 24556 20804
rect 24612 20748 26908 20804
rect 27346 20748 27356 20804
rect 27412 20748 28252 20804
rect 28308 20748 28318 20804
rect 29474 20748 29484 20804
rect 29540 20748 30380 20804
rect 30436 20748 30446 20804
rect 3154 20636 3164 20692
rect 3220 20636 5516 20692
rect 5572 20636 5582 20692
rect 6178 20636 6188 20692
rect 6244 20636 6748 20692
rect 6804 20636 6814 20692
rect 9314 20636 9324 20692
rect 9380 20636 10332 20692
rect 10388 20636 10398 20692
rect 24770 20636 24780 20692
rect 24836 20636 25340 20692
rect 25396 20636 25406 20692
rect 29586 20636 29596 20692
rect 29652 20636 31836 20692
rect 31892 20636 32732 20692
rect 32788 20636 32798 20692
rect 5058 20524 5068 20580
rect 5124 20524 6636 20580
rect 6692 20524 6702 20580
rect 8754 20524 8764 20580
rect 8820 20524 9548 20580
rect 9604 20524 9614 20580
rect 12338 20524 12348 20580
rect 12404 20524 13804 20580
rect 13860 20524 14140 20580
rect 14196 20524 14588 20580
rect 14644 20524 14654 20580
rect 23650 20524 23660 20580
rect 23716 20524 29708 20580
rect 29764 20524 29774 20580
rect 13998 20356 14008 20412
rect 14064 20356 14112 20412
rect 14168 20356 14216 20412
rect 14272 20356 14320 20412
rect 14376 20356 14424 20412
rect 14480 20356 14528 20412
rect 14584 20356 14632 20412
rect 14688 20356 14736 20412
rect 14792 20356 14840 20412
rect 14896 20356 14944 20412
rect 15000 20356 15048 20412
rect 15104 20356 15152 20412
rect 15208 20356 15218 20412
rect 33998 20356 34008 20412
rect 34064 20356 34112 20412
rect 34168 20356 34216 20412
rect 34272 20356 34320 20412
rect 34376 20356 34424 20412
rect 34480 20356 34528 20412
rect 34584 20356 34632 20412
rect 34688 20356 34736 20412
rect 34792 20356 34840 20412
rect 34896 20356 34944 20412
rect 35000 20356 35048 20412
rect 35104 20356 35152 20412
rect 35208 20356 35218 20412
rect 0 20244 800 20272
rect 0 20188 2492 20244
rect 2548 20188 2558 20244
rect 6150 20188 6188 20244
rect 6244 20188 6254 20244
rect 13122 20188 13132 20244
rect 13188 20188 14028 20244
rect 14084 20188 14094 20244
rect 25302 20188 25340 20244
rect 25396 20188 25406 20244
rect 0 20160 800 20188
rect 9650 20076 9660 20132
rect 9716 20076 10332 20132
rect 10388 20076 10398 20132
rect 10546 20076 10556 20132
rect 10612 20076 11564 20132
rect 11620 20076 11630 20132
rect 11778 20076 11788 20132
rect 11844 20076 12572 20132
rect 12628 20076 13692 20132
rect 13748 20076 15148 20132
rect 15586 20076 15596 20132
rect 15652 20076 16044 20132
rect 16100 20076 18284 20132
rect 18340 20076 18732 20132
rect 18788 20076 18798 20132
rect 20290 20076 20300 20132
rect 20356 20076 25452 20132
rect 25508 20076 30268 20132
rect 30324 20076 30334 20132
rect 30818 20076 30828 20132
rect 30884 20076 31948 20132
rect 32004 20076 33628 20132
rect 33684 20076 33694 20132
rect 15092 20020 15148 20076
rect 8866 19964 8876 20020
rect 8932 19964 9884 20020
rect 9940 19964 9950 20020
rect 13458 19964 13468 20020
rect 13524 19964 13916 20020
rect 13972 19964 14812 20020
rect 14868 19964 14878 20020
rect 15092 19964 16492 20020
rect 16548 19964 16558 20020
rect 22530 19964 22540 20020
rect 22596 19964 23212 20020
rect 23268 19964 23660 20020
rect 23716 19964 25564 20020
rect 25620 19964 25630 20020
rect 28018 19964 28028 20020
rect 28084 19964 30156 20020
rect 30212 19964 30222 20020
rect 14242 19852 14252 19908
rect 14308 19852 15708 19908
rect 15764 19852 15774 19908
rect 16594 19852 16604 19908
rect 16660 19852 23548 19908
rect 23604 19852 23614 19908
rect 29810 19852 29820 19908
rect 29876 19852 30940 19908
rect 30996 19852 31006 19908
rect 21410 19740 21420 19796
rect 21476 19740 23772 19796
rect 23828 19740 23838 19796
rect 28466 19740 28476 19796
rect 28532 19740 29932 19796
rect 29988 19740 29998 19796
rect 30258 19740 30268 19796
rect 30324 19740 32284 19796
rect 32340 19740 32350 19796
rect 25666 19628 25676 19684
rect 25732 19628 27244 19684
rect 27300 19628 27310 19684
rect 27458 19628 27468 19684
rect 27524 19628 31500 19684
rect 31556 19628 31566 19684
rect 3998 19572 4008 19628
rect 4064 19572 4112 19628
rect 4168 19572 4216 19628
rect 4272 19572 4320 19628
rect 4376 19572 4424 19628
rect 4480 19572 4528 19628
rect 4584 19572 4632 19628
rect 4688 19572 4736 19628
rect 4792 19572 4840 19628
rect 4896 19572 4944 19628
rect 5000 19572 5048 19628
rect 5104 19572 5152 19628
rect 5208 19572 5218 19628
rect 23998 19572 24008 19628
rect 24064 19572 24112 19628
rect 24168 19572 24216 19628
rect 24272 19572 24320 19628
rect 24376 19572 24424 19628
rect 24480 19572 24528 19628
rect 24584 19572 24632 19628
rect 24688 19572 24736 19628
rect 24792 19572 24840 19628
rect 24896 19572 24944 19628
rect 25000 19572 25048 19628
rect 25104 19572 25152 19628
rect 25208 19572 25218 19628
rect 20514 19404 20524 19460
rect 20580 19404 21420 19460
rect 21476 19404 21486 19460
rect 26898 19404 26908 19460
rect 26964 19404 27804 19460
rect 27860 19404 27870 19460
rect 14578 19292 14588 19348
rect 14644 19292 15820 19348
rect 15876 19292 15886 19348
rect 2482 19180 2492 19236
rect 2548 19180 2558 19236
rect 2818 19180 2828 19236
rect 2884 19180 3612 19236
rect 3668 19180 3678 19236
rect 13356 19180 14700 19236
rect 14756 19180 14766 19236
rect 18946 19180 18956 19236
rect 19012 19180 20524 19236
rect 20580 19180 20590 19236
rect 25106 19180 25116 19236
rect 25172 19180 25340 19236
rect 25396 19180 25406 19236
rect 27122 19180 27132 19236
rect 27188 19180 27468 19236
rect 27524 19180 27534 19236
rect 28354 19180 28364 19236
rect 28420 19180 29148 19236
rect 29204 19180 29214 19236
rect 30034 19180 30044 19236
rect 30100 19180 32732 19236
rect 32788 19180 32798 19236
rect 0 19124 800 19152
rect 2492 19124 2548 19180
rect 13356 19124 13412 19180
rect 0 19068 2548 19124
rect 13346 19068 13356 19124
rect 13412 19068 13422 19124
rect 13682 19068 13692 19124
rect 13748 19068 14364 19124
rect 14420 19068 14430 19124
rect 16380 19068 18508 19124
rect 18564 19068 18574 19124
rect 19506 19068 19516 19124
rect 19572 19068 20300 19124
rect 20356 19068 20366 19124
rect 26450 19068 26460 19124
rect 26516 19068 28476 19124
rect 28532 19068 28542 19124
rect 0 19040 800 19068
rect 16380 19012 16436 19068
rect 14242 18956 14252 19012
rect 14308 18956 16380 19012
rect 16436 18956 16446 19012
rect 18050 18956 18060 19012
rect 18116 18956 19628 19012
rect 19684 18956 19694 19012
rect 13998 18788 14008 18844
rect 14064 18788 14112 18844
rect 14168 18788 14216 18844
rect 14272 18788 14320 18844
rect 14376 18788 14424 18844
rect 14480 18788 14528 18844
rect 14584 18788 14632 18844
rect 14688 18788 14736 18844
rect 14792 18788 14840 18844
rect 14896 18788 14944 18844
rect 15000 18788 15048 18844
rect 15104 18788 15152 18844
rect 15208 18788 15218 18844
rect 33998 18788 34008 18844
rect 34064 18788 34112 18844
rect 34168 18788 34216 18844
rect 34272 18788 34320 18844
rect 34376 18788 34424 18844
rect 34480 18788 34528 18844
rect 34584 18788 34632 18844
rect 34688 18788 34736 18844
rect 34792 18788 34840 18844
rect 34896 18788 34944 18844
rect 35000 18788 35048 18844
rect 35104 18788 35152 18844
rect 35208 18788 35218 18844
rect 6402 18732 6412 18788
rect 6468 18732 7420 18788
rect 7476 18732 7486 18788
rect 23762 18620 23772 18676
rect 23828 18620 25788 18676
rect 25844 18620 25854 18676
rect 27122 18620 27132 18676
rect 27188 18620 27916 18676
rect 27972 18620 27982 18676
rect 28130 18620 28140 18676
rect 28196 18620 29596 18676
rect 29652 18620 30604 18676
rect 30660 18620 30670 18676
rect 12226 18508 12236 18564
rect 12292 18508 13916 18564
rect 13972 18508 13982 18564
rect 26338 18508 26348 18564
rect 26404 18508 26796 18564
rect 26852 18508 29036 18564
rect 29092 18508 30828 18564
rect 30884 18508 30894 18564
rect 16706 18396 16716 18452
rect 16772 18396 21196 18452
rect 21252 18396 21262 18452
rect 12562 18284 12572 18340
rect 12628 18284 13020 18340
rect 13076 18284 14812 18340
rect 14868 18284 14878 18340
rect 15810 18284 15820 18340
rect 15876 18284 16604 18340
rect 16660 18284 16670 18340
rect 28354 18284 28364 18340
rect 28420 18284 30156 18340
rect 30212 18284 30222 18340
rect 19282 18172 19292 18228
rect 19348 18172 21084 18228
rect 21140 18172 22652 18228
rect 22708 18172 22718 18228
rect 22418 18060 22428 18116
rect 22484 18060 23212 18116
rect 23268 18060 23278 18116
rect 0 17920 800 18032
rect 3998 18004 4008 18060
rect 4064 18004 4112 18060
rect 4168 18004 4216 18060
rect 4272 18004 4320 18060
rect 4376 18004 4424 18060
rect 4480 18004 4528 18060
rect 4584 18004 4632 18060
rect 4688 18004 4736 18060
rect 4792 18004 4840 18060
rect 4896 18004 4944 18060
rect 5000 18004 5048 18060
rect 5104 18004 5152 18060
rect 5208 18004 5218 18060
rect 23998 18004 24008 18060
rect 24064 18004 24112 18060
rect 24168 18004 24216 18060
rect 24272 18004 24320 18060
rect 24376 18004 24424 18060
rect 24480 18004 24528 18060
rect 24584 18004 24632 18060
rect 24688 18004 24736 18060
rect 24792 18004 24840 18060
rect 24896 18004 24944 18060
rect 25000 18004 25048 18060
rect 25104 18004 25152 18060
rect 25208 18004 25218 18060
rect 12002 17948 12012 18004
rect 12068 17948 12684 18004
rect 12740 17948 13804 18004
rect 13860 17948 13870 18004
rect 3266 17836 3276 17892
rect 3332 17836 4172 17892
rect 4228 17836 4238 17892
rect 3826 17724 3836 17780
rect 3892 17724 17948 17780
rect 18004 17724 18014 17780
rect 8530 17612 8540 17668
rect 8596 17612 9996 17668
rect 10052 17612 10062 17668
rect 10882 17612 10892 17668
rect 10948 17612 11900 17668
rect 11956 17612 11966 17668
rect 19394 17612 19404 17668
rect 19460 17612 20412 17668
rect 20468 17612 21532 17668
rect 21588 17612 21598 17668
rect 22306 17612 22316 17668
rect 22372 17612 23100 17668
rect 23156 17612 23166 17668
rect 9996 17556 10052 17612
rect 4946 17500 4956 17556
rect 5012 17500 7084 17556
rect 7140 17500 9212 17556
rect 9268 17500 9660 17556
rect 9716 17500 9726 17556
rect 9996 17500 13804 17556
rect 13860 17500 14420 17556
rect 18610 17500 18620 17556
rect 18676 17500 19292 17556
rect 19348 17500 19358 17556
rect 21858 17500 21868 17556
rect 21924 17500 22764 17556
rect 22820 17500 22830 17556
rect 26198 17500 26236 17556
rect 26292 17500 26796 17556
rect 26852 17500 26862 17556
rect 14364 17444 14420 17500
rect 8642 17388 8652 17444
rect 8708 17388 10780 17444
rect 10836 17388 10846 17444
rect 11106 17388 11116 17444
rect 11172 17388 11564 17444
rect 11620 17388 12348 17444
rect 12404 17388 12908 17444
rect 12964 17388 12974 17444
rect 14354 17388 14364 17444
rect 14420 17388 18060 17444
rect 18116 17388 18126 17444
rect 18498 17388 18508 17444
rect 18564 17388 23548 17444
rect 23604 17388 24892 17444
rect 24948 17388 24958 17444
rect 26852 17388 28252 17444
rect 28308 17388 29708 17444
rect 29764 17388 29774 17444
rect 11218 17276 11228 17332
rect 11284 17276 12572 17332
rect 12628 17276 12638 17332
rect 22418 17276 22428 17332
rect 22484 17276 23884 17332
rect 23940 17276 25340 17332
rect 25396 17276 25406 17332
rect 13998 17220 14008 17276
rect 14064 17220 14112 17276
rect 14168 17220 14216 17276
rect 14272 17220 14320 17276
rect 14376 17220 14424 17276
rect 14480 17220 14528 17276
rect 14584 17220 14632 17276
rect 14688 17220 14736 17276
rect 14792 17220 14840 17276
rect 14896 17220 14944 17276
rect 15000 17220 15048 17276
rect 15104 17220 15152 17276
rect 15208 17220 15218 17276
rect 26852 17220 26908 17388
rect 33998 17220 34008 17276
rect 34064 17220 34112 17276
rect 34168 17220 34216 17276
rect 34272 17220 34320 17276
rect 34376 17220 34424 17276
rect 34480 17220 34528 17276
rect 34584 17220 34632 17276
rect 34688 17220 34736 17276
rect 34792 17220 34840 17276
rect 34896 17220 34944 17276
rect 35000 17220 35048 17276
rect 35104 17220 35152 17276
rect 35208 17220 35218 17276
rect 15362 17164 15372 17220
rect 15428 17164 16492 17220
rect 16548 17164 18508 17220
rect 18564 17164 22484 17220
rect 23314 17164 23324 17220
rect 23380 17164 24220 17220
rect 24276 17164 24286 17220
rect 25218 17164 25228 17220
rect 25284 17164 26572 17220
rect 26628 17164 26908 17220
rect 22428 17108 22484 17164
rect 2482 17052 2492 17108
rect 2548 17052 3052 17108
rect 3108 17052 3118 17108
rect 14914 17052 14924 17108
rect 14980 17052 15372 17108
rect 15428 17052 15438 17108
rect 20066 17052 20076 17108
rect 20132 17052 20860 17108
rect 20916 17052 20926 17108
rect 21410 17052 21420 17108
rect 21476 17052 22204 17108
rect 22260 17052 22270 17108
rect 22428 17052 23940 17108
rect 24098 17052 24108 17108
rect 24164 17052 26684 17108
rect 26740 17052 26750 17108
rect 23884 16996 23940 17052
rect 1922 16940 1932 16996
rect 1988 16940 2940 16996
rect 2996 16940 3388 16996
rect 3444 16940 3454 16996
rect 8418 16940 8428 16996
rect 8484 16940 10444 16996
rect 10500 16940 10510 16996
rect 10994 16940 11004 16996
rect 11060 16940 11788 16996
rect 11844 16940 12348 16996
rect 12404 16940 12414 16996
rect 15092 16940 15484 16996
rect 15540 16940 15550 16996
rect 15698 16940 15708 16996
rect 15764 16940 16268 16996
rect 16324 16940 18172 16996
rect 18228 16940 18238 16996
rect 22530 16940 22540 16996
rect 22596 16940 23212 16996
rect 23268 16940 23660 16996
rect 23716 16940 23726 16996
rect 23884 16940 27020 16996
rect 27076 16940 27086 16996
rect 0 16800 800 16912
rect 4610 16828 4620 16884
rect 4676 16828 5404 16884
rect 5460 16828 5740 16884
rect 5796 16828 5806 16884
rect 6178 16828 6188 16884
rect 6244 16828 6972 16884
rect 7028 16828 9548 16884
rect 9604 16828 9614 16884
rect 3266 16716 3276 16772
rect 3332 16716 3948 16772
rect 4004 16716 4014 16772
rect 6066 16716 6076 16772
rect 6132 16716 6860 16772
rect 6916 16716 6926 16772
rect 8082 16716 8092 16772
rect 8148 16716 8596 16772
rect 11218 16716 11228 16772
rect 11284 16716 12124 16772
rect 12180 16716 13244 16772
rect 13300 16716 13310 16772
rect 4722 16604 4732 16660
rect 4788 16604 5852 16660
rect 5908 16604 5918 16660
rect 7746 16604 7756 16660
rect 7812 16604 8316 16660
rect 8372 16604 8382 16660
rect 8540 16548 8596 16716
rect 15092 16660 15148 16940
rect 15586 16828 15596 16884
rect 15652 16828 17052 16884
rect 17108 16828 17612 16884
rect 17668 16828 17678 16884
rect 20402 16828 20412 16884
rect 20468 16828 21644 16884
rect 21700 16828 21710 16884
rect 22642 16828 22652 16884
rect 22708 16828 23324 16884
rect 23380 16828 23772 16884
rect 23828 16828 25452 16884
rect 25508 16828 25518 16884
rect 19282 16716 19292 16772
rect 19348 16716 20188 16772
rect 20244 16716 20254 16772
rect 21074 16716 21084 16772
rect 21140 16716 22316 16772
rect 22372 16716 22382 16772
rect 12674 16604 12684 16660
rect 12740 16604 13580 16660
rect 13636 16604 15148 16660
rect 19506 16604 19516 16660
rect 19572 16604 20748 16660
rect 20804 16604 20814 16660
rect 23734 16604 23772 16660
rect 23828 16604 23838 16660
rect 8540 16492 15148 16548
rect 3998 16436 4008 16492
rect 4064 16436 4112 16492
rect 4168 16436 4216 16492
rect 4272 16436 4320 16492
rect 4376 16436 4424 16492
rect 4480 16436 4528 16492
rect 4584 16436 4632 16492
rect 4688 16436 4736 16492
rect 4792 16436 4840 16492
rect 4896 16436 4944 16492
rect 5000 16436 5048 16492
rect 5104 16436 5152 16492
rect 5208 16436 5218 16492
rect 7410 16380 7420 16436
rect 7476 16380 7868 16436
rect 7924 16380 7934 16436
rect 13318 16380 13356 16436
rect 13412 16380 13422 16436
rect 15092 16324 15148 16492
rect 23998 16436 24008 16492
rect 24064 16436 24112 16492
rect 24168 16436 24216 16492
rect 24272 16436 24320 16492
rect 24376 16436 24424 16492
rect 24480 16436 24528 16492
rect 24584 16436 24632 16492
rect 24688 16436 24736 16492
rect 24792 16436 24840 16492
rect 24896 16436 24944 16492
rect 25000 16436 25048 16492
rect 25104 16436 25152 16492
rect 25208 16436 25218 16492
rect 5954 16268 5964 16324
rect 6020 16268 6030 16324
rect 13458 16268 13468 16324
rect 13524 16268 14028 16324
rect 14084 16268 14094 16324
rect 15092 16268 25788 16324
rect 25844 16268 29372 16324
rect 29428 16268 30380 16324
rect 30436 16268 30446 16324
rect 3938 16156 3948 16212
rect 4004 16156 4732 16212
rect 4788 16156 5404 16212
rect 5460 16156 5470 16212
rect 2594 16044 2604 16100
rect 2660 16044 2670 16100
rect 0 15764 800 15792
rect 2604 15764 2660 16044
rect 4162 15932 4172 15988
rect 4228 15932 5292 15988
rect 5348 15932 5740 15988
rect 5796 15932 5806 15988
rect 0 15708 2660 15764
rect 5964 15764 6020 16268
rect 8642 16156 8652 16212
rect 8708 16156 11228 16212
rect 11284 16156 11294 16212
rect 13234 16156 13244 16212
rect 13300 16156 14700 16212
rect 14756 16156 14766 16212
rect 23762 16156 23772 16212
rect 23828 16156 24556 16212
rect 24612 16156 24622 16212
rect 16706 16044 16716 16100
rect 16772 16044 17612 16100
rect 17668 16044 26796 16100
rect 26852 16044 26862 16100
rect 14018 15932 14028 15988
rect 14084 15932 14588 15988
rect 14644 15932 14654 15988
rect 18050 15932 18060 15988
rect 18116 15932 21644 15988
rect 21700 15932 21710 15988
rect 25106 15932 25116 15988
rect 25172 15932 26684 15988
rect 26740 15932 26750 15988
rect 12226 15820 12236 15876
rect 12292 15820 13132 15876
rect 13188 15820 14140 15876
rect 14196 15820 14206 15876
rect 22642 15820 22652 15876
rect 22708 15820 23884 15876
rect 23940 15820 23950 15876
rect 25302 15820 25340 15876
rect 25396 15820 29036 15876
rect 29092 15820 29102 15876
rect 5964 15708 10500 15764
rect 0 15680 800 15708
rect 4722 15596 4732 15652
rect 4788 15596 6188 15652
rect 6244 15596 6254 15652
rect 10444 15540 10500 15708
rect 13998 15652 14008 15708
rect 14064 15652 14112 15708
rect 14168 15652 14216 15708
rect 14272 15652 14320 15708
rect 14376 15652 14424 15708
rect 14480 15652 14528 15708
rect 14584 15652 14632 15708
rect 14688 15652 14736 15708
rect 14792 15652 14840 15708
rect 14896 15652 14944 15708
rect 15000 15652 15048 15708
rect 15104 15652 15152 15708
rect 15208 15652 15218 15708
rect 33998 15652 34008 15708
rect 34064 15652 34112 15708
rect 34168 15652 34216 15708
rect 34272 15652 34320 15708
rect 34376 15652 34424 15708
rect 34480 15652 34528 15708
rect 34584 15652 34632 15708
rect 34688 15652 34736 15708
rect 34792 15652 34840 15708
rect 34896 15652 34944 15708
rect 35000 15652 35048 15708
rect 35104 15652 35152 15708
rect 35208 15652 35218 15708
rect 5842 15484 5852 15540
rect 5908 15484 6412 15540
rect 6468 15484 7308 15540
rect 7364 15484 7374 15540
rect 7522 15484 7532 15540
rect 7588 15484 9660 15540
rect 9716 15484 9726 15540
rect 10444 15484 22204 15540
rect 22260 15484 22988 15540
rect 23044 15484 23054 15540
rect 28466 15484 28476 15540
rect 28532 15484 29260 15540
rect 29316 15484 29326 15540
rect 6066 15372 6076 15428
rect 6132 15372 7196 15428
rect 7252 15372 7262 15428
rect 9538 15372 9548 15428
rect 9604 15372 11564 15428
rect 11620 15372 11630 15428
rect 13906 15372 13916 15428
rect 13972 15372 15708 15428
rect 15764 15372 15774 15428
rect 18722 15260 18732 15316
rect 18788 15260 22316 15316
rect 22372 15260 22382 15316
rect 25554 15260 25564 15316
rect 25620 15260 27580 15316
rect 27636 15260 28252 15316
rect 28308 15260 29932 15316
rect 29988 15260 29998 15316
rect 1810 15148 1820 15204
rect 1876 15148 5628 15204
rect 5684 15148 5694 15204
rect 13458 15148 13468 15204
rect 13524 15148 14364 15204
rect 14420 15148 14430 15204
rect 20514 15148 20524 15204
rect 20580 15148 21756 15204
rect 21812 15148 22204 15204
rect 22260 15148 22270 15204
rect 6962 15036 6972 15092
rect 7028 15036 8764 15092
rect 8820 15036 8830 15092
rect 23772 15036 24220 15092
rect 24276 15036 24286 15092
rect 24434 15036 24444 15092
rect 24500 15036 26908 15092
rect 26964 15036 26974 15092
rect 23772 14980 23828 15036
rect 8866 14924 8876 14980
rect 8932 14924 9100 14980
rect 9156 14924 10556 14980
rect 10612 14924 11452 14980
rect 11508 14924 12348 14980
rect 12404 14924 12796 14980
rect 12852 14924 13356 14980
rect 13412 14924 16716 14980
rect 16772 14924 16782 14980
rect 23762 14924 23772 14980
rect 23828 14924 23838 14980
rect 3998 14868 4008 14924
rect 4064 14868 4112 14924
rect 4168 14868 4216 14924
rect 4272 14868 4320 14924
rect 4376 14868 4424 14924
rect 4480 14868 4528 14924
rect 4584 14868 4632 14924
rect 4688 14868 4736 14924
rect 4792 14868 4840 14924
rect 4896 14868 4944 14924
rect 5000 14868 5048 14924
rect 5104 14868 5152 14924
rect 5208 14868 5218 14924
rect 23998 14868 24008 14924
rect 24064 14868 24112 14924
rect 24168 14868 24216 14924
rect 24272 14868 24320 14924
rect 24376 14868 24424 14924
rect 24480 14868 24528 14924
rect 24584 14868 24632 14924
rect 24688 14868 24736 14924
rect 24792 14868 24840 14924
rect 24896 14868 24944 14924
rect 25000 14868 25048 14924
rect 25104 14868 25152 14924
rect 25208 14868 25218 14924
rect 3154 14700 3164 14756
rect 3220 14700 4060 14756
rect 4116 14700 4126 14756
rect 6514 14700 6524 14756
rect 6580 14700 15148 14756
rect 17154 14700 17164 14756
rect 17220 14700 18172 14756
rect 18228 14700 20692 14756
rect 0 14644 800 14672
rect 15092 14644 15148 14700
rect 20636 14644 20692 14700
rect 0 14588 1708 14644
rect 1764 14588 1774 14644
rect 11442 14588 11452 14644
rect 11508 14588 13132 14644
rect 13188 14588 13198 14644
rect 15092 14588 18620 14644
rect 18676 14588 19852 14644
rect 19908 14588 19918 14644
rect 20626 14588 20636 14644
rect 20692 14588 21980 14644
rect 22036 14588 23212 14644
rect 23268 14588 23278 14644
rect 0 14560 800 14588
rect 5954 14476 5964 14532
rect 6020 14476 8428 14532
rect 8484 14476 8494 14532
rect 9986 14476 9996 14532
rect 10052 14476 10556 14532
rect 10612 14476 11116 14532
rect 11172 14476 11900 14532
rect 11956 14476 12348 14532
rect 12404 14476 15372 14532
rect 15428 14476 15438 14532
rect 4722 14364 4732 14420
rect 4788 14364 6412 14420
rect 6468 14364 6478 14420
rect 7186 14364 7196 14420
rect 7252 14364 8204 14420
rect 8260 14364 8270 14420
rect 8754 14364 8764 14420
rect 8820 14364 9548 14420
rect 9604 14364 9614 14420
rect 17602 14364 17612 14420
rect 17668 14364 18956 14420
rect 19012 14364 19022 14420
rect 5730 14252 5740 14308
rect 5796 14252 6188 14308
rect 6244 14252 6254 14308
rect 19506 14252 19516 14308
rect 19572 14252 20972 14308
rect 21028 14252 21038 14308
rect 27906 14252 27916 14308
rect 27972 14252 28476 14308
rect 28532 14252 28542 14308
rect 13998 14084 14008 14140
rect 14064 14084 14112 14140
rect 14168 14084 14216 14140
rect 14272 14084 14320 14140
rect 14376 14084 14424 14140
rect 14480 14084 14528 14140
rect 14584 14084 14632 14140
rect 14688 14084 14736 14140
rect 14792 14084 14840 14140
rect 14896 14084 14944 14140
rect 15000 14084 15048 14140
rect 15104 14084 15152 14140
rect 15208 14084 15218 14140
rect 33998 14084 34008 14140
rect 34064 14084 34112 14140
rect 34168 14084 34216 14140
rect 34272 14084 34320 14140
rect 34376 14084 34424 14140
rect 34480 14084 34528 14140
rect 34584 14084 34632 14140
rect 34688 14084 34736 14140
rect 34792 14084 34840 14140
rect 34896 14084 34944 14140
rect 35000 14084 35048 14140
rect 35104 14084 35152 14140
rect 35208 14084 35218 14140
rect 3602 13916 3612 13972
rect 3668 13916 3836 13972
rect 3892 13916 3902 13972
rect 9090 13916 9100 13972
rect 9156 13916 9884 13972
rect 9940 13916 11228 13972
rect 11284 13916 11294 13972
rect 11732 13916 12348 13972
rect 12404 13916 13468 13972
rect 13524 13916 13534 13972
rect 9538 13804 9548 13860
rect 9604 13804 10780 13860
rect 10836 13804 10846 13860
rect 6962 13692 6972 13748
rect 7028 13692 7196 13748
rect 7252 13692 7756 13748
rect 7812 13692 8596 13748
rect 8540 13636 8596 13692
rect 11732 13636 11788 13916
rect 16818 13804 16828 13860
rect 16884 13804 18060 13860
rect 18116 13804 20188 13860
rect 20244 13804 21196 13860
rect 21252 13804 22428 13860
rect 22484 13804 22494 13860
rect 12450 13692 12460 13748
rect 12516 13692 13244 13748
rect 13300 13692 14252 13748
rect 14308 13692 14318 13748
rect 14802 13692 14812 13748
rect 14868 13692 15372 13748
rect 15428 13692 15438 13748
rect 24658 13692 24668 13748
rect 24724 13692 26908 13748
rect 26964 13692 27916 13748
rect 27972 13692 27982 13748
rect 7074 13580 7084 13636
rect 7140 13580 8204 13636
rect 8260 13580 8270 13636
rect 8530 13580 8540 13636
rect 8596 13580 9212 13636
rect 9268 13580 9548 13636
rect 9604 13580 11452 13636
rect 11508 13580 11788 13636
rect 26114 13580 26124 13636
rect 26180 13580 26684 13636
rect 26740 13580 26750 13636
rect 0 13524 800 13552
rect 0 13468 1932 13524
rect 1988 13468 1998 13524
rect 10098 13468 10108 13524
rect 10164 13468 15260 13524
rect 15316 13468 16044 13524
rect 16100 13468 16110 13524
rect 26450 13468 26460 13524
rect 26516 13468 26796 13524
rect 26852 13468 26862 13524
rect 0 13440 800 13468
rect 3998 13300 4008 13356
rect 4064 13300 4112 13356
rect 4168 13300 4216 13356
rect 4272 13300 4320 13356
rect 4376 13300 4424 13356
rect 4480 13300 4528 13356
rect 4584 13300 4632 13356
rect 4688 13300 4736 13356
rect 4792 13300 4840 13356
rect 4896 13300 4944 13356
rect 5000 13300 5048 13356
rect 5104 13300 5152 13356
rect 5208 13300 5218 13356
rect 23998 13300 24008 13356
rect 24064 13300 24112 13356
rect 24168 13300 24216 13356
rect 24272 13300 24320 13356
rect 24376 13300 24424 13356
rect 24480 13300 24528 13356
rect 24584 13300 24632 13356
rect 24688 13300 24736 13356
rect 24792 13300 24840 13356
rect 24896 13300 24944 13356
rect 25000 13300 25048 13356
rect 25104 13300 25152 13356
rect 25208 13300 25218 13356
rect 14914 13132 14924 13188
rect 14980 13132 15820 13188
rect 15876 13132 15886 13188
rect 23762 13132 23772 13188
rect 23828 13132 24556 13188
rect 24612 13132 24622 13188
rect 26852 13132 27356 13188
rect 27412 13132 27422 13188
rect 26852 13076 26908 13132
rect 4274 13020 4284 13076
rect 4340 13020 4844 13076
rect 4900 13020 5404 13076
rect 5460 13020 5470 13076
rect 6514 13020 6524 13076
rect 6580 13020 7196 13076
rect 7252 13020 10444 13076
rect 10500 13020 11676 13076
rect 11732 13020 11742 13076
rect 22418 13020 22428 13076
rect 22484 13020 23436 13076
rect 23492 13020 23502 13076
rect 26562 13020 26572 13076
rect 26628 13020 26908 13076
rect 15586 12908 15596 12964
rect 15652 12908 16380 12964
rect 16436 12908 16446 12964
rect 21746 12908 21756 12964
rect 21812 12908 23212 12964
rect 23268 12908 24444 12964
rect 24500 12908 24510 12964
rect 8754 12796 8764 12852
rect 8820 12796 9772 12852
rect 9828 12796 9838 12852
rect 12898 12796 12908 12852
rect 12964 12796 13692 12852
rect 13748 12796 14364 12852
rect 14420 12796 14430 12852
rect 23986 12796 23996 12852
rect 24052 12796 25788 12852
rect 25844 12796 25854 12852
rect 8194 12684 8204 12740
rect 8260 12684 9100 12740
rect 9156 12684 9166 12740
rect 13804 12684 14588 12740
rect 14644 12684 14654 12740
rect 15250 12684 15260 12740
rect 15316 12684 15596 12740
rect 15652 12684 15662 12740
rect 19170 12684 19180 12740
rect 19236 12684 20300 12740
rect 20356 12684 21308 12740
rect 21364 12684 21374 12740
rect 0 12320 800 12432
rect 13804 12404 13860 12684
rect 13998 12516 14008 12572
rect 14064 12516 14112 12572
rect 14168 12516 14216 12572
rect 14272 12516 14320 12572
rect 14376 12516 14424 12572
rect 14480 12516 14528 12572
rect 14584 12516 14632 12572
rect 14688 12516 14736 12572
rect 14792 12516 14840 12572
rect 14896 12516 14944 12572
rect 15000 12516 15048 12572
rect 15104 12516 15152 12572
rect 15208 12516 15218 12572
rect 33998 12516 34008 12572
rect 34064 12516 34112 12572
rect 34168 12516 34216 12572
rect 34272 12516 34320 12572
rect 34376 12516 34424 12572
rect 34480 12516 34528 12572
rect 34584 12516 34632 12572
rect 34688 12516 34736 12572
rect 34792 12516 34840 12572
rect 34896 12516 34944 12572
rect 35000 12516 35048 12572
rect 35104 12516 35152 12572
rect 35208 12516 35218 12572
rect 4834 12348 4844 12404
rect 4900 12348 5740 12404
rect 5796 12348 5806 12404
rect 6066 12348 6076 12404
rect 6132 12348 6748 12404
rect 6804 12348 6814 12404
rect 8978 12348 8988 12404
rect 9044 12348 10332 12404
rect 10388 12348 10892 12404
rect 10948 12348 10958 12404
rect 13804 12348 14588 12404
rect 14644 12348 14654 12404
rect 16706 12348 16716 12404
rect 16772 12348 17500 12404
rect 17556 12348 17566 12404
rect 27346 12348 27356 12404
rect 27412 12348 28252 12404
rect 28308 12348 28318 12404
rect 6850 12236 6860 12292
rect 6916 12236 7420 12292
rect 7476 12236 7486 12292
rect 4050 12124 4060 12180
rect 4116 12124 5292 12180
rect 5348 12124 10220 12180
rect 10276 12124 10286 12180
rect 19842 12124 19852 12180
rect 19908 12124 22540 12180
rect 22596 12124 22606 12180
rect 5506 12012 5516 12068
rect 5572 12012 7084 12068
rect 7140 12012 7150 12068
rect 7298 12012 7308 12068
rect 7364 12012 8988 12068
rect 9044 12012 9054 12068
rect 17938 12012 17948 12068
rect 18004 12012 19180 12068
rect 19236 12012 19246 12068
rect 6962 11900 6972 11956
rect 7028 11900 8316 11956
rect 8372 11900 8382 11956
rect 13570 11788 13580 11844
rect 13636 11788 15484 11844
rect 15540 11788 15550 11844
rect 3998 11732 4008 11788
rect 4064 11732 4112 11788
rect 4168 11732 4216 11788
rect 4272 11732 4320 11788
rect 4376 11732 4424 11788
rect 4480 11732 4528 11788
rect 4584 11732 4632 11788
rect 4688 11732 4736 11788
rect 4792 11732 4840 11788
rect 4896 11732 4944 11788
rect 5000 11732 5048 11788
rect 5104 11732 5152 11788
rect 5208 11732 5218 11788
rect 23998 11732 24008 11788
rect 24064 11732 24112 11788
rect 24168 11732 24216 11788
rect 24272 11732 24320 11788
rect 24376 11732 24424 11788
rect 24480 11732 24528 11788
rect 24584 11732 24632 11788
rect 24688 11732 24736 11788
rect 24792 11732 24840 11788
rect 24896 11732 24944 11788
rect 25000 11732 25048 11788
rect 25104 11732 25152 11788
rect 25208 11732 25218 11788
rect 2370 11564 2380 11620
rect 2436 11564 3388 11620
rect 3444 11564 3454 11620
rect 13234 11564 13244 11620
rect 13300 11564 13916 11620
rect 13972 11564 13982 11620
rect 4386 11452 4396 11508
rect 4452 11452 5068 11508
rect 5124 11452 5404 11508
rect 5460 11452 5470 11508
rect 25442 11452 25452 11508
rect 25508 11452 26124 11508
rect 26180 11452 26684 11508
rect 26740 11452 26750 11508
rect 4498 11340 4508 11396
rect 4564 11340 5404 11396
rect 5460 11340 6860 11396
rect 6916 11340 6926 11396
rect 0 11200 800 11312
rect 16370 11228 16380 11284
rect 16436 11228 17836 11284
rect 17892 11228 17902 11284
rect 5730 11116 5740 11172
rect 5796 11116 7980 11172
rect 8036 11116 8876 11172
rect 8932 11116 9660 11172
rect 9716 11116 12012 11172
rect 12068 11116 12078 11172
rect 14578 11116 14588 11172
rect 14644 11116 17052 11172
rect 17108 11116 17118 11172
rect 10882 11004 10892 11060
rect 10948 11004 12460 11060
rect 12516 11004 13244 11060
rect 13300 11004 13310 11060
rect 13998 10948 14008 11004
rect 14064 10948 14112 11004
rect 14168 10948 14216 11004
rect 14272 10948 14320 11004
rect 14376 10948 14424 11004
rect 14480 10948 14528 11004
rect 14584 10948 14632 11004
rect 14688 10948 14736 11004
rect 14792 10948 14840 11004
rect 14896 10948 14944 11004
rect 15000 10948 15048 11004
rect 15104 10948 15152 11004
rect 15208 10948 15218 11004
rect 15372 10836 15428 11116
rect 33998 10948 34008 11004
rect 34064 10948 34112 11004
rect 34168 10948 34216 11004
rect 34272 10948 34320 11004
rect 34376 10948 34424 11004
rect 34480 10948 34528 11004
rect 34584 10948 34632 11004
rect 34688 10948 34736 11004
rect 34792 10948 34840 11004
rect 34896 10948 34944 11004
rect 35000 10948 35048 11004
rect 35104 10948 35152 11004
rect 35208 10948 35218 11004
rect 4722 10780 4732 10836
rect 4788 10780 5964 10836
rect 6020 10780 6030 10836
rect 13234 10780 13244 10836
rect 13300 10780 14588 10836
rect 14644 10780 14654 10836
rect 15138 10780 15148 10836
rect 15204 10780 15428 10836
rect 22530 10780 22540 10836
rect 22596 10780 23660 10836
rect 23716 10780 25004 10836
rect 25060 10780 25070 10836
rect 14588 10388 14644 10780
rect 19730 10668 19740 10724
rect 19796 10668 22316 10724
rect 22372 10668 23996 10724
rect 24052 10668 26572 10724
rect 26628 10668 26638 10724
rect 14588 10332 15596 10388
rect 15652 10332 16380 10388
rect 16436 10332 16446 10388
rect 0 10080 800 10192
rect 3998 10164 4008 10220
rect 4064 10164 4112 10220
rect 4168 10164 4216 10220
rect 4272 10164 4320 10220
rect 4376 10164 4424 10220
rect 4480 10164 4528 10220
rect 4584 10164 4632 10220
rect 4688 10164 4736 10220
rect 4792 10164 4840 10220
rect 4896 10164 4944 10220
rect 5000 10164 5048 10220
rect 5104 10164 5152 10220
rect 5208 10164 5218 10220
rect 23998 10164 24008 10220
rect 24064 10164 24112 10220
rect 24168 10164 24216 10220
rect 24272 10164 24320 10220
rect 24376 10164 24424 10220
rect 24480 10164 24528 10220
rect 24584 10164 24632 10220
rect 24688 10164 24736 10220
rect 24792 10164 24840 10220
rect 24896 10164 24944 10220
rect 25000 10164 25048 10220
rect 25104 10164 25152 10220
rect 25208 10164 25218 10220
rect 9202 10108 9212 10164
rect 9268 10108 10892 10164
rect 10948 10108 10958 10164
rect 25778 9884 25788 9940
rect 25844 9884 27020 9940
rect 27076 9884 27086 9940
rect 25890 9660 25900 9716
rect 25956 9660 28028 9716
rect 28084 9660 28094 9716
rect 13998 9380 14008 9436
rect 14064 9380 14112 9436
rect 14168 9380 14216 9436
rect 14272 9380 14320 9436
rect 14376 9380 14424 9436
rect 14480 9380 14528 9436
rect 14584 9380 14632 9436
rect 14688 9380 14736 9436
rect 14792 9380 14840 9436
rect 14896 9380 14944 9436
rect 15000 9380 15048 9436
rect 15104 9380 15152 9436
rect 15208 9380 15218 9436
rect 33998 9380 34008 9436
rect 34064 9380 34112 9436
rect 34168 9380 34216 9436
rect 34272 9380 34320 9436
rect 34376 9380 34424 9436
rect 34480 9380 34528 9436
rect 34584 9380 34632 9436
rect 34688 9380 34736 9436
rect 34792 9380 34840 9436
rect 34896 9380 34944 9436
rect 35000 9380 35048 9436
rect 35104 9380 35152 9436
rect 35208 9380 35218 9436
rect 28242 9100 28252 9156
rect 28308 9100 29036 9156
rect 29092 9100 29102 9156
rect 0 8960 800 9072
rect 25330 8988 25340 9044
rect 25396 8988 28364 9044
rect 28420 8988 29596 9044
rect 29652 8988 29662 9044
rect 3998 8596 4008 8652
rect 4064 8596 4112 8652
rect 4168 8596 4216 8652
rect 4272 8596 4320 8652
rect 4376 8596 4424 8652
rect 4480 8596 4528 8652
rect 4584 8596 4632 8652
rect 4688 8596 4736 8652
rect 4792 8596 4840 8652
rect 4896 8596 4944 8652
rect 5000 8596 5048 8652
rect 5104 8596 5152 8652
rect 5208 8596 5218 8652
rect 23998 8596 24008 8652
rect 24064 8596 24112 8652
rect 24168 8596 24216 8652
rect 24272 8596 24320 8652
rect 24376 8596 24424 8652
rect 24480 8596 24528 8652
rect 24584 8596 24632 8652
rect 24688 8596 24736 8652
rect 24792 8596 24840 8652
rect 24896 8596 24944 8652
rect 25000 8596 25048 8652
rect 25104 8596 25152 8652
rect 25208 8596 25218 8652
rect 17602 8428 17612 8484
rect 17668 8428 19404 8484
rect 19460 8428 19470 8484
rect 6066 8316 6076 8372
rect 6132 8316 7308 8372
rect 7364 8316 7980 8372
rect 8036 8316 9212 8372
rect 9268 8316 9278 8372
rect 18946 8316 18956 8372
rect 19012 8316 19740 8372
rect 19796 8316 19806 8372
rect 18610 8204 18620 8260
rect 18676 8204 19516 8260
rect 19572 8204 21196 8260
rect 21252 8204 21262 8260
rect 18050 8092 18060 8148
rect 18116 8092 18732 8148
rect 18788 8092 19964 8148
rect 20020 8092 20030 8148
rect 3490 7980 3500 8036
rect 3556 7980 5404 8036
rect 5460 7980 5852 8036
rect 5908 7980 6636 8036
rect 6692 7980 6702 8036
rect 19506 7980 19516 8036
rect 19572 7980 20300 8036
rect 20356 7980 20366 8036
rect 0 7840 800 7952
rect 13998 7812 14008 7868
rect 14064 7812 14112 7868
rect 14168 7812 14216 7868
rect 14272 7812 14320 7868
rect 14376 7812 14424 7868
rect 14480 7812 14528 7868
rect 14584 7812 14632 7868
rect 14688 7812 14736 7868
rect 14792 7812 14840 7868
rect 14896 7812 14944 7868
rect 15000 7812 15048 7868
rect 15104 7812 15152 7868
rect 15208 7812 15218 7868
rect 33998 7812 34008 7868
rect 34064 7812 34112 7868
rect 34168 7812 34216 7868
rect 34272 7812 34320 7868
rect 34376 7812 34424 7868
rect 34480 7812 34528 7868
rect 34584 7812 34632 7868
rect 34688 7812 34736 7868
rect 34792 7812 34840 7868
rect 34896 7812 34944 7868
rect 35000 7812 35048 7868
rect 35104 7812 35152 7868
rect 35208 7812 35218 7868
rect 25330 7756 25340 7812
rect 25396 7756 26348 7812
rect 26404 7756 26908 7812
rect 26964 7756 27580 7812
rect 27636 7756 28140 7812
rect 28196 7756 28206 7812
rect 4722 7644 4732 7700
rect 4788 7644 6076 7700
rect 6132 7644 6142 7700
rect 16818 7644 16828 7700
rect 16884 7644 19292 7700
rect 19348 7644 19358 7700
rect 19730 7644 19740 7700
rect 19796 7644 21420 7700
rect 21476 7644 21486 7700
rect 20066 7532 20076 7588
rect 20132 7532 20636 7588
rect 20692 7532 26012 7588
rect 26068 7532 26078 7588
rect 6738 7420 6748 7476
rect 6804 7420 7532 7476
rect 7588 7420 7980 7476
rect 8036 7420 8046 7476
rect 13570 7420 13580 7476
rect 13636 7420 14588 7476
rect 14644 7420 15148 7476
rect 15204 7420 15214 7476
rect 5506 7308 5516 7364
rect 5572 7308 6636 7364
rect 6692 7308 6702 7364
rect 6850 7308 6860 7364
rect 6916 7308 7644 7364
rect 7700 7308 7710 7364
rect 7970 7196 7980 7252
rect 8036 7196 8428 7252
rect 8484 7196 8494 7252
rect 24658 7196 24668 7252
rect 24724 7196 25676 7252
rect 25732 7196 25742 7252
rect 3998 7028 4008 7084
rect 4064 7028 4112 7084
rect 4168 7028 4216 7084
rect 4272 7028 4320 7084
rect 4376 7028 4424 7084
rect 4480 7028 4528 7084
rect 4584 7028 4632 7084
rect 4688 7028 4736 7084
rect 4792 7028 4840 7084
rect 4896 7028 4944 7084
rect 5000 7028 5048 7084
rect 5104 7028 5152 7084
rect 5208 7028 5218 7084
rect 23998 7028 24008 7084
rect 24064 7028 24112 7084
rect 24168 7028 24216 7084
rect 24272 7028 24320 7084
rect 24376 7028 24424 7084
rect 24480 7028 24528 7084
rect 24584 7028 24632 7084
rect 24688 7028 24736 7084
rect 24792 7028 24840 7084
rect 24896 7028 24944 7084
rect 25000 7028 25048 7084
rect 25104 7028 25152 7084
rect 25208 7028 25218 7084
rect 3332 6860 3500 6916
rect 3556 6860 3566 6916
rect 4162 6860 4172 6916
rect 4228 6860 5628 6916
rect 5684 6860 5694 6916
rect 8082 6860 8092 6916
rect 8148 6860 8540 6916
rect 8596 6860 8606 6916
rect 8754 6860 8764 6916
rect 8820 6860 9772 6916
rect 9828 6860 9838 6916
rect 20290 6860 20300 6916
rect 20356 6860 21308 6916
rect 21364 6860 21374 6916
rect 0 6720 800 6832
rect 3332 6692 3388 6860
rect 3602 6748 3612 6804
rect 3668 6748 4508 6804
rect 4564 6748 4574 6804
rect 4722 6748 4732 6804
rect 4788 6748 6300 6804
rect 6356 6748 6366 6804
rect 14242 6748 14252 6804
rect 14308 6748 15036 6804
rect 15092 6748 15102 6804
rect 2482 6636 2492 6692
rect 2548 6636 3388 6692
rect 4050 6636 4060 6692
rect 4116 6636 5292 6692
rect 5348 6636 5358 6692
rect 6738 6636 6748 6692
rect 6804 6636 7756 6692
rect 7812 6636 7822 6692
rect 9986 6636 9996 6692
rect 10052 6636 13244 6692
rect 13300 6636 16716 6692
rect 16772 6636 16782 6692
rect 21074 6636 21084 6692
rect 21140 6636 22092 6692
rect 22148 6636 25340 6692
rect 25396 6636 25406 6692
rect 3042 6412 3052 6468
rect 3108 6412 3118 6468
rect 3052 6356 3108 6412
rect 4060 6356 4116 6636
rect 6402 6524 6412 6580
rect 6468 6524 7980 6580
rect 8036 6524 8316 6580
rect 8372 6524 8382 6580
rect 13010 6524 13020 6580
rect 13076 6524 13916 6580
rect 13972 6524 13982 6580
rect 16818 6524 16828 6580
rect 16884 6524 18060 6580
rect 18116 6524 18126 6580
rect 25554 6524 25564 6580
rect 25620 6524 27804 6580
rect 27860 6524 27870 6580
rect 5730 6412 5740 6468
rect 5796 6412 7532 6468
rect 7588 6412 7598 6468
rect 16482 6412 16492 6468
rect 16548 6412 17500 6468
rect 17556 6412 17566 6468
rect 26002 6412 26012 6468
rect 26068 6412 29820 6468
rect 29876 6412 29886 6468
rect 3052 6300 4116 6356
rect 13998 6244 14008 6300
rect 14064 6244 14112 6300
rect 14168 6244 14216 6300
rect 14272 6244 14320 6300
rect 14376 6244 14424 6300
rect 14480 6244 14528 6300
rect 14584 6244 14632 6300
rect 14688 6244 14736 6300
rect 14792 6244 14840 6300
rect 14896 6244 14944 6300
rect 15000 6244 15048 6300
rect 15104 6244 15152 6300
rect 15208 6244 15218 6300
rect 33998 6244 34008 6300
rect 34064 6244 34112 6300
rect 34168 6244 34216 6300
rect 34272 6244 34320 6300
rect 34376 6244 34424 6300
rect 34480 6244 34528 6300
rect 34584 6244 34632 6300
rect 34688 6244 34736 6300
rect 34792 6244 34840 6300
rect 34896 6244 34944 6300
rect 35000 6244 35048 6300
rect 35104 6244 35152 6300
rect 35208 6244 35218 6300
rect 8530 6076 8540 6132
rect 8596 6076 8932 6132
rect 18610 6076 18620 6132
rect 18676 6076 20188 6132
rect 20244 6076 20748 6132
rect 20804 6076 21532 6132
rect 21588 6076 21598 6132
rect 27010 6076 27020 6132
rect 27076 6076 28812 6132
rect 28868 6076 28878 6132
rect 2146 5964 2156 6020
rect 2212 5964 3500 6020
rect 3556 5964 3566 6020
rect 8876 5908 8932 6076
rect 6738 5852 6748 5908
rect 6804 5852 8428 5908
rect 8484 5852 8494 5908
rect 8866 5852 8876 5908
rect 8932 5852 8942 5908
rect 9090 5852 9100 5908
rect 9156 5852 9996 5908
rect 10052 5852 10062 5908
rect 16370 5852 16380 5908
rect 16436 5852 17276 5908
rect 17332 5852 17342 5908
rect 24322 5852 24332 5908
rect 24388 5852 26012 5908
rect 26068 5852 26078 5908
rect 3602 5740 3612 5796
rect 3668 5740 5964 5796
rect 6020 5740 6030 5796
rect 7522 5740 7532 5796
rect 7588 5740 8540 5796
rect 8596 5740 11116 5796
rect 11172 5740 11182 5796
rect 0 5684 800 5712
rect 0 5628 2044 5684
rect 2100 5628 2828 5684
rect 2884 5628 2894 5684
rect 8306 5628 8316 5684
rect 8372 5628 8764 5684
rect 8820 5628 8830 5684
rect 9202 5628 9212 5684
rect 9268 5628 10108 5684
rect 10164 5628 13132 5684
rect 13188 5628 13198 5684
rect 0 5600 800 5628
rect 3998 5460 4008 5516
rect 4064 5460 4112 5516
rect 4168 5460 4216 5516
rect 4272 5460 4320 5516
rect 4376 5460 4424 5516
rect 4480 5460 4528 5516
rect 4584 5460 4632 5516
rect 4688 5460 4736 5516
rect 4792 5460 4840 5516
rect 4896 5460 4944 5516
rect 5000 5460 5048 5516
rect 5104 5460 5152 5516
rect 5208 5460 5218 5516
rect 23998 5460 24008 5516
rect 24064 5460 24112 5516
rect 24168 5460 24216 5516
rect 24272 5460 24320 5516
rect 24376 5460 24424 5516
rect 24480 5460 24528 5516
rect 24584 5460 24632 5516
rect 24688 5460 24736 5516
rect 24792 5460 24840 5516
rect 24896 5460 24944 5516
rect 25000 5460 25048 5516
rect 25104 5460 25152 5516
rect 25208 5460 25218 5516
rect 9100 5180 11340 5236
rect 11396 5180 11900 5236
rect 11956 5180 13580 5236
rect 13636 5180 14028 5236
rect 14084 5180 14094 5236
rect 5282 5068 5292 5124
rect 5348 5068 6076 5124
rect 6132 5068 6142 5124
rect 9100 5012 9156 5180
rect 9314 5068 9324 5124
rect 9380 5068 10332 5124
rect 10388 5068 10892 5124
rect 10948 5068 10958 5124
rect 20402 5068 20412 5124
rect 20468 5068 22316 5124
rect 22372 5068 22382 5124
rect 4722 4956 4732 5012
rect 4788 4956 6636 5012
rect 6692 4956 7308 5012
rect 7364 4956 7532 5012
rect 7588 4956 9156 5012
rect 13234 4956 13244 5012
rect 13300 4956 15372 5012
rect 15428 4956 16828 5012
rect 16884 4956 16894 5012
rect 13794 4844 13804 4900
rect 13860 4844 16436 4900
rect 13998 4676 14008 4732
rect 14064 4676 14112 4732
rect 14168 4676 14216 4732
rect 14272 4676 14320 4732
rect 14376 4676 14424 4732
rect 14480 4676 14528 4732
rect 14584 4676 14632 4732
rect 14688 4676 14736 4732
rect 14792 4676 14840 4732
rect 14896 4676 14944 4732
rect 15000 4676 15048 4732
rect 15104 4676 15152 4732
rect 15208 4676 15218 4732
rect 0 4480 800 4592
rect 16380 4564 16436 4844
rect 33998 4676 34008 4732
rect 34064 4676 34112 4732
rect 34168 4676 34216 4732
rect 34272 4676 34320 4732
rect 34376 4676 34424 4732
rect 34480 4676 34528 4732
rect 34584 4676 34632 4732
rect 34688 4676 34736 4732
rect 34792 4676 34840 4732
rect 34896 4676 34944 4732
rect 35000 4676 35048 4732
rect 35104 4676 35152 4732
rect 35208 4676 35218 4732
rect 12562 4508 12572 4564
rect 12628 4508 13804 4564
rect 13860 4508 13870 4564
rect 16370 4508 16380 4564
rect 16436 4508 20076 4564
rect 20132 4508 20142 4564
rect 18050 4396 18060 4452
rect 18116 4396 19068 4452
rect 19124 4396 23996 4452
rect 24052 4396 24062 4452
rect 24770 4396 24780 4452
rect 24836 4396 25900 4452
rect 25956 4396 25966 4452
rect 1922 4284 1932 4340
rect 1988 4284 3836 4340
rect 3892 4284 5964 4340
rect 6020 4284 6030 4340
rect 9650 4284 9660 4340
rect 9716 4284 13244 4340
rect 13300 4284 13310 4340
rect 13122 4060 13132 4116
rect 13188 4060 17948 4116
rect 18004 4060 18014 4116
rect 25442 4060 25452 4116
rect 25508 4060 26572 4116
rect 26628 4060 26638 4116
rect 16930 3948 16940 4004
rect 16996 3948 18172 4004
rect 18228 3948 19852 4004
rect 19908 3948 19918 4004
rect 3998 3892 4008 3948
rect 4064 3892 4112 3948
rect 4168 3892 4216 3948
rect 4272 3892 4320 3948
rect 4376 3892 4424 3948
rect 4480 3892 4528 3948
rect 4584 3892 4632 3948
rect 4688 3892 4736 3948
rect 4792 3892 4840 3948
rect 4896 3892 4944 3948
rect 5000 3892 5048 3948
rect 5104 3892 5152 3948
rect 5208 3892 5218 3948
rect 23998 3892 24008 3948
rect 24064 3892 24112 3948
rect 24168 3892 24216 3948
rect 24272 3892 24320 3948
rect 24376 3892 24424 3948
rect 24480 3892 24528 3948
rect 24584 3892 24632 3948
rect 24688 3892 24736 3948
rect 24792 3892 24840 3948
rect 24896 3892 24944 3948
rect 25000 3892 25048 3948
rect 25104 3892 25152 3948
rect 25208 3892 25218 3948
rect 17266 3724 17276 3780
rect 17332 3724 20860 3780
rect 20916 3724 20926 3780
rect 5954 3612 5964 3668
rect 6020 3612 8316 3668
rect 8372 3612 9324 3668
rect 9380 3612 9390 3668
rect 13906 3612 13916 3668
rect 13972 3612 16940 3668
rect 16996 3612 17006 3668
rect 15092 3500 25452 3556
rect 25508 3500 25518 3556
rect 15092 3444 15148 3500
rect 9874 3388 9884 3444
rect 9940 3388 13244 3444
rect 13300 3388 13692 3444
rect 13748 3388 15148 3444
rect 16146 3388 16156 3444
rect 16212 3388 18732 3444
rect 18788 3388 18798 3444
rect 13998 3108 14008 3164
rect 14064 3108 14112 3164
rect 14168 3108 14216 3164
rect 14272 3108 14320 3164
rect 14376 3108 14424 3164
rect 14480 3108 14528 3164
rect 14584 3108 14632 3164
rect 14688 3108 14736 3164
rect 14792 3108 14840 3164
rect 14896 3108 14944 3164
rect 15000 3108 15048 3164
rect 15104 3108 15152 3164
rect 15208 3108 15218 3164
rect 33998 3108 34008 3164
rect 34064 3108 34112 3164
rect 34168 3108 34216 3164
rect 34272 3108 34320 3164
rect 34376 3108 34424 3164
rect 34480 3108 34528 3164
rect 34584 3108 34632 3164
rect 34688 3108 34736 3164
rect 34792 3108 34840 3164
rect 34896 3108 34944 3164
rect 35000 3108 35048 3164
rect 35104 3108 35152 3164
rect 35208 3108 35218 3164
<< via3 >>
rect 4008 96404 4064 96460
rect 4112 96404 4168 96460
rect 4216 96404 4272 96460
rect 4320 96404 4376 96460
rect 4424 96404 4480 96460
rect 4528 96404 4584 96460
rect 4632 96404 4688 96460
rect 4736 96404 4792 96460
rect 4840 96404 4896 96460
rect 4944 96404 5000 96460
rect 5048 96404 5104 96460
rect 5152 96404 5208 96460
rect 24008 96404 24064 96460
rect 24112 96404 24168 96460
rect 24216 96404 24272 96460
rect 24320 96404 24376 96460
rect 24424 96404 24480 96460
rect 24528 96404 24584 96460
rect 24632 96404 24688 96460
rect 24736 96404 24792 96460
rect 24840 96404 24896 96460
rect 24944 96404 25000 96460
rect 25048 96404 25104 96460
rect 25152 96404 25208 96460
rect 14008 95620 14064 95676
rect 14112 95620 14168 95676
rect 14216 95620 14272 95676
rect 14320 95620 14376 95676
rect 14424 95620 14480 95676
rect 14528 95620 14584 95676
rect 14632 95620 14688 95676
rect 14736 95620 14792 95676
rect 14840 95620 14896 95676
rect 14944 95620 15000 95676
rect 15048 95620 15104 95676
rect 15152 95620 15208 95676
rect 34008 95620 34064 95676
rect 34112 95620 34168 95676
rect 34216 95620 34272 95676
rect 34320 95620 34376 95676
rect 34424 95620 34480 95676
rect 34528 95620 34584 95676
rect 34632 95620 34688 95676
rect 34736 95620 34792 95676
rect 34840 95620 34896 95676
rect 34944 95620 35000 95676
rect 35048 95620 35104 95676
rect 35152 95620 35208 95676
rect 4008 94836 4064 94892
rect 4112 94836 4168 94892
rect 4216 94836 4272 94892
rect 4320 94836 4376 94892
rect 4424 94836 4480 94892
rect 4528 94836 4584 94892
rect 4632 94836 4688 94892
rect 4736 94836 4792 94892
rect 4840 94836 4896 94892
rect 4944 94836 5000 94892
rect 5048 94836 5104 94892
rect 5152 94836 5208 94892
rect 24008 94836 24064 94892
rect 24112 94836 24168 94892
rect 24216 94836 24272 94892
rect 24320 94836 24376 94892
rect 24424 94836 24480 94892
rect 24528 94836 24584 94892
rect 24632 94836 24688 94892
rect 24736 94836 24792 94892
rect 24840 94836 24896 94892
rect 24944 94836 25000 94892
rect 25048 94836 25104 94892
rect 25152 94836 25208 94892
rect 14008 94052 14064 94108
rect 14112 94052 14168 94108
rect 14216 94052 14272 94108
rect 14320 94052 14376 94108
rect 14424 94052 14480 94108
rect 14528 94052 14584 94108
rect 14632 94052 14688 94108
rect 14736 94052 14792 94108
rect 14840 94052 14896 94108
rect 14944 94052 15000 94108
rect 15048 94052 15104 94108
rect 15152 94052 15208 94108
rect 34008 94052 34064 94108
rect 34112 94052 34168 94108
rect 34216 94052 34272 94108
rect 34320 94052 34376 94108
rect 34424 94052 34480 94108
rect 34528 94052 34584 94108
rect 34632 94052 34688 94108
rect 34736 94052 34792 94108
rect 34840 94052 34896 94108
rect 34944 94052 35000 94108
rect 35048 94052 35104 94108
rect 35152 94052 35208 94108
rect 4008 93268 4064 93324
rect 4112 93268 4168 93324
rect 4216 93268 4272 93324
rect 4320 93268 4376 93324
rect 4424 93268 4480 93324
rect 4528 93268 4584 93324
rect 4632 93268 4688 93324
rect 4736 93268 4792 93324
rect 4840 93268 4896 93324
rect 4944 93268 5000 93324
rect 5048 93268 5104 93324
rect 5152 93268 5208 93324
rect 24008 93268 24064 93324
rect 24112 93268 24168 93324
rect 24216 93268 24272 93324
rect 24320 93268 24376 93324
rect 24424 93268 24480 93324
rect 24528 93268 24584 93324
rect 24632 93268 24688 93324
rect 24736 93268 24792 93324
rect 24840 93268 24896 93324
rect 24944 93268 25000 93324
rect 25048 93268 25104 93324
rect 25152 93268 25208 93324
rect 14008 92484 14064 92540
rect 14112 92484 14168 92540
rect 14216 92484 14272 92540
rect 14320 92484 14376 92540
rect 14424 92484 14480 92540
rect 14528 92484 14584 92540
rect 14632 92484 14688 92540
rect 14736 92484 14792 92540
rect 14840 92484 14896 92540
rect 14944 92484 15000 92540
rect 15048 92484 15104 92540
rect 15152 92484 15208 92540
rect 34008 92484 34064 92540
rect 34112 92484 34168 92540
rect 34216 92484 34272 92540
rect 34320 92484 34376 92540
rect 34424 92484 34480 92540
rect 34528 92484 34584 92540
rect 34632 92484 34688 92540
rect 34736 92484 34792 92540
rect 34840 92484 34896 92540
rect 34944 92484 35000 92540
rect 35048 92484 35104 92540
rect 35152 92484 35208 92540
rect 4008 91700 4064 91756
rect 4112 91700 4168 91756
rect 4216 91700 4272 91756
rect 4320 91700 4376 91756
rect 4424 91700 4480 91756
rect 4528 91700 4584 91756
rect 4632 91700 4688 91756
rect 4736 91700 4792 91756
rect 4840 91700 4896 91756
rect 4944 91700 5000 91756
rect 5048 91700 5104 91756
rect 5152 91700 5208 91756
rect 24008 91700 24064 91756
rect 24112 91700 24168 91756
rect 24216 91700 24272 91756
rect 24320 91700 24376 91756
rect 24424 91700 24480 91756
rect 24528 91700 24584 91756
rect 24632 91700 24688 91756
rect 24736 91700 24792 91756
rect 24840 91700 24896 91756
rect 24944 91700 25000 91756
rect 25048 91700 25104 91756
rect 25152 91700 25208 91756
rect 14008 90916 14064 90972
rect 14112 90916 14168 90972
rect 14216 90916 14272 90972
rect 14320 90916 14376 90972
rect 14424 90916 14480 90972
rect 14528 90916 14584 90972
rect 14632 90916 14688 90972
rect 14736 90916 14792 90972
rect 14840 90916 14896 90972
rect 14944 90916 15000 90972
rect 15048 90916 15104 90972
rect 15152 90916 15208 90972
rect 34008 90916 34064 90972
rect 34112 90916 34168 90972
rect 34216 90916 34272 90972
rect 34320 90916 34376 90972
rect 34424 90916 34480 90972
rect 34528 90916 34584 90972
rect 34632 90916 34688 90972
rect 34736 90916 34792 90972
rect 34840 90916 34896 90972
rect 34944 90916 35000 90972
rect 35048 90916 35104 90972
rect 35152 90916 35208 90972
rect 4008 90132 4064 90188
rect 4112 90132 4168 90188
rect 4216 90132 4272 90188
rect 4320 90132 4376 90188
rect 4424 90132 4480 90188
rect 4528 90132 4584 90188
rect 4632 90132 4688 90188
rect 4736 90132 4792 90188
rect 4840 90132 4896 90188
rect 4944 90132 5000 90188
rect 5048 90132 5104 90188
rect 5152 90132 5208 90188
rect 24008 90132 24064 90188
rect 24112 90132 24168 90188
rect 24216 90132 24272 90188
rect 24320 90132 24376 90188
rect 24424 90132 24480 90188
rect 24528 90132 24584 90188
rect 24632 90132 24688 90188
rect 24736 90132 24792 90188
rect 24840 90132 24896 90188
rect 24944 90132 25000 90188
rect 25048 90132 25104 90188
rect 25152 90132 25208 90188
rect 14008 89348 14064 89404
rect 14112 89348 14168 89404
rect 14216 89348 14272 89404
rect 14320 89348 14376 89404
rect 14424 89348 14480 89404
rect 14528 89348 14584 89404
rect 14632 89348 14688 89404
rect 14736 89348 14792 89404
rect 14840 89348 14896 89404
rect 14944 89348 15000 89404
rect 15048 89348 15104 89404
rect 15152 89348 15208 89404
rect 34008 89348 34064 89404
rect 34112 89348 34168 89404
rect 34216 89348 34272 89404
rect 34320 89348 34376 89404
rect 34424 89348 34480 89404
rect 34528 89348 34584 89404
rect 34632 89348 34688 89404
rect 34736 89348 34792 89404
rect 34840 89348 34896 89404
rect 34944 89348 35000 89404
rect 35048 89348 35104 89404
rect 35152 89348 35208 89404
rect 4008 88564 4064 88620
rect 4112 88564 4168 88620
rect 4216 88564 4272 88620
rect 4320 88564 4376 88620
rect 4424 88564 4480 88620
rect 4528 88564 4584 88620
rect 4632 88564 4688 88620
rect 4736 88564 4792 88620
rect 4840 88564 4896 88620
rect 4944 88564 5000 88620
rect 5048 88564 5104 88620
rect 5152 88564 5208 88620
rect 24008 88564 24064 88620
rect 24112 88564 24168 88620
rect 24216 88564 24272 88620
rect 24320 88564 24376 88620
rect 24424 88564 24480 88620
rect 24528 88564 24584 88620
rect 24632 88564 24688 88620
rect 24736 88564 24792 88620
rect 24840 88564 24896 88620
rect 24944 88564 25000 88620
rect 25048 88564 25104 88620
rect 25152 88564 25208 88620
rect 14008 87780 14064 87836
rect 14112 87780 14168 87836
rect 14216 87780 14272 87836
rect 14320 87780 14376 87836
rect 14424 87780 14480 87836
rect 14528 87780 14584 87836
rect 14632 87780 14688 87836
rect 14736 87780 14792 87836
rect 14840 87780 14896 87836
rect 14944 87780 15000 87836
rect 15048 87780 15104 87836
rect 15152 87780 15208 87836
rect 34008 87780 34064 87836
rect 34112 87780 34168 87836
rect 34216 87780 34272 87836
rect 34320 87780 34376 87836
rect 34424 87780 34480 87836
rect 34528 87780 34584 87836
rect 34632 87780 34688 87836
rect 34736 87780 34792 87836
rect 34840 87780 34896 87836
rect 34944 87780 35000 87836
rect 35048 87780 35104 87836
rect 35152 87780 35208 87836
rect 4008 86996 4064 87052
rect 4112 86996 4168 87052
rect 4216 86996 4272 87052
rect 4320 86996 4376 87052
rect 4424 86996 4480 87052
rect 4528 86996 4584 87052
rect 4632 86996 4688 87052
rect 4736 86996 4792 87052
rect 4840 86996 4896 87052
rect 4944 86996 5000 87052
rect 5048 86996 5104 87052
rect 5152 86996 5208 87052
rect 24008 86996 24064 87052
rect 24112 86996 24168 87052
rect 24216 86996 24272 87052
rect 24320 86996 24376 87052
rect 24424 86996 24480 87052
rect 24528 86996 24584 87052
rect 24632 86996 24688 87052
rect 24736 86996 24792 87052
rect 24840 86996 24896 87052
rect 24944 86996 25000 87052
rect 25048 86996 25104 87052
rect 25152 86996 25208 87052
rect 13804 86604 13860 86660
rect 14008 86212 14064 86268
rect 14112 86212 14168 86268
rect 14216 86212 14272 86268
rect 14320 86212 14376 86268
rect 14424 86212 14480 86268
rect 14528 86212 14584 86268
rect 14632 86212 14688 86268
rect 14736 86212 14792 86268
rect 14840 86212 14896 86268
rect 14944 86212 15000 86268
rect 15048 86212 15104 86268
rect 15152 86212 15208 86268
rect 34008 86212 34064 86268
rect 34112 86212 34168 86268
rect 34216 86212 34272 86268
rect 34320 86212 34376 86268
rect 34424 86212 34480 86268
rect 34528 86212 34584 86268
rect 34632 86212 34688 86268
rect 34736 86212 34792 86268
rect 34840 86212 34896 86268
rect 34944 86212 35000 86268
rect 35048 86212 35104 86268
rect 35152 86212 35208 86268
rect 13804 85820 13860 85876
rect 4008 85428 4064 85484
rect 4112 85428 4168 85484
rect 4216 85428 4272 85484
rect 4320 85428 4376 85484
rect 4424 85428 4480 85484
rect 4528 85428 4584 85484
rect 4632 85428 4688 85484
rect 4736 85428 4792 85484
rect 4840 85428 4896 85484
rect 4944 85428 5000 85484
rect 5048 85428 5104 85484
rect 5152 85428 5208 85484
rect 24008 85428 24064 85484
rect 24112 85428 24168 85484
rect 24216 85428 24272 85484
rect 24320 85428 24376 85484
rect 24424 85428 24480 85484
rect 24528 85428 24584 85484
rect 24632 85428 24688 85484
rect 24736 85428 24792 85484
rect 24840 85428 24896 85484
rect 24944 85428 25000 85484
rect 25048 85428 25104 85484
rect 25152 85428 25208 85484
rect 15372 85148 15428 85204
rect 13692 84924 13748 84980
rect 14008 84644 14064 84700
rect 14112 84644 14168 84700
rect 14216 84644 14272 84700
rect 14320 84644 14376 84700
rect 14424 84644 14480 84700
rect 14528 84644 14584 84700
rect 14632 84644 14688 84700
rect 14736 84644 14792 84700
rect 14840 84644 14896 84700
rect 14944 84644 15000 84700
rect 15048 84644 15104 84700
rect 15152 84644 15208 84700
rect 34008 84644 34064 84700
rect 34112 84644 34168 84700
rect 34216 84644 34272 84700
rect 34320 84644 34376 84700
rect 34424 84644 34480 84700
rect 34528 84644 34584 84700
rect 34632 84644 34688 84700
rect 34736 84644 34792 84700
rect 34840 84644 34896 84700
rect 34944 84644 35000 84700
rect 35048 84644 35104 84700
rect 35152 84644 35208 84700
rect 13580 84028 13636 84084
rect 19292 84028 19348 84084
rect 4008 83860 4064 83916
rect 4112 83860 4168 83916
rect 4216 83860 4272 83916
rect 4320 83860 4376 83916
rect 4424 83860 4480 83916
rect 4528 83860 4584 83916
rect 4632 83860 4688 83916
rect 4736 83860 4792 83916
rect 4840 83860 4896 83916
rect 4944 83860 5000 83916
rect 5048 83860 5104 83916
rect 5152 83860 5208 83916
rect 24008 83860 24064 83916
rect 24112 83860 24168 83916
rect 24216 83860 24272 83916
rect 24320 83860 24376 83916
rect 24424 83860 24480 83916
rect 24528 83860 24584 83916
rect 24632 83860 24688 83916
rect 24736 83860 24792 83916
rect 24840 83860 24896 83916
rect 24944 83860 25000 83916
rect 25048 83860 25104 83916
rect 25152 83860 25208 83916
rect 13804 83244 13860 83300
rect 13692 83132 13748 83188
rect 14008 83076 14064 83132
rect 14112 83076 14168 83132
rect 14216 83076 14272 83132
rect 14320 83076 14376 83132
rect 14424 83076 14480 83132
rect 14528 83076 14584 83132
rect 14632 83076 14688 83132
rect 14736 83076 14792 83132
rect 14840 83076 14896 83132
rect 14944 83076 15000 83132
rect 15048 83076 15104 83132
rect 15152 83076 15208 83132
rect 34008 83076 34064 83132
rect 34112 83076 34168 83132
rect 34216 83076 34272 83132
rect 34320 83076 34376 83132
rect 34424 83076 34480 83132
rect 34528 83076 34584 83132
rect 34632 83076 34688 83132
rect 34736 83076 34792 83132
rect 34840 83076 34896 83132
rect 34944 83076 35000 83132
rect 35048 83076 35104 83132
rect 35152 83076 35208 83132
rect 13804 82684 13860 82740
rect 10220 82460 10276 82516
rect 4008 82292 4064 82348
rect 4112 82292 4168 82348
rect 4216 82292 4272 82348
rect 4320 82292 4376 82348
rect 4424 82292 4480 82348
rect 4528 82292 4584 82348
rect 4632 82292 4688 82348
rect 4736 82292 4792 82348
rect 4840 82292 4896 82348
rect 4944 82292 5000 82348
rect 5048 82292 5104 82348
rect 5152 82292 5208 82348
rect 24008 82292 24064 82348
rect 24112 82292 24168 82348
rect 24216 82292 24272 82348
rect 24320 82292 24376 82348
rect 24424 82292 24480 82348
rect 24528 82292 24584 82348
rect 24632 82292 24688 82348
rect 24736 82292 24792 82348
rect 24840 82292 24896 82348
rect 24944 82292 25000 82348
rect 25048 82292 25104 82348
rect 25152 82292 25208 82348
rect 11004 82124 11060 82180
rect 13804 81900 13860 81956
rect 15484 81788 15540 81844
rect 10220 81452 10276 81508
rect 14008 81508 14064 81564
rect 14112 81508 14168 81564
rect 14216 81508 14272 81564
rect 14320 81508 14376 81564
rect 14424 81508 14480 81564
rect 14528 81508 14584 81564
rect 14632 81508 14688 81564
rect 14736 81508 14792 81564
rect 14840 81508 14896 81564
rect 14944 81508 15000 81564
rect 15048 81508 15104 81564
rect 15152 81508 15208 81564
rect 34008 81508 34064 81564
rect 34112 81508 34168 81564
rect 34216 81508 34272 81564
rect 34320 81508 34376 81564
rect 34424 81508 34480 81564
rect 34528 81508 34584 81564
rect 34632 81508 34688 81564
rect 34736 81508 34792 81564
rect 34840 81508 34896 81564
rect 34944 81508 35000 81564
rect 35048 81508 35104 81564
rect 35152 81508 35208 81564
rect 13804 81004 13860 81060
rect 4008 80724 4064 80780
rect 4112 80724 4168 80780
rect 4216 80724 4272 80780
rect 4320 80724 4376 80780
rect 4424 80724 4480 80780
rect 4528 80724 4584 80780
rect 4632 80724 4688 80780
rect 4736 80724 4792 80780
rect 4840 80724 4896 80780
rect 4944 80724 5000 80780
rect 5048 80724 5104 80780
rect 5152 80724 5208 80780
rect 24008 80724 24064 80780
rect 24112 80724 24168 80780
rect 24216 80724 24272 80780
rect 24320 80724 24376 80780
rect 24424 80724 24480 80780
rect 24528 80724 24584 80780
rect 24632 80724 24688 80780
rect 24736 80724 24792 80780
rect 24840 80724 24896 80780
rect 24944 80724 25000 80780
rect 25048 80724 25104 80780
rect 25152 80724 25208 80780
rect 15484 80556 15540 80612
rect 11004 80444 11060 80500
rect 14008 79940 14064 79996
rect 14112 79940 14168 79996
rect 14216 79940 14272 79996
rect 14320 79940 14376 79996
rect 14424 79940 14480 79996
rect 14528 79940 14584 79996
rect 14632 79940 14688 79996
rect 14736 79940 14792 79996
rect 14840 79940 14896 79996
rect 14944 79940 15000 79996
rect 15048 79940 15104 79996
rect 15152 79940 15208 79996
rect 34008 79940 34064 79996
rect 34112 79940 34168 79996
rect 34216 79940 34272 79996
rect 34320 79940 34376 79996
rect 34424 79940 34480 79996
rect 34528 79940 34584 79996
rect 34632 79940 34688 79996
rect 34736 79940 34792 79996
rect 34840 79940 34896 79996
rect 34944 79940 35000 79996
rect 35048 79940 35104 79996
rect 35152 79940 35208 79996
rect 5292 79772 5348 79828
rect 4008 79156 4064 79212
rect 4112 79156 4168 79212
rect 4216 79156 4272 79212
rect 4320 79156 4376 79212
rect 4424 79156 4480 79212
rect 4528 79156 4584 79212
rect 4632 79156 4688 79212
rect 4736 79156 4792 79212
rect 4840 79156 4896 79212
rect 4944 79156 5000 79212
rect 5048 79156 5104 79212
rect 5152 79156 5208 79212
rect 24008 79156 24064 79212
rect 24112 79156 24168 79212
rect 24216 79156 24272 79212
rect 24320 79156 24376 79212
rect 24424 79156 24480 79212
rect 24528 79156 24584 79212
rect 24632 79156 24688 79212
rect 24736 79156 24792 79212
rect 24840 79156 24896 79212
rect 24944 79156 25000 79212
rect 25048 79156 25104 79212
rect 25152 79156 25208 79212
rect 13692 78988 13748 79044
rect 15484 78652 15540 78708
rect 11004 78540 11060 78596
rect 14008 78372 14064 78428
rect 14112 78372 14168 78428
rect 14216 78372 14272 78428
rect 14320 78372 14376 78428
rect 14424 78372 14480 78428
rect 14528 78372 14584 78428
rect 14632 78372 14688 78428
rect 14736 78372 14792 78428
rect 14840 78372 14896 78428
rect 14944 78372 15000 78428
rect 15048 78372 15104 78428
rect 15152 78372 15208 78428
rect 34008 78372 34064 78428
rect 34112 78372 34168 78428
rect 34216 78372 34272 78428
rect 34320 78372 34376 78428
rect 34424 78372 34480 78428
rect 34528 78372 34584 78428
rect 34632 78372 34688 78428
rect 34736 78372 34792 78428
rect 34840 78372 34896 78428
rect 34944 78372 35000 78428
rect 35048 78372 35104 78428
rect 35152 78372 35208 78428
rect 5292 78204 5348 78260
rect 13692 78092 13748 78148
rect 15484 77980 15540 78036
rect 4008 77588 4064 77644
rect 4112 77588 4168 77644
rect 4216 77588 4272 77644
rect 4320 77588 4376 77644
rect 4424 77588 4480 77644
rect 4528 77588 4584 77644
rect 4632 77588 4688 77644
rect 4736 77588 4792 77644
rect 4840 77588 4896 77644
rect 4944 77588 5000 77644
rect 5048 77588 5104 77644
rect 5152 77588 5208 77644
rect 24008 77588 24064 77644
rect 24112 77588 24168 77644
rect 24216 77588 24272 77644
rect 24320 77588 24376 77644
rect 24424 77588 24480 77644
rect 24528 77588 24584 77644
rect 24632 77588 24688 77644
rect 24736 77588 24792 77644
rect 24840 77588 24896 77644
rect 24944 77588 25000 77644
rect 25048 77588 25104 77644
rect 25152 77588 25208 77644
rect 13804 77308 13860 77364
rect 14008 76804 14064 76860
rect 14112 76804 14168 76860
rect 14216 76804 14272 76860
rect 14320 76804 14376 76860
rect 14424 76804 14480 76860
rect 14528 76804 14584 76860
rect 14632 76804 14688 76860
rect 14736 76804 14792 76860
rect 14840 76804 14896 76860
rect 14944 76804 15000 76860
rect 15048 76804 15104 76860
rect 15152 76804 15208 76860
rect 34008 76804 34064 76860
rect 34112 76804 34168 76860
rect 34216 76804 34272 76860
rect 34320 76804 34376 76860
rect 34424 76804 34480 76860
rect 34528 76804 34584 76860
rect 34632 76804 34688 76860
rect 34736 76804 34792 76860
rect 34840 76804 34896 76860
rect 34944 76804 35000 76860
rect 35048 76804 35104 76860
rect 35152 76804 35208 76860
rect 3836 76636 3892 76692
rect 19292 76300 19348 76356
rect 4008 76020 4064 76076
rect 4112 76020 4168 76076
rect 4216 76020 4272 76076
rect 4320 76020 4376 76076
rect 4424 76020 4480 76076
rect 4528 76020 4584 76076
rect 4632 76020 4688 76076
rect 4736 76020 4792 76076
rect 4840 76020 4896 76076
rect 4944 76020 5000 76076
rect 5048 76020 5104 76076
rect 5152 76020 5208 76076
rect 24008 76020 24064 76076
rect 24112 76020 24168 76076
rect 24216 76020 24272 76076
rect 24320 76020 24376 76076
rect 24424 76020 24480 76076
rect 24528 76020 24584 76076
rect 24632 76020 24688 76076
rect 24736 76020 24792 76076
rect 24840 76020 24896 76076
rect 24944 76020 25000 76076
rect 25048 76020 25104 76076
rect 25152 76020 25208 76076
rect 13692 75516 13748 75572
rect 14008 75236 14064 75292
rect 14112 75236 14168 75292
rect 14216 75236 14272 75292
rect 14320 75236 14376 75292
rect 14424 75236 14480 75292
rect 14528 75236 14584 75292
rect 14632 75236 14688 75292
rect 14736 75236 14792 75292
rect 14840 75236 14896 75292
rect 14944 75236 15000 75292
rect 15048 75236 15104 75292
rect 15152 75236 15208 75292
rect 34008 75236 34064 75292
rect 34112 75236 34168 75292
rect 34216 75236 34272 75292
rect 34320 75236 34376 75292
rect 34424 75236 34480 75292
rect 34528 75236 34584 75292
rect 34632 75236 34688 75292
rect 34736 75236 34792 75292
rect 34840 75236 34896 75292
rect 34944 75236 35000 75292
rect 35048 75236 35104 75292
rect 35152 75236 35208 75292
rect 13804 75068 13860 75124
rect 15372 75068 15428 75124
rect 4008 74452 4064 74508
rect 4112 74452 4168 74508
rect 4216 74452 4272 74508
rect 4320 74452 4376 74508
rect 4424 74452 4480 74508
rect 4528 74452 4584 74508
rect 4632 74452 4688 74508
rect 4736 74452 4792 74508
rect 4840 74452 4896 74508
rect 4944 74452 5000 74508
rect 5048 74452 5104 74508
rect 5152 74452 5208 74508
rect 24008 74452 24064 74508
rect 24112 74452 24168 74508
rect 24216 74452 24272 74508
rect 24320 74452 24376 74508
rect 24424 74452 24480 74508
rect 24528 74452 24584 74508
rect 24632 74452 24688 74508
rect 24736 74452 24792 74508
rect 24840 74452 24896 74508
rect 24944 74452 25000 74508
rect 25048 74452 25104 74508
rect 25152 74452 25208 74508
rect 3836 74060 3892 74116
rect 13580 73948 13636 74004
rect 13692 73836 13748 73892
rect 14008 73668 14064 73724
rect 14112 73668 14168 73724
rect 14216 73668 14272 73724
rect 14320 73668 14376 73724
rect 14424 73668 14480 73724
rect 14528 73668 14584 73724
rect 14632 73668 14688 73724
rect 14736 73668 14792 73724
rect 14840 73668 14896 73724
rect 14944 73668 15000 73724
rect 15048 73668 15104 73724
rect 15152 73668 15208 73724
rect 34008 73668 34064 73724
rect 34112 73668 34168 73724
rect 34216 73668 34272 73724
rect 34320 73668 34376 73724
rect 34424 73668 34480 73724
rect 34528 73668 34584 73724
rect 34632 73668 34688 73724
rect 34736 73668 34792 73724
rect 34840 73668 34896 73724
rect 34944 73668 35000 73724
rect 35048 73668 35104 73724
rect 35152 73668 35208 73724
rect 13692 73500 13748 73556
rect 4008 72884 4064 72940
rect 4112 72884 4168 72940
rect 4216 72884 4272 72940
rect 4320 72884 4376 72940
rect 4424 72884 4480 72940
rect 4528 72884 4584 72940
rect 4632 72884 4688 72940
rect 4736 72884 4792 72940
rect 4840 72884 4896 72940
rect 4944 72884 5000 72940
rect 5048 72884 5104 72940
rect 5152 72884 5208 72940
rect 24008 72884 24064 72940
rect 24112 72884 24168 72940
rect 24216 72884 24272 72940
rect 24320 72884 24376 72940
rect 24424 72884 24480 72940
rect 24528 72884 24584 72940
rect 24632 72884 24688 72940
rect 24736 72884 24792 72940
rect 24840 72884 24896 72940
rect 24944 72884 25000 72940
rect 25048 72884 25104 72940
rect 25152 72884 25208 72940
rect 14008 72100 14064 72156
rect 14112 72100 14168 72156
rect 14216 72100 14272 72156
rect 14320 72100 14376 72156
rect 14424 72100 14480 72156
rect 14528 72100 14584 72156
rect 14632 72100 14688 72156
rect 14736 72100 14792 72156
rect 14840 72100 14896 72156
rect 14944 72100 15000 72156
rect 15048 72100 15104 72156
rect 15152 72100 15208 72156
rect 34008 72100 34064 72156
rect 34112 72100 34168 72156
rect 34216 72100 34272 72156
rect 34320 72100 34376 72156
rect 34424 72100 34480 72156
rect 34528 72100 34584 72156
rect 34632 72100 34688 72156
rect 34736 72100 34792 72156
rect 34840 72100 34896 72156
rect 34944 72100 35000 72156
rect 35048 72100 35104 72156
rect 35152 72100 35208 72156
rect 35308 71484 35364 71540
rect 4008 71316 4064 71372
rect 4112 71316 4168 71372
rect 4216 71316 4272 71372
rect 4320 71316 4376 71372
rect 4424 71316 4480 71372
rect 4528 71316 4584 71372
rect 4632 71316 4688 71372
rect 4736 71316 4792 71372
rect 4840 71316 4896 71372
rect 4944 71316 5000 71372
rect 5048 71316 5104 71372
rect 5152 71316 5208 71372
rect 24008 71316 24064 71372
rect 24112 71316 24168 71372
rect 24216 71316 24272 71372
rect 24320 71316 24376 71372
rect 24424 71316 24480 71372
rect 24528 71316 24584 71372
rect 24632 71316 24688 71372
rect 24736 71316 24792 71372
rect 24840 71316 24896 71372
rect 24944 71316 25000 71372
rect 25048 71316 25104 71372
rect 25152 71316 25208 71372
rect 13468 70588 13524 70644
rect 14008 70532 14064 70588
rect 14112 70532 14168 70588
rect 14216 70532 14272 70588
rect 14320 70532 14376 70588
rect 14424 70532 14480 70588
rect 14528 70532 14584 70588
rect 14632 70532 14688 70588
rect 14736 70532 14792 70588
rect 14840 70532 14896 70588
rect 14944 70532 15000 70588
rect 15048 70532 15104 70588
rect 15152 70532 15208 70588
rect 34008 70532 34064 70588
rect 34112 70532 34168 70588
rect 34216 70532 34272 70588
rect 34320 70532 34376 70588
rect 34424 70532 34480 70588
rect 34528 70532 34584 70588
rect 34632 70532 34688 70588
rect 34736 70532 34792 70588
rect 34840 70532 34896 70588
rect 34944 70532 35000 70588
rect 35048 70532 35104 70588
rect 35152 70532 35208 70588
rect 35308 70364 35364 70420
rect 4008 69748 4064 69804
rect 4112 69748 4168 69804
rect 4216 69748 4272 69804
rect 4320 69748 4376 69804
rect 4424 69748 4480 69804
rect 4528 69748 4584 69804
rect 4632 69748 4688 69804
rect 4736 69748 4792 69804
rect 4840 69748 4896 69804
rect 4944 69748 5000 69804
rect 5048 69748 5104 69804
rect 5152 69748 5208 69804
rect 24008 69748 24064 69804
rect 24112 69748 24168 69804
rect 24216 69748 24272 69804
rect 24320 69748 24376 69804
rect 24424 69748 24480 69804
rect 24528 69748 24584 69804
rect 24632 69748 24688 69804
rect 24736 69748 24792 69804
rect 24840 69748 24896 69804
rect 24944 69748 25000 69804
rect 25048 69748 25104 69804
rect 25152 69748 25208 69804
rect 13692 69692 13748 69748
rect 15372 69468 15428 69524
rect 19404 69132 19460 69188
rect 14008 68964 14064 69020
rect 14112 68964 14168 69020
rect 14216 68964 14272 69020
rect 14320 68964 14376 69020
rect 14424 68964 14480 69020
rect 14528 68964 14584 69020
rect 14632 68964 14688 69020
rect 14736 68964 14792 69020
rect 14840 68964 14896 69020
rect 14944 68964 15000 69020
rect 15048 68964 15104 69020
rect 15152 68964 15208 69020
rect 13580 68796 13636 68852
rect 34008 68964 34064 69020
rect 34112 68964 34168 69020
rect 34216 68964 34272 69020
rect 34320 68964 34376 69020
rect 34424 68964 34480 69020
rect 34528 68964 34584 69020
rect 34632 68964 34688 69020
rect 34736 68964 34792 69020
rect 34840 68964 34896 69020
rect 34944 68964 35000 69020
rect 35048 68964 35104 69020
rect 35152 68964 35208 69020
rect 4008 68180 4064 68236
rect 4112 68180 4168 68236
rect 4216 68180 4272 68236
rect 4320 68180 4376 68236
rect 4424 68180 4480 68236
rect 4528 68180 4584 68236
rect 4632 68180 4688 68236
rect 4736 68180 4792 68236
rect 4840 68180 4896 68236
rect 4944 68180 5000 68236
rect 5048 68180 5104 68236
rect 5152 68180 5208 68236
rect 24008 68180 24064 68236
rect 24112 68180 24168 68236
rect 24216 68180 24272 68236
rect 24320 68180 24376 68236
rect 24424 68180 24480 68236
rect 24528 68180 24584 68236
rect 24632 68180 24688 68236
rect 24736 68180 24792 68236
rect 24840 68180 24896 68236
rect 24944 68180 25000 68236
rect 25048 68180 25104 68236
rect 25152 68180 25208 68236
rect 15372 67788 15428 67844
rect 6524 67340 6580 67396
rect 14008 67396 14064 67452
rect 14112 67396 14168 67452
rect 14216 67396 14272 67452
rect 14320 67396 14376 67452
rect 14424 67396 14480 67452
rect 14528 67396 14584 67452
rect 14632 67396 14688 67452
rect 14736 67396 14792 67452
rect 14840 67396 14896 67452
rect 14944 67396 15000 67452
rect 15048 67396 15104 67452
rect 15152 67396 15208 67452
rect 34008 67396 34064 67452
rect 34112 67396 34168 67452
rect 34216 67396 34272 67452
rect 34320 67396 34376 67452
rect 34424 67396 34480 67452
rect 34528 67396 34584 67452
rect 34632 67396 34688 67452
rect 34736 67396 34792 67452
rect 34840 67396 34896 67452
rect 34944 67396 35000 67452
rect 35048 67396 35104 67452
rect 35152 67396 35208 67452
rect 25340 66892 25396 66948
rect 4008 66612 4064 66668
rect 4112 66612 4168 66668
rect 4216 66612 4272 66668
rect 4320 66612 4376 66668
rect 4424 66612 4480 66668
rect 4528 66612 4584 66668
rect 4632 66612 4688 66668
rect 4736 66612 4792 66668
rect 4840 66612 4896 66668
rect 4944 66612 5000 66668
rect 5048 66612 5104 66668
rect 5152 66612 5208 66668
rect 24008 66612 24064 66668
rect 24112 66612 24168 66668
rect 24216 66612 24272 66668
rect 24320 66612 24376 66668
rect 24424 66612 24480 66668
rect 24528 66612 24584 66668
rect 24632 66612 24688 66668
rect 24736 66612 24792 66668
rect 24840 66612 24896 66668
rect 24944 66612 25000 66668
rect 25048 66612 25104 66668
rect 25152 66612 25208 66668
rect 19180 66220 19236 66276
rect 14008 65828 14064 65884
rect 14112 65828 14168 65884
rect 14216 65828 14272 65884
rect 14320 65828 14376 65884
rect 14424 65828 14480 65884
rect 14528 65828 14584 65884
rect 14632 65828 14688 65884
rect 14736 65828 14792 65884
rect 14840 65828 14896 65884
rect 14944 65828 15000 65884
rect 15048 65828 15104 65884
rect 15152 65828 15208 65884
rect 34008 65828 34064 65884
rect 34112 65828 34168 65884
rect 34216 65828 34272 65884
rect 34320 65828 34376 65884
rect 34424 65828 34480 65884
rect 34528 65828 34584 65884
rect 34632 65828 34688 65884
rect 34736 65828 34792 65884
rect 34840 65828 34896 65884
rect 34944 65828 35000 65884
rect 35048 65828 35104 65884
rect 35152 65828 35208 65884
rect 5292 65548 5348 65604
rect 13580 65324 13636 65380
rect 25340 65324 25396 65380
rect 13804 65100 13860 65156
rect 15484 65100 15540 65156
rect 4008 65044 4064 65100
rect 4112 65044 4168 65100
rect 4216 65044 4272 65100
rect 4320 65044 4376 65100
rect 4424 65044 4480 65100
rect 4528 65044 4584 65100
rect 4632 65044 4688 65100
rect 4736 65044 4792 65100
rect 4840 65044 4896 65100
rect 4944 65044 5000 65100
rect 5048 65044 5104 65100
rect 5152 65044 5208 65100
rect 24008 65044 24064 65100
rect 24112 65044 24168 65100
rect 24216 65044 24272 65100
rect 24320 65044 24376 65100
rect 24424 65044 24480 65100
rect 24528 65044 24584 65100
rect 24632 65044 24688 65100
rect 24736 65044 24792 65100
rect 24840 65044 24896 65100
rect 24944 65044 25000 65100
rect 25048 65044 25104 65100
rect 25152 65044 25208 65100
rect 15372 64764 15428 64820
rect 19180 64428 19236 64484
rect 14008 64260 14064 64316
rect 14112 64260 14168 64316
rect 14216 64260 14272 64316
rect 14320 64260 14376 64316
rect 14424 64260 14480 64316
rect 14528 64260 14584 64316
rect 14632 64260 14688 64316
rect 14736 64260 14792 64316
rect 14840 64260 14896 64316
rect 14944 64260 15000 64316
rect 15048 64260 15104 64316
rect 15152 64260 15208 64316
rect 34008 64260 34064 64316
rect 34112 64260 34168 64316
rect 34216 64260 34272 64316
rect 34320 64260 34376 64316
rect 34424 64260 34480 64316
rect 34528 64260 34584 64316
rect 34632 64260 34688 64316
rect 34736 64260 34792 64316
rect 34840 64260 34896 64316
rect 34944 64260 35000 64316
rect 35048 64260 35104 64316
rect 35152 64260 35208 64316
rect 13692 64092 13748 64148
rect 15372 64092 15428 64148
rect 5404 63980 5460 64036
rect 19964 63980 20020 64036
rect 4008 63476 4064 63532
rect 4112 63476 4168 63532
rect 4216 63476 4272 63532
rect 4320 63476 4376 63532
rect 4424 63476 4480 63532
rect 4528 63476 4584 63532
rect 4632 63476 4688 63532
rect 4736 63476 4792 63532
rect 4840 63476 4896 63532
rect 4944 63476 5000 63532
rect 5048 63476 5104 63532
rect 5152 63476 5208 63532
rect 13804 63644 13860 63700
rect 13692 63532 13748 63588
rect 24008 63476 24064 63532
rect 24112 63476 24168 63532
rect 24216 63476 24272 63532
rect 24320 63476 24376 63532
rect 24424 63476 24480 63532
rect 24528 63476 24584 63532
rect 24632 63476 24688 63532
rect 24736 63476 24792 63532
rect 24840 63476 24896 63532
rect 24944 63476 25000 63532
rect 25048 63476 25104 63532
rect 25152 63476 25208 63532
rect 13692 63308 13748 63364
rect 33852 63196 33908 63252
rect 15484 62972 15540 63028
rect 25340 62972 25396 63028
rect 19964 62860 20020 62916
rect 14008 62692 14064 62748
rect 14112 62692 14168 62748
rect 14216 62692 14272 62748
rect 14320 62692 14376 62748
rect 14424 62692 14480 62748
rect 14528 62692 14584 62748
rect 14632 62692 14688 62748
rect 14736 62692 14792 62748
rect 14840 62692 14896 62748
rect 14944 62692 15000 62748
rect 15048 62692 15104 62748
rect 15152 62692 15208 62748
rect 34008 62692 34064 62748
rect 34112 62692 34168 62748
rect 34216 62692 34272 62748
rect 34320 62692 34376 62748
rect 34424 62692 34480 62748
rect 34528 62692 34584 62748
rect 34632 62692 34688 62748
rect 34736 62692 34792 62748
rect 34840 62692 34896 62748
rect 34944 62692 35000 62748
rect 35048 62692 35104 62748
rect 35152 62692 35208 62748
rect 13804 62636 13860 62692
rect 19404 62524 19460 62580
rect 13580 62412 13636 62468
rect 33852 62412 33908 62468
rect 5292 62300 5348 62356
rect 4008 61908 4064 61964
rect 4112 61908 4168 61964
rect 4216 61908 4272 61964
rect 4320 61908 4376 61964
rect 4424 61908 4480 61964
rect 4528 61908 4584 61964
rect 4632 61908 4688 61964
rect 4736 61908 4792 61964
rect 4840 61908 4896 61964
rect 4944 61908 5000 61964
rect 5048 61908 5104 61964
rect 5152 61908 5208 61964
rect 24008 61908 24064 61964
rect 24112 61908 24168 61964
rect 24216 61908 24272 61964
rect 24320 61908 24376 61964
rect 24424 61908 24480 61964
rect 24528 61908 24584 61964
rect 24632 61908 24688 61964
rect 24736 61908 24792 61964
rect 24840 61908 24896 61964
rect 24944 61908 25000 61964
rect 25048 61908 25104 61964
rect 25152 61908 25208 61964
rect 13804 61628 13860 61684
rect 19292 61516 19348 61572
rect 5292 61404 5348 61460
rect 25340 61404 25396 61460
rect 5404 61292 5460 61348
rect 13692 61292 13748 61348
rect 14008 61124 14064 61180
rect 14112 61124 14168 61180
rect 14216 61124 14272 61180
rect 14320 61124 14376 61180
rect 14424 61124 14480 61180
rect 14528 61124 14584 61180
rect 14632 61124 14688 61180
rect 14736 61124 14792 61180
rect 14840 61124 14896 61180
rect 14944 61124 15000 61180
rect 15048 61124 15104 61180
rect 15152 61124 15208 61180
rect 34008 61124 34064 61180
rect 34112 61124 34168 61180
rect 34216 61124 34272 61180
rect 34320 61124 34376 61180
rect 34424 61124 34480 61180
rect 34528 61124 34584 61180
rect 34632 61124 34688 61180
rect 34736 61124 34792 61180
rect 34840 61124 34896 61180
rect 34944 61124 35000 61180
rect 35048 61124 35104 61180
rect 35152 61124 35208 61180
rect 4008 60340 4064 60396
rect 4112 60340 4168 60396
rect 4216 60340 4272 60396
rect 4320 60340 4376 60396
rect 4424 60340 4480 60396
rect 4528 60340 4584 60396
rect 4632 60340 4688 60396
rect 4736 60340 4792 60396
rect 4840 60340 4896 60396
rect 4944 60340 5000 60396
rect 5048 60340 5104 60396
rect 5152 60340 5208 60396
rect 24008 60340 24064 60396
rect 24112 60340 24168 60396
rect 24216 60340 24272 60396
rect 24320 60340 24376 60396
rect 24424 60340 24480 60396
rect 24528 60340 24584 60396
rect 24632 60340 24688 60396
rect 24736 60340 24792 60396
rect 24840 60340 24896 60396
rect 24944 60340 25000 60396
rect 25048 60340 25104 60396
rect 25152 60340 25208 60396
rect 6524 59724 6580 59780
rect 14008 59556 14064 59612
rect 14112 59556 14168 59612
rect 14216 59556 14272 59612
rect 14320 59556 14376 59612
rect 14424 59556 14480 59612
rect 14528 59556 14584 59612
rect 14632 59556 14688 59612
rect 14736 59556 14792 59612
rect 14840 59556 14896 59612
rect 14944 59556 15000 59612
rect 15048 59556 15104 59612
rect 15152 59556 15208 59612
rect 34008 59556 34064 59612
rect 34112 59556 34168 59612
rect 34216 59556 34272 59612
rect 34320 59556 34376 59612
rect 34424 59556 34480 59612
rect 34528 59556 34584 59612
rect 34632 59556 34688 59612
rect 34736 59556 34792 59612
rect 34840 59556 34896 59612
rect 34944 59556 35000 59612
rect 35048 59556 35104 59612
rect 35152 59556 35208 59612
rect 19068 59500 19124 59556
rect 13804 58940 13860 58996
rect 19292 58828 19348 58884
rect 4008 58772 4064 58828
rect 4112 58772 4168 58828
rect 4216 58772 4272 58828
rect 4320 58772 4376 58828
rect 4424 58772 4480 58828
rect 4528 58772 4584 58828
rect 4632 58772 4688 58828
rect 4736 58772 4792 58828
rect 4840 58772 4896 58828
rect 4944 58772 5000 58828
rect 5048 58772 5104 58828
rect 5152 58772 5208 58828
rect 24008 58772 24064 58828
rect 24112 58772 24168 58828
rect 24216 58772 24272 58828
rect 24320 58772 24376 58828
rect 24424 58772 24480 58828
rect 24528 58772 24584 58828
rect 24632 58772 24688 58828
rect 24736 58772 24792 58828
rect 24840 58772 24896 58828
rect 24944 58772 25000 58828
rect 25048 58772 25104 58828
rect 25152 58772 25208 58828
rect 13468 58716 13524 58772
rect 19740 58716 19796 58772
rect 7420 58604 7476 58660
rect 18508 58604 18564 58660
rect 19628 58604 19684 58660
rect 15372 58156 15428 58212
rect 14008 57988 14064 58044
rect 14112 57988 14168 58044
rect 14216 57988 14272 58044
rect 14320 57988 14376 58044
rect 14424 57988 14480 58044
rect 14528 57988 14584 58044
rect 14632 57988 14688 58044
rect 14736 57988 14792 58044
rect 14840 57988 14896 58044
rect 14944 57988 15000 58044
rect 15048 57988 15104 58044
rect 15152 57988 15208 58044
rect 13692 57932 13748 57988
rect 34008 57988 34064 58044
rect 34112 57988 34168 58044
rect 34216 57988 34272 58044
rect 34320 57988 34376 58044
rect 34424 57988 34480 58044
rect 34528 57988 34584 58044
rect 34632 57988 34688 58044
rect 34736 57988 34792 58044
rect 34840 57988 34896 58044
rect 34944 57988 35000 58044
rect 35048 57988 35104 58044
rect 35152 57988 35208 58044
rect 19292 57372 19348 57428
rect 19740 57372 19796 57428
rect 4008 57204 4064 57260
rect 4112 57204 4168 57260
rect 4216 57204 4272 57260
rect 4320 57204 4376 57260
rect 4424 57204 4480 57260
rect 4528 57204 4584 57260
rect 4632 57204 4688 57260
rect 4736 57204 4792 57260
rect 4840 57204 4896 57260
rect 4944 57204 5000 57260
rect 5048 57204 5104 57260
rect 5152 57204 5208 57260
rect 24008 57204 24064 57260
rect 24112 57204 24168 57260
rect 24216 57204 24272 57260
rect 24320 57204 24376 57260
rect 24424 57204 24480 57260
rect 24528 57204 24584 57260
rect 24632 57204 24688 57260
rect 24736 57204 24792 57260
rect 24840 57204 24896 57260
rect 24944 57204 25000 57260
rect 25048 57204 25104 57260
rect 25152 57204 25208 57260
rect 13804 56812 13860 56868
rect 13468 56700 13524 56756
rect 5292 56588 5348 56644
rect 14008 56420 14064 56476
rect 14112 56420 14168 56476
rect 14216 56420 14272 56476
rect 14320 56420 14376 56476
rect 14424 56420 14480 56476
rect 14528 56420 14584 56476
rect 14632 56420 14688 56476
rect 14736 56420 14792 56476
rect 14840 56420 14896 56476
rect 14944 56420 15000 56476
rect 15048 56420 15104 56476
rect 15152 56420 15208 56476
rect 34008 56420 34064 56476
rect 34112 56420 34168 56476
rect 34216 56420 34272 56476
rect 34320 56420 34376 56476
rect 34424 56420 34480 56476
rect 34528 56420 34584 56476
rect 34632 56420 34688 56476
rect 34736 56420 34792 56476
rect 34840 56420 34896 56476
rect 34944 56420 35000 56476
rect 35048 56420 35104 56476
rect 35152 56420 35208 56476
rect 18508 56252 18564 56308
rect 13580 56140 13636 56196
rect 13804 55692 13860 55748
rect 4008 55636 4064 55692
rect 4112 55636 4168 55692
rect 4216 55636 4272 55692
rect 4320 55636 4376 55692
rect 4424 55636 4480 55692
rect 4528 55636 4584 55692
rect 4632 55636 4688 55692
rect 4736 55636 4792 55692
rect 4840 55636 4896 55692
rect 4944 55636 5000 55692
rect 5048 55636 5104 55692
rect 5152 55636 5208 55692
rect 24008 55636 24064 55692
rect 24112 55636 24168 55692
rect 24216 55636 24272 55692
rect 24320 55636 24376 55692
rect 24424 55636 24480 55692
rect 24528 55636 24584 55692
rect 24632 55636 24688 55692
rect 24736 55636 24792 55692
rect 24840 55636 24896 55692
rect 24944 55636 25000 55692
rect 25048 55636 25104 55692
rect 25152 55636 25208 55692
rect 10108 55468 10164 55524
rect 13468 55356 13524 55412
rect 19068 55356 19124 55412
rect 13804 55132 13860 55188
rect 14008 54852 14064 54908
rect 14112 54852 14168 54908
rect 14216 54852 14272 54908
rect 14320 54852 14376 54908
rect 14424 54852 14480 54908
rect 14528 54852 14584 54908
rect 14632 54852 14688 54908
rect 14736 54852 14792 54908
rect 14840 54852 14896 54908
rect 14944 54852 15000 54908
rect 15048 54852 15104 54908
rect 15152 54852 15208 54908
rect 34008 54852 34064 54908
rect 34112 54852 34168 54908
rect 34216 54852 34272 54908
rect 34320 54852 34376 54908
rect 34424 54852 34480 54908
rect 34528 54852 34584 54908
rect 34632 54852 34688 54908
rect 34736 54852 34792 54908
rect 34840 54852 34896 54908
rect 34944 54852 35000 54908
rect 35048 54852 35104 54908
rect 35152 54852 35208 54908
rect 6300 54572 6356 54628
rect 4008 54068 4064 54124
rect 4112 54068 4168 54124
rect 4216 54068 4272 54124
rect 4320 54068 4376 54124
rect 4424 54068 4480 54124
rect 4528 54068 4584 54124
rect 4632 54068 4688 54124
rect 4736 54068 4792 54124
rect 4840 54068 4896 54124
rect 4944 54068 5000 54124
rect 5048 54068 5104 54124
rect 5152 54068 5208 54124
rect 24008 54068 24064 54124
rect 24112 54068 24168 54124
rect 24216 54068 24272 54124
rect 24320 54068 24376 54124
rect 24424 54068 24480 54124
rect 24528 54068 24584 54124
rect 24632 54068 24688 54124
rect 24736 54068 24792 54124
rect 24840 54068 24896 54124
rect 24944 54068 25000 54124
rect 25048 54068 25104 54124
rect 25152 54068 25208 54124
rect 15372 53900 15428 53956
rect 11900 53564 11956 53620
rect 15372 53452 15428 53508
rect 14008 53284 14064 53340
rect 14112 53284 14168 53340
rect 14216 53284 14272 53340
rect 14320 53284 14376 53340
rect 14424 53284 14480 53340
rect 14528 53284 14584 53340
rect 14632 53284 14688 53340
rect 14736 53284 14792 53340
rect 14840 53284 14896 53340
rect 14944 53284 15000 53340
rect 15048 53284 15104 53340
rect 15152 53284 15208 53340
rect 34008 53284 34064 53340
rect 34112 53284 34168 53340
rect 34216 53284 34272 53340
rect 34320 53284 34376 53340
rect 34424 53284 34480 53340
rect 34528 53284 34584 53340
rect 34632 53284 34688 53340
rect 34736 53284 34792 53340
rect 34840 53284 34896 53340
rect 34944 53284 35000 53340
rect 35048 53284 35104 53340
rect 35152 53284 35208 53340
rect 3500 53116 3556 53172
rect 7420 53116 7476 53172
rect 6300 53004 6356 53060
rect 5292 52780 5348 52836
rect 4008 52500 4064 52556
rect 4112 52500 4168 52556
rect 4216 52500 4272 52556
rect 4320 52500 4376 52556
rect 4424 52500 4480 52556
rect 4528 52500 4584 52556
rect 4632 52500 4688 52556
rect 4736 52500 4792 52556
rect 4840 52500 4896 52556
rect 4944 52500 5000 52556
rect 5048 52500 5104 52556
rect 5152 52500 5208 52556
rect 24008 52500 24064 52556
rect 24112 52500 24168 52556
rect 24216 52500 24272 52556
rect 24320 52500 24376 52556
rect 24424 52500 24480 52556
rect 24528 52500 24584 52556
rect 24632 52500 24688 52556
rect 24736 52500 24792 52556
rect 24840 52500 24896 52556
rect 24944 52500 25000 52556
rect 25048 52500 25104 52556
rect 25152 52500 25208 52556
rect 13468 52444 13524 52500
rect 11900 52108 11956 52164
rect 14008 51716 14064 51772
rect 14112 51716 14168 51772
rect 14216 51716 14272 51772
rect 14320 51716 14376 51772
rect 14424 51716 14480 51772
rect 14528 51716 14584 51772
rect 14632 51716 14688 51772
rect 14736 51716 14792 51772
rect 14840 51716 14896 51772
rect 14944 51716 15000 51772
rect 15048 51716 15104 51772
rect 15152 51716 15208 51772
rect 34008 51716 34064 51772
rect 34112 51716 34168 51772
rect 34216 51716 34272 51772
rect 34320 51716 34376 51772
rect 34424 51716 34480 51772
rect 34528 51716 34584 51772
rect 34632 51716 34688 51772
rect 34736 51716 34792 51772
rect 34840 51716 34896 51772
rect 34944 51716 35000 51772
rect 35048 51716 35104 51772
rect 35152 51716 35208 51772
rect 3500 51660 3556 51716
rect 5292 51660 5348 51716
rect 13804 51660 13860 51716
rect 13580 51548 13636 51604
rect 4008 50932 4064 50988
rect 4112 50932 4168 50988
rect 4216 50932 4272 50988
rect 4320 50932 4376 50988
rect 4424 50932 4480 50988
rect 4528 50932 4584 50988
rect 4632 50932 4688 50988
rect 4736 50932 4792 50988
rect 4840 50932 4896 50988
rect 4944 50932 5000 50988
rect 5048 50932 5104 50988
rect 5152 50932 5208 50988
rect 24008 50932 24064 50988
rect 24112 50932 24168 50988
rect 24216 50932 24272 50988
rect 24320 50932 24376 50988
rect 24424 50932 24480 50988
rect 24528 50932 24584 50988
rect 24632 50932 24688 50988
rect 24736 50932 24792 50988
rect 24840 50932 24896 50988
rect 24944 50932 25000 50988
rect 25048 50932 25104 50988
rect 25152 50932 25208 50988
rect 19628 50652 19684 50708
rect 13804 50540 13860 50596
rect 33852 50428 33908 50484
rect 14008 50148 14064 50204
rect 14112 50148 14168 50204
rect 14216 50148 14272 50204
rect 14320 50148 14376 50204
rect 14424 50148 14480 50204
rect 14528 50148 14584 50204
rect 14632 50148 14688 50204
rect 14736 50148 14792 50204
rect 14840 50148 14896 50204
rect 14944 50148 15000 50204
rect 15048 50148 15104 50204
rect 15152 50148 15208 50204
rect 34008 50148 34064 50204
rect 34112 50148 34168 50204
rect 34216 50148 34272 50204
rect 34320 50148 34376 50204
rect 34424 50148 34480 50204
rect 34528 50148 34584 50204
rect 34632 50148 34688 50204
rect 34736 50148 34792 50204
rect 34840 50148 34896 50204
rect 34944 50148 35000 50204
rect 35048 50148 35104 50204
rect 35152 50148 35208 50204
rect 4008 49364 4064 49420
rect 4112 49364 4168 49420
rect 4216 49364 4272 49420
rect 4320 49364 4376 49420
rect 4424 49364 4480 49420
rect 4528 49364 4584 49420
rect 4632 49364 4688 49420
rect 4736 49364 4792 49420
rect 4840 49364 4896 49420
rect 4944 49364 5000 49420
rect 5048 49364 5104 49420
rect 5152 49364 5208 49420
rect 24008 49364 24064 49420
rect 24112 49364 24168 49420
rect 24216 49364 24272 49420
rect 24320 49364 24376 49420
rect 24424 49364 24480 49420
rect 24528 49364 24584 49420
rect 24632 49364 24688 49420
rect 24736 49364 24792 49420
rect 24840 49364 24896 49420
rect 24944 49364 25000 49420
rect 25048 49364 25104 49420
rect 25152 49364 25208 49420
rect 13804 48972 13860 49028
rect 33852 48748 33908 48804
rect 14008 48580 14064 48636
rect 14112 48580 14168 48636
rect 14216 48580 14272 48636
rect 14320 48580 14376 48636
rect 14424 48580 14480 48636
rect 14528 48580 14584 48636
rect 14632 48580 14688 48636
rect 14736 48580 14792 48636
rect 14840 48580 14896 48636
rect 14944 48580 15000 48636
rect 15048 48580 15104 48636
rect 15152 48580 15208 48636
rect 34008 48580 34064 48636
rect 34112 48580 34168 48636
rect 34216 48580 34272 48636
rect 34320 48580 34376 48636
rect 34424 48580 34480 48636
rect 34528 48580 34584 48636
rect 34632 48580 34688 48636
rect 34736 48580 34792 48636
rect 34840 48580 34896 48636
rect 34944 48580 35000 48636
rect 35048 48580 35104 48636
rect 35152 48580 35208 48636
rect 5292 48076 5348 48132
rect 4008 47796 4064 47852
rect 4112 47796 4168 47852
rect 4216 47796 4272 47852
rect 4320 47796 4376 47852
rect 4424 47796 4480 47852
rect 4528 47796 4584 47852
rect 4632 47796 4688 47852
rect 4736 47796 4792 47852
rect 4840 47796 4896 47852
rect 4944 47796 5000 47852
rect 5048 47796 5104 47852
rect 5152 47796 5208 47852
rect 24008 47796 24064 47852
rect 24112 47796 24168 47852
rect 24216 47796 24272 47852
rect 24320 47796 24376 47852
rect 24424 47796 24480 47852
rect 24528 47796 24584 47852
rect 24632 47796 24688 47852
rect 24736 47796 24792 47852
rect 24840 47796 24896 47852
rect 24944 47796 25000 47852
rect 25048 47796 25104 47852
rect 25152 47796 25208 47852
rect 3388 47516 3444 47572
rect 10108 47404 10164 47460
rect 13804 47404 13860 47460
rect 5292 47068 5348 47124
rect 14008 47012 14064 47068
rect 14112 47012 14168 47068
rect 14216 47012 14272 47068
rect 14320 47012 14376 47068
rect 14424 47012 14480 47068
rect 14528 47012 14584 47068
rect 14632 47012 14688 47068
rect 14736 47012 14792 47068
rect 14840 47012 14896 47068
rect 14944 47012 15000 47068
rect 15048 47012 15104 47068
rect 15152 47012 15208 47068
rect 34008 47012 34064 47068
rect 34112 47012 34168 47068
rect 34216 47012 34272 47068
rect 34320 47012 34376 47068
rect 34424 47012 34480 47068
rect 34528 47012 34584 47068
rect 34632 47012 34688 47068
rect 34736 47012 34792 47068
rect 34840 47012 34896 47068
rect 34944 47012 35000 47068
rect 35048 47012 35104 47068
rect 35152 47012 35208 47068
rect 15372 46956 15428 47012
rect 17612 46508 17668 46564
rect 4008 46228 4064 46284
rect 4112 46228 4168 46284
rect 4216 46228 4272 46284
rect 4320 46228 4376 46284
rect 4424 46228 4480 46284
rect 4528 46228 4584 46284
rect 4632 46228 4688 46284
rect 4736 46228 4792 46284
rect 4840 46228 4896 46284
rect 4944 46228 5000 46284
rect 5048 46228 5104 46284
rect 5152 46228 5208 46284
rect 24008 46228 24064 46284
rect 24112 46228 24168 46284
rect 24216 46228 24272 46284
rect 24320 46228 24376 46284
rect 24424 46228 24480 46284
rect 24528 46228 24584 46284
rect 24632 46228 24688 46284
rect 24736 46228 24792 46284
rect 24840 46228 24896 46284
rect 24944 46228 25000 46284
rect 25048 46228 25104 46284
rect 25152 46228 25208 46284
rect 25788 45948 25844 46004
rect 17612 45724 17668 45780
rect 14008 45444 14064 45500
rect 14112 45444 14168 45500
rect 14216 45444 14272 45500
rect 14320 45444 14376 45500
rect 14424 45444 14480 45500
rect 14528 45444 14584 45500
rect 14632 45444 14688 45500
rect 14736 45444 14792 45500
rect 14840 45444 14896 45500
rect 14944 45444 15000 45500
rect 15048 45444 15104 45500
rect 15152 45444 15208 45500
rect 34008 45444 34064 45500
rect 34112 45444 34168 45500
rect 34216 45444 34272 45500
rect 34320 45444 34376 45500
rect 34424 45444 34480 45500
rect 34528 45444 34584 45500
rect 34632 45444 34688 45500
rect 34736 45444 34792 45500
rect 34840 45444 34896 45500
rect 34944 45444 35000 45500
rect 35048 45444 35104 45500
rect 35152 45444 35208 45500
rect 13692 45276 13748 45332
rect 5964 44828 6020 44884
rect 4008 44660 4064 44716
rect 4112 44660 4168 44716
rect 4216 44660 4272 44716
rect 4320 44660 4376 44716
rect 4424 44660 4480 44716
rect 4528 44660 4584 44716
rect 4632 44660 4688 44716
rect 4736 44660 4792 44716
rect 4840 44660 4896 44716
rect 4944 44660 5000 44716
rect 5048 44660 5104 44716
rect 5152 44660 5208 44716
rect 3836 44492 3892 44548
rect 24008 44660 24064 44716
rect 24112 44660 24168 44716
rect 24216 44660 24272 44716
rect 24320 44660 24376 44716
rect 24424 44660 24480 44716
rect 24528 44660 24584 44716
rect 24632 44660 24688 44716
rect 24736 44660 24792 44716
rect 24840 44660 24896 44716
rect 24944 44660 25000 44716
rect 25048 44660 25104 44716
rect 25152 44660 25208 44716
rect 23772 44380 23828 44436
rect 33516 44268 33572 44324
rect 33628 44044 33684 44100
rect 3388 43932 3444 43988
rect 14008 43876 14064 43932
rect 14112 43876 14168 43932
rect 14216 43876 14272 43932
rect 14320 43876 14376 43932
rect 14424 43876 14480 43932
rect 14528 43876 14584 43932
rect 14632 43876 14688 43932
rect 14736 43876 14792 43932
rect 14840 43876 14896 43932
rect 14944 43876 15000 43932
rect 15048 43876 15104 43932
rect 15152 43876 15208 43932
rect 34008 43876 34064 43932
rect 34112 43876 34168 43932
rect 34216 43876 34272 43932
rect 34320 43876 34376 43932
rect 34424 43876 34480 43932
rect 34528 43876 34584 43932
rect 34632 43876 34688 43932
rect 34736 43876 34792 43932
rect 34840 43876 34896 43932
rect 34944 43876 35000 43932
rect 35048 43876 35104 43932
rect 35152 43876 35208 43932
rect 3388 43596 3444 43652
rect 33516 43372 33572 43428
rect 4008 43092 4064 43148
rect 4112 43092 4168 43148
rect 4216 43092 4272 43148
rect 4320 43092 4376 43148
rect 4424 43092 4480 43148
rect 4528 43092 4584 43148
rect 4632 43092 4688 43148
rect 4736 43092 4792 43148
rect 4840 43092 4896 43148
rect 4944 43092 5000 43148
rect 5048 43092 5104 43148
rect 5152 43092 5208 43148
rect 24008 43092 24064 43148
rect 24112 43092 24168 43148
rect 24216 43092 24272 43148
rect 24320 43092 24376 43148
rect 24424 43092 24480 43148
rect 24528 43092 24584 43148
rect 24632 43092 24688 43148
rect 24736 43092 24792 43148
rect 24840 43092 24896 43148
rect 24944 43092 25000 43148
rect 25048 43092 25104 43148
rect 25152 43092 25208 43148
rect 33404 43036 33460 43092
rect 23548 42812 23604 42868
rect 33628 42812 33684 42868
rect 14008 42308 14064 42364
rect 14112 42308 14168 42364
rect 14216 42308 14272 42364
rect 14320 42308 14376 42364
rect 14424 42308 14480 42364
rect 14528 42308 14584 42364
rect 14632 42308 14688 42364
rect 14736 42308 14792 42364
rect 14840 42308 14896 42364
rect 14944 42308 15000 42364
rect 15048 42308 15104 42364
rect 15152 42308 15208 42364
rect 34008 42308 34064 42364
rect 34112 42308 34168 42364
rect 34216 42308 34272 42364
rect 34320 42308 34376 42364
rect 34424 42308 34480 42364
rect 34528 42308 34584 42364
rect 34632 42308 34688 42364
rect 34736 42308 34792 42364
rect 34840 42308 34896 42364
rect 34944 42308 35000 42364
rect 35048 42308 35104 42364
rect 35152 42308 35208 42364
rect 4008 41524 4064 41580
rect 4112 41524 4168 41580
rect 4216 41524 4272 41580
rect 4320 41524 4376 41580
rect 4424 41524 4480 41580
rect 4528 41524 4584 41580
rect 4632 41524 4688 41580
rect 4736 41524 4792 41580
rect 4840 41524 4896 41580
rect 4944 41524 5000 41580
rect 5048 41524 5104 41580
rect 5152 41524 5208 41580
rect 24008 41524 24064 41580
rect 24112 41524 24168 41580
rect 24216 41524 24272 41580
rect 24320 41524 24376 41580
rect 24424 41524 24480 41580
rect 24528 41524 24584 41580
rect 24632 41524 24688 41580
rect 24736 41524 24792 41580
rect 24840 41524 24896 41580
rect 24944 41524 25000 41580
rect 25048 41524 25104 41580
rect 25152 41524 25208 41580
rect 33740 41468 33796 41524
rect 33852 41020 33908 41076
rect 14008 40740 14064 40796
rect 14112 40740 14168 40796
rect 14216 40740 14272 40796
rect 14320 40740 14376 40796
rect 14424 40740 14480 40796
rect 14528 40740 14584 40796
rect 14632 40740 14688 40796
rect 14736 40740 14792 40796
rect 14840 40740 14896 40796
rect 14944 40740 15000 40796
rect 15048 40740 15104 40796
rect 15152 40740 15208 40796
rect 34008 40740 34064 40796
rect 34112 40740 34168 40796
rect 34216 40740 34272 40796
rect 34320 40740 34376 40796
rect 34424 40740 34480 40796
rect 34528 40740 34584 40796
rect 34632 40740 34688 40796
rect 34736 40740 34792 40796
rect 34840 40740 34896 40796
rect 34944 40740 35000 40796
rect 35048 40740 35104 40796
rect 35152 40740 35208 40796
rect 23660 40684 23716 40740
rect 33740 40572 33796 40628
rect 25788 40348 25844 40404
rect 4008 39956 4064 40012
rect 4112 39956 4168 40012
rect 4216 39956 4272 40012
rect 4320 39956 4376 40012
rect 4424 39956 4480 40012
rect 4528 39956 4584 40012
rect 4632 39956 4688 40012
rect 4736 39956 4792 40012
rect 4840 39956 4896 40012
rect 4944 39956 5000 40012
rect 5048 39956 5104 40012
rect 5152 39956 5208 40012
rect 24008 39956 24064 40012
rect 24112 39956 24168 40012
rect 24216 39956 24272 40012
rect 24320 39956 24376 40012
rect 24424 39956 24480 40012
rect 24528 39956 24584 40012
rect 24632 39956 24688 40012
rect 24736 39956 24792 40012
rect 24840 39956 24896 40012
rect 24944 39956 25000 40012
rect 25048 39956 25104 40012
rect 25152 39956 25208 40012
rect 23548 39676 23604 39732
rect 33628 39676 33684 39732
rect 3836 39564 3892 39620
rect 23100 39564 23156 39620
rect 23660 39564 23716 39620
rect 5964 39452 6020 39508
rect 14008 39172 14064 39228
rect 14112 39172 14168 39228
rect 14216 39172 14272 39228
rect 14320 39172 14376 39228
rect 14424 39172 14480 39228
rect 14528 39172 14584 39228
rect 14632 39172 14688 39228
rect 14736 39172 14792 39228
rect 14840 39172 14896 39228
rect 14944 39172 15000 39228
rect 15048 39172 15104 39228
rect 15152 39172 15208 39228
rect 34008 39172 34064 39228
rect 34112 39172 34168 39228
rect 34216 39172 34272 39228
rect 34320 39172 34376 39228
rect 34424 39172 34480 39228
rect 34528 39172 34584 39228
rect 34632 39172 34688 39228
rect 34736 39172 34792 39228
rect 34840 39172 34896 39228
rect 34944 39172 35000 39228
rect 35048 39172 35104 39228
rect 35152 39172 35208 39228
rect 33852 39004 33908 39060
rect 17612 38444 17668 38500
rect 33516 38444 33572 38500
rect 33852 38444 33908 38500
rect 4008 38388 4064 38444
rect 4112 38388 4168 38444
rect 4216 38388 4272 38444
rect 4320 38388 4376 38444
rect 4424 38388 4480 38444
rect 4528 38388 4584 38444
rect 4632 38388 4688 38444
rect 4736 38388 4792 38444
rect 4840 38388 4896 38444
rect 4944 38388 5000 38444
rect 5048 38388 5104 38444
rect 5152 38388 5208 38444
rect 24008 38388 24064 38444
rect 24112 38388 24168 38444
rect 24216 38388 24272 38444
rect 24320 38388 24376 38444
rect 24424 38388 24480 38444
rect 24528 38388 24584 38444
rect 24632 38388 24688 38444
rect 24736 38388 24792 38444
rect 24840 38388 24896 38444
rect 24944 38388 25000 38444
rect 25048 38388 25104 38444
rect 25152 38388 25208 38444
rect 33404 37660 33460 37716
rect 14008 37604 14064 37660
rect 14112 37604 14168 37660
rect 14216 37604 14272 37660
rect 14320 37604 14376 37660
rect 14424 37604 14480 37660
rect 14528 37604 14584 37660
rect 14632 37604 14688 37660
rect 14736 37604 14792 37660
rect 14840 37604 14896 37660
rect 14944 37604 15000 37660
rect 15048 37604 15104 37660
rect 15152 37604 15208 37660
rect 34008 37604 34064 37660
rect 34112 37604 34168 37660
rect 34216 37604 34272 37660
rect 34320 37604 34376 37660
rect 34424 37604 34480 37660
rect 34528 37604 34584 37660
rect 34632 37604 34688 37660
rect 34736 37604 34792 37660
rect 34840 37604 34896 37660
rect 34944 37604 35000 37660
rect 35048 37604 35104 37660
rect 35152 37604 35208 37660
rect 23772 37324 23828 37380
rect 27020 37324 27076 37380
rect 4008 36820 4064 36876
rect 4112 36820 4168 36876
rect 4216 36820 4272 36876
rect 4320 36820 4376 36876
rect 4424 36820 4480 36876
rect 4528 36820 4584 36876
rect 4632 36820 4688 36876
rect 4736 36820 4792 36876
rect 4840 36820 4896 36876
rect 4944 36820 5000 36876
rect 5048 36820 5104 36876
rect 5152 36820 5208 36876
rect 24008 36820 24064 36876
rect 24112 36820 24168 36876
rect 24216 36820 24272 36876
rect 24320 36820 24376 36876
rect 24424 36820 24480 36876
rect 24528 36820 24584 36876
rect 24632 36820 24688 36876
rect 24736 36820 24792 36876
rect 24840 36820 24896 36876
rect 24944 36820 25000 36876
rect 25048 36820 25104 36876
rect 25152 36820 25208 36876
rect 23100 36204 23156 36260
rect 14008 36036 14064 36092
rect 14112 36036 14168 36092
rect 14216 36036 14272 36092
rect 14320 36036 14376 36092
rect 14424 36036 14480 36092
rect 14528 36036 14584 36092
rect 14632 36036 14688 36092
rect 14736 36036 14792 36092
rect 14840 36036 14896 36092
rect 14944 36036 15000 36092
rect 15048 36036 15104 36092
rect 15152 36036 15208 36092
rect 34008 36036 34064 36092
rect 34112 36036 34168 36092
rect 34216 36036 34272 36092
rect 34320 36036 34376 36092
rect 34424 36036 34480 36092
rect 34528 36036 34584 36092
rect 34632 36036 34688 36092
rect 34736 36036 34792 36092
rect 34840 36036 34896 36092
rect 34944 36036 35000 36092
rect 35048 36036 35104 36092
rect 35152 36036 35208 36092
rect 4008 35252 4064 35308
rect 4112 35252 4168 35308
rect 4216 35252 4272 35308
rect 4320 35252 4376 35308
rect 4424 35252 4480 35308
rect 4528 35252 4584 35308
rect 4632 35252 4688 35308
rect 4736 35252 4792 35308
rect 4840 35252 4896 35308
rect 4944 35252 5000 35308
rect 5048 35252 5104 35308
rect 5152 35252 5208 35308
rect 24008 35252 24064 35308
rect 24112 35252 24168 35308
rect 24216 35252 24272 35308
rect 24320 35252 24376 35308
rect 24424 35252 24480 35308
rect 24528 35252 24584 35308
rect 24632 35252 24688 35308
rect 24736 35252 24792 35308
rect 24840 35252 24896 35308
rect 24944 35252 25000 35308
rect 25048 35252 25104 35308
rect 25152 35252 25208 35308
rect 13804 35084 13860 35140
rect 7308 34972 7364 35028
rect 13692 34972 13748 35028
rect 33628 34860 33684 34916
rect 33852 34636 33908 34692
rect 14008 34468 14064 34524
rect 14112 34468 14168 34524
rect 14216 34468 14272 34524
rect 14320 34468 14376 34524
rect 14424 34468 14480 34524
rect 14528 34468 14584 34524
rect 14632 34468 14688 34524
rect 14736 34468 14792 34524
rect 14840 34468 14896 34524
rect 14944 34468 15000 34524
rect 15048 34468 15104 34524
rect 15152 34468 15208 34524
rect 34008 34468 34064 34524
rect 34112 34468 34168 34524
rect 34216 34468 34272 34524
rect 34320 34468 34376 34524
rect 34424 34468 34480 34524
rect 34528 34468 34584 34524
rect 34632 34468 34688 34524
rect 34736 34468 34792 34524
rect 34840 34468 34896 34524
rect 34944 34468 35000 34524
rect 35048 34468 35104 34524
rect 35152 34468 35208 34524
rect 33628 34188 33684 34244
rect 4008 33684 4064 33740
rect 4112 33684 4168 33740
rect 4216 33684 4272 33740
rect 4320 33684 4376 33740
rect 4424 33684 4480 33740
rect 4528 33684 4584 33740
rect 4632 33684 4688 33740
rect 4736 33684 4792 33740
rect 4840 33684 4896 33740
rect 4944 33684 5000 33740
rect 5048 33684 5104 33740
rect 5152 33684 5208 33740
rect 24008 33684 24064 33740
rect 24112 33684 24168 33740
rect 24216 33684 24272 33740
rect 24320 33684 24376 33740
rect 24424 33684 24480 33740
rect 24528 33684 24584 33740
rect 24632 33684 24688 33740
rect 24736 33684 24792 33740
rect 24840 33684 24896 33740
rect 24944 33684 25000 33740
rect 25048 33684 25104 33740
rect 25152 33684 25208 33740
rect 3500 33628 3556 33684
rect 5292 33516 5348 33572
rect 27020 32956 27076 33012
rect 33740 32956 33796 33012
rect 14008 32900 14064 32956
rect 14112 32900 14168 32956
rect 14216 32900 14272 32956
rect 14320 32900 14376 32956
rect 14424 32900 14480 32956
rect 14528 32900 14584 32956
rect 14632 32900 14688 32956
rect 14736 32900 14792 32956
rect 14840 32900 14896 32956
rect 14944 32900 15000 32956
rect 15048 32900 15104 32956
rect 15152 32900 15208 32956
rect 34008 32900 34064 32956
rect 34112 32900 34168 32956
rect 34216 32900 34272 32956
rect 34320 32900 34376 32956
rect 34424 32900 34480 32956
rect 34528 32900 34584 32956
rect 34632 32900 34688 32956
rect 34736 32900 34792 32956
rect 34840 32900 34896 32956
rect 34944 32900 35000 32956
rect 35048 32900 35104 32956
rect 35152 32900 35208 32956
rect 15484 32732 15540 32788
rect 1820 32508 1876 32564
rect 4008 32116 4064 32172
rect 4112 32116 4168 32172
rect 4216 32116 4272 32172
rect 4320 32116 4376 32172
rect 4424 32116 4480 32172
rect 4528 32116 4584 32172
rect 4632 32116 4688 32172
rect 4736 32116 4792 32172
rect 4840 32116 4896 32172
rect 4944 32116 5000 32172
rect 5048 32116 5104 32172
rect 5152 32116 5208 32172
rect 24008 32116 24064 32172
rect 24112 32116 24168 32172
rect 24216 32116 24272 32172
rect 24320 32116 24376 32172
rect 24424 32116 24480 32172
rect 24528 32116 24584 32172
rect 24632 32116 24688 32172
rect 24736 32116 24792 32172
rect 24840 32116 24896 32172
rect 24944 32116 25000 32172
rect 25048 32116 25104 32172
rect 25152 32116 25208 32172
rect 3836 32060 3892 32116
rect 15372 31612 15428 31668
rect 26572 31500 26628 31556
rect 14008 31332 14064 31388
rect 14112 31332 14168 31388
rect 14216 31332 14272 31388
rect 14320 31332 14376 31388
rect 14424 31332 14480 31388
rect 14528 31332 14584 31388
rect 14632 31332 14688 31388
rect 14736 31332 14792 31388
rect 14840 31332 14896 31388
rect 14944 31332 15000 31388
rect 15048 31332 15104 31388
rect 15152 31332 15208 31388
rect 34008 31332 34064 31388
rect 34112 31332 34168 31388
rect 34216 31332 34272 31388
rect 34320 31332 34376 31388
rect 34424 31332 34480 31388
rect 34528 31332 34584 31388
rect 34632 31332 34688 31388
rect 34736 31332 34792 31388
rect 34840 31332 34896 31388
rect 34944 31332 35000 31388
rect 35048 31332 35104 31388
rect 35152 31332 35208 31388
rect 4008 30548 4064 30604
rect 4112 30548 4168 30604
rect 4216 30548 4272 30604
rect 4320 30548 4376 30604
rect 4424 30548 4480 30604
rect 4528 30548 4584 30604
rect 4632 30548 4688 30604
rect 4736 30548 4792 30604
rect 4840 30548 4896 30604
rect 4944 30548 5000 30604
rect 5048 30548 5104 30604
rect 5152 30548 5208 30604
rect 24008 30548 24064 30604
rect 24112 30548 24168 30604
rect 24216 30548 24272 30604
rect 24320 30548 24376 30604
rect 24424 30548 24480 30604
rect 24528 30548 24584 30604
rect 24632 30548 24688 30604
rect 24736 30548 24792 30604
rect 24840 30548 24896 30604
rect 24944 30548 25000 30604
rect 25048 30548 25104 30604
rect 25152 30548 25208 30604
rect 3164 30156 3220 30212
rect 5292 30156 5348 30212
rect 13468 29932 13524 29988
rect 14008 29764 14064 29820
rect 14112 29764 14168 29820
rect 14216 29764 14272 29820
rect 14320 29764 14376 29820
rect 14424 29764 14480 29820
rect 14528 29764 14584 29820
rect 14632 29764 14688 29820
rect 14736 29764 14792 29820
rect 14840 29764 14896 29820
rect 14944 29764 15000 29820
rect 15048 29764 15104 29820
rect 15152 29764 15208 29820
rect 34008 29764 34064 29820
rect 34112 29764 34168 29820
rect 34216 29764 34272 29820
rect 34320 29764 34376 29820
rect 34424 29764 34480 29820
rect 34528 29764 34584 29820
rect 34632 29764 34688 29820
rect 34736 29764 34792 29820
rect 34840 29764 34896 29820
rect 34944 29764 35000 29820
rect 35048 29764 35104 29820
rect 35152 29764 35208 29820
rect 15484 29596 15540 29652
rect 4008 28980 4064 29036
rect 4112 28980 4168 29036
rect 4216 28980 4272 29036
rect 4320 28980 4376 29036
rect 4424 28980 4480 29036
rect 4528 28980 4584 29036
rect 4632 28980 4688 29036
rect 4736 28980 4792 29036
rect 4840 28980 4896 29036
rect 4944 28980 5000 29036
rect 5048 28980 5104 29036
rect 5152 28980 5208 29036
rect 24008 28980 24064 29036
rect 24112 28980 24168 29036
rect 24216 28980 24272 29036
rect 24320 28980 24376 29036
rect 24424 28980 24480 29036
rect 24528 28980 24584 29036
rect 24632 28980 24688 29036
rect 24736 28980 24792 29036
rect 24840 28980 24896 29036
rect 24944 28980 25000 29036
rect 25048 28980 25104 29036
rect 25152 28980 25208 29036
rect 3612 28812 3668 28868
rect 3836 28588 3892 28644
rect 6076 28476 6132 28532
rect 3612 28364 3668 28420
rect 13468 28252 13524 28308
rect 14008 28196 14064 28252
rect 14112 28196 14168 28252
rect 14216 28196 14272 28252
rect 14320 28196 14376 28252
rect 14424 28196 14480 28252
rect 14528 28196 14584 28252
rect 14632 28196 14688 28252
rect 14736 28196 14792 28252
rect 14840 28196 14896 28252
rect 14944 28196 15000 28252
rect 15048 28196 15104 28252
rect 15152 28196 15208 28252
rect 34008 28196 34064 28252
rect 34112 28196 34168 28252
rect 34216 28196 34272 28252
rect 34320 28196 34376 28252
rect 34424 28196 34480 28252
rect 34528 28196 34584 28252
rect 34632 28196 34688 28252
rect 34736 28196 34792 28252
rect 34840 28196 34896 28252
rect 34944 28196 35000 28252
rect 35048 28196 35104 28252
rect 35152 28196 35208 28252
rect 4008 27412 4064 27468
rect 4112 27412 4168 27468
rect 4216 27412 4272 27468
rect 4320 27412 4376 27468
rect 4424 27412 4480 27468
rect 4528 27412 4584 27468
rect 4632 27412 4688 27468
rect 4736 27412 4792 27468
rect 4840 27412 4896 27468
rect 4944 27412 5000 27468
rect 5048 27412 5104 27468
rect 5152 27412 5208 27468
rect 24008 27412 24064 27468
rect 24112 27412 24168 27468
rect 24216 27412 24272 27468
rect 24320 27412 24376 27468
rect 24424 27412 24480 27468
rect 24528 27412 24584 27468
rect 24632 27412 24688 27468
rect 24736 27412 24792 27468
rect 24840 27412 24896 27468
rect 24944 27412 25000 27468
rect 25048 27412 25104 27468
rect 25152 27412 25208 27468
rect 5964 27356 6020 27412
rect 3276 27020 3332 27076
rect 6188 27020 6244 27076
rect 13804 27020 13860 27076
rect 3388 26908 3444 26964
rect 7308 26908 7364 26964
rect 5964 26796 6020 26852
rect 14008 26628 14064 26684
rect 14112 26628 14168 26684
rect 14216 26628 14272 26684
rect 14320 26628 14376 26684
rect 14424 26628 14480 26684
rect 14528 26628 14584 26684
rect 14632 26628 14688 26684
rect 14736 26628 14792 26684
rect 14840 26628 14896 26684
rect 14944 26628 15000 26684
rect 15048 26628 15104 26684
rect 15152 26628 15208 26684
rect 34008 26628 34064 26684
rect 34112 26628 34168 26684
rect 34216 26628 34272 26684
rect 34320 26628 34376 26684
rect 34424 26628 34480 26684
rect 34528 26628 34584 26684
rect 34632 26628 34688 26684
rect 34736 26628 34792 26684
rect 34840 26628 34896 26684
rect 34944 26628 35000 26684
rect 35048 26628 35104 26684
rect 35152 26628 35208 26684
rect 1820 26572 1876 26628
rect 6076 26572 6132 26628
rect 3836 26460 3892 26516
rect 4008 25844 4064 25900
rect 4112 25844 4168 25900
rect 4216 25844 4272 25900
rect 4320 25844 4376 25900
rect 4424 25844 4480 25900
rect 4528 25844 4584 25900
rect 4632 25844 4688 25900
rect 4736 25844 4792 25900
rect 4840 25844 4896 25900
rect 4944 25844 5000 25900
rect 5048 25844 5104 25900
rect 5152 25844 5208 25900
rect 24008 25844 24064 25900
rect 24112 25844 24168 25900
rect 24216 25844 24272 25900
rect 24320 25844 24376 25900
rect 24424 25844 24480 25900
rect 24528 25844 24584 25900
rect 24632 25844 24688 25900
rect 24736 25844 24792 25900
rect 24840 25844 24896 25900
rect 24944 25844 25000 25900
rect 25048 25844 25104 25900
rect 25152 25844 25208 25900
rect 3164 25788 3220 25844
rect 3500 25676 3556 25732
rect 3836 25564 3892 25620
rect 13692 25564 13748 25620
rect 5292 25340 5348 25396
rect 26572 25116 26628 25172
rect 14008 25060 14064 25116
rect 14112 25060 14168 25116
rect 14216 25060 14272 25116
rect 14320 25060 14376 25116
rect 14424 25060 14480 25116
rect 14528 25060 14584 25116
rect 14632 25060 14688 25116
rect 14736 25060 14792 25116
rect 14840 25060 14896 25116
rect 14944 25060 15000 25116
rect 15048 25060 15104 25116
rect 15152 25060 15208 25116
rect 34008 25060 34064 25116
rect 34112 25060 34168 25116
rect 34216 25060 34272 25116
rect 34320 25060 34376 25116
rect 34424 25060 34480 25116
rect 34528 25060 34584 25116
rect 34632 25060 34688 25116
rect 34736 25060 34792 25116
rect 34840 25060 34896 25116
rect 34944 25060 35000 25116
rect 35048 25060 35104 25116
rect 35152 25060 35208 25116
rect 6188 24892 6244 24948
rect 3164 24668 3220 24724
rect 4008 24276 4064 24332
rect 4112 24276 4168 24332
rect 4216 24276 4272 24332
rect 4320 24276 4376 24332
rect 4424 24276 4480 24332
rect 4528 24276 4584 24332
rect 4632 24276 4688 24332
rect 4736 24276 4792 24332
rect 4840 24276 4896 24332
rect 4944 24276 5000 24332
rect 5048 24276 5104 24332
rect 5152 24276 5208 24332
rect 24008 24276 24064 24332
rect 24112 24276 24168 24332
rect 24216 24276 24272 24332
rect 24320 24276 24376 24332
rect 24424 24276 24480 24332
rect 24528 24276 24584 24332
rect 24632 24276 24688 24332
rect 24736 24276 24792 24332
rect 24840 24276 24896 24332
rect 24944 24276 25000 24332
rect 25048 24276 25104 24332
rect 25152 24276 25208 24332
rect 13804 23772 13860 23828
rect 3276 23660 3332 23716
rect 14008 23492 14064 23548
rect 14112 23492 14168 23548
rect 14216 23492 14272 23548
rect 14320 23492 14376 23548
rect 14424 23492 14480 23548
rect 14528 23492 14584 23548
rect 14632 23492 14688 23548
rect 14736 23492 14792 23548
rect 14840 23492 14896 23548
rect 14944 23492 15000 23548
rect 15048 23492 15104 23548
rect 15152 23492 15208 23548
rect 34008 23492 34064 23548
rect 34112 23492 34168 23548
rect 34216 23492 34272 23548
rect 34320 23492 34376 23548
rect 34424 23492 34480 23548
rect 34528 23492 34584 23548
rect 34632 23492 34688 23548
rect 34736 23492 34792 23548
rect 34840 23492 34896 23548
rect 34944 23492 35000 23548
rect 35048 23492 35104 23548
rect 35152 23492 35208 23548
rect 3052 23436 3108 23492
rect 13692 23436 13748 23492
rect 3836 23212 3892 23268
rect 13804 23100 13860 23156
rect 5292 22876 5348 22932
rect 13692 22876 13748 22932
rect 4008 22708 4064 22764
rect 4112 22708 4168 22764
rect 4216 22708 4272 22764
rect 4320 22708 4376 22764
rect 4424 22708 4480 22764
rect 4528 22708 4584 22764
rect 4632 22708 4688 22764
rect 4736 22708 4792 22764
rect 4840 22708 4896 22764
rect 4944 22708 5000 22764
rect 5048 22708 5104 22764
rect 5152 22708 5208 22764
rect 24008 22708 24064 22764
rect 24112 22708 24168 22764
rect 24216 22708 24272 22764
rect 24320 22708 24376 22764
rect 24424 22708 24480 22764
rect 24528 22708 24584 22764
rect 24632 22708 24688 22764
rect 24736 22708 24792 22764
rect 24840 22708 24896 22764
rect 24944 22708 25000 22764
rect 25048 22708 25104 22764
rect 25152 22708 25208 22764
rect 13804 22652 13860 22708
rect 13692 22540 13748 22596
rect 13692 22204 13748 22260
rect 25340 22204 25396 22260
rect 14008 21924 14064 21980
rect 14112 21924 14168 21980
rect 14216 21924 14272 21980
rect 14320 21924 14376 21980
rect 14424 21924 14480 21980
rect 14528 21924 14584 21980
rect 14632 21924 14688 21980
rect 14736 21924 14792 21980
rect 14840 21924 14896 21980
rect 14944 21924 15000 21980
rect 15048 21924 15104 21980
rect 15152 21924 15208 21980
rect 34008 21924 34064 21980
rect 34112 21924 34168 21980
rect 34216 21924 34272 21980
rect 34320 21924 34376 21980
rect 34424 21924 34480 21980
rect 34528 21924 34584 21980
rect 34632 21924 34688 21980
rect 34736 21924 34792 21980
rect 34840 21924 34896 21980
rect 34944 21924 35000 21980
rect 35048 21924 35104 21980
rect 35152 21924 35208 21980
rect 6188 21756 6244 21812
rect 5404 21420 5460 21476
rect 4008 21140 4064 21196
rect 4112 21140 4168 21196
rect 4216 21140 4272 21196
rect 4320 21140 4376 21196
rect 4424 21140 4480 21196
rect 4528 21140 4584 21196
rect 4632 21140 4688 21196
rect 4736 21140 4792 21196
rect 4840 21140 4896 21196
rect 4944 21140 5000 21196
rect 5048 21140 5104 21196
rect 5152 21140 5208 21196
rect 24008 21140 24064 21196
rect 24112 21140 24168 21196
rect 24216 21140 24272 21196
rect 24320 21140 24376 21196
rect 24424 21140 24480 21196
rect 24528 21140 24584 21196
rect 24632 21140 24688 21196
rect 24736 21140 24792 21196
rect 24840 21140 24896 21196
rect 24944 21140 25000 21196
rect 25048 21140 25104 21196
rect 25152 21140 25208 21196
rect 5292 20972 5348 21028
rect 13692 20972 13748 21028
rect 26236 20860 26292 20916
rect 25340 20636 25396 20692
rect 13804 20524 13860 20580
rect 14008 20356 14064 20412
rect 14112 20356 14168 20412
rect 14216 20356 14272 20412
rect 14320 20356 14376 20412
rect 14424 20356 14480 20412
rect 14528 20356 14584 20412
rect 14632 20356 14688 20412
rect 14736 20356 14792 20412
rect 14840 20356 14896 20412
rect 14944 20356 15000 20412
rect 15048 20356 15104 20412
rect 15152 20356 15208 20412
rect 34008 20356 34064 20412
rect 34112 20356 34168 20412
rect 34216 20356 34272 20412
rect 34320 20356 34376 20412
rect 34424 20356 34480 20412
rect 34528 20356 34584 20412
rect 34632 20356 34688 20412
rect 34736 20356 34792 20412
rect 34840 20356 34896 20412
rect 34944 20356 35000 20412
rect 35048 20356 35104 20412
rect 35152 20356 35208 20412
rect 6188 20188 6244 20244
rect 25340 20188 25396 20244
rect 13468 19964 13524 20020
rect 4008 19572 4064 19628
rect 4112 19572 4168 19628
rect 4216 19572 4272 19628
rect 4320 19572 4376 19628
rect 4424 19572 4480 19628
rect 4528 19572 4584 19628
rect 4632 19572 4688 19628
rect 4736 19572 4792 19628
rect 4840 19572 4896 19628
rect 4944 19572 5000 19628
rect 5048 19572 5104 19628
rect 5152 19572 5208 19628
rect 24008 19572 24064 19628
rect 24112 19572 24168 19628
rect 24216 19572 24272 19628
rect 24320 19572 24376 19628
rect 24424 19572 24480 19628
rect 24528 19572 24584 19628
rect 24632 19572 24688 19628
rect 24736 19572 24792 19628
rect 24840 19572 24896 19628
rect 24944 19572 25000 19628
rect 25048 19572 25104 19628
rect 25152 19572 25208 19628
rect 25340 19180 25396 19236
rect 13356 19068 13412 19124
rect 14008 18788 14064 18844
rect 14112 18788 14168 18844
rect 14216 18788 14272 18844
rect 14320 18788 14376 18844
rect 14424 18788 14480 18844
rect 14528 18788 14584 18844
rect 14632 18788 14688 18844
rect 14736 18788 14792 18844
rect 14840 18788 14896 18844
rect 14944 18788 15000 18844
rect 15048 18788 15104 18844
rect 15152 18788 15208 18844
rect 34008 18788 34064 18844
rect 34112 18788 34168 18844
rect 34216 18788 34272 18844
rect 34320 18788 34376 18844
rect 34424 18788 34480 18844
rect 34528 18788 34584 18844
rect 34632 18788 34688 18844
rect 34736 18788 34792 18844
rect 34840 18788 34896 18844
rect 34944 18788 35000 18844
rect 35048 18788 35104 18844
rect 35152 18788 35208 18844
rect 4008 18004 4064 18060
rect 4112 18004 4168 18060
rect 4216 18004 4272 18060
rect 4320 18004 4376 18060
rect 4424 18004 4480 18060
rect 4528 18004 4584 18060
rect 4632 18004 4688 18060
rect 4736 18004 4792 18060
rect 4840 18004 4896 18060
rect 4944 18004 5000 18060
rect 5048 18004 5104 18060
rect 5152 18004 5208 18060
rect 24008 18004 24064 18060
rect 24112 18004 24168 18060
rect 24216 18004 24272 18060
rect 24320 18004 24376 18060
rect 24424 18004 24480 18060
rect 24528 18004 24584 18060
rect 24632 18004 24688 18060
rect 24736 18004 24792 18060
rect 24840 18004 24896 18060
rect 24944 18004 25000 18060
rect 25048 18004 25104 18060
rect 25152 18004 25208 18060
rect 13804 17500 13860 17556
rect 26236 17500 26292 17556
rect 25340 17276 25396 17332
rect 14008 17220 14064 17276
rect 14112 17220 14168 17276
rect 14216 17220 14272 17276
rect 14320 17220 14376 17276
rect 14424 17220 14480 17276
rect 14528 17220 14584 17276
rect 14632 17220 14688 17276
rect 14736 17220 14792 17276
rect 14840 17220 14896 17276
rect 14944 17220 15000 17276
rect 15048 17220 15104 17276
rect 15152 17220 15208 17276
rect 34008 17220 34064 17276
rect 34112 17220 34168 17276
rect 34216 17220 34272 17276
rect 34320 17220 34376 17276
rect 34424 17220 34480 17276
rect 34528 17220 34584 17276
rect 34632 17220 34688 17276
rect 34736 17220 34792 17276
rect 34840 17220 34896 17276
rect 34944 17220 35000 17276
rect 35048 17220 35104 17276
rect 35152 17220 35208 17276
rect 3052 17052 3108 17108
rect 15372 17052 15428 17108
rect 3388 16940 3444 16996
rect 23772 16604 23828 16660
rect 4008 16436 4064 16492
rect 4112 16436 4168 16492
rect 4216 16436 4272 16492
rect 4320 16436 4376 16492
rect 4424 16436 4480 16492
rect 4528 16436 4584 16492
rect 4632 16436 4688 16492
rect 4736 16436 4792 16492
rect 4840 16436 4896 16492
rect 4944 16436 5000 16492
rect 5048 16436 5104 16492
rect 5152 16436 5208 16492
rect 13356 16380 13412 16436
rect 24008 16436 24064 16492
rect 24112 16436 24168 16492
rect 24216 16436 24272 16492
rect 24320 16436 24376 16492
rect 24424 16436 24480 16492
rect 24528 16436 24584 16492
rect 24632 16436 24688 16492
rect 24736 16436 24792 16492
rect 24840 16436 24896 16492
rect 24944 16436 25000 16492
rect 25048 16436 25104 16492
rect 25152 16436 25208 16492
rect 13468 16268 13524 16324
rect 5404 16156 5460 16212
rect 23772 16156 23828 16212
rect 25340 15820 25396 15876
rect 6188 15596 6244 15652
rect 14008 15652 14064 15708
rect 14112 15652 14168 15708
rect 14216 15652 14272 15708
rect 14320 15652 14376 15708
rect 14424 15652 14480 15708
rect 14528 15652 14584 15708
rect 14632 15652 14688 15708
rect 14736 15652 14792 15708
rect 14840 15652 14896 15708
rect 14944 15652 15000 15708
rect 15048 15652 15104 15708
rect 15152 15652 15208 15708
rect 34008 15652 34064 15708
rect 34112 15652 34168 15708
rect 34216 15652 34272 15708
rect 34320 15652 34376 15708
rect 34424 15652 34480 15708
rect 34528 15652 34584 15708
rect 34632 15652 34688 15708
rect 34736 15652 34792 15708
rect 34840 15652 34896 15708
rect 34944 15652 35000 15708
rect 35048 15652 35104 15708
rect 35152 15652 35208 15708
rect 13468 15148 13524 15204
rect 4008 14868 4064 14924
rect 4112 14868 4168 14924
rect 4216 14868 4272 14924
rect 4320 14868 4376 14924
rect 4424 14868 4480 14924
rect 4528 14868 4584 14924
rect 4632 14868 4688 14924
rect 4736 14868 4792 14924
rect 4840 14868 4896 14924
rect 4944 14868 5000 14924
rect 5048 14868 5104 14924
rect 5152 14868 5208 14924
rect 24008 14868 24064 14924
rect 24112 14868 24168 14924
rect 24216 14868 24272 14924
rect 24320 14868 24376 14924
rect 24424 14868 24480 14924
rect 24528 14868 24584 14924
rect 24632 14868 24688 14924
rect 24736 14868 24792 14924
rect 24840 14868 24896 14924
rect 24944 14868 25000 14924
rect 25048 14868 25104 14924
rect 25152 14868 25208 14924
rect 6188 14252 6244 14308
rect 14008 14084 14064 14140
rect 14112 14084 14168 14140
rect 14216 14084 14272 14140
rect 14320 14084 14376 14140
rect 14424 14084 14480 14140
rect 14528 14084 14584 14140
rect 14632 14084 14688 14140
rect 14736 14084 14792 14140
rect 14840 14084 14896 14140
rect 14944 14084 15000 14140
rect 15048 14084 15104 14140
rect 15152 14084 15208 14140
rect 34008 14084 34064 14140
rect 34112 14084 34168 14140
rect 34216 14084 34272 14140
rect 34320 14084 34376 14140
rect 34424 14084 34480 14140
rect 34528 14084 34584 14140
rect 34632 14084 34688 14140
rect 34736 14084 34792 14140
rect 34840 14084 34896 14140
rect 34944 14084 35000 14140
rect 35048 14084 35104 14140
rect 35152 14084 35208 14140
rect 3836 13916 3892 13972
rect 13468 13916 13524 13972
rect 4008 13300 4064 13356
rect 4112 13300 4168 13356
rect 4216 13300 4272 13356
rect 4320 13300 4376 13356
rect 4424 13300 4480 13356
rect 4528 13300 4584 13356
rect 4632 13300 4688 13356
rect 4736 13300 4792 13356
rect 4840 13300 4896 13356
rect 4944 13300 5000 13356
rect 5048 13300 5104 13356
rect 5152 13300 5208 13356
rect 24008 13300 24064 13356
rect 24112 13300 24168 13356
rect 24216 13300 24272 13356
rect 24320 13300 24376 13356
rect 24424 13300 24480 13356
rect 24528 13300 24584 13356
rect 24632 13300 24688 13356
rect 24736 13300 24792 13356
rect 24840 13300 24896 13356
rect 24944 13300 25000 13356
rect 25048 13300 25104 13356
rect 25152 13300 25208 13356
rect 5404 13020 5460 13076
rect 13692 12796 13748 12852
rect 14008 12516 14064 12572
rect 14112 12516 14168 12572
rect 14216 12516 14272 12572
rect 14320 12516 14376 12572
rect 14424 12516 14480 12572
rect 14528 12516 14584 12572
rect 14632 12516 14688 12572
rect 14736 12516 14792 12572
rect 14840 12516 14896 12572
rect 14944 12516 15000 12572
rect 15048 12516 15104 12572
rect 15152 12516 15208 12572
rect 34008 12516 34064 12572
rect 34112 12516 34168 12572
rect 34216 12516 34272 12572
rect 34320 12516 34376 12572
rect 34424 12516 34480 12572
rect 34528 12516 34584 12572
rect 34632 12516 34688 12572
rect 34736 12516 34792 12572
rect 34840 12516 34896 12572
rect 34944 12516 35000 12572
rect 35048 12516 35104 12572
rect 35152 12516 35208 12572
rect 4008 11732 4064 11788
rect 4112 11732 4168 11788
rect 4216 11732 4272 11788
rect 4320 11732 4376 11788
rect 4424 11732 4480 11788
rect 4528 11732 4584 11788
rect 4632 11732 4688 11788
rect 4736 11732 4792 11788
rect 4840 11732 4896 11788
rect 4944 11732 5000 11788
rect 5048 11732 5104 11788
rect 5152 11732 5208 11788
rect 24008 11732 24064 11788
rect 24112 11732 24168 11788
rect 24216 11732 24272 11788
rect 24320 11732 24376 11788
rect 24424 11732 24480 11788
rect 24528 11732 24584 11788
rect 24632 11732 24688 11788
rect 24736 11732 24792 11788
rect 24840 11732 24896 11788
rect 24944 11732 25000 11788
rect 25048 11732 25104 11788
rect 25152 11732 25208 11788
rect 5404 11452 5460 11508
rect 14008 10948 14064 11004
rect 14112 10948 14168 11004
rect 14216 10948 14272 11004
rect 14320 10948 14376 11004
rect 14424 10948 14480 11004
rect 14528 10948 14584 11004
rect 14632 10948 14688 11004
rect 14736 10948 14792 11004
rect 14840 10948 14896 11004
rect 14944 10948 15000 11004
rect 15048 10948 15104 11004
rect 15152 10948 15208 11004
rect 34008 10948 34064 11004
rect 34112 10948 34168 11004
rect 34216 10948 34272 11004
rect 34320 10948 34376 11004
rect 34424 10948 34480 11004
rect 34528 10948 34584 11004
rect 34632 10948 34688 11004
rect 34736 10948 34792 11004
rect 34840 10948 34896 11004
rect 34944 10948 35000 11004
rect 35048 10948 35104 11004
rect 35152 10948 35208 11004
rect 4008 10164 4064 10220
rect 4112 10164 4168 10220
rect 4216 10164 4272 10220
rect 4320 10164 4376 10220
rect 4424 10164 4480 10220
rect 4528 10164 4584 10220
rect 4632 10164 4688 10220
rect 4736 10164 4792 10220
rect 4840 10164 4896 10220
rect 4944 10164 5000 10220
rect 5048 10164 5104 10220
rect 5152 10164 5208 10220
rect 24008 10164 24064 10220
rect 24112 10164 24168 10220
rect 24216 10164 24272 10220
rect 24320 10164 24376 10220
rect 24424 10164 24480 10220
rect 24528 10164 24584 10220
rect 24632 10164 24688 10220
rect 24736 10164 24792 10220
rect 24840 10164 24896 10220
rect 24944 10164 25000 10220
rect 25048 10164 25104 10220
rect 25152 10164 25208 10220
rect 14008 9380 14064 9436
rect 14112 9380 14168 9436
rect 14216 9380 14272 9436
rect 14320 9380 14376 9436
rect 14424 9380 14480 9436
rect 14528 9380 14584 9436
rect 14632 9380 14688 9436
rect 14736 9380 14792 9436
rect 14840 9380 14896 9436
rect 14944 9380 15000 9436
rect 15048 9380 15104 9436
rect 15152 9380 15208 9436
rect 34008 9380 34064 9436
rect 34112 9380 34168 9436
rect 34216 9380 34272 9436
rect 34320 9380 34376 9436
rect 34424 9380 34480 9436
rect 34528 9380 34584 9436
rect 34632 9380 34688 9436
rect 34736 9380 34792 9436
rect 34840 9380 34896 9436
rect 34944 9380 35000 9436
rect 35048 9380 35104 9436
rect 35152 9380 35208 9436
rect 4008 8596 4064 8652
rect 4112 8596 4168 8652
rect 4216 8596 4272 8652
rect 4320 8596 4376 8652
rect 4424 8596 4480 8652
rect 4528 8596 4584 8652
rect 4632 8596 4688 8652
rect 4736 8596 4792 8652
rect 4840 8596 4896 8652
rect 4944 8596 5000 8652
rect 5048 8596 5104 8652
rect 5152 8596 5208 8652
rect 24008 8596 24064 8652
rect 24112 8596 24168 8652
rect 24216 8596 24272 8652
rect 24320 8596 24376 8652
rect 24424 8596 24480 8652
rect 24528 8596 24584 8652
rect 24632 8596 24688 8652
rect 24736 8596 24792 8652
rect 24840 8596 24896 8652
rect 24944 8596 25000 8652
rect 25048 8596 25104 8652
rect 25152 8596 25208 8652
rect 14008 7812 14064 7868
rect 14112 7812 14168 7868
rect 14216 7812 14272 7868
rect 14320 7812 14376 7868
rect 14424 7812 14480 7868
rect 14528 7812 14584 7868
rect 14632 7812 14688 7868
rect 14736 7812 14792 7868
rect 14840 7812 14896 7868
rect 14944 7812 15000 7868
rect 15048 7812 15104 7868
rect 15152 7812 15208 7868
rect 34008 7812 34064 7868
rect 34112 7812 34168 7868
rect 34216 7812 34272 7868
rect 34320 7812 34376 7868
rect 34424 7812 34480 7868
rect 34528 7812 34584 7868
rect 34632 7812 34688 7868
rect 34736 7812 34792 7868
rect 34840 7812 34896 7868
rect 34944 7812 35000 7868
rect 35048 7812 35104 7868
rect 35152 7812 35208 7868
rect 4008 7028 4064 7084
rect 4112 7028 4168 7084
rect 4216 7028 4272 7084
rect 4320 7028 4376 7084
rect 4424 7028 4480 7084
rect 4528 7028 4584 7084
rect 4632 7028 4688 7084
rect 4736 7028 4792 7084
rect 4840 7028 4896 7084
rect 4944 7028 5000 7084
rect 5048 7028 5104 7084
rect 5152 7028 5208 7084
rect 24008 7028 24064 7084
rect 24112 7028 24168 7084
rect 24216 7028 24272 7084
rect 24320 7028 24376 7084
rect 24424 7028 24480 7084
rect 24528 7028 24584 7084
rect 24632 7028 24688 7084
rect 24736 7028 24792 7084
rect 24840 7028 24896 7084
rect 24944 7028 25000 7084
rect 25048 7028 25104 7084
rect 25152 7028 25208 7084
rect 14008 6244 14064 6300
rect 14112 6244 14168 6300
rect 14216 6244 14272 6300
rect 14320 6244 14376 6300
rect 14424 6244 14480 6300
rect 14528 6244 14584 6300
rect 14632 6244 14688 6300
rect 14736 6244 14792 6300
rect 14840 6244 14896 6300
rect 14944 6244 15000 6300
rect 15048 6244 15104 6300
rect 15152 6244 15208 6300
rect 34008 6244 34064 6300
rect 34112 6244 34168 6300
rect 34216 6244 34272 6300
rect 34320 6244 34376 6300
rect 34424 6244 34480 6300
rect 34528 6244 34584 6300
rect 34632 6244 34688 6300
rect 34736 6244 34792 6300
rect 34840 6244 34896 6300
rect 34944 6244 35000 6300
rect 35048 6244 35104 6300
rect 35152 6244 35208 6300
rect 4008 5460 4064 5516
rect 4112 5460 4168 5516
rect 4216 5460 4272 5516
rect 4320 5460 4376 5516
rect 4424 5460 4480 5516
rect 4528 5460 4584 5516
rect 4632 5460 4688 5516
rect 4736 5460 4792 5516
rect 4840 5460 4896 5516
rect 4944 5460 5000 5516
rect 5048 5460 5104 5516
rect 5152 5460 5208 5516
rect 24008 5460 24064 5516
rect 24112 5460 24168 5516
rect 24216 5460 24272 5516
rect 24320 5460 24376 5516
rect 24424 5460 24480 5516
rect 24528 5460 24584 5516
rect 24632 5460 24688 5516
rect 24736 5460 24792 5516
rect 24840 5460 24896 5516
rect 24944 5460 25000 5516
rect 25048 5460 25104 5516
rect 25152 5460 25208 5516
rect 14008 4676 14064 4732
rect 14112 4676 14168 4732
rect 14216 4676 14272 4732
rect 14320 4676 14376 4732
rect 14424 4676 14480 4732
rect 14528 4676 14584 4732
rect 14632 4676 14688 4732
rect 14736 4676 14792 4732
rect 14840 4676 14896 4732
rect 14944 4676 15000 4732
rect 15048 4676 15104 4732
rect 15152 4676 15208 4732
rect 34008 4676 34064 4732
rect 34112 4676 34168 4732
rect 34216 4676 34272 4732
rect 34320 4676 34376 4732
rect 34424 4676 34480 4732
rect 34528 4676 34584 4732
rect 34632 4676 34688 4732
rect 34736 4676 34792 4732
rect 34840 4676 34896 4732
rect 34944 4676 35000 4732
rect 35048 4676 35104 4732
rect 35152 4676 35208 4732
rect 4008 3892 4064 3948
rect 4112 3892 4168 3948
rect 4216 3892 4272 3948
rect 4320 3892 4376 3948
rect 4424 3892 4480 3948
rect 4528 3892 4584 3948
rect 4632 3892 4688 3948
rect 4736 3892 4792 3948
rect 4840 3892 4896 3948
rect 4944 3892 5000 3948
rect 5048 3892 5104 3948
rect 5152 3892 5208 3948
rect 24008 3892 24064 3948
rect 24112 3892 24168 3948
rect 24216 3892 24272 3948
rect 24320 3892 24376 3948
rect 24424 3892 24480 3948
rect 24528 3892 24584 3948
rect 24632 3892 24688 3948
rect 24736 3892 24792 3948
rect 24840 3892 24896 3948
rect 24944 3892 25000 3948
rect 25048 3892 25104 3948
rect 25152 3892 25208 3948
rect 14008 3108 14064 3164
rect 14112 3108 14168 3164
rect 14216 3108 14272 3164
rect 14320 3108 14376 3164
rect 14424 3108 14480 3164
rect 14528 3108 14584 3164
rect 14632 3108 14688 3164
rect 14736 3108 14792 3164
rect 14840 3108 14896 3164
rect 14944 3108 15000 3164
rect 15048 3108 15104 3164
rect 15152 3108 15208 3164
rect 34008 3108 34064 3164
rect 34112 3108 34168 3164
rect 34216 3108 34272 3164
rect 34320 3108 34376 3164
rect 34424 3108 34480 3164
rect 34528 3108 34584 3164
rect 34632 3108 34688 3164
rect 34736 3108 34792 3164
rect 34840 3108 34896 3164
rect 34944 3108 35000 3164
rect 35048 3108 35104 3164
rect 35152 3108 35208 3164
<< metal4 >>
rect 3988 96460 5228 96492
rect 3988 96404 4008 96460
rect 4064 96404 4112 96460
rect 4168 96404 4216 96460
rect 4272 96404 4320 96460
rect 4376 96404 4424 96460
rect 4480 96404 4528 96460
rect 4584 96404 4632 96460
rect 4688 96404 4736 96460
rect 4792 96404 4840 96460
rect 4896 96404 4944 96460
rect 5000 96404 5048 96460
rect 5104 96404 5152 96460
rect 5208 96404 5228 96460
rect 3988 94892 5228 96404
rect 3988 94836 4008 94892
rect 4064 94836 4112 94892
rect 4168 94836 4216 94892
rect 4272 94836 4320 94892
rect 4376 94836 4424 94892
rect 4480 94836 4528 94892
rect 4584 94836 4632 94892
rect 4688 94836 4736 94892
rect 4792 94836 4840 94892
rect 4896 94836 4944 94892
rect 5000 94836 5048 94892
rect 5104 94836 5152 94892
rect 5208 94836 5228 94892
rect 3988 93324 5228 94836
rect 3988 93268 4008 93324
rect 4064 93268 4112 93324
rect 4168 93268 4216 93324
rect 4272 93268 4320 93324
rect 4376 93268 4424 93324
rect 4480 93268 4528 93324
rect 4584 93268 4632 93324
rect 4688 93268 4736 93324
rect 4792 93268 4840 93324
rect 4896 93268 4944 93324
rect 5000 93268 5048 93324
rect 5104 93268 5152 93324
rect 5208 93268 5228 93324
rect 3988 91756 5228 93268
rect 3988 91700 4008 91756
rect 4064 91700 4112 91756
rect 4168 91700 4216 91756
rect 4272 91700 4320 91756
rect 4376 91700 4424 91756
rect 4480 91700 4528 91756
rect 4584 91700 4632 91756
rect 4688 91700 4736 91756
rect 4792 91700 4840 91756
rect 4896 91700 4944 91756
rect 5000 91700 5048 91756
rect 5104 91700 5152 91756
rect 5208 91700 5228 91756
rect 3988 90188 5228 91700
rect 3988 90132 4008 90188
rect 4064 90132 4112 90188
rect 4168 90132 4216 90188
rect 4272 90132 4320 90188
rect 4376 90132 4424 90188
rect 4480 90132 4528 90188
rect 4584 90132 4632 90188
rect 4688 90132 4736 90188
rect 4792 90132 4840 90188
rect 4896 90132 4944 90188
rect 5000 90132 5048 90188
rect 5104 90132 5152 90188
rect 5208 90132 5228 90188
rect 3988 88620 5228 90132
rect 3988 88564 4008 88620
rect 4064 88564 4112 88620
rect 4168 88564 4216 88620
rect 4272 88564 4320 88620
rect 4376 88564 4424 88620
rect 4480 88564 4528 88620
rect 4584 88564 4632 88620
rect 4688 88564 4736 88620
rect 4792 88564 4840 88620
rect 4896 88564 4944 88620
rect 5000 88564 5048 88620
rect 5104 88564 5152 88620
rect 5208 88564 5228 88620
rect 3988 87052 5228 88564
rect 3988 86996 4008 87052
rect 4064 86996 4112 87052
rect 4168 86996 4216 87052
rect 4272 86996 4320 87052
rect 4376 86996 4424 87052
rect 4480 86996 4528 87052
rect 4584 86996 4632 87052
rect 4688 86996 4736 87052
rect 4792 86996 4840 87052
rect 4896 86996 4944 87052
rect 5000 86996 5048 87052
rect 5104 86996 5152 87052
rect 5208 86996 5228 87052
rect 3988 85484 5228 86996
rect 13988 95676 15228 96492
rect 13988 95620 14008 95676
rect 14064 95620 14112 95676
rect 14168 95620 14216 95676
rect 14272 95620 14320 95676
rect 14376 95620 14424 95676
rect 14480 95620 14528 95676
rect 14584 95620 14632 95676
rect 14688 95620 14736 95676
rect 14792 95620 14840 95676
rect 14896 95620 14944 95676
rect 15000 95620 15048 95676
rect 15104 95620 15152 95676
rect 15208 95620 15228 95676
rect 13988 94108 15228 95620
rect 13988 94052 14008 94108
rect 14064 94052 14112 94108
rect 14168 94052 14216 94108
rect 14272 94052 14320 94108
rect 14376 94052 14424 94108
rect 14480 94052 14528 94108
rect 14584 94052 14632 94108
rect 14688 94052 14736 94108
rect 14792 94052 14840 94108
rect 14896 94052 14944 94108
rect 15000 94052 15048 94108
rect 15104 94052 15152 94108
rect 15208 94052 15228 94108
rect 13988 92540 15228 94052
rect 13988 92484 14008 92540
rect 14064 92484 14112 92540
rect 14168 92484 14216 92540
rect 14272 92484 14320 92540
rect 14376 92484 14424 92540
rect 14480 92484 14528 92540
rect 14584 92484 14632 92540
rect 14688 92484 14736 92540
rect 14792 92484 14840 92540
rect 14896 92484 14944 92540
rect 15000 92484 15048 92540
rect 15104 92484 15152 92540
rect 15208 92484 15228 92540
rect 13988 90972 15228 92484
rect 13988 90916 14008 90972
rect 14064 90916 14112 90972
rect 14168 90916 14216 90972
rect 14272 90916 14320 90972
rect 14376 90916 14424 90972
rect 14480 90916 14528 90972
rect 14584 90916 14632 90972
rect 14688 90916 14736 90972
rect 14792 90916 14840 90972
rect 14896 90916 14944 90972
rect 15000 90916 15048 90972
rect 15104 90916 15152 90972
rect 15208 90916 15228 90972
rect 13988 89404 15228 90916
rect 13988 89348 14008 89404
rect 14064 89348 14112 89404
rect 14168 89348 14216 89404
rect 14272 89348 14320 89404
rect 14376 89348 14424 89404
rect 14480 89348 14528 89404
rect 14584 89348 14632 89404
rect 14688 89348 14736 89404
rect 14792 89348 14840 89404
rect 14896 89348 14944 89404
rect 15000 89348 15048 89404
rect 15104 89348 15152 89404
rect 15208 89348 15228 89404
rect 13988 87836 15228 89348
rect 13988 87780 14008 87836
rect 14064 87780 14112 87836
rect 14168 87780 14216 87836
rect 14272 87780 14320 87836
rect 14376 87780 14424 87836
rect 14480 87780 14528 87836
rect 14584 87780 14632 87836
rect 14688 87780 14736 87836
rect 14792 87780 14840 87836
rect 14896 87780 14944 87836
rect 15000 87780 15048 87836
rect 15104 87780 15152 87836
rect 15208 87780 15228 87836
rect 13804 86660 13860 86670
rect 13804 85876 13860 86604
rect 13804 85810 13860 85820
rect 13988 86268 15228 87780
rect 13988 86212 14008 86268
rect 14064 86212 14112 86268
rect 14168 86212 14216 86268
rect 14272 86212 14320 86268
rect 14376 86212 14424 86268
rect 14480 86212 14528 86268
rect 14584 86212 14632 86268
rect 14688 86212 14736 86268
rect 14792 86212 14840 86268
rect 14896 86212 14944 86268
rect 15000 86212 15048 86268
rect 15104 86212 15152 86268
rect 15208 86212 15228 86268
rect 3988 85428 4008 85484
rect 4064 85428 4112 85484
rect 4168 85428 4216 85484
rect 4272 85428 4320 85484
rect 4376 85428 4424 85484
rect 4480 85428 4528 85484
rect 4584 85428 4632 85484
rect 4688 85428 4736 85484
rect 4792 85428 4840 85484
rect 4896 85428 4944 85484
rect 5000 85428 5048 85484
rect 5104 85428 5152 85484
rect 5208 85428 5228 85484
rect 3988 83916 5228 85428
rect 13692 84980 13748 84990
rect 3988 83860 4008 83916
rect 4064 83860 4112 83916
rect 4168 83860 4216 83916
rect 4272 83860 4320 83916
rect 4376 83860 4424 83916
rect 4480 83860 4528 83916
rect 4584 83860 4632 83916
rect 4688 83860 4736 83916
rect 4792 83860 4840 83916
rect 4896 83860 4944 83916
rect 5000 83860 5048 83916
rect 5104 83860 5152 83916
rect 5208 83860 5228 83916
rect 3988 82348 5228 83860
rect 13580 84084 13636 84094
rect 3988 82292 4008 82348
rect 4064 82292 4112 82348
rect 4168 82292 4216 82348
rect 4272 82292 4320 82348
rect 4376 82292 4424 82348
rect 4480 82292 4528 82348
rect 4584 82292 4632 82348
rect 4688 82292 4736 82348
rect 4792 82292 4840 82348
rect 4896 82292 4944 82348
rect 5000 82292 5048 82348
rect 5104 82292 5152 82348
rect 5208 82292 5228 82348
rect 3988 80780 5228 82292
rect 10220 82516 10276 82526
rect 10220 81508 10276 82460
rect 10220 81442 10276 81452
rect 11004 82180 11060 82190
rect 3988 80724 4008 80780
rect 4064 80724 4112 80780
rect 4168 80724 4216 80780
rect 4272 80724 4320 80780
rect 4376 80724 4424 80780
rect 4480 80724 4528 80780
rect 4584 80724 4632 80780
rect 4688 80724 4736 80780
rect 4792 80724 4840 80780
rect 4896 80724 4944 80780
rect 5000 80724 5048 80780
rect 5104 80724 5152 80780
rect 5208 80724 5228 80780
rect 3988 79212 5228 80724
rect 11004 80500 11060 82124
rect 3988 79156 4008 79212
rect 4064 79156 4112 79212
rect 4168 79156 4216 79212
rect 4272 79156 4320 79212
rect 4376 79156 4424 79212
rect 4480 79156 4528 79212
rect 4584 79156 4632 79212
rect 4688 79156 4736 79212
rect 4792 79156 4840 79212
rect 4896 79156 4944 79212
rect 5000 79156 5048 79212
rect 5104 79156 5152 79212
rect 5208 79156 5228 79212
rect 3988 77644 5228 79156
rect 5292 79828 5348 79838
rect 5292 78260 5348 79772
rect 11004 78596 11060 80444
rect 11004 78530 11060 78540
rect 5292 78194 5348 78204
rect 3988 77588 4008 77644
rect 4064 77588 4112 77644
rect 4168 77588 4216 77644
rect 4272 77588 4320 77644
rect 4376 77588 4424 77644
rect 4480 77588 4528 77644
rect 4584 77588 4632 77644
rect 4688 77588 4736 77644
rect 4792 77588 4840 77644
rect 4896 77588 4944 77644
rect 5000 77588 5048 77644
rect 5104 77588 5152 77644
rect 5208 77588 5228 77644
rect 3836 76692 3892 76702
rect 3836 74116 3892 76636
rect 3836 74050 3892 74060
rect 3988 76076 5228 77588
rect 3988 76020 4008 76076
rect 4064 76020 4112 76076
rect 4168 76020 4216 76076
rect 4272 76020 4320 76076
rect 4376 76020 4424 76076
rect 4480 76020 4528 76076
rect 4584 76020 4632 76076
rect 4688 76020 4736 76076
rect 4792 76020 4840 76076
rect 4896 76020 4944 76076
rect 5000 76020 5048 76076
rect 5104 76020 5152 76076
rect 5208 76020 5228 76076
rect 3988 74508 5228 76020
rect 3988 74452 4008 74508
rect 4064 74452 4112 74508
rect 4168 74452 4216 74508
rect 4272 74452 4320 74508
rect 4376 74452 4424 74508
rect 4480 74452 4528 74508
rect 4584 74452 4632 74508
rect 4688 74452 4736 74508
rect 4792 74452 4840 74508
rect 4896 74452 4944 74508
rect 5000 74452 5048 74508
rect 5104 74452 5152 74508
rect 5208 74452 5228 74508
rect 3988 72940 5228 74452
rect 3988 72884 4008 72940
rect 4064 72884 4112 72940
rect 4168 72884 4216 72940
rect 4272 72884 4320 72940
rect 4376 72884 4424 72940
rect 4480 72884 4528 72940
rect 4584 72884 4632 72940
rect 4688 72884 4736 72940
rect 4792 72884 4840 72940
rect 4896 72884 4944 72940
rect 5000 72884 5048 72940
rect 5104 72884 5152 72940
rect 5208 72884 5228 72940
rect 3988 71372 5228 72884
rect 3988 71316 4008 71372
rect 4064 71316 4112 71372
rect 4168 71316 4216 71372
rect 4272 71316 4320 71372
rect 4376 71316 4424 71372
rect 4480 71316 4528 71372
rect 4584 71316 4632 71372
rect 4688 71316 4736 71372
rect 4792 71316 4840 71372
rect 4896 71316 4944 71372
rect 5000 71316 5048 71372
rect 5104 71316 5152 71372
rect 5208 71316 5228 71372
rect 3988 69804 5228 71316
rect 13580 74004 13636 84028
rect 13692 83188 13748 84924
rect 13988 84700 15228 86212
rect 23988 96460 25228 96492
rect 23988 96404 24008 96460
rect 24064 96404 24112 96460
rect 24168 96404 24216 96460
rect 24272 96404 24320 96460
rect 24376 96404 24424 96460
rect 24480 96404 24528 96460
rect 24584 96404 24632 96460
rect 24688 96404 24736 96460
rect 24792 96404 24840 96460
rect 24896 96404 24944 96460
rect 25000 96404 25048 96460
rect 25104 96404 25152 96460
rect 25208 96404 25228 96460
rect 23988 94892 25228 96404
rect 23988 94836 24008 94892
rect 24064 94836 24112 94892
rect 24168 94836 24216 94892
rect 24272 94836 24320 94892
rect 24376 94836 24424 94892
rect 24480 94836 24528 94892
rect 24584 94836 24632 94892
rect 24688 94836 24736 94892
rect 24792 94836 24840 94892
rect 24896 94836 24944 94892
rect 25000 94836 25048 94892
rect 25104 94836 25152 94892
rect 25208 94836 25228 94892
rect 23988 93324 25228 94836
rect 23988 93268 24008 93324
rect 24064 93268 24112 93324
rect 24168 93268 24216 93324
rect 24272 93268 24320 93324
rect 24376 93268 24424 93324
rect 24480 93268 24528 93324
rect 24584 93268 24632 93324
rect 24688 93268 24736 93324
rect 24792 93268 24840 93324
rect 24896 93268 24944 93324
rect 25000 93268 25048 93324
rect 25104 93268 25152 93324
rect 25208 93268 25228 93324
rect 23988 91756 25228 93268
rect 23988 91700 24008 91756
rect 24064 91700 24112 91756
rect 24168 91700 24216 91756
rect 24272 91700 24320 91756
rect 24376 91700 24424 91756
rect 24480 91700 24528 91756
rect 24584 91700 24632 91756
rect 24688 91700 24736 91756
rect 24792 91700 24840 91756
rect 24896 91700 24944 91756
rect 25000 91700 25048 91756
rect 25104 91700 25152 91756
rect 25208 91700 25228 91756
rect 23988 90188 25228 91700
rect 23988 90132 24008 90188
rect 24064 90132 24112 90188
rect 24168 90132 24216 90188
rect 24272 90132 24320 90188
rect 24376 90132 24424 90188
rect 24480 90132 24528 90188
rect 24584 90132 24632 90188
rect 24688 90132 24736 90188
rect 24792 90132 24840 90188
rect 24896 90132 24944 90188
rect 25000 90132 25048 90188
rect 25104 90132 25152 90188
rect 25208 90132 25228 90188
rect 23988 88620 25228 90132
rect 23988 88564 24008 88620
rect 24064 88564 24112 88620
rect 24168 88564 24216 88620
rect 24272 88564 24320 88620
rect 24376 88564 24424 88620
rect 24480 88564 24528 88620
rect 24584 88564 24632 88620
rect 24688 88564 24736 88620
rect 24792 88564 24840 88620
rect 24896 88564 24944 88620
rect 25000 88564 25048 88620
rect 25104 88564 25152 88620
rect 25208 88564 25228 88620
rect 23988 87052 25228 88564
rect 23988 86996 24008 87052
rect 24064 86996 24112 87052
rect 24168 86996 24216 87052
rect 24272 86996 24320 87052
rect 24376 86996 24424 87052
rect 24480 86996 24528 87052
rect 24584 86996 24632 87052
rect 24688 86996 24736 87052
rect 24792 86996 24840 87052
rect 24896 86996 24944 87052
rect 25000 86996 25048 87052
rect 25104 86996 25152 87052
rect 25208 86996 25228 87052
rect 23988 85484 25228 86996
rect 23988 85428 24008 85484
rect 24064 85428 24112 85484
rect 24168 85428 24216 85484
rect 24272 85428 24320 85484
rect 24376 85428 24424 85484
rect 24480 85428 24528 85484
rect 24584 85428 24632 85484
rect 24688 85428 24736 85484
rect 24792 85428 24840 85484
rect 24896 85428 24944 85484
rect 25000 85428 25048 85484
rect 25104 85428 25152 85484
rect 25208 85428 25228 85484
rect 13988 84644 14008 84700
rect 14064 84644 14112 84700
rect 14168 84644 14216 84700
rect 14272 84644 14320 84700
rect 14376 84644 14424 84700
rect 14480 84644 14528 84700
rect 14584 84644 14632 84700
rect 14688 84644 14736 84700
rect 14792 84644 14840 84700
rect 14896 84644 14944 84700
rect 15000 84644 15048 84700
rect 15104 84644 15152 84700
rect 15208 84644 15228 84700
rect 13692 83122 13748 83132
rect 13804 83300 13860 83310
rect 13804 82740 13860 83244
rect 13804 82674 13860 82684
rect 13988 83132 15228 84644
rect 13988 83076 14008 83132
rect 14064 83076 14112 83132
rect 14168 83076 14216 83132
rect 14272 83076 14320 83132
rect 14376 83076 14424 83132
rect 14480 83076 14528 83132
rect 14584 83076 14632 83132
rect 14688 83076 14736 83132
rect 14792 83076 14840 83132
rect 14896 83076 14944 83132
rect 15000 83076 15048 83132
rect 15104 83076 15152 83132
rect 15208 83076 15228 83132
rect 13804 81956 13860 81966
rect 13804 81060 13860 81900
rect 13804 80994 13860 81004
rect 13988 81564 15228 83076
rect 13988 81508 14008 81564
rect 14064 81508 14112 81564
rect 14168 81508 14216 81564
rect 14272 81508 14320 81564
rect 14376 81508 14424 81564
rect 14480 81508 14528 81564
rect 14584 81508 14632 81564
rect 14688 81508 14736 81564
rect 14792 81508 14840 81564
rect 14896 81508 14944 81564
rect 15000 81508 15048 81564
rect 15104 81508 15152 81564
rect 15208 81508 15228 81564
rect 13988 79996 15228 81508
rect 13988 79940 14008 79996
rect 14064 79940 14112 79996
rect 14168 79940 14216 79996
rect 14272 79940 14320 79996
rect 14376 79940 14424 79996
rect 14480 79940 14528 79996
rect 14584 79940 14632 79996
rect 14688 79940 14736 79996
rect 14792 79940 14840 79996
rect 14896 79940 14944 79996
rect 15000 79940 15048 79996
rect 15104 79940 15152 79996
rect 15208 79940 15228 79996
rect 13692 79044 13748 79054
rect 13692 78148 13748 78988
rect 13692 78082 13748 78092
rect 13988 78428 15228 79940
rect 13988 78372 14008 78428
rect 14064 78372 14112 78428
rect 14168 78372 14216 78428
rect 14272 78372 14320 78428
rect 14376 78372 14424 78428
rect 14480 78372 14528 78428
rect 14584 78372 14632 78428
rect 14688 78372 14736 78428
rect 14792 78372 14840 78428
rect 14896 78372 14944 78428
rect 15000 78372 15048 78428
rect 15104 78372 15152 78428
rect 15208 78372 15228 78428
rect 13804 77364 13860 77374
rect 3988 69748 4008 69804
rect 4064 69748 4112 69804
rect 4168 69748 4216 69804
rect 4272 69748 4320 69804
rect 4376 69748 4424 69804
rect 4480 69748 4528 69804
rect 4584 69748 4632 69804
rect 4688 69748 4736 69804
rect 4792 69748 4840 69804
rect 4896 69748 4944 69804
rect 5000 69748 5048 69804
rect 5104 69748 5152 69804
rect 5208 69748 5228 69804
rect 3988 68236 5228 69748
rect 3988 68180 4008 68236
rect 4064 68180 4112 68236
rect 4168 68180 4216 68236
rect 4272 68180 4320 68236
rect 4376 68180 4424 68236
rect 4480 68180 4528 68236
rect 4584 68180 4632 68236
rect 4688 68180 4736 68236
rect 4792 68180 4840 68236
rect 4896 68180 4944 68236
rect 5000 68180 5048 68236
rect 5104 68180 5152 68236
rect 5208 68180 5228 68236
rect 3988 66668 5228 68180
rect 13468 70644 13524 70654
rect 3988 66612 4008 66668
rect 4064 66612 4112 66668
rect 4168 66612 4216 66668
rect 4272 66612 4320 66668
rect 4376 66612 4424 66668
rect 4480 66612 4528 66668
rect 4584 66612 4632 66668
rect 4688 66612 4736 66668
rect 4792 66612 4840 66668
rect 4896 66612 4944 66668
rect 5000 66612 5048 66668
rect 5104 66612 5152 66668
rect 5208 66612 5228 66668
rect 3988 65100 5228 66612
rect 6524 67396 6580 67406
rect 3988 65044 4008 65100
rect 4064 65044 4112 65100
rect 4168 65044 4216 65100
rect 4272 65044 4320 65100
rect 4376 65044 4424 65100
rect 4480 65044 4528 65100
rect 4584 65044 4632 65100
rect 4688 65044 4736 65100
rect 4792 65044 4840 65100
rect 4896 65044 4944 65100
rect 5000 65044 5048 65100
rect 5104 65044 5152 65100
rect 5208 65044 5228 65100
rect 3988 63532 5228 65044
rect 3988 63476 4008 63532
rect 4064 63476 4112 63532
rect 4168 63476 4216 63532
rect 4272 63476 4320 63532
rect 4376 63476 4424 63532
rect 4480 63476 4528 63532
rect 4584 63476 4632 63532
rect 4688 63476 4736 63532
rect 4792 63476 4840 63532
rect 4896 63476 4944 63532
rect 5000 63476 5048 63532
rect 5104 63476 5152 63532
rect 5208 63476 5228 63532
rect 3988 61964 5228 63476
rect 3988 61908 4008 61964
rect 4064 61908 4112 61964
rect 4168 61908 4216 61964
rect 4272 61908 4320 61964
rect 4376 61908 4424 61964
rect 4480 61908 4528 61964
rect 4584 61908 4632 61964
rect 4688 61908 4736 61964
rect 4792 61908 4840 61964
rect 4896 61908 4944 61964
rect 5000 61908 5048 61964
rect 5104 61908 5152 61964
rect 5208 61908 5228 61964
rect 3988 60396 5228 61908
rect 5292 65604 5348 65614
rect 5292 62356 5348 65548
rect 5292 61460 5348 62300
rect 5292 61394 5348 61404
rect 5404 64036 5460 64046
rect 5404 61348 5460 63980
rect 5404 61282 5460 61292
rect 3988 60340 4008 60396
rect 4064 60340 4112 60396
rect 4168 60340 4216 60396
rect 4272 60340 4320 60396
rect 4376 60340 4424 60396
rect 4480 60340 4528 60396
rect 4584 60340 4632 60396
rect 4688 60340 4736 60396
rect 4792 60340 4840 60396
rect 4896 60340 4944 60396
rect 5000 60340 5048 60396
rect 5104 60340 5152 60396
rect 5208 60340 5228 60396
rect 3988 58828 5228 60340
rect 6524 59780 6580 67340
rect 6524 59714 6580 59724
rect 3988 58772 4008 58828
rect 4064 58772 4112 58828
rect 4168 58772 4216 58828
rect 4272 58772 4320 58828
rect 4376 58772 4424 58828
rect 4480 58772 4528 58828
rect 4584 58772 4632 58828
rect 4688 58772 4736 58828
rect 4792 58772 4840 58828
rect 4896 58772 4944 58828
rect 5000 58772 5048 58828
rect 5104 58772 5152 58828
rect 5208 58772 5228 58828
rect 3988 57260 5228 58772
rect 13468 58772 13524 70588
rect 13580 68852 13636 73948
rect 13692 75572 13748 75582
rect 13692 73892 13748 75516
rect 13804 75124 13860 77308
rect 13804 75058 13860 75068
rect 13988 76860 15228 78372
rect 13988 76804 14008 76860
rect 14064 76804 14112 76860
rect 14168 76804 14216 76860
rect 14272 76804 14320 76860
rect 14376 76804 14424 76860
rect 14480 76804 14528 76860
rect 14584 76804 14632 76860
rect 14688 76804 14736 76860
rect 14792 76804 14840 76860
rect 14896 76804 14944 76860
rect 15000 76804 15048 76860
rect 15104 76804 15152 76860
rect 15208 76804 15228 76860
rect 13988 75292 15228 76804
rect 13988 75236 14008 75292
rect 14064 75236 14112 75292
rect 14168 75236 14216 75292
rect 14272 75236 14320 75292
rect 14376 75236 14424 75292
rect 14480 75236 14528 75292
rect 14584 75236 14632 75292
rect 14688 75236 14736 75292
rect 14792 75236 14840 75292
rect 14896 75236 14944 75292
rect 15000 75236 15048 75292
rect 15104 75236 15152 75292
rect 15208 75236 15228 75292
rect 13692 73556 13748 73836
rect 13692 73490 13748 73500
rect 13988 73724 15228 75236
rect 15372 85204 15428 85214
rect 15372 75124 15428 85148
rect 19292 84084 19348 84094
rect 15484 81844 15540 81854
rect 15484 80612 15540 81788
rect 15484 78708 15540 80556
rect 15484 78036 15540 78652
rect 15484 77970 15540 77980
rect 15372 75058 15428 75068
rect 19292 76356 19348 84028
rect 13988 73668 14008 73724
rect 14064 73668 14112 73724
rect 14168 73668 14216 73724
rect 14272 73668 14320 73724
rect 14376 73668 14424 73724
rect 14480 73668 14528 73724
rect 14584 73668 14632 73724
rect 14688 73668 14736 73724
rect 14792 73668 14840 73724
rect 14896 73668 14944 73724
rect 15000 73668 15048 73724
rect 15104 73668 15152 73724
rect 15208 73668 15228 73724
rect 13988 72156 15228 73668
rect 13988 72100 14008 72156
rect 14064 72100 14112 72156
rect 14168 72100 14216 72156
rect 14272 72100 14320 72156
rect 14376 72100 14424 72156
rect 14480 72100 14528 72156
rect 14584 72100 14632 72156
rect 14688 72100 14736 72156
rect 14792 72100 14840 72156
rect 14896 72100 14944 72156
rect 15000 72100 15048 72156
rect 15104 72100 15152 72156
rect 15208 72100 15228 72156
rect 13988 70588 15228 72100
rect 13988 70532 14008 70588
rect 14064 70532 14112 70588
rect 14168 70532 14216 70588
rect 14272 70532 14320 70588
rect 14376 70532 14424 70588
rect 14480 70532 14528 70588
rect 14584 70532 14632 70588
rect 14688 70532 14736 70588
rect 14792 70532 14840 70588
rect 14896 70532 14944 70588
rect 15000 70532 15048 70588
rect 15104 70532 15152 70588
rect 15208 70532 15228 70588
rect 13580 68786 13636 68796
rect 13692 69748 13748 69758
rect 13580 65380 13636 65390
rect 13580 62468 13636 65324
rect 13692 64148 13748 69692
rect 13988 69020 15228 70532
rect 13988 68964 14008 69020
rect 14064 68964 14112 69020
rect 14168 68964 14216 69020
rect 14272 68964 14320 69020
rect 14376 68964 14424 69020
rect 14480 68964 14528 69020
rect 14584 68964 14632 69020
rect 14688 68964 14736 69020
rect 14792 68964 14840 69020
rect 14896 68964 14944 69020
rect 15000 68964 15048 69020
rect 15104 68964 15152 69020
rect 15208 68964 15228 69020
rect 13988 67452 15228 68964
rect 15372 69524 15428 69534
rect 15372 67844 15428 69468
rect 15372 67778 15428 67788
rect 13988 67396 14008 67452
rect 14064 67396 14112 67452
rect 14168 67396 14216 67452
rect 14272 67396 14320 67452
rect 14376 67396 14424 67452
rect 14480 67396 14528 67452
rect 14584 67396 14632 67452
rect 14688 67396 14736 67452
rect 14792 67396 14840 67452
rect 14896 67396 14944 67452
rect 15000 67396 15048 67452
rect 15104 67396 15152 67452
rect 15208 67396 15228 67452
rect 13988 65884 15228 67396
rect 13988 65828 14008 65884
rect 14064 65828 14112 65884
rect 14168 65828 14216 65884
rect 14272 65828 14320 65884
rect 14376 65828 14424 65884
rect 14480 65828 14528 65884
rect 14584 65828 14632 65884
rect 14688 65828 14736 65884
rect 14792 65828 14840 65884
rect 14896 65828 14944 65884
rect 15000 65828 15048 65884
rect 15104 65828 15152 65884
rect 15208 65828 15228 65884
rect 13692 63588 13748 64092
rect 13692 63522 13748 63532
rect 13804 65156 13860 65166
rect 13804 63700 13860 65100
rect 13580 62402 13636 62412
rect 13692 63364 13748 63374
rect 13692 61348 13748 63308
rect 13804 62692 13860 63644
rect 13804 62626 13860 62636
rect 13988 64316 15228 65828
rect 19180 66276 19236 66286
rect 15484 65156 15540 65166
rect 13988 64260 14008 64316
rect 14064 64260 14112 64316
rect 14168 64260 14216 64316
rect 14272 64260 14320 64316
rect 14376 64260 14424 64316
rect 14480 64260 14528 64316
rect 14584 64260 14632 64316
rect 14688 64260 14736 64316
rect 14792 64260 14840 64316
rect 14896 64260 14944 64316
rect 15000 64260 15048 64316
rect 15104 64260 15152 64316
rect 15208 64260 15228 64316
rect 13988 62748 15228 64260
rect 15372 64820 15428 64830
rect 15372 64148 15428 64764
rect 15372 64082 15428 64092
rect 15484 63028 15540 65100
rect 19180 64484 19236 66220
rect 19180 64418 19236 64428
rect 15484 62962 15540 62972
rect 13988 62692 14008 62748
rect 14064 62692 14112 62748
rect 14168 62692 14216 62748
rect 14272 62692 14320 62748
rect 14376 62692 14424 62748
rect 14480 62692 14528 62748
rect 14584 62692 14632 62748
rect 14688 62692 14736 62748
rect 14792 62692 14840 62748
rect 14896 62692 14944 62748
rect 15000 62692 15048 62748
rect 15104 62692 15152 62748
rect 15208 62692 15228 62748
rect 13692 61282 13748 61292
rect 13804 61684 13860 61694
rect 13804 58996 13860 61628
rect 13804 58930 13860 58940
rect 13988 61180 15228 62692
rect 19292 61572 19348 76300
rect 23988 83916 25228 85428
rect 23988 83860 24008 83916
rect 24064 83860 24112 83916
rect 24168 83860 24216 83916
rect 24272 83860 24320 83916
rect 24376 83860 24424 83916
rect 24480 83860 24528 83916
rect 24584 83860 24632 83916
rect 24688 83860 24736 83916
rect 24792 83860 24840 83916
rect 24896 83860 24944 83916
rect 25000 83860 25048 83916
rect 25104 83860 25152 83916
rect 25208 83860 25228 83916
rect 23988 82348 25228 83860
rect 23988 82292 24008 82348
rect 24064 82292 24112 82348
rect 24168 82292 24216 82348
rect 24272 82292 24320 82348
rect 24376 82292 24424 82348
rect 24480 82292 24528 82348
rect 24584 82292 24632 82348
rect 24688 82292 24736 82348
rect 24792 82292 24840 82348
rect 24896 82292 24944 82348
rect 25000 82292 25048 82348
rect 25104 82292 25152 82348
rect 25208 82292 25228 82348
rect 23988 80780 25228 82292
rect 23988 80724 24008 80780
rect 24064 80724 24112 80780
rect 24168 80724 24216 80780
rect 24272 80724 24320 80780
rect 24376 80724 24424 80780
rect 24480 80724 24528 80780
rect 24584 80724 24632 80780
rect 24688 80724 24736 80780
rect 24792 80724 24840 80780
rect 24896 80724 24944 80780
rect 25000 80724 25048 80780
rect 25104 80724 25152 80780
rect 25208 80724 25228 80780
rect 23988 79212 25228 80724
rect 23988 79156 24008 79212
rect 24064 79156 24112 79212
rect 24168 79156 24216 79212
rect 24272 79156 24320 79212
rect 24376 79156 24424 79212
rect 24480 79156 24528 79212
rect 24584 79156 24632 79212
rect 24688 79156 24736 79212
rect 24792 79156 24840 79212
rect 24896 79156 24944 79212
rect 25000 79156 25048 79212
rect 25104 79156 25152 79212
rect 25208 79156 25228 79212
rect 23988 77644 25228 79156
rect 23988 77588 24008 77644
rect 24064 77588 24112 77644
rect 24168 77588 24216 77644
rect 24272 77588 24320 77644
rect 24376 77588 24424 77644
rect 24480 77588 24528 77644
rect 24584 77588 24632 77644
rect 24688 77588 24736 77644
rect 24792 77588 24840 77644
rect 24896 77588 24944 77644
rect 25000 77588 25048 77644
rect 25104 77588 25152 77644
rect 25208 77588 25228 77644
rect 23988 76076 25228 77588
rect 23988 76020 24008 76076
rect 24064 76020 24112 76076
rect 24168 76020 24216 76076
rect 24272 76020 24320 76076
rect 24376 76020 24424 76076
rect 24480 76020 24528 76076
rect 24584 76020 24632 76076
rect 24688 76020 24736 76076
rect 24792 76020 24840 76076
rect 24896 76020 24944 76076
rect 25000 76020 25048 76076
rect 25104 76020 25152 76076
rect 25208 76020 25228 76076
rect 23988 74508 25228 76020
rect 23988 74452 24008 74508
rect 24064 74452 24112 74508
rect 24168 74452 24216 74508
rect 24272 74452 24320 74508
rect 24376 74452 24424 74508
rect 24480 74452 24528 74508
rect 24584 74452 24632 74508
rect 24688 74452 24736 74508
rect 24792 74452 24840 74508
rect 24896 74452 24944 74508
rect 25000 74452 25048 74508
rect 25104 74452 25152 74508
rect 25208 74452 25228 74508
rect 23988 72940 25228 74452
rect 23988 72884 24008 72940
rect 24064 72884 24112 72940
rect 24168 72884 24216 72940
rect 24272 72884 24320 72940
rect 24376 72884 24424 72940
rect 24480 72884 24528 72940
rect 24584 72884 24632 72940
rect 24688 72884 24736 72940
rect 24792 72884 24840 72940
rect 24896 72884 24944 72940
rect 25000 72884 25048 72940
rect 25104 72884 25152 72940
rect 25208 72884 25228 72940
rect 23988 71372 25228 72884
rect 23988 71316 24008 71372
rect 24064 71316 24112 71372
rect 24168 71316 24216 71372
rect 24272 71316 24320 71372
rect 24376 71316 24424 71372
rect 24480 71316 24528 71372
rect 24584 71316 24632 71372
rect 24688 71316 24736 71372
rect 24792 71316 24840 71372
rect 24896 71316 24944 71372
rect 25000 71316 25048 71372
rect 25104 71316 25152 71372
rect 25208 71316 25228 71372
rect 23988 69804 25228 71316
rect 23988 69748 24008 69804
rect 24064 69748 24112 69804
rect 24168 69748 24216 69804
rect 24272 69748 24320 69804
rect 24376 69748 24424 69804
rect 24480 69748 24528 69804
rect 24584 69748 24632 69804
rect 24688 69748 24736 69804
rect 24792 69748 24840 69804
rect 24896 69748 24944 69804
rect 25000 69748 25048 69804
rect 25104 69748 25152 69804
rect 25208 69748 25228 69804
rect 19404 69188 19460 69198
rect 19404 62580 19460 69132
rect 23988 68236 25228 69748
rect 23988 68180 24008 68236
rect 24064 68180 24112 68236
rect 24168 68180 24216 68236
rect 24272 68180 24320 68236
rect 24376 68180 24424 68236
rect 24480 68180 24528 68236
rect 24584 68180 24632 68236
rect 24688 68180 24736 68236
rect 24792 68180 24840 68236
rect 24896 68180 24944 68236
rect 25000 68180 25048 68236
rect 25104 68180 25152 68236
rect 25208 68180 25228 68236
rect 23988 66668 25228 68180
rect 33988 95676 35228 96492
rect 33988 95620 34008 95676
rect 34064 95620 34112 95676
rect 34168 95620 34216 95676
rect 34272 95620 34320 95676
rect 34376 95620 34424 95676
rect 34480 95620 34528 95676
rect 34584 95620 34632 95676
rect 34688 95620 34736 95676
rect 34792 95620 34840 95676
rect 34896 95620 34944 95676
rect 35000 95620 35048 95676
rect 35104 95620 35152 95676
rect 35208 95620 35228 95676
rect 33988 94108 35228 95620
rect 33988 94052 34008 94108
rect 34064 94052 34112 94108
rect 34168 94052 34216 94108
rect 34272 94052 34320 94108
rect 34376 94052 34424 94108
rect 34480 94052 34528 94108
rect 34584 94052 34632 94108
rect 34688 94052 34736 94108
rect 34792 94052 34840 94108
rect 34896 94052 34944 94108
rect 35000 94052 35048 94108
rect 35104 94052 35152 94108
rect 35208 94052 35228 94108
rect 33988 92540 35228 94052
rect 33988 92484 34008 92540
rect 34064 92484 34112 92540
rect 34168 92484 34216 92540
rect 34272 92484 34320 92540
rect 34376 92484 34424 92540
rect 34480 92484 34528 92540
rect 34584 92484 34632 92540
rect 34688 92484 34736 92540
rect 34792 92484 34840 92540
rect 34896 92484 34944 92540
rect 35000 92484 35048 92540
rect 35104 92484 35152 92540
rect 35208 92484 35228 92540
rect 33988 90972 35228 92484
rect 33988 90916 34008 90972
rect 34064 90916 34112 90972
rect 34168 90916 34216 90972
rect 34272 90916 34320 90972
rect 34376 90916 34424 90972
rect 34480 90916 34528 90972
rect 34584 90916 34632 90972
rect 34688 90916 34736 90972
rect 34792 90916 34840 90972
rect 34896 90916 34944 90972
rect 35000 90916 35048 90972
rect 35104 90916 35152 90972
rect 35208 90916 35228 90972
rect 33988 89404 35228 90916
rect 33988 89348 34008 89404
rect 34064 89348 34112 89404
rect 34168 89348 34216 89404
rect 34272 89348 34320 89404
rect 34376 89348 34424 89404
rect 34480 89348 34528 89404
rect 34584 89348 34632 89404
rect 34688 89348 34736 89404
rect 34792 89348 34840 89404
rect 34896 89348 34944 89404
rect 35000 89348 35048 89404
rect 35104 89348 35152 89404
rect 35208 89348 35228 89404
rect 33988 87836 35228 89348
rect 33988 87780 34008 87836
rect 34064 87780 34112 87836
rect 34168 87780 34216 87836
rect 34272 87780 34320 87836
rect 34376 87780 34424 87836
rect 34480 87780 34528 87836
rect 34584 87780 34632 87836
rect 34688 87780 34736 87836
rect 34792 87780 34840 87836
rect 34896 87780 34944 87836
rect 35000 87780 35048 87836
rect 35104 87780 35152 87836
rect 35208 87780 35228 87836
rect 33988 86268 35228 87780
rect 33988 86212 34008 86268
rect 34064 86212 34112 86268
rect 34168 86212 34216 86268
rect 34272 86212 34320 86268
rect 34376 86212 34424 86268
rect 34480 86212 34528 86268
rect 34584 86212 34632 86268
rect 34688 86212 34736 86268
rect 34792 86212 34840 86268
rect 34896 86212 34944 86268
rect 35000 86212 35048 86268
rect 35104 86212 35152 86268
rect 35208 86212 35228 86268
rect 33988 84700 35228 86212
rect 33988 84644 34008 84700
rect 34064 84644 34112 84700
rect 34168 84644 34216 84700
rect 34272 84644 34320 84700
rect 34376 84644 34424 84700
rect 34480 84644 34528 84700
rect 34584 84644 34632 84700
rect 34688 84644 34736 84700
rect 34792 84644 34840 84700
rect 34896 84644 34944 84700
rect 35000 84644 35048 84700
rect 35104 84644 35152 84700
rect 35208 84644 35228 84700
rect 33988 83132 35228 84644
rect 33988 83076 34008 83132
rect 34064 83076 34112 83132
rect 34168 83076 34216 83132
rect 34272 83076 34320 83132
rect 34376 83076 34424 83132
rect 34480 83076 34528 83132
rect 34584 83076 34632 83132
rect 34688 83076 34736 83132
rect 34792 83076 34840 83132
rect 34896 83076 34944 83132
rect 35000 83076 35048 83132
rect 35104 83076 35152 83132
rect 35208 83076 35228 83132
rect 33988 81564 35228 83076
rect 33988 81508 34008 81564
rect 34064 81508 34112 81564
rect 34168 81508 34216 81564
rect 34272 81508 34320 81564
rect 34376 81508 34424 81564
rect 34480 81508 34528 81564
rect 34584 81508 34632 81564
rect 34688 81508 34736 81564
rect 34792 81508 34840 81564
rect 34896 81508 34944 81564
rect 35000 81508 35048 81564
rect 35104 81508 35152 81564
rect 35208 81508 35228 81564
rect 33988 79996 35228 81508
rect 33988 79940 34008 79996
rect 34064 79940 34112 79996
rect 34168 79940 34216 79996
rect 34272 79940 34320 79996
rect 34376 79940 34424 79996
rect 34480 79940 34528 79996
rect 34584 79940 34632 79996
rect 34688 79940 34736 79996
rect 34792 79940 34840 79996
rect 34896 79940 34944 79996
rect 35000 79940 35048 79996
rect 35104 79940 35152 79996
rect 35208 79940 35228 79996
rect 33988 78428 35228 79940
rect 33988 78372 34008 78428
rect 34064 78372 34112 78428
rect 34168 78372 34216 78428
rect 34272 78372 34320 78428
rect 34376 78372 34424 78428
rect 34480 78372 34528 78428
rect 34584 78372 34632 78428
rect 34688 78372 34736 78428
rect 34792 78372 34840 78428
rect 34896 78372 34944 78428
rect 35000 78372 35048 78428
rect 35104 78372 35152 78428
rect 35208 78372 35228 78428
rect 33988 76860 35228 78372
rect 33988 76804 34008 76860
rect 34064 76804 34112 76860
rect 34168 76804 34216 76860
rect 34272 76804 34320 76860
rect 34376 76804 34424 76860
rect 34480 76804 34528 76860
rect 34584 76804 34632 76860
rect 34688 76804 34736 76860
rect 34792 76804 34840 76860
rect 34896 76804 34944 76860
rect 35000 76804 35048 76860
rect 35104 76804 35152 76860
rect 35208 76804 35228 76860
rect 33988 75292 35228 76804
rect 33988 75236 34008 75292
rect 34064 75236 34112 75292
rect 34168 75236 34216 75292
rect 34272 75236 34320 75292
rect 34376 75236 34424 75292
rect 34480 75236 34528 75292
rect 34584 75236 34632 75292
rect 34688 75236 34736 75292
rect 34792 75236 34840 75292
rect 34896 75236 34944 75292
rect 35000 75236 35048 75292
rect 35104 75236 35152 75292
rect 35208 75236 35228 75292
rect 33988 73724 35228 75236
rect 33988 73668 34008 73724
rect 34064 73668 34112 73724
rect 34168 73668 34216 73724
rect 34272 73668 34320 73724
rect 34376 73668 34424 73724
rect 34480 73668 34528 73724
rect 34584 73668 34632 73724
rect 34688 73668 34736 73724
rect 34792 73668 34840 73724
rect 34896 73668 34944 73724
rect 35000 73668 35048 73724
rect 35104 73668 35152 73724
rect 35208 73668 35228 73724
rect 33988 72156 35228 73668
rect 33988 72100 34008 72156
rect 34064 72100 34112 72156
rect 34168 72100 34216 72156
rect 34272 72100 34320 72156
rect 34376 72100 34424 72156
rect 34480 72100 34528 72156
rect 34584 72100 34632 72156
rect 34688 72100 34736 72156
rect 34792 72100 34840 72156
rect 34896 72100 34944 72156
rect 35000 72100 35048 72156
rect 35104 72100 35152 72156
rect 35208 72100 35228 72156
rect 33988 70588 35228 72100
rect 33988 70532 34008 70588
rect 34064 70532 34112 70588
rect 34168 70532 34216 70588
rect 34272 70532 34320 70588
rect 34376 70532 34424 70588
rect 34480 70532 34528 70588
rect 34584 70532 34632 70588
rect 34688 70532 34736 70588
rect 34792 70532 34840 70588
rect 34896 70532 34944 70588
rect 35000 70532 35048 70588
rect 35104 70532 35152 70588
rect 35208 70532 35228 70588
rect 33988 69020 35228 70532
rect 35308 71540 35364 71550
rect 35308 70420 35364 71484
rect 35308 70354 35364 70364
rect 33988 68964 34008 69020
rect 34064 68964 34112 69020
rect 34168 68964 34216 69020
rect 34272 68964 34320 69020
rect 34376 68964 34424 69020
rect 34480 68964 34528 69020
rect 34584 68964 34632 69020
rect 34688 68964 34736 69020
rect 34792 68964 34840 69020
rect 34896 68964 34944 69020
rect 35000 68964 35048 69020
rect 35104 68964 35152 69020
rect 35208 68964 35228 69020
rect 33988 67452 35228 68964
rect 33988 67396 34008 67452
rect 34064 67396 34112 67452
rect 34168 67396 34216 67452
rect 34272 67396 34320 67452
rect 34376 67396 34424 67452
rect 34480 67396 34528 67452
rect 34584 67396 34632 67452
rect 34688 67396 34736 67452
rect 34792 67396 34840 67452
rect 34896 67396 34944 67452
rect 35000 67396 35048 67452
rect 35104 67396 35152 67452
rect 35208 67396 35228 67452
rect 23988 66612 24008 66668
rect 24064 66612 24112 66668
rect 24168 66612 24216 66668
rect 24272 66612 24320 66668
rect 24376 66612 24424 66668
rect 24480 66612 24528 66668
rect 24584 66612 24632 66668
rect 24688 66612 24736 66668
rect 24792 66612 24840 66668
rect 24896 66612 24944 66668
rect 25000 66612 25048 66668
rect 25104 66612 25152 66668
rect 25208 66612 25228 66668
rect 23988 65100 25228 66612
rect 23988 65044 24008 65100
rect 24064 65044 24112 65100
rect 24168 65044 24216 65100
rect 24272 65044 24320 65100
rect 24376 65044 24424 65100
rect 24480 65044 24528 65100
rect 24584 65044 24632 65100
rect 24688 65044 24736 65100
rect 24792 65044 24840 65100
rect 24896 65044 24944 65100
rect 25000 65044 25048 65100
rect 25104 65044 25152 65100
rect 25208 65044 25228 65100
rect 19964 64036 20020 64046
rect 19964 62916 20020 63980
rect 19964 62850 20020 62860
rect 23988 63532 25228 65044
rect 23988 63476 24008 63532
rect 24064 63476 24112 63532
rect 24168 63476 24216 63532
rect 24272 63476 24320 63532
rect 24376 63476 24424 63532
rect 24480 63476 24528 63532
rect 24584 63476 24632 63532
rect 24688 63476 24736 63532
rect 24792 63476 24840 63532
rect 24896 63476 24944 63532
rect 25000 63476 25048 63532
rect 25104 63476 25152 63532
rect 25208 63476 25228 63532
rect 19404 62514 19460 62524
rect 19292 61506 19348 61516
rect 23988 61964 25228 63476
rect 23988 61908 24008 61964
rect 24064 61908 24112 61964
rect 24168 61908 24216 61964
rect 24272 61908 24320 61964
rect 24376 61908 24424 61964
rect 24480 61908 24528 61964
rect 24584 61908 24632 61964
rect 24688 61908 24736 61964
rect 24792 61908 24840 61964
rect 24896 61908 24944 61964
rect 25000 61908 25048 61964
rect 25104 61908 25152 61964
rect 25208 61908 25228 61964
rect 13988 61124 14008 61180
rect 14064 61124 14112 61180
rect 14168 61124 14216 61180
rect 14272 61124 14320 61180
rect 14376 61124 14424 61180
rect 14480 61124 14528 61180
rect 14584 61124 14632 61180
rect 14688 61124 14736 61180
rect 14792 61124 14840 61180
rect 14896 61124 14944 61180
rect 15000 61124 15048 61180
rect 15104 61124 15152 61180
rect 15208 61124 15228 61180
rect 13988 59612 15228 61124
rect 13988 59556 14008 59612
rect 14064 59556 14112 59612
rect 14168 59556 14216 59612
rect 14272 59556 14320 59612
rect 14376 59556 14424 59612
rect 14480 59556 14528 59612
rect 14584 59556 14632 59612
rect 14688 59556 14736 59612
rect 14792 59556 14840 59612
rect 14896 59556 14944 59612
rect 15000 59556 15048 59612
rect 15104 59556 15152 59612
rect 15208 59556 15228 59612
rect 23988 60396 25228 61908
rect 25340 66948 25396 66958
rect 25340 65380 25396 66892
rect 25340 63028 25396 65324
rect 33988 65884 35228 67396
rect 33988 65828 34008 65884
rect 34064 65828 34112 65884
rect 34168 65828 34216 65884
rect 34272 65828 34320 65884
rect 34376 65828 34424 65884
rect 34480 65828 34528 65884
rect 34584 65828 34632 65884
rect 34688 65828 34736 65884
rect 34792 65828 34840 65884
rect 34896 65828 34944 65884
rect 35000 65828 35048 65884
rect 35104 65828 35152 65884
rect 35208 65828 35228 65884
rect 33988 64316 35228 65828
rect 33988 64260 34008 64316
rect 34064 64260 34112 64316
rect 34168 64260 34216 64316
rect 34272 64260 34320 64316
rect 34376 64260 34424 64316
rect 34480 64260 34528 64316
rect 34584 64260 34632 64316
rect 34688 64260 34736 64316
rect 34792 64260 34840 64316
rect 34896 64260 34944 64316
rect 35000 64260 35048 64316
rect 35104 64260 35152 64316
rect 35208 64260 35228 64316
rect 25340 61460 25396 62972
rect 33852 63252 33908 63262
rect 33852 62468 33908 63196
rect 33852 62402 33908 62412
rect 33988 62748 35228 64260
rect 33988 62692 34008 62748
rect 34064 62692 34112 62748
rect 34168 62692 34216 62748
rect 34272 62692 34320 62748
rect 34376 62692 34424 62748
rect 34480 62692 34528 62748
rect 34584 62692 34632 62748
rect 34688 62692 34736 62748
rect 34792 62692 34840 62748
rect 34896 62692 34944 62748
rect 35000 62692 35048 62748
rect 35104 62692 35152 62748
rect 35208 62692 35228 62748
rect 25340 61394 25396 61404
rect 23988 60340 24008 60396
rect 24064 60340 24112 60396
rect 24168 60340 24216 60396
rect 24272 60340 24320 60396
rect 24376 60340 24424 60396
rect 24480 60340 24528 60396
rect 24584 60340 24632 60396
rect 24688 60340 24736 60396
rect 24792 60340 24840 60396
rect 24896 60340 24944 60396
rect 25000 60340 25048 60396
rect 25104 60340 25152 60396
rect 25208 60340 25228 60396
rect 13468 58706 13524 58716
rect 3988 57204 4008 57260
rect 4064 57204 4112 57260
rect 4168 57204 4216 57260
rect 4272 57204 4320 57260
rect 4376 57204 4424 57260
rect 4480 57204 4528 57260
rect 4584 57204 4632 57260
rect 4688 57204 4736 57260
rect 4792 57204 4840 57260
rect 4896 57204 4944 57260
rect 5000 57204 5048 57260
rect 5104 57204 5152 57260
rect 5208 57204 5228 57260
rect 3988 55692 5228 57204
rect 7420 58660 7476 58670
rect 3988 55636 4008 55692
rect 4064 55636 4112 55692
rect 4168 55636 4216 55692
rect 4272 55636 4320 55692
rect 4376 55636 4424 55692
rect 4480 55636 4528 55692
rect 4584 55636 4632 55692
rect 4688 55636 4736 55692
rect 4792 55636 4840 55692
rect 4896 55636 4944 55692
rect 5000 55636 5048 55692
rect 5104 55636 5152 55692
rect 5208 55636 5228 55692
rect 3988 54124 5228 55636
rect 3988 54068 4008 54124
rect 4064 54068 4112 54124
rect 4168 54068 4216 54124
rect 4272 54068 4320 54124
rect 4376 54068 4424 54124
rect 4480 54068 4528 54124
rect 4584 54068 4632 54124
rect 4688 54068 4736 54124
rect 4792 54068 4840 54124
rect 4896 54068 4944 54124
rect 5000 54068 5048 54124
rect 5104 54068 5152 54124
rect 5208 54068 5228 54124
rect 3500 53172 3556 53182
rect 3500 51716 3556 53116
rect 3500 51650 3556 51660
rect 3988 52556 5228 54068
rect 3988 52500 4008 52556
rect 4064 52500 4112 52556
rect 4168 52500 4216 52556
rect 4272 52500 4320 52556
rect 4376 52500 4424 52556
rect 4480 52500 4528 52556
rect 4584 52500 4632 52556
rect 4688 52500 4736 52556
rect 4792 52500 4840 52556
rect 4896 52500 4944 52556
rect 5000 52500 5048 52556
rect 5104 52500 5152 52556
rect 5208 52500 5228 52556
rect 3988 50988 5228 52500
rect 5292 56644 5348 56654
rect 5292 52836 5348 56588
rect 6300 54628 6356 54638
rect 6300 53060 6356 54572
rect 7420 53172 7476 58604
rect 13988 58044 15228 59556
rect 19068 59556 19124 59566
rect 18508 58660 18564 58670
rect 13692 57988 13748 57998
rect 13468 56756 13524 56766
rect 7420 53106 7476 53116
rect 10108 55524 10164 55534
rect 6300 52994 6356 53004
rect 5292 51716 5348 52780
rect 5292 51650 5348 51660
rect 3988 50932 4008 50988
rect 4064 50932 4112 50988
rect 4168 50932 4216 50988
rect 4272 50932 4320 50988
rect 4376 50932 4424 50988
rect 4480 50932 4528 50988
rect 4584 50932 4632 50988
rect 4688 50932 4736 50988
rect 4792 50932 4840 50988
rect 4896 50932 4944 50988
rect 5000 50932 5048 50988
rect 5104 50932 5152 50988
rect 5208 50932 5228 50988
rect 3988 49420 5228 50932
rect 3988 49364 4008 49420
rect 4064 49364 4112 49420
rect 4168 49364 4216 49420
rect 4272 49364 4320 49420
rect 4376 49364 4424 49420
rect 4480 49364 4528 49420
rect 4584 49364 4632 49420
rect 4688 49364 4736 49420
rect 4792 49364 4840 49420
rect 4896 49364 4944 49420
rect 5000 49364 5048 49420
rect 5104 49364 5152 49420
rect 5208 49364 5228 49420
rect 3988 47852 5228 49364
rect 3988 47796 4008 47852
rect 4064 47796 4112 47852
rect 4168 47796 4216 47852
rect 4272 47796 4320 47852
rect 4376 47796 4424 47852
rect 4480 47796 4528 47852
rect 4584 47796 4632 47852
rect 4688 47796 4736 47852
rect 4792 47796 4840 47852
rect 4896 47796 4944 47852
rect 5000 47796 5048 47852
rect 5104 47796 5152 47852
rect 5208 47796 5228 47852
rect 3388 47572 3444 47582
rect 3388 43988 3444 47516
rect 3988 46284 5228 47796
rect 5292 48132 5348 48142
rect 5292 47124 5348 48076
rect 10108 47460 10164 55468
rect 13468 55412 13524 56700
rect 11900 53620 11956 53630
rect 11900 52164 11956 53564
rect 13468 52500 13524 55356
rect 13468 52434 13524 52444
rect 13580 56196 13636 56206
rect 11900 52098 11956 52108
rect 13580 51604 13636 56140
rect 13580 51538 13636 51548
rect 10108 47394 10164 47404
rect 5292 47058 5348 47068
rect 3988 46228 4008 46284
rect 4064 46228 4112 46284
rect 4168 46228 4216 46284
rect 4272 46228 4320 46284
rect 4376 46228 4424 46284
rect 4480 46228 4528 46284
rect 4584 46228 4632 46284
rect 4688 46228 4736 46284
rect 4792 46228 4840 46284
rect 4896 46228 4944 46284
rect 5000 46228 5048 46284
rect 5104 46228 5152 46284
rect 5208 46228 5228 46284
rect 3988 44716 5228 46228
rect 13692 45332 13748 57932
rect 13988 57988 14008 58044
rect 14064 57988 14112 58044
rect 14168 57988 14216 58044
rect 14272 57988 14320 58044
rect 14376 57988 14424 58044
rect 14480 57988 14528 58044
rect 14584 57988 14632 58044
rect 14688 57988 14736 58044
rect 14792 57988 14840 58044
rect 14896 57988 14944 58044
rect 15000 57988 15048 58044
rect 15104 57988 15152 58044
rect 15208 57988 15228 58044
rect 13804 56868 13860 56878
rect 13804 55748 13860 56812
rect 13804 55682 13860 55692
rect 13988 56476 15228 57988
rect 13988 56420 14008 56476
rect 14064 56420 14112 56476
rect 14168 56420 14216 56476
rect 14272 56420 14320 56476
rect 14376 56420 14424 56476
rect 14480 56420 14528 56476
rect 14584 56420 14632 56476
rect 14688 56420 14736 56476
rect 14792 56420 14840 56476
rect 14896 56420 14944 56476
rect 15000 56420 15048 56476
rect 15104 56420 15152 56476
rect 15208 56420 15228 56476
rect 13804 55188 13860 55198
rect 13804 51716 13860 55132
rect 13804 50596 13860 51660
rect 13804 50530 13860 50540
rect 13988 54908 15228 56420
rect 13988 54852 14008 54908
rect 14064 54852 14112 54908
rect 14168 54852 14216 54908
rect 14272 54852 14320 54908
rect 14376 54852 14424 54908
rect 14480 54852 14528 54908
rect 14584 54852 14632 54908
rect 14688 54852 14736 54908
rect 14792 54852 14840 54908
rect 14896 54852 14944 54908
rect 15000 54852 15048 54908
rect 15104 54852 15152 54908
rect 15208 54852 15228 54908
rect 13988 53340 15228 54852
rect 15372 58212 15428 58222
rect 15372 53956 15428 58156
rect 18508 56308 18564 58604
rect 18508 56242 18564 56252
rect 19068 55412 19124 59500
rect 19292 58884 19348 58894
rect 19292 57428 19348 58828
rect 23988 58828 25228 60340
rect 19740 58772 19796 58782
rect 19292 57362 19348 57372
rect 19628 58660 19684 58670
rect 19068 55346 19124 55356
rect 15372 53890 15428 53900
rect 13988 53284 14008 53340
rect 14064 53284 14112 53340
rect 14168 53284 14216 53340
rect 14272 53284 14320 53340
rect 14376 53284 14424 53340
rect 14480 53284 14528 53340
rect 14584 53284 14632 53340
rect 14688 53284 14736 53340
rect 14792 53284 14840 53340
rect 14896 53284 14944 53340
rect 15000 53284 15048 53340
rect 15104 53284 15152 53340
rect 15208 53284 15228 53340
rect 13988 51772 15228 53284
rect 13988 51716 14008 51772
rect 14064 51716 14112 51772
rect 14168 51716 14216 51772
rect 14272 51716 14320 51772
rect 14376 51716 14424 51772
rect 14480 51716 14528 51772
rect 14584 51716 14632 51772
rect 14688 51716 14736 51772
rect 14792 51716 14840 51772
rect 14896 51716 14944 51772
rect 15000 51716 15048 51772
rect 15104 51716 15152 51772
rect 15208 51716 15228 51772
rect 13988 50204 15228 51716
rect 13988 50148 14008 50204
rect 14064 50148 14112 50204
rect 14168 50148 14216 50204
rect 14272 50148 14320 50204
rect 14376 50148 14424 50204
rect 14480 50148 14528 50204
rect 14584 50148 14632 50204
rect 14688 50148 14736 50204
rect 14792 50148 14840 50204
rect 14896 50148 14944 50204
rect 15000 50148 15048 50204
rect 15104 50148 15152 50204
rect 15208 50148 15228 50204
rect 13804 49028 13860 49038
rect 13804 47460 13860 48972
rect 13804 47394 13860 47404
rect 13988 48636 15228 50148
rect 13988 48580 14008 48636
rect 14064 48580 14112 48636
rect 14168 48580 14216 48636
rect 14272 48580 14320 48636
rect 14376 48580 14424 48636
rect 14480 48580 14528 48636
rect 14584 48580 14632 48636
rect 14688 48580 14736 48636
rect 14792 48580 14840 48636
rect 14896 48580 14944 48636
rect 15000 48580 15048 48636
rect 15104 48580 15152 48636
rect 15208 48580 15228 48636
rect 13692 45266 13748 45276
rect 13988 47068 15228 48580
rect 13988 47012 14008 47068
rect 14064 47012 14112 47068
rect 14168 47012 14216 47068
rect 14272 47012 14320 47068
rect 14376 47012 14424 47068
rect 14480 47012 14528 47068
rect 14584 47012 14632 47068
rect 14688 47012 14736 47068
rect 14792 47012 14840 47068
rect 14896 47012 14944 47068
rect 15000 47012 15048 47068
rect 15104 47012 15152 47068
rect 15208 47012 15228 47068
rect 13988 45500 15228 47012
rect 15372 53508 15428 53518
rect 15372 47012 15428 53452
rect 19628 50708 19684 58604
rect 19740 57428 19796 58716
rect 19740 57362 19796 57372
rect 23988 58772 24008 58828
rect 24064 58772 24112 58828
rect 24168 58772 24216 58828
rect 24272 58772 24320 58828
rect 24376 58772 24424 58828
rect 24480 58772 24528 58828
rect 24584 58772 24632 58828
rect 24688 58772 24736 58828
rect 24792 58772 24840 58828
rect 24896 58772 24944 58828
rect 25000 58772 25048 58828
rect 25104 58772 25152 58828
rect 25208 58772 25228 58828
rect 19628 50642 19684 50652
rect 23988 57260 25228 58772
rect 23988 57204 24008 57260
rect 24064 57204 24112 57260
rect 24168 57204 24216 57260
rect 24272 57204 24320 57260
rect 24376 57204 24424 57260
rect 24480 57204 24528 57260
rect 24584 57204 24632 57260
rect 24688 57204 24736 57260
rect 24792 57204 24840 57260
rect 24896 57204 24944 57260
rect 25000 57204 25048 57260
rect 25104 57204 25152 57260
rect 25208 57204 25228 57260
rect 23988 55692 25228 57204
rect 23988 55636 24008 55692
rect 24064 55636 24112 55692
rect 24168 55636 24216 55692
rect 24272 55636 24320 55692
rect 24376 55636 24424 55692
rect 24480 55636 24528 55692
rect 24584 55636 24632 55692
rect 24688 55636 24736 55692
rect 24792 55636 24840 55692
rect 24896 55636 24944 55692
rect 25000 55636 25048 55692
rect 25104 55636 25152 55692
rect 25208 55636 25228 55692
rect 23988 54124 25228 55636
rect 23988 54068 24008 54124
rect 24064 54068 24112 54124
rect 24168 54068 24216 54124
rect 24272 54068 24320 54124
rect 24376 54068 24424 54124
rect 24480 54068 24528 54124
rect 24584 54068 24632 54124
rect 24688 54068 24736 54124
rect 24792 54068 24840 54124
rect 24896 54068 24944 54124
rect 25000 54068 25048 54124
rect 25104 54068 25152 54124
rect 25208 54068 25228 54124
rect 23988 52556 25228 54068
rect 23988 52500 24008 52556
rect 24064 52500 24112 52556
rect 24168 52500 24216 52556
rect 24272 52500 24320 52556
rect 24376 52500 24424 52556
rect 24480 52500 24528 52556
rect 24584 52500 24632 52556
rect 24688 52500 24736 52556
rect 24792 52500 24840 52556
rect 24896 52500 24944 52556
rect 25000 52500 25048 52556
rect 25104 52500 25152 52556
rect 25208 52500 25228 52556
rect 23988 50988 25228 52500
rect 23988 50932 24008 50988
rect 24064 50932 24112 50988
rect 24168 50932 24216 50988
rect 24272 50932 24320 50988
rect 24376 50932 24424 50988
rect 24480 50932 24528 50988
rect 24584 50932 24632 50988
rect 24688 50932 24736 50988
rect 24792 50932 24840 50988
rect 24896 50932 24944 50988
rect 25000 50932 25048 50988
rect 25104 50932 25152 50988
rect 25208 50932 25228 50988
rect 15372 46946 15428 46956
rect 23988 49420 25228 50932
rect 33988 61180 35228 62692
rect 33988 61124 34008 61180
rect 34064 61124 34112 61180
rect 34168 61124 34216 61180
rect 34272 61124 34320 61180
rect 34376 61124 34424 61180
rect 34480 61124 34528 61180
rect 34584 61124 34632 61180
rect 34688 61124 34736 61180
rect 34792 61124 34840 61180
rect 34896 61124 34944 61180
rect 35000 61124 35048 61180
rect 35104 61124 35152 61180
rect 35208 61124 35228 61180
rect 33988 59612 35228 61124
rect 33988 59556 34008 59612
rect 34064 59556 34112 59612
rect 34168 59556 34216 59612
rect 34272 59556 34320 59612
rect 34376 59556 34424 59612
rect 34480 59556 34528 59612
rect 34584 59556 34632 59612
rect 34688 59556 34736 59612
rect 34792 59556 34840 59612
rect 34896 59556 34944 59612
rect 35000 59556 35048 59612
rect 35104 59556 35152 59612
rect 35208 59556 35228 59612
rect 33988 58044 35228 59556
rect 33988 57988 34008 58044
rect 34064 57988 34112 58044
rect 34168 57988 34216 58044
rect 34272 57988 34320 58044
rect 34376 57988 34424 58044
rect 34480 57988 34528 58044
rect 34584 57988 34632 58044
rect 34688 57988 34736 58044
rect 34792 57988 34840 58044
rect 34896 57988 34944 58044
rect 35000 57988 35048 58044
rect 35104 57988 35152 58044
rect 35208 57988 35228 58044
rect 33988 56476 35228 57988
rect 33988 56420 34008 56476
rect 34064 56420 34112 56476
rect 34168 56420 34216 56476
rect 34272 56420 34320 56476
rect 34376 56420 34424 56476
rect 34480 56420 34528 56476
rect 34584 56420 34632 56476
rect 34688 56420 34736 56476
rect 34792 56420 34840 56476
rect 34896 56420 34944 56476
rect 35000 56420 35048 56476
rect 35104 56420 35152 56476
rect 35208 56420 35228 56476
rect 33988 54908 35228 56420
rect 33988 54852 34008 54908
rect 34064 54852 34112 54908
rect 34168 54852 34216 54908
rect 34272 54852 34320 54908
rect 34376 54852 34424 54908
rect 34480 54852 34528 54908
rect 34584 54852 34632 54908
rect 34688 54852 34736 54908
rect 34792 54852 34840 54908
rect 34896 54852 34944 54908
rect 35000 54852 35048 54908
rect 35104 54852 35152 54908
rect 35208 54852 35228 54908
rect 33988 53340 35228 54852
rect 33988 53284 34008 53340
rect 34064 53284 34112 53340
rect 34168 53284 34216 53340
rect 34272 53284 34320 53340
rect 34376 53284 34424 53340
rect 34480 53284 34528 53340
rect 34584 53284 34632 53340
rect 34688 53284 34736 53340
rect 34792 53284 34840 53340
rect 34896 53284 34944 53340
rect 35000 53284 35048 53340
rect 35104 53284 35152 53340
rect 35208 53284 35228 53340
rect 33988 51772 35228 53284
rect 33988 51716 34008 51772
rect 34064 51716 34112 51772
rect 34168 51716 34216 51772
rect 34272 51716 34320 51772
rect 34376 51716 34424 51772
rect 34480 51716 34528 51772
rect 34584 51716 34632 51772
rect 34688 51716 34736 51772
rect 34792 51716 34840 51772
rect 34896 51716 34944 51772
rect 35000 51716 35048 51772
rect 35104 51716 35152 51772
rect 35208 51716 35228 51772
rect 23988 49364 24008 49420
rect 24064 49364 24112 49420
rect 24168 49364 24216 49420
rect 24272 49364 24320 49420
rect 24376 49364 24424 49420
rect 24480 49364 24528 49420
rect 24584 49364 24632 49420
rect 24688 49364 24736 49420
rect 24792 49364 24840 49420
rect 24896 49364 24944 49420
rect 25000 49364 25048 49420
rect 25104 49364 25152 49420
rect 25208 49364 25228 49420
rect 23988 47852 25228 49364
rect 33852 50484 33908 50494
rect 33852 48804 33908 50428
rect 33852 48738 33908 48748
rect 33988 50204 35228 51716
rect 33988 50148 34008 50204
rect 34064 50148 34112 50204
rect 34168 50148 34216 50204
rect 34272 50148 34320 50204
rect 34376 50148 34424 50204
rect 34480 50148 34528 50204
rect 34584 50148 34632 50204
rect 34688 50148 34736 50204
rect 34792 50148 34840 50204
rect 34896 50148 34944 50204
rect 35000 50148 35048 50204
rect 35104 50148 35152 50204
rect 35208 50148 35228 50204
rect 23988 47796 24008 47852
rect 24064 47796 24112 47852
rect 24168 47796 24216 47852
rect 24272 47796 24320 47852
rect 24376 47796 24424 47852
rect 24480 47796 24528 47852
rect 24584 47796 24632 47852
rect 24688 47796 24736 47852
rect 24792 47796 24840 47852
rect 24896 47796 24944 47852
rect 25000 47796 25048 47852
rect 25104 47796 25152 47852
rect 25208 47796 25228 47852
rect 13988 45444 14008 45500
rect 14064 45444 14112 45500
rect 14168 45444 14216 45500
rect 14272 45444 14320 45500
rect 14376 45444 14424 45500
rect 14480 45444 14528 45500
rect 14584 45444 14632 45500
rect 14688 45444 14736 45500
rect 14792 45444 14840 45500
rect 14896 45444 14944 45500
rect 15000 45444 15048 45500
rect 15104 45444 15152 45500
rect 15208 45444 15228 45500
rect 3988 44660 4008 44716
rect 4064 44660 4112 44716
rect 4168 44660 4216 44716
rect 4272 44660 4320 44716
rect 4376 44660 4424 44716
rect 4480 44660 4528 44716
rect 4584 44660 4632 44716
rect 4688 44660 4736 44716
rect 4792 44660 4840 44716
rect 4896 44660 4944 44716
rect 5000 44660 5048 44716
rect 5104 44660 5152 44716
rect 5208 44660 5228 44716
rect 3388 43652 3444 43932
rect 3388 43586 3444 43596
rect 3836 44548 3892 44558
rect 3836 39620 3892 44492
rect 3836 39554 3892 39564
rect 3988 43148 5228 44660
rect 3988 43092 4008 43148
rect 4064 43092 4112 43148
rect 4168 43092 4216 43148
rect 4272 43092 4320 43148
rect 4376 43092 4424 43148
rect 4480 43092 4528 43148
rect 4584 43092 4632 43148
rect 4688 43092 4736 43148
rect 4792 43092 4840 43148
rect 4896 43092 4944 43148
rect 5000 43092 5048 43148
rect 5104 43092 5152 43148
rect 5208 43092 5228 43148
rect 3988 41580 5228 43092
rect 3988 41524 4008 41580
rect 4064 41524 4112 41580
rect 4168 41524 4216 41580
rect 4272 41524 4320 41580
rect 4376 41524 4424 41580
rect 4480 41524 4528 41580
rect 4584 41524 4632 41580
rect 4688 41524 4736 41580
rect 4792 41524 4840 41580
rect 4896 41524 4944 41580
rect 5000 41524 5048 41580
rect 5104 41524 5152 41580
rect 5208 41524 5228 41580
rect 3988 40012 5228 41524
rect 3988 39956 4008 40012
rect 4064 39956 4112 40012
rect 4168 39956 4216 40012
rect 4272 39956 4320 40012
rect 4376 39956 4424 40012
rect 4480 39956 4528 40012
rect 4584 39956 4632 40012
rect 4688 39956 4736 40012
rect 4792 39956 4840 40012
rect 4896 39956 4944 40012
rect 5000 39956 5048 40012
rect 5104 39956 5152 40012
rect 5208 39956 5228 40012
rect 3988 38444 5228 39956
rect 5964 44884 6020 44894
rect 5964 39508 6020 44828
rect 5964 39442 6020 39452
rect 13988 43932 15228 45444
rect 13988 43876 14008 43932
rect 14064 43876 14112 43932
rect 14168 43876 14216 43932
rect 14272 43876 14320 43932
rect 14376 43876 14424 43932
rect 14480 43876 14528 43932
rect 14584 43876 14632 43932
rect 14688 43876 14736 43932
rect 14792 43876 14840 43932
rect 14896 43876 14944 43932
rect 15000 43876 15048 43932
rect 15104 43876 15152 43932
rect 15208 43876 15228 43932
rect 13988 42364 15228 43876
rect 13988 42308 14008 42364
rect 14064 42308 14112 42364
rect 14168 42308 14216 42364
rect 14272 42308 14320 42364
rect 14376 42308 14424 42364
rect 14480 42308 14528 42364
rect 14584 42308 14632 42364
rect 14688 42308 14736 42364
rect 14792 42308 14840 42364
rect 14896 42308 14944 42364
rect 15000 42308 15048 42364
rect 15104 42308 15152 42364
rect 15208 42308 15228 42364
rect 13988 40796 15228 42308
rect 13988 40740 14008 40796
rect 14064 40740 14112 40796
rect 14168 40740 14216 40796
rect 14272 40740 14320 40796
rect 14376 40740 14424 40796
rect 14480 40740 14528 40796
rect 14584 40740 14632 40796
rect 14688 40740 14736 40796
rect 14792 40740 14840 40796
rect 14896 40740 14944 40796
rect 15000 40740 15048 40796
rect 15104 40740 15152 40796
rect 15208 40740 15228 40796
rect 3988 38388 4008 38444
rect 4064 38388 4112 38444
rect 4168 38388 4216 38444
rect 4272 38388 4320 38444
rect 4376 38388 4424 38444
rect 4480 38388 4528 38444
rect 4584 38388 4632 38444
rect 4688 38388 4736 38444
rect 4792 38388 4840 38444
rect 4896 38388 4944 38444
rect 5000 38388 5048 38444
rect 5104 38388 5152 38444
rect 5208 38388 5228 38444
rect 3988 36876 5228 38388
rect 3988 36820 4008 36876
rect 4064 36820 4112 36876
rect 4168 36820 4216 36876
rect 4272 36820 4320 36876
rect 4376 36820 4424 36876
rect 4480 36820 4528 36876
rect 4584 36820 4632 36876
rect 4688 36820 4736 36876
rect 4792 36820 4840 36876
rect 4896 36820 4944 36876
rect 5000 36820 5048 36876
rect 5104 36820 5152 36876
rect 5208 36820 5228 36876
rect 3988 35308 5228 36820
rect 3988 35252 4008 35308
rect 4064 35252 4112 35308
rect 4168 35252 4216 35308
rect 4272 35252 4320 35308
rect 4376 35252 4424 35308
rect 4480 35252 4528 35308
rect 4584 35252 4632 35308
rect 4688 35252 4736 35308
rect 4792 35252 4840 35308
rect 4896 35252 4944 35308
rect 5000 35252 5048 35308
rect 5104 35252 5152 35308
rect 5208 35252 5228 35308
rect 3988 33740 5228 35252
rect 13988 39228 15228 40740
rect 13988 39172 14008 39228
rect 14064 39172 14112 39228
rect 14168 39172 14216 39228
rect 14272 39172 14320 39228
rect 14376 39172 14424 39228
rect 14480 39172 14528 39228
rect 14584 39172 14632 39228
rect 14688 39172 14736 39228
rect 14792 39172 14840 39228
rect 14896 39172 14944 39228
rect 15000 39172 15048 39228
rect 15104 39172 15152 39228
rect 15208 39172 15228 39228
rect 13988 37660 15228 39172
rect 17612 46564 17668 46574
rect 17612 45780 17668 46508
rect 17612 38500 17668 45724
rect 23988 46284 25228 47796
rect 23988 46228 24008 46284
rect 24064 46228 24112 46284
rect 24168 46228 24216 46284
rect 24272 46228 24320 46284
rect 24376 46228 24424 46284
rect 24480 46228 24528 46284
rect 24584 46228 24632 46284
rect 24688 46228 24736 46284
rect 24792 46228 24840 46284
rect 24896 46228 24944 46284
rect 25000 46228 25048 46284
rect 25104 46228 25152 46284
rect 25208 46228 25228 46284
rect 23988 44716 25228 46228
rect 33988 48636 35228 50148
rect 33988 48580 34008 48636
rect 34064 48580 34112 48636
rect 34168 48580 34216 48636
rect 34272 48580 34320 48636
rect 34376 48580 34424 48636
rect 34480 48580 34528 48636
rect 34584 48580 34632 48636
rect 34688 48580 34736 48636
rect 34792 48580 34840 48636
rect 34896 48580 34944 48636
rect 35000 48580 35048 48636
rect 35104 48580 35152 48636
rect 35208 48580 35228 48636
rect 33988 47068 35228 48580
rect 33988 47012 34008 47068
rect 34064 47012 34112 47068
rect 34168 47012 34216 47068
rect 34272 47012 34320 47068
rect 34376 47012 34424 47068
rect 34480 47012 34528 47068
rect 34584 47012 34632 47068
rect 34688 47012 34736 47068
rect 34792 47012 34840 47068
rect 34896 47012 34944 47068
rect 35000 47012 35048 47068
rect 35104 47012 35152 47068
rect 35208 47012 35228 47068
rect 23988 44660 24008 44716
rect 24064 44660 24112 44716
rect 24168 44660 24216 44716
rect 24272 44660 24320 44716
rect 24376 44660 24424 44716
rect 24480 44660 24528 44716
rect 24584 44660 24632 44716
rect 24688 44660 24736 44716
rect 24792 44660 24840 44716
rect 24896 44660 24944 44716
rect 25000 44660 25048 44716
rect 25104 44660 25152 44716
rect 25208 44660 25228 44716
rect 23772 44436 23828 44446
rect 23548 42868 23604 42878
rect 23548 39732 23604 42812
rect 23548 39666 23604 39676
rect 23660 40740 23716 40750
rect 17612 38434 17668 38444
rect 23100 39620 23156 39630
rect 13988 37604 14008 37660
rect 14064 37604 14112 37660
rect 14168 37604 14216 37660
rect 14272 37604 14320 37660
rect 14376 37604 14424 37660
rect 14480 37604 14528 37660
rect 14584 37604 14632 37660
rect 14688 37604 14736 37660
rect 14792 37604 14840 37660
rect 14896 37604 14944 37660
rect 15000 37604 15048 37660
rect 15104 37604 15152 37660
rect 15208 37604 15228 37660
rect 13988 36092 15228 37604
rect 23100 36260 23156 39564
rect 23660 39620 23716 40684
rect 23660 39554 23716 39564
rect 23772 37380 23828 44380
rect 23772 37314 23828 37324
rect 23988 43148 25228 44660
rect 23988 43092 24008 43148
rect 24064 43092 24112 43148
rect 24168 43092 24216 43148
rect 24272 43092 24320 43148
rect 24376 43092 24424 43148
rect 24480 43092 24528 43148
rect 24584 43092 24632 43148
rect 24688 43092 24736 43148
rect 24792 43092 24840 43148
rect 24896 43092 24944 43148
rect 25000 43092 25048 43148
rect 25104 43092 25152 43148
rect 25208 43092 25228 43148
rect 23988 41580 25228 43092
rect 23988 41524 24008 41580
rect 24064 41524 24112 41580
rect 24168 41524 24216 41580
rect 24272 41524 24320 41580
rect 24376 41524 24424 41580
rect 24480 41524 24528 41580
rect 24584 41524 24632 41580
rect 24688 41524 24736 41580
rect 24792 41524 24840 41580
rect 24896 41524 24944 41580
rect 25000 41524 25048 41580
rect 25104 41524 25152 41580
rect 25208 41524 25228 41580
rect 23988 40012 25228 41524
rect 25788 46004 25844 46014
rect 25788 40404 25844 45948
rect 33988 45500 35228 47012
rect 33988 45444 34008 45500
rect 34064 45444 34112 45500
rect 34168 45444 34216 45500
rect 34272 45444 34320 45500
rect 34376 45444 34424 45500
rect 34480 45444 34528 45500
rect 34584 45444 34632 45500
rect 34688 45444 34736 45500
rect 34792 45444 34840 45500
rect 34896 45444 34944 45500
rect 35000 45444 35048 45500
rect 35104 45444 35152 45500
rect 35208 45444 35228 45500
rect 33516 44324 33572 44334
rect 33516 43428 33572 44268
rect 25788 40338 25844 40348
rect 33404 43092 33460 43102
rect 23988 39956 24008 40012
rect 24064 39956 24112 40012
rect 24168 39956 24216 40012
rect 24272 39956 24320 40012
rect 24376 39956 24424 40012
rect 24480 39956 24528 40012
rect 24584 39956 24632 40012
rect 24688 39956 24736 40012
rect 24792 39956 24840 40012
rect 24896 39956 24944 40012
rect 25000 39956 25048 40012
rect 25104 39956 25152 40012
rect 25208 39956 25228 40012
rect 23988 38444 25228 39956
rect 23988 38388 24008 38444
rect 24064 38388 24112 38444
rect 24168 38388 24216 38444
rect 24272 38388 24320 38444
rect 24376 38388 24424 38444
rect 24480 38388 24528 38444
rect 24584 38388 24632 38444
rect 24688 38388 24736 38444
rect 24792 38388 24840 38444
rect 24896 38388 24944 38444
rect 25000 38388 25048 38444
rect 25104 38388 25152 38444
rect 25208 38388 25228 38444
rect 23100 36194 23156 36204
rect 23988 36876 25228 38388
rect 33404 37716 33460 43036
rect 33516 38500 33572 43372
rect 33628 44100 33684 44110
rect 33628 42868 33684 44044
rect 33628 39732 33684 42812
rect 33988 43932 35228 45444
rect 33988 43876 34008 43932
rect 34064 43876 34112 43932
rect 34168 43876 34216 43932
rect 34272 43876 34320 43932
rect 34376 43876 34424 43932
rect 34480 43876 34528 43932
rect 34584 43876 34632 43932
rect 34688 43876 34736 43932
rect 34792 43876 34840 43932
rect 34896 43876 34944 43932
rect 35000 43876 35048 43932
rect 35104 43876 35152 43932
rect 35208 43876 35228 43932
rect 33988 42364 35228 43876
rect 33988 42308 34008 42364
rect 34064 42308 34112 42364
rect 34168 42308 34216 42364
rect 34272 42308 34320 42364
rect 34376 42308 34424 42364
rect 34480 42308 34528 42364
rect 34584 42308 34632 42364
rect 34688 42308 34736 42364
rect 34792 42308 34840 42364
rect 34896 42308 34944 42364
rect 35000 42308 35048 42364
rect 35104 42308 35152 42364
rect 35208 42308 35228 42364
rect 33740 41524 33796 41534
rect 33740 40628 33796 41468
rect 33740 40562 33796 40572
rect 33852 41076 33908 41086
rect 33628 39666 33684 39676
rect 33852 39060 33908 41020
rect 33852 38668 33908 39004
rect 33516 38434 33572 38444
rect 33740 38612 33908 38668
rect 33988 40796 35228 42308
rect 33988 40740 34008 40796
rect 34064 40740 34112 40796
rect 34168 40740 34216 40796
rect 34272 40740 34320 40796
rect 34376 40740 34424 40796
rect 34480 40740 34528 40796
rect 34584 40740 34632 40796
rect 34688 40740 34736 40796
rect 34792 40740 34840 40796
rect 34896 40740 34944 40796
rect 35000 40740 35048 40796
rect 35104 40740 35152 40796
rect 35208 40740 35228 40796
rect 33988 39228 35228 40740
rect 33988 39172 34008 39228
rect 34064 39172 34112 39228
rect 34168 39172 34216 39228
rect 34272 39172 34320 39228
rect 34376 39172 34424 39228
rect 34480 39172 34528 39228
rect 34584 39172 34632 39228
rect 34688 39172 34736 39228
rect 34792 39172 34840 39228
rect 34896 39172 34944 39228
rect 35000 39172 35048 39228
rect 35104 39172 35152 39228
rect 35208 39172 35228 39228
rect 33404 37650 33460 37660
rect 23988 36820 24008 36876
rect 24064 36820 24112 36876
rect 24168 36820 24216 36876
rect 24272 36820 24320 36876
rect 24376 36820 24424 36876
rect 24480 36820 24528 36876
rect 24584 36820 24632 36876
rect 24688 36820 24736 36876
rect 24792 36820 24840 36876
rect 24896 36820 24944 36876
rect 25000 36820 25048 36876
rect 25104 36820 25152 36876
rect 25208 36820 25228 36876
rect 13988 36036 14008 36092
rect 14064 36036 14112 36092
rect 14168 36036 14216 36092
rect 14272 36036 14320 36092
rect 14376 36036 14424 36092
rect 14480 36036 14528 36092
rect 14584 36036 14632 36092
rect 14688 36036 14736 36092
rect 14792 36036 14840 36092
rect 14896 36036 14944 36092
rect 15000 36036 15048 36092
rect 15104 36036 15152 36092
rect 15208 36036 15228 36092
rect 13804 35140 13860 35150
rect 3500 33684 3556 33694
rect 1820 32564 1876 32574
rect 1820 26628 1876 32508
rect 1820 26562 1876 26572
rect 3164 30212 3220 30222
rect 3164 25844 3220 30156
rect 3164 24724 3220 25788
rect 3164 24658 3220 24668
rect 3276 27076 3332 27086
rect 3276 23716 3332 27020
rect 3276 23650 3332 23660
rect 3388 26964 3444 26974
rect 3052 23492 3108 23502
rect 3052 17108 3108 23436
rect 3052 17042 3108 17052
rect 3388 16996 3444 26908
rect 3500 25732 3556 33628
rect 3988 33684 4008 33740
rect 4064 33684 4112 33740
rect 4168 33684 4216 33740
rect 4272 33684 4320 33740
rect 4376 33684 4424 33740
rect 4480 33684 4528 33740
rect 4584 33684 4632 33740
rect 4688 33684 4736 33740
rect 4792 33684 4840 33740
rect 4896 33684 4944 33740
rect 5000 33684 5048 33740
rect 5104 33684 5152 33740
rect 5208 33684 5228 33740
rect 3988 32172 5228 33684
rect 7308 35028 7364 35038
rect 3836 32116 3892 32126
rect 3612 28868 3668 28878
rect 3612 28420 3668 28812
rect 3836 28644 3892 32060
rect 3836 28578 3892 28588
rect 3988 32116 4008 32172
rect 4064 32116 4112 32172
rect 4168 32116 4216 32172
rect 4272 32116 4320 32172
rect 4376 32116 4424 32172
rect 4480 32116 4528 32172
rect 4584 32116 4632 32172
rect 4688 32116 4736 32172
rect 4792 32116 4840 32172
rect 4896 32116 4944 32172
rect 5000 32116 5048 32172
rect 5104 32116 5152 32172
rect 5208 32116 5228 32172
rect 3988 30604 5228 32116
rect 3988 30548 4008 30604
rect 4064 30548 4112 30604
rect 4168 30548 4216 30604
rect 4272 30548 4320 30604
rect 4376 30548 4424 30604
rect 4480 30548 4528 30604
rect 4584 30548 4632 30604
rect 4688 30548 4736 30604
rect 4792 30548 4840 30604
rect 4896 30548 4944 30604
rect 5000 30548 5048 30604
rect 5104 30548 5152 30604
rect 5208 30548 5228 30604
rect 3988 29036 5228 30548
rect 3988 28980 4008 29036
rect 4064 28980 4112 29036
rect 4168 28980 4216 29036
rect 4272 28980 4320 29036
rect 4376 28980 4424 29036
rect 4480 28980 4528 29036
rect 4584 28980 4632 29036
rect 4688 28980 4736 29036
rect 4792 28980 4840 29036
rect 4896 28980 4944 29036
rect 5000 28980 5048 29036
rect 5104 28980 5152 29036
rect 5208 28980 5228 29036
rect 3612 28354 3668 28364
rect 3988 27468 5228 28980
rect 3988 27412 4008 27468
rect 4064 27412 4112 27468
rect 4168 27412 4216 27468
rect 4272 27412 4320 27468
rect 4376 27412 4424 27468
rect 4480 27412 4528 27468
rect 4584 27412 4632 27468
rect 4688 27412 4736 27468
rect 4792 27412 4840 27468
rect 4896 27412 4944 27468
rect 5000 27412 5048 27468
rect 5104 27412 5152 27468
rect 5208 27412 5228 27468
rect 3500 25666 3556 25676
rect 3836 26516 3892 26526
rect 3836 25620 3892 26460
rect 3836 25554 3892 25564
rect 3988 25900 5228 27412
rect 3988 25844 4008 25900
rect 4064 25844 4112 25900
rect 4168 25844 4216 25900
rect 4272 25844 4320 25900
rect 4376 25844 4424 25900
rect 4480 25844 4528 25900
rect 4584 25844 4632 25900
rect 4688 25844 4736 25900
rect 4792 25844 4840 25900
rect 4896 25844 4944 25900
rect 5000 25844 5048 25900
rect 5104 25844 5152 25900
rect 5208 25844 5228 25900
rect 3988 24332 5228 25844
rect 5292 33572 5348 33582
rect 5292 30212 5348 33516
rect 5292 25396 5348 30156
rect 6076 28532 6132 28542
rect 5964 27412 6020 27422
rect 5964 26852 6020 27356
rect 5964 26786 6020 26796
rect 6076 26628 6132 28476
rect 6076 26562 6132 26572
rect 6188 27076 6244 27086
rect 5292 25330 5348 25340
rect 6188 24948 6244 27020
rect 7308 26964 7364 34972
rect 13692 35028 13748 35038
rect 13468 29988 13524 29998
rect 13468 28308 13524 29932
rect 13468 28242 13524 28252
rect 7308 26898 7364 26908
rect 13692 25620 13748 34972
rect 13804 27076 13860 35084
rect 13804 27010 13860 27020
rect 13988 34524 15228 36036
rect 13988 34468 14008 34524
rect 14064 34468 14112 34524
rect 14168 34468 14216 34524
rect 14272 34468 14320 34524
rect 14376 34468 14424 34524
rect 14480 34468 14528 34524
rect 14584 34468 14632 34524
rect 14688 34468 14736 34524
rect 14792 34468 14840 34524
rect 14896 34468 14944 34524
rect 15000 34468 15048 34524
rect 15104 34468 15152 34524
rect 15208 34468 15228 34524
rect 13988 32956 15228 34468
rect 13988 32900 14008 32956
rect 14064 32900 14112 32956
rect 14168 32900 14216 32956
rect 14272 32900 14320 32956
rect 14376 32900 14424 32956
rect 14480 32900 14528 32956
rect 14584 32900 14632 32956
rect 14688 32900 14736 32956
rect 14792 32900 14840 32956
rect 14896 32900 14944 32956
rect 15000 32900 15048 32956
rect 15104 32900 15152 32956
rect 15208 32900 15228 32956
rect 13988 31388 15228 32900
rect 23988 35308 25228 36820
rect 23988 35252 24008 35308
rect 24064 35252 24112 35308
rect 24168 35252 24216 35308
rect 24272 35252 24320 35308
rect 24376 35252 24424 35308
rect 24480 35252 24528 35308
rect 24584 35252 24632 35308
rect 24688 35252 24736 35308
rect 24792 35252 24840 35308
rect 24896 35252 24944 35308
rect 25000 35252 25048 35308
rect 25104 35252 25152 35308
rect 25208 35252 25228 35308
rect 23988 33740 25228 35252
rect 23988 33684 24008 33740
rect 24064 33684 24112 33740
rect 24168 33684 24216 33740
rect 24272 33684 24320 33740
rect 24376 33684 24424 33740
rect 24480 33684 24528 33740
rect 24584 33684 24632 33740
rect 24688 33684 24736 33740
rect 24792 33684 24840 33740
rect 24896 33684 24944 33740
rect 25000 33684 25048 33740
rect 25104 33684 25152 33740
rect 25208 33684 25228 33740
rect 15484 32788 15540 32798
rect 13988 31332 14008 31388
rect 14064 31332 14112 31388
rect 14168 31332 14216 31388
rect 14272 31332 14320 31388
rect 14376 31332 14424 31388
rect 14480 31332 14528 31388
rect 14584 31332 14632 31388
rect 14688 31332 14736 31388
rect 14792 31332 14840 31388
rect 14896 31332 14944 31388
rect 15000 31332 15048 31388
rect 15104 31332 15152 31388
rect 15208 31332 15228 31388
rect 13988 29820 15228 31332
rect 13988 29764 14008 29820
rect 14064 29764 14112 29820
rect 14168 29764 14216 29820
rect 14272 29764 14320 29820
rect 14376 29764 14424 29820
rect 14480 29764 14528 29820
rect 14584 29764 14632 29820
rect 14688 29764 14736 29820
rect 14792 29764 14840 29820
rect 14896 29764 14944 29820
rect 15000 29764 15048 29820
rect 15104 29764 15152 29820
rect 15208 29764 15228 29820
rect 13988 28252 15228 29764
rect 13988 28196 14008 28252
rect 14064 28196 14112 28252
rect 14168 28196 14216 28252
rect 14272 28196 14320 28252
rect 14376 28196 14424 28252
rect 14480 28196 14528 28252
rect 14584 28196 14632 28252
rect 14688 28196 14736 28252
rect 14792 28196 14840 28252
rect 14896 28196 14944 28252
rect 15000 28196 15048 28252
rect 15104 28196 15152 28252
rect 15208 28196 15228 28252
rect 13692 25554 13748 25564
rect 13988 26684 15228 28196
rect 13988 26628 14008 26684
rect 14064 26628 14112 26684
rect 14168 26628 14216 26684
rect 14272 26628 14320 26684
rect 14376 26628 14424 26684
rect 14480 26628 14528 26684
rect 14584 26628 14632 26684
rect 14688 26628 14736 26684
rect 14792 26628 14840 26684
rect 14896 26628 14944 26684
rect 15000 26628 15048 26684
rect 15104 26628 15152 26684
rect 15208 26628 15228 26684
rect 6188 24882 6244 24892
rect 13988 25116 15228 26628
rect 13988 25060 14008 25116
rect 14064 25060 14112 25116
rect 14168 25060 14216 25116
rect 14272 25060 14320 25116
rect 14376 25060 14424 25116
rect 14480 25060 14528 25116
rect 14584 25060 14632 25116
rect 14688 25060 14736 25116
rect 14792 25060 14840 25116
rect 14896 25060 14944 25116
rect 15000 25060 15048 25116
rect 15104 25060 15152 25116
rect 15208 25060 15228 25116
rect 3988 24276 4008 24332
rect 4064 24276 4112 24332
rect 4168 24276 4216 24332
rect 4272 24276 4320 24332
rect 4376 24276 4424 24332
rect 4480 24276 4528 24332
rect 4584 24276 4632 24332
rect 4688 24276 4736 24332
rect 4792 24276 4840 24332
rect 4896 24276 4944 24332
rect 5000 24276 5048 24332
rect 5104 24276 5152 24332
rect 5208 24276 5228 24332
rect 3388 16930 3444 16940
rect 3836 23268 3892 23278
rect 3836 13972 3892 23212
rect 3836 13906 3892 13916
rect 3988 22764 5228 24276
rect 13804 23828 13860 23838
rect 13692 23492 13748 23502
rect 3988 22708 4008 22764
rect 4064 22708 4112 22764
rect 4168 22708 4216 22764
rect 4272 22708 4320 22764
rect 4376 22708 4424 22764
rect 4480 22708 4528 22764
rect 4584 22708 4632 22764
rect 4688 22708 4736 22764
rect 4792 22708 4840 22764
rect 4896 22708 4944 22764
rect 5000 22708 5048 22764
rect 5104 22708 5152 22764
rect 5208 22708 5228 22764
rect 3988 21196 5228 22708
rect 3988 21140 4008 21196
rect 4064 21140 4112 21196
rect 4168 21140 4216 21196
rect 4272 21140 4320 21196
rect 4376 21140 4424 21196
rect 4480 21140 4528 21196
rect 4584 21140 4632 21196
rect 4688 21140 4736 21196
rect 4792 21140 4840 21196
rect 4896 21140 4944 21196
rect 5000 21140 5048 21196
rect 5104 21140 5152 21196
rect 5208 21140 5228 21196
rect 3988 19628 5228 21140
rect 5292 22932 5348 22942
rect 5292 21028 5348 22876
rect 13692 22932 13748 23436
rect 13804 23156 13860 23772
rect 13804 23090 13860 23100
rect 13988 23548 15228 25060
rect 13988 23492 14008 23548
rect 14064 23492 14112 23548
rect 14168 23492 14216 23548
rect 14272 23492 14320 23548
rect 14376 23492 14424 23548
rect 14480 23492 14528 23548
rect 14584 23492 14632 23548
rect 14688 23492 14736 23548
rect 14792 23492 14840 23548
rect 14896 23492 14944 23548
rect 15000 23492 15048 23548
rect 15104 23492 15152 23548
rect 15208 23492 15228 23548
rect 13692 22866 13748 22876
rect 13804 22708 13860 22718
rect 13692 22596 13748 22606
rect 13692 22260 13748 22540
rect 6188 21812 6244 21822
rect 5292 20962 5348 20972
rect 5404 21476 5460 21486
rect 3988 19572 4008 19628
rect 4064 19572 4112 19628
rect 4168 19572 4216 19628
rect 4272 19572 4320 19628
rect 4376 19572 4424 19628
rect 4480 19572 4528 19628
rect 4584 19572 4632 19628
rect 4688 19572 4736 19628
rect 4792 19572 4840 19628
rect 4896 19572 4944 19628
rect 5000 19572 5048 19628
rect 5104 19572 5152 19628
rect 5208 19572 5228 19628
rect 3988 18060 5228 19572
rect 3988 18004 4008 18060
rect 4064 18004 4112 18060
rect 4168 18004 4216 18060
rect 4272 18004 4320 18060
rect 4376 18004 4424 18060
rect 4480 18004 4528 18060
rect 4584 18004 4632 18060
rect 4688 18004 4736 18060
rect 4792 18004 4840 18060
rect 4896 18004 4944 18060
rect 5000 18004 5048 18060
rect 5104 18004 5152 18060
rect 5208 18004 5228 18060
rect 3988 16492 5228 18004
rect 3988 16436 4008 16492
rect 4064 16436 4112 16492
rect 4168 16436 4216 16492
rect 4272 16436 4320 16492
rect 4376 16436 4424 16492
rect 4480 16436 4528 16492
rect 4584 16436 4632 16492
rect 4688 16436 4736 16492
rect 4792 16436 4840 16492
rect 4896 16436 4944 16492
rect 5000 16436 5048 16492
rect 5104 16436 5152 16492
rect 5208 16436 5228 16492
rect 3988 14924 5228 16436
rect 3988 14868 4008 14924
rect 4064 14868 4112 14924
rect 4168 14868 4216 14924
rect 4272 14868 4320 14924
rect 4376 14868 4424 14924
rect 4480 14868 4528 14924
rect 4584 14868 4632 14924
rect 4688 14868 4736 14924
rect 4792 14868 4840 14924
rect 4896 14868 4944 14924
rect 5000 14868 5048 14924
rect 5104 14868 5152 14924
rect 5208 14868 5228 14924
rect 3988 13356 5228 14868
rect 3988 13300 4008 13356
rect 4064 13300 4112 13356
rect 4168 13300 4216 13356
rect 4272 13300 4320 13356
rect 4376 13300 4424 13356
rect 4480 13300 4528 13356
rect 4584 13300 4632 13356
rect 4688 13300 4736 13356
rect 4792 13300 4840 13356
rect 4896 13300 4944 13356
rect 5000 13300 5048 13356
rect 5104 13300 5152 13356
rect 5208 13300 5228 13356
rect 3988 11788 5228 13300
rect 3988 11732 4008 11788
rect 4064 11732 4112 11788
rect 4168 11732 4216 11788
rect 4272 11732 4320 11788
rect 4376 11732 4424 11788
rect 4480 11732 4528 11788
rect 4584 11732 4632 11788
rect 4688 11732 4736 11788
rect 4792 11732 4840 11788
rect 4896 11732 4944 11788
rect 5000 11732 5048 11788
rect 5104 11732 5152 11788
rect 5208 11732 5228 11788
rect 3988 10220 5228 11732
rect 5404 16212 5460 21420
rect 5404 13076 5460 16156
rect 6188 20244 6244 21756
rect 6188 15652 6244 20188
rect 13692 21028 13748 22204
rect 13468 20020 13524 20030
rect 13356 19124 13412 19134
rect 13356 16436 13412 19068
rect 13356 16370 13412 16380
rect 6188 14308 6244 15596
rect 6188 14242 6244 14252
rect 13468 16324 13524 19964
rect 13468 15204 13524 16268
rect 13468 13972 13524 15148
rect 13468 13906 13524 13916
rect 5404 11508 5460 13020
rect 13692 12852 13748 20972
rect 13804 20580 13860 22652
rect 13804 17556 13860 20524
rect 13804 17490 13860 17500
rect 13988 21980 15228 23492
rect 13988 21924 14008 21980
rect 14064 21924 14112 21980
rect 14168 21924 14216 21980
rect 14272 21924 14320 21980
rect 14376 21924 14424 21980
rect 14480 21924 14528 21980
rect 14584 21924 14632 21980
rect 14688 21924 14736 21980
rect 14792 21924 14840 21980
rect 14896 21924 14944 21980
rect 15000 21924 15048 21980
rect 15104 21924 15152 21980
rect 15208 21924 15228 21980
rect 13988 20412 15228 21924
rect 13988 20356 14008 20412
rect 14064 20356 14112 20412
rect 14168 20356 14216 20412
rect 14272 20356 14320 20412
rect 14376 20356 14424 20412
rect 14480 20356 14528 20412
rect 14584 20356 14632 20412
rect 14688 20356 14736 20412
rect 14792 20356 14840 20412
rect 14896 20356 14944 20412
rect 15000 20356 15048 20412
rect 15104 20356 15152 20412
rect 15208 20356 15228 20412
rect 13988 18844 15228 20356
rect 13988 18788 14008 18844
rect 14064 18788 14112 18844
rect 14168 18788 14216 18844
rect 14272 18788 14320 18844
rect 14376 18788 14424 18844
rect 14480 18788 14528 18844
rect 14584 18788 14632 18844
rect 14688 18788 14736 18844
rect 14792 18788 14840 18844
rect 14896 18788 14944 18844
rect 15000 18788 15048 18844
rect 15104 18788 15152 18844
rect 15208 18788 15228 18844
rect 13692 12786 13748 12796
rect 13988 17276 15228 18788
rect 13988 17220 14008 17276
rect 14064 17220 14112 17276
rect 14168 17220 14216 17276
rect 14272 17220 14320 17276
rect 14376 17220 14424 17276
rect 14480 17220 14528 17276
rect 14584 17220 14632 17276
rect 14688 17220 14736 17276
rect 14792 17220 14840 17276
rect 14896 17220 14944 17276
rect 15000 17220 15048 17276
rect 15104 17220 15152 17276
rect 15208 17220 15228 17276
rect 13988 15708 15228 17220
rect 15372 31668 15428 31678
rect 15372 17108 15428 31612
rect 15484 29652 15540 32732
rect 15484 29586 15540 29596
rect 23988 32172 25228 33684
rect 27020 37380 27076 37390
rect 27020 33012 27076 37324
rect 33628 34916 33684 34926
rect 33628 34244 33684 34860
rect 33628 34178 33684 34188
rect 27020 32946 27076 32956
rect 33740 33012 33796 38612
rect 33852 38500 33908 38510
rect 33852 34692 33908 38444
rect 33852 34626 33908 34636
rect 33988 37660 35228 39172
rect 33988 37604 34008 37660
rect 34064 37604 34112 37660
rect 34168 37604 34216 37660
rect 34272 37604 34320 37660
rect 34376 37604 34424 37660
rect 34480 37604 34528 37660
rect 34584 37604 34632 37660
rect 34688 37604 34736 37660
rect 34792 37604 34840 37660
rect 34896 37604 34944 37660
rect 35000 37604 35048 37660
rect 35104 37604 35152 37660
rect 35208 37604 35228 37660
rect 33988 36092 35228 37604
rect 33988 36036 34008 36092
rect 34064 36036 34112 36092
rect 34168 36036 34216 36092
rect 34272 36036 34320 36092
rect 34376 36036 34424 36092
rect 34480 36036 34528 36092
rect 34584 36036 34632 36092
rect 34688 36036 34736 36092
rect 34792 36036 34840 36092
rect 34896 36036 34944 36092
rect 35000 36036 35048 36092
rect 35104 36036 35152 36092
rect 35208 36036 35228 36092
rect 33740 32946 33796 32956
rect 33988 34524 35228 36036
rect 33988 34468 34008 34524
rect 34064 34468 34112 34524
rect 34168 34468 34216 34524
rect 34272 34468 34320 34524
rect 34376 34468 34424 34524
rect 34480 34468 34528 34524
rect 34584 34468 34632 34524
rect 34688 34468 34736 34524
rect 34792 34468 34840 34524
rect 34896 34468 34944 34524
rect 35000 34468 35048 34524
rect 35104 34468 35152 34524
rect 35208 34468 35228 34524
rect 33988 32956 35228 34468
rect 23988 32116 24008 32172
rect 24064 32116 24112 32172
rect 24168 32116 24216 32172
rect 24272 32116 24320 32172
rect 24376 32116 24424 32172
rect 24480 32116 24528 32172
rect 24584 32116 24632 32172
rect 24688 32116 24736 32172
rect 24792 32116 24840 32172
rect 24896 32116 24944 32172
rect 25000 32116 25048 32172
rect 25104 32116 25152 32172
rect 25208 32116 25228 32172
rect 23988 30604 25228 32116
rect 33988 32900 34008 32956
rect 34064 32900 34112 32956
rect 34168 32900 34216 32956
rect 34272 32900 34320 32956
rect 34376 32900 34424 32956
rect 34480 32900 34528 32956
rect 34584 32900 34632 32956
rect 34688 32900 34736 32956
rect 34792 32900 34840 32956
rect 34896 32900 34944 32956
rect 35000 32900 35048 32956
rect 35104 32900 35152 32956
rect 35208 32900 35228 32956
rect 23988 30548 24008 30604
rect 24064 30548 24112 30604
rect 24168 30548 24216 30604
rect 24272 30548 24320 30604
rect 24376 30548 24424 30604
rect 24480 30548 24528 30604
rect 24584 30548 24632 30604
rect 24688 30548 24736 30604
rect 24792 30548 24840 30604
rect 24896 30548 24944 30604
rect 25000 30548 25048 30604
rect 25104 30548 25152 30604
rect 25208 30548 25228 30604
rect 15372 17042 15428 17052
rect 23988 29036 25228 30548
rect 23988 28980 24008 29036
rect 24064 28980 24112 29036
rect 24168 28980 24216 29036
rect 24272 28980 24320 29036
rect 24376 28980 24424 29036
rect 24480 28980 24528 29036
rect 24584 28980 24632 29036
rect 24688 28980 24736 29036
rect 24792 28980 24840 29036
rect 24896 28980 24944 29036
rect 25000 28980 25048 29036
rect 25104 28980 25152 29036
rect 25208 28980 25228 29036
rect 23988 27468 25228 28980
rect 23988 27412 24008 27468
rect 24064 27412 24112 27468
rect 24168 27412 24216 27468
rect 24272 27412 24320 27468
rect 24376 27412 24424 27468
rect 24480 27412 24528 27468
rect 24584 27412 24632 27468
rect 24688 27412 24736 27468
rect 24792 27412 24840 27468
rect 24896 27412 24944 27468
rect 25000 27412 25048 27468
rect 25104 27412 25152 27468
rect 25208 27412 25228 27468
rect 23988 25900 25228 27412
rect 23988 25844 24008 25900
rect 24064 25844 24112 25900
rect 24168 25844 24216 25900
rect 24272 25844 24320 25900
rect 24376 25844 24424 25900
rect 24480 25844 24528 25900
rect 24584 25844 24632 25900
rect 24688 25844 24736 25900
rect 24792 25844 24840 25900
rect 24896 25844 24944 25900
rect 25000 25844 25048 25900
rect 25104 25844 25152 25900
rect 25208 25844 25228 25900
rect 23988 24332 25228 25844
rect 26572 31556 26628 31566
rect 26572 25172 26628 31500
rect 26572 25106 26628 25116
rect 33988 31388 35228 32900
rect 33988 31332 34008 31388
rect 34064 31332 34112 31388
rect 34168 31332 34216 31388
rect 34272 31332 34320 31388
rect 34376 31332 34424 31388
rect 34480 31332 34528 31388
rect 34584 31332 34632 31388
rect 34688 31332 34736 31388
rect 34792 31332 34840 31388
rect 34896 31332 34944 31388
rect 35000 31332 35048 31388
rect 35104 31332 35152 31388
rect 35208 31332 35228 31388
rect 33988 29820 35228 31332
rect 33988 29764 34008 29820
rect 34064 29764 34112 29820
rect 34168 29764 34216 29820
rect 34272 29764 34320 29820
rect 34376 29764 34424 29820
rect 34480 29764 34528 29820
rect 34584 29764 34632 29820
rect 34688 29764 34736 29820
rect 34792 29764 34840 29820
rect 34896 29764 34944 29820
rect 35000 29764 35048 29820
rect 35104 29764 35152 29820
rect 35208 29764 35228 29820
rect 33988 28252 35228 29764
rect 33988 28196 34008 28252
rect 34064 28196 34112 28252
rect 34168 28196 34216 28252
rect 34272 28196 34320 28252
rect 34376 28196 34424 28252
rect 34480 28196 34528 28252
rect 34584 28196 34632 28252
rect 34688 28196 34736 28252
rect 34792 28196 34840 28252
rect 34896 28196 34944 28252
rect 35000 28196 35048 28252
rect 35104 28196 35152 28252
rect 35208 28196 35228 28252
rect 33988 26684 35228 28196
rect 33988 26628 34008 26684
rect 34064 26628 34112 26684
rect 34168 26628 34216 26684
rect 34272 26628 34320 26684
rect 34376 26628 34424 26684
rect 34480 26628 34528 26684
rect 34584 26628 34632 26684
rect 34688 26628 34736 26684
rect 34792 26628 34840 26684
rect 34896 26628 34944 26684
rect 35000 26628 35048 26684
rect 35104 26628 35152 26684
rect 35208 26628 35228 26684
rect 33988 25116 35228 26628
rect 23988 24276 24008 24332
rect 24064 24276 24112 24332
rect 24168 24276 24216 24332
rect 24272 24276 24320 24332
rect 24376 24276 24424 24332
rect 24480 24276 24528 24332
rect 24584 24276 24632 24332
rect 24688 24276 24736 24332
rect 24792 24276 24840 24332
rect 24896 24276 24944 24332
rect 25000 24276 25048 24332
rect 25104 24276 25152 24332
rect 25208 24276 25228 24332
rect 23988 22764 25228 24276
rect 23988 22708 24008 22764
rect 24064 22708 24112 22764
rect 24168 22708 24216 22764
rect 24272 22708 24320 22764
rect 24376 22708 24424 22764
rect 24480 22708 24528 22764
rect 24584 22708 24632 22764
rect 24688 22708 24736 22764
rect 24792 22708 24840 22764
rect 24896 22708 24944 22764
rect 25000 22708 25048 22764
rect 25104 22708 25152 22764
rect 25208 22708 25228 22764
rect 23988 21196 25228 22708
rect 33988 25060 34008 25116
rect 34064 25060 34112 25116
rect 34168 25060 34216 25116
rect 34272 25060 34320 25116
rect 34376 25060 34424 25116
rect 34480 25060 34528 25116
rect 34584 25060 34632 25116
rect 34688 25060 34736 25116
rect 34792 25060 34840 25116
rect 34896 25060 34944 25116
rect 35000 25060 35048 25116
rect 35104 25060 35152 25116
rect 35208 25060 35228 25116
rect 33988 23548 35228 25060
rect 33988 23492 34008 23548
rect 34064 23492 34112 23548
rect 34168 23492 34216 23548
rect 34272 23492 34320 23548
rect 34376 23492 34424 23548
rect 34480 23492 34528 23548
rect 34584 23492 34632 23548
rect 34688 23492 34736 23548
rect 34792 23492 34840 23548
rect 34896 23492 34944 23548
rect 35000 23492 35048 23548
rect 35104 23492 35152 23548
rect 35208 23492 35228 23548
rect 23988 21140 24008 21196
rect 24064 21140 24112 21196
rect 24168 21140 24216 21196
rect 24272 21140 24320 21196
rect 24376 21140 24424 21196
rect 24480 21140 24528 21196
rect 24584 21140 24632 21196
rect 24688 21140 24736 21196
rect 24792 21140 24840 21196
rect 24896 21140 24944 21196
rect 25000 21140 25048 21196
rect 25104 21140 25152 21196
rect 25208 21140 25228 21196
rect 23988 19628 25228 21140
rect 25340 22260 25396 22270
rect 25340 20692 25396 22204
rect 33988 21980 35228 23492
rect 33988 21924 34008 21980
rect 34064 21924 34112 21980
rect 34168 21924 34216 21980
rect 34272 21924 34320 21980
rect 34376 21924 34424 21980
rect 34480 21924 34528 21980
rect 34584 21924 34632 21980
rect 34688 21924 34736 21980
rect 34792 21924 34840 21980
rect 34896 21924 34944 21980
rect 35000 21924 35048 21980
rect 35104 21924 35152 21980
rect 35208 21924 35228 21980
rect 25340 20626 25396 20636
rect 26236 20916 26292 20926
rect 23988 19572 24008 19628
rect 24064 19572 24112 19628
rect 24168 19572 24216 19628
rect 24272 19572 24320 19628
rect 24376 19572 24424 19628
rect 24480 19572 24528 19628
rect 24584 19572 24632 19628
rect 24688 19572 24736 19628
rect 24792 19572 24840 19628
rect 24896 19572 24944 19628
rect 25000 19572 25048 19628
rect 25104 19572 25152 19628
rect 25208 19572 25228 19628
rect 23988 18060 25228 19572
rect 25340 20244 25396 20254
rect 25340 19236 25396 20188
rect 25340 19170 25396 19180
rect 23988 18004 24008 18060
rect 24064 18004 24112 18060
rect 24168 18004 24216 18060
rect 24272 18004 24320 18060
rect 24376 18004 24424 18060
rect 24480 18004 24528 18060
rect 24584 18004 24632 18060
rect 24688 18004 24736 18060
rect 24792 18004 24840 18060
rect 24896 18004 24944 18060
rect 25000 18004 25048 18060
rect 25104 18004 25152 18060
rect 25208 18004 25228 18060
rect 23772 16660 23828 16670
rect 23772 16212 23828 16604
rect 23772 16146 23828 16156
rect 23988 16492 25228 18004
rect 26236 17556 26292 20860
rect 26236 17490 26292 17500
rect 33988 20412 35228 21924
rect 33988 20356 34008 20412
rect 34064 20356 34112 20412
rect 34168 20356 34216 20412
rect 34272 20356 34320 20412
rect 34376 20356 34424 20412
rect 34480 20356 34528 20412
rect 34584 20356 34632 20412
rect 34688 20356 34736 20412
rect 34792 20356 34840 20412
rect 34896 20356 34944 20412
rect 35000 20356 35048 20412
rect 35104 20356 35152 20412
rect 35208 20356 35228 20412
rect 33988 18844 35228 20356
rect 33988 18788 34008 18844
rect 34064 18788 34112 18844
rect 34168 18788 34216 18844
rect 34272 18788 34320 18844
rect 34376 18788 34424 18844
rect 34480 18788 34528 18844
rect 34584 18788 34632 18844
rect 34688 18788 34736 18844
rect 34792 18788 34840 18844
rect 34896 18788 34944 18844
rect 35000 18788 35048 18844
rect 35104 18788 35152 18844
rect 35208 18788 35228 18844
rect 23988 16436 24008 16492
rect 24064 16436 24112 16492
rect 24168 16436 24216 16492
rect 24272 16436 24320 16492
rect 24376 16436 24424 16492
rect 24480 16436 24528 16492
rect 24584 16436 24632 16492
rect 24688 16436 24736 16492
rect 24792 16436 24840 16492
rect 24896 16436 24944 16492
rect 25000 16436 25048 16492
rect 25104 16436 25152 16492
rect 25208 16436 25228 16492
rect 13988 15652 14008 15708
rect 14064 15652 14112 15708
rect 14168 15652 14216 15708
rect 14272 15652 14320 15708
rect 14376 15652 14424 15708
rect 14480 15652 14528 15708
rect 14584 15652 14632 15708
rect 14688 15652 14736 15708
rect 14792 15652 14840 15708
rect 14896 15652 14944 15708
rect 15000 15652 15048 15708
rect 15104 15652 15152 15708
rect 15208 15652 15228 15708
rect 13988 14140 15228 15652
rect 13988 14084 14008 14140
rect 14064 14084 14112 14140
rect 14168 14084 14216 14140
rect 14272 14084 14320 14140
rect 14376 14084 14424 14140
rect 14480 14084 14528 14140
rect 14584 14084 14632 14140
rect 14688 14084 14736 14140
rect 14792 14084 14840 14140
rect 14896 14084 14944 14140
rect 15000 14084 15048 14140
rect 15104 14084 15152 14140
rect 15208 14084 15228 14140
rect 5404 11442 5460 11452
rect 13988 12572 15228 14084
rect 13988 12516 14008 12572
rect 14064 12516 14112 12572
rect 14168 12516 14216 12572
rect 14272 12516 14320 12572
rect 14376 12516 14424 12572
rect 14480 12516 14528 12572
rect 14584 12516 14632 12572
rect 14688 12516 14736 12572
rect 14792 12516 14840 12572
rect 14896 12516 14944 12572
rect 15000 12516 15048 12572
rect 15104 12516 15152 12572
rect 15208 12516 15228 12572
rect 3988 10164 4008 10220
rect 4064 10164 4112 10220
rect 4168 10164 4216 10220
rect 4272 10164 4320 10220
rect 4376 10164 4424 10220
rect 4480 10164 4528 10220
rect 4584 10164 4632 10220
rect 4688 10164 4736 10220
rect 4792 10164 4840 10220
rect 4896 10164 4944 10220
rect 5000 10164 5048 10220
rect 5104 10164 5152 10220
rect 5208 10164 5228 10220
rect 3988 8652 5228 10164
rect 3988 8596 4008 8652
rect 4064 8596 4112 8652
rect 4168 8596 4216 8652
rect 4272 8596 4320 8652
rect 4376 8596 4424 8652
rect 4480 8596 4528 8652
rect 4584 8596 4632 8652
rect 4688 8596 4736 8652
rect 4792 8596 4840 8652
rect 4896 8596 4944 8652
rect 5000 8596 5048 8652
rect 5104 8596 5152 8652
rect 5208 8596 5228 8652
rect 3988 7084 5228 8596
rect 3988 7028 4008 7084
rect 4064 7028 4112 7084
rect 4168 7028 4216 7084
rect 4272 7028 4320 7084
rect 4376 7028 4424 7084
rect 4480 7028 4528 7084
rect 4584 7028 4632 7084
rect 4688 7028 4736 7084
rect 4792 7028 4840 7084
rect 4896 7028 4944 7084
rect 5000 7028 5048 7084
rect 5104 7028 5152 7084
rect 5208 7028 5228 7084
rect 3988 5516 5228 7028
rect 3988 5460 4008 5516
rect 4064 5460 4112 5516
rect 4168 5460 4216 5516
rect 4272 5460 4320 5516
rect 4376 5460 4424 5516
rect 4480 5460 4528 5516
rect 4584 5460 4632 5516
rect 4688 5460 4736 5516
rect 4792 5460 4840 5516
rect 4896 5460 4944 5516
rect 5000 5460 5048 5516
rect 5104 5460 5152 5516
rect 5208 5460 5228 5516
rect 3988 3948 5228 5460
rect 3988 3892 4008 3948
rect 4064 3892 4112 3948
rect 4168 3892 4216 3948
rect 4272 3892 4320 3948
rect 4376 3892 4424 3948
rect 4480 3892 4528 3948
rect 4584 3892 4632 3948
rect 4688 3892 4736 3948
rect 4792 3892 4840 3948
rect 4896 3892 4944 3948
rect 5000 3892 5048 3948
rect 5104 3892 5152 3948
rect 5208 3892 5228 3948
rect 3988 3076 5228 3892
rect 13988 11004 15228 12516
rect 13988 10948 14008 11004
rect 14064 10948 14112 11004
rect 14168 10948 14216 11004
rect 14272 10948 14320 11004
rect 14376 10948 14424 11004
rect 14480 10948 14528 11004
rect 14584 10948 14632 11004
rect 14688 10948 14736 11004
rect 14792 10948 14840 11004
rect 14896 10948 14944 11004
rect 15000 10948 15048 11004
rect 15104 10948 15152 11004
rect 15208 10948 15228 11004
rect 13988 9436 15228 10948
rect 13988 9380 14008 9436
rect 14064 9380 14112 9436
rect 14168 9380 14216 9436
rect 14272 9380 14320 9436
rect 14376 9380 14424 9436
rect 14480 9380 14528 9436
rect 14584 9380 14632 9436
rect 14688 9380 14736 9436
rect 14792 9380 14840 9436
rect 14896 9380 14944 9436
rect 15000 9380 15048 9436
rect 15104 9380 15152 9436
rect 15208 9380 15228 9436
rect 13988 7868 15228 9380
rect 13988 7812 14008 7868
rect 14064 7812 14112 7868
rect 14168 7812 14216 7868
rect 14272 7812 14320 7868
rect 14376 7812 14424 7868
rect 14480 7812 14528 7868
rect 14584 7812 14632 7868
rect 14688 7812 14736 7868
rect 14792 7812 14840 7868
rect 14896 7812 14944 7868
rect 15000 7812 15048 7868
rect 15104 7812 15152 7868
rect 15208 7812 15228 7868
rect 13988 6300 15228 7812
rect 13988 6244 14008 6300
rect 14064 6244 14112 6300
rect 14168 6244 14216 6300
rect 14272 6244 14320 6300
rect 14376 6244 14424 6300
rect 14480 6244 14528 6300
rect 14584 6244 14632 6300
rect 14688 6244 14736 6300
rect 14792 6244 14840 6300
rect 14896 6244 14944 6300
rect 15000 6244 15048 6300
rect 15104 6244 15152 6300
rect 15208 6244 15228 6300
rect 13988 4732 15228 6244
rect 13988 4676 14008 4732
rect 14064 4676 14112 4732
rect 14168 4676 14216 4732
rect 14272 4676 14320 4732
rect 14376 4676 14424 4732
rect 14480 4676 14528 4732
rect 14584 4676 14632 4732
rect 14688 4676 14736 4732
rect 14792 4676 14840 4732
rect 14896 4676 14944 4732
rect 15000 4676 15048 4732
rect 15104 4676 15152 4732
rect 15208 4676 15228 4732
rect 13988 3164 15228 4676
rect 13988 3108 14008 3164
rect 14064 3108 14112 3164
rect 14168 3108 14216 3164
rect 14272 3108 14320 3164
rect 14376 3108 14424 3164
rect 14480 3108 14528 3164
rect 14584 3108 14632 3164
rect 14688 3108 14736 3164
rect 14792 3108 14840 3164
rect 14896 3108 14944 3164
rect 15000 3108 15048 3164
rect 15104 3108 15152 3164
rect 15208 3108 15228 3164
rect 13988 3076 15228 3108
rect 23988 14924 25228 16436
rect 25340 17332 25396 17342
rect 25340 15876 25396 17276
rect 25340 15810 25396 15820
rect 33988 17276 35228 18788
rect 33988 17220 34008 17276
rect 34064 17220 34112 17276
rect 34168 17220 34216 17276
rect 34272 17220 34320 17276
rect 34376 17220 34424 17276
rect 34480 17220 34528 17276
rect 34584 17220 34632 17276
rect 34688 17220 34736 17276
rect 34792 17220 34840 17276
rect 34896 17220 34944 17276
rect 35000 17220 35048 17276
rect 35104 17220 35152 17276
rect 35208 17220 35228 17276
rect 23988 14868 24008 14924
rect 24064 14868 24112 14924
rect 24168 14868 24216 14924
rect 24272 14868 24320 14924
rect 24376 14868 24424 14924
rect 24480 14868 24528 14924
rect 24584 14868 24632 14924
rect 24688 14868 24736 14924
rect 24792 14868 24840 14924
rect 24896 14868 24944 14924
rect 25000 14868 25048 14924
rect 25104 14868 25152 14924
rect 25208 14868 25228 14924
rect 23988 13356 25228 14868
rect 23988 13300 24008 13356
rect 24064 13300 24112 13356
rect 24168 13300 24216 13356
rect 24272 13300 24320 13356
rect 24376 13300 24424 13356
rect 24480 13300 24528 13356
rect 24584 13300 24632 13356
rect 24688 13300 24736 13356
rect 24792 13300 24840 13356
rect 24896 13300 24944 13356
rect 25000 13300 25048 13356
rect 25104 13300 25152 13356
rect 25208 13300 25228 13356
rect 23988 11788 25228 13300
rect 23988 11732 24008 11788
rect 24064 11732 24112 11788
rect 24168 11732 24216 11788
rect 24272 11732 24320 11788
rect 24376 11732 24424 11788
rect 24480 11732 24528 11788
rect 24584 11732 24632 11788
rect 24688 11732 24736 11788
rect 24792 11732 24840 11788
rect 24896 11732 24944 11788
rect 25000 11732 25048 11788
rect 25104 11732 25152 11788
rect 25208 11732 25228 11788
rect 23988 10220 25228 11732
rect 23988 10164 24008 10220
rect 24064 10164 24112 10220
rect 24168 10164 24216 10220
rect 24272 10164 24320 10220
rect 24376 10164 24424 10220
rect 24480 10164 24528 10220
rect 24584 10164 24632 10220
rect 24688 10164 24736 10220
rect 24792 10164 24840 10220
rect 24896 10164 24944 10220
rect 25000 10164 25048 10220
rect 25104 10164 25152 10220
rect 25208 10164 25228 10220
rect 23988 8652 25228 10164
rect 23988 8596 24008 8652
rect 24064 8596 24112 8652
rect 24168 8596 24216 8652
rect 24272 8596 24320 8652
rect 24376 8596 24424 8652
rect 24480 8596 24528 8652
rect 24584 8596 24632 8652
rect 24688 8596 24736 8652
rect 24792 8596 24840 8652
rect 24896 8596 24944 8652
rect 25000 8596 25048 8652
rect 25104 8596 25152 8652
rect 25208 8596 25228 8652
rect 23988 7084 25228 8596
rect 23988 7028 24008 7084
rect 24064 7028 24112 7084
rect 24168 7028 24216 7084
rect 24272 7028 24320 7084
rect 24376 7028 24424 7084
rect 24480 7028 24528 7084
rect 24584 7028 24632 7084
rect 24688 7028 24736 7084
rect 24792 7028 24840 7084
rect 24896 7028 24944 7084
rect 25000 7028 25048 7084
rect 25104 7028 25152 7084
rect 25208 7028 25228 7084
rect 23988 5516 25228 7028
rect 23988 5460 24008 5516
rect 24064 5460 24112 5516
rect 24168 5460 24216 5516
rect 24272 5460 24320 5516
rect 24376 5460 24424 5516
rect 24480 5460 24528 5516
rect 24584 5460 24632 5516
rect 24688 5460 24736 5516
rect 24792 5460 24840 5516
rect 24896 5460 24944 5516
rect 25000 5460 25048 5516
rect 25104 5460 25152 5516
rect 25208 5460 25228 5516
rect 23988 3948 25228 5460
rect 23988 3892 24008 3948
rect 24064 3892 24112 3948
rect 24168 3892 24216 3948
rect 24272 3892 24320 3948
rect 24376 3892 24424 3948
rect 24480 3892 24528 3948
rect 24584 3892 24632 3948
rect 24688 3892 24736 3948
rect 24792 3892 24840 3948
rect 24896 3892 24944 3948
rect 25000 3892 25048 3948
rect 25104 3892 25152 3948
rect 25208 3892 25228 3948
rect 23988 3076 25228 3892
rect 33988 15708 35228 17220
rect 33988 15652 34008 15708
rect 34064 15652 34112 15708
rect 34168 15652 34216 15708
rect 34272 15652 34320 15708
rect 34376 15652 34424 15708
rect 34480 15652 34528 15708
rect 34584 15652 34632 15708
rect 34688 15652 34736 15708
rect 34792 15652 34840 15708
rect 34896 15652 34944 15708
rect 35000 15652 35048 15708
rect 35104 15652 35152 15708
rect 35208 15652 35228 15708
rect 33988 14140 35228 15652
rect 33988 14084 34008 14140
rect 34064 14084 34112 14140
rect 34168 14084 34216 14140
rect 34272 14084 34320 14140
rect 34376 14084 34424 14140
rect 34480 14084 34528 14140
rect 34584 14084 34632 14140
rect 34688 14084 34736 14140
rect 34792 14084 34840 14140
rect 34896 14084 34944 14140
rect 35000 14084 35048 14140
rect 35104 14084 35152 14140
rect 35208 14084 35228 14140
rect 33988 12572 35228 14084
rect 33988 12516 34008 12572
rect 34064 12516 34112 12572
rect 34168 12516 34216 12572
rect 34272 12516 34320 12572
rect 34376 12516 34424 12572
rect 34480 12516 34528 12572
rect 34584 12516 34632 12572
rect 34688 12516 34736 12572
rect 34792 12516 34840 12572
rect 34896 12516 34944 12572
rect 35000 12516 35048 12572
rect 35104 12516 35152 12572
rect 35208 12516 35228 12572
rect 33988 11004 35228 12516
rect 33988 10948 34008 11004
rect 34064 10948 34112 11004
rect 34168 10948 34216 11004
rect 34272 10948 34320 11004
rect 34376 10948 34424 11004
rect 34480 10948 34528 11004
rect 34584 10948 34632 11004
rect 34688 10948 34736 11004
rect 34792 10948 34840 11004
rect 34896 10948 34944 11004
rect 35000 10948 35048 11004
rect 35104 10948 35152 11004
rect 35208 10948 35228 11004
rect 33988 9436 35228 10948
rect 33988 9380 34008 9436
rect 34064 9380 34112 9436
rect 34168 9380 34216 9436
rect 34272 9380 34320 9436
rect 34376 9380 34424 9436
rect 34480 9380 34528 9436
rect 34584 9380 34632 9436
rect 34688 9380 34736 9436
rect 34792 9380 34840 9436
rect 34896 9380 34944 9436
rect 35000 9380 35048 9436
rect 35104 9380 35152 9436
rect 35208 9380 35228 9436
rect 33988 7868 35228 9380
rect 33988 7812 34008 7868
rect 34064 7812 34112 7868
rect 34168 7812 34216 7868
rect 34272 7812 34320 7868
rect 34376 7812 34424 7868
rect 34480 7812 34528 7868
rect 34584 7812 34632 7868
rect 34688 7812 34736 7868
rect 34792 7812 34840 7868
rect 34896 7812 34944 7868
rect 35000 7812 35048 7868
rect 35104 7812 35152 7868
rect 35208 7812 35228 7868
rect 33988 6300 35228 7812
rect 33988 6244 34008 6300
rect 34064 6244 34112 6300
rect 34168 6244 34216 6300
rect 34272 6244 34320 6300
rect 34376 6244 34424 6300
rect 34480 6244 34528 6300
rect 34584 6244 34632 6300
rect 34688 6244 34736 6300
rect 34792 6244 34840 6300
rect 34896 6244 34944 6300
rect 35000 6244 35048 6300
rect 35104 6244 35152 6300
rect 35208 6244 35228 6300
rect 33988 4732 35228 6244
rect 33988 4676 34008 4732
rect 34064 4676 34112 4732
rect 34168 4676 34216 4732
rect 34272 4676 34320 4732
rect 34376 4676 34424 4732
rect 34480 4676 34528 4732
rect 34584 4676 34632 4732
rect 34688 4676 34736 4732
rect 34792 4676 34840 4732
rect 34896 4676 34944 4732
rect 35000 4676 35048 4732
rect 35104 4676 35152 4732
rect 35208 4676 35228 4732
rect 33988 3164 35228 4676
rect 33988 3108 34008 3164
rect 34064 3108 34112 3164
rect 34168 3108 34216 3164
rect 34272 3108 34320 3164
rect 34376 3108 34424 3164
rect 34480 3108 34528 3164
rect 34584 3108 34632 3164
rect 34688 3108 34736 3164
rect 34792 3108 34840 3164
rect 34896 3108 34944 3164
rect 35000 3108 35048 3164
rect 35104 3108 35152 3164
rect 35208 3108 35228 3164
rect 33988 3076 35228 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_mclk_I open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_rtc_clk_I
timestamp 1698431365
transform 1 0 18928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_rtc_clk_I
timestamp 1698431365
transform -1 0 11312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_rtc_clk_I
timestamp 1698431365
transform -1 0 14784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_rtc_clk_I
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_rtc_clk_I
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_rtc_clk_I
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_rtc_clk_I
timestamp 1698431365
transform 1 0 24080 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_rtc_clk_I
timestamp 1698431365
transform 1 0 24080 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_rtc_clk_I
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_rtc_clk_I
timestamp 1698431365
transform 1 0 9968 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_rtc_clk_I
timestamp 1698431365
transform 1 0 13552 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_rtc_clk_I
timestamp 1698431365
transform 1 0 9744 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_rtc_clk_I
timestamp 1698431365
transform -1 0 16464 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_rtc_clk_I
timestamp 1698431365
transform 1 0 23408 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_rtc_clk_I
timestamp 1698431365
transform 1 0 26656 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_rtc_clk_I
timestamp 1698431365
transform 1 0 24192 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_rtc_clk_I
timestamp 1698431365
transform 1 0 27440 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout2_I
timestamp 1698431365
transform 1 0 8512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout4_I
timestamp 1698431365
transform 1 0 9296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout5_I
timestamp 1698431365
transform 1 0 8960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout6_I
timestamp 1698431365
transform 1 0 22400 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout7_I
timestamp 1698431365
transform 1 0 28224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout8_I
timestamp 1698431365
transform 1 0 21280 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout9_I
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout10_I
timestamp 1698431365
transform 1 0 26656 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout11_I
timestamp 1698431365
transform 1 0 29568 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout12_I
timestamp 1698431365
transform 1 0 17584 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout13_I
timestamp 1698431365
transform 1 0 24304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout14_I
timestamp 1698431365
transform 1 0 27104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout16_I
timestamp 1698431365
transform -1 0 29456 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout17_I
timestamp 1698431365
transform 1 0 13328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout18_I
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout19_I
timestamp 1698431365
transform 1 0 5600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout20_I
timestamp 1698431365
transform 1 0 8512 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_hold7_I
timestamp 1698431365
transform 1 0 13216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output1_I
timestamp 1698431365
transform -1 0 29904 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rst_sync.u_buf.genblk1.u_mux_I1
timestamp 1698431365
transform -1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._102__A2
timestamp 1698431365
transform -1 0 6160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._107__A3
timestamp 1698431365
transform 1 0 5824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._110__A1
timestamp 1698431365
transform 1 0 7504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._185__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._185__RN
timestamp 1698431365
transform 1 0 13552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._186__CLK
timestamp 1698431365
transform 1 0 15120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._186__RN
timestamp 1698431365
transform 1 0 15568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._189__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._189__RN
timestamp 1698431365
transform 1 0 6048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._190__CLK
timestamp 1698431365
transform -1 0 8400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._190__RN
timestamp 1698431365
transform 1 0 7952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._191__CLK
timestamp 1698431365
transform 1 0 10864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._191__RN
timestamp 1698431365
transform 1 0 11312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._192__CLK
timestamp 1698431365
transform 1 0 10080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._192__RN
timestamp 1698431365
transform 1 0 14000 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._231__I
timestamp 1698431365
transform -1 0 2688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._232__I
timestamp 1698431365
transform 1 0 1792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._233__I
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._234__I
timestamp 1698431365
transform -1 0 2016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._235__I
timestamp 1698431365
transform 1 0 1792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._236__I
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._237__I
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._238__I
timestamp 1698431365
transform 1 0 2464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._239__I
timestamp 1698431365
transform -1 0 2688 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._240__I
timestamp 1698431365
transform 1 0 2352 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._241__I
timestamp 1698431365
transform -1 0 2688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._242__I
timestamp 1698431365
transform 1 0 2464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._243__I
timestamp 1698431365
transform 1 0 2016 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._244__I
timestamp 1698431365
transform -1 0 2688 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._245__I
timestamp 1698431365
transform -1 0 2688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._246__I
timestamp 1698431365
transform 1 0 2464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._247__I
timestamp 1698431365
transform 1 0 2464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._248__I
timestamp 1698431365
transform -1 0 2240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._249__I
timestamp 1698431365
transform 1 0 2464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._250__I
timestamp 1698431365
transform 1 0 2464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._251__I
timestamp 1698431365
transform -1 0 2688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._252__I
timestamp 1698431365
transform 1 0 2464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._253__I
timestamp 1698431365
transform -1 0 2688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._254__I
timestamp 1698431365
transform -1 0 2688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._255__I
timestamp 1698431365
transform -1 0 2576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._256__I
timestamp 1698431365
transform 1 0 2464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._257__I
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._258__I
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._259__I
timestamp 1698431365
transform -1 0 2688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._260__I
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._261__I
timestamp 1698431365
transform -1 0 2016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._262__I
timestamp 1698431365
transform -1 0 2240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._263__I
timestamp 1698431365
transform -1 0 2688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._264__I
timestamp 1698431365
transform -1 0 2240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._265__I
timestamp 1698431365
transform 1 0 1792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._266__I
timestamp 1698431365
transform -1 0 2016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._267__I
timestamp 1698431365
transform -1 0 2688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._268__I
timestamp 1698431365
transform 1 0 2016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._269__I
timestamp 1698431365
transform -1 0 2016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_async_reg_bus._270__I
timestamp 1698431365
transform 1 0 2016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._405__I
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._406__I
timestamp 1698431365
transform 1 0 37968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._407__I
timestamp 1698431365
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._408__I
timestamp 1698431365
transform 1 0 37072 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._409__I
timestamp 1698431365
transform 1 0 33600 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._414__I
timestamp 1698431365
transform 1 0 30128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._415__I
timestamp 1698431365
transform 1 0 33712 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._423__I
timestamp 1698431365
transform 1 0 14336 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._432__I1
timestamp 1698431365
transform -1 0 31920 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._434__A3
timestamp 1698431365
transform 1 0 17472 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._438__A1
timestamp 1698431365
transform 1 0 7840 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._438__A2
timestamp 1698431365
transform 1 0 9184 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._439__A2
timestamp 1698431365
transform 1 0 20384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._441__A2
timestamp 1698431365
transform 1 0 6832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._441__A3
timestamp 1698431365
transform 1 0 8960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._443__A1
timestamp 1698431365
transform 1 0 8736 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._445__A1
timestamp 1698431365
transform -1 0 10752 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._448__A1
timestamp 1698431365
transform 1 0 10752 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._450__B
timestamp 1698431365
transform -1 0 11200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._451__A1
timestamp 1698431365
transform 1 0 9968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._451__B
timestamp 1698431365
transform 1 0 8176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._453__A1
timestamp 1698431365
transform 1 0 13776 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._453__A2
timestamp 1698431365
transform 1 0 8400 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._457__I
timestamp 1698431365
transform 1 0 12096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._458__I0
timestamp 1698431365
transform 1 0 27440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._458__I1
timestamp 1698431365
transform 1 0 29568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._460__A3
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._465__A2
timestamp 1698431365
transform -1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._466__A2
timestamp 1698431365
transform 1 0 31472 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._469__A3
timestamp 1698431365
transform 1 0 31808 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._473__A1
timestamp 1698431365
transform 1 0 37520 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._473__A2
timestamp 1698431365
transform 1 0 33824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._474__A1
timestamp 1698431365
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._474__A2
timestamp 1698431365
transform 1 0 37520 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._481__A1
timestamp 1698431365
transform 1 0 32256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._482__A2
timestamp 1698431365
transform 1 0 32704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._483__A3
timestamp 1698431365
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._487__A2
timestamp 1698431365
transform 1 0 34160 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._493__A3
timestamp 1698431365
transform 1 0 37856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._496__A1
timestamp 1698431365
transform 1 0 37520 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._496__A3
timestamp 1698431365
transform 1 0 37968 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._497__C
timestamp 1698431365
transform -1 0 37296 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._498__A3
timestamp 1698431365
transform 1 0 33264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._501__A2
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._502__A2
timestamp 1698431365
transform 1 0 37408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._514__B
timestamp 1698431365
transform 1 0 14784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._521__A2
timestamp 1698431365
transform -1 0 35280 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._522__A2
timestamp 1698431365
transform 1 0 34608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._523__S
timestamp 1698431365
transform -1 0 33936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._541__I
timestamp 1698431365
transform 1 0 31472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._542__A2
timestamp 1698431365
transform 1 0 31808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._546__A2
timestamp 1698431365
transform -1 0 28000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._549__A1
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._550__I
timestamp 1698431365
transform 1 0 11872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._554__A1
timestamp 1698431365
transform 1 0 31248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._555__A1
timestamp 1698431365
transform 1 0 28560 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._556__A1
timestamp 1698431365
transform 1 0 32704 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._568__A1
timestamp 1698431365
transform 1 0 29792 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._570__A1
timestamp 1698431365
transform 1 0 30912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._571__A1
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._573__B
timestamp 1698431365
transform 1 0 31024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._574__A1
timestamp 1698431365
transform 1 0 30800 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._575__A1
timestamp 1698431365
transform 1 0 26992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._580__S
timestamp 1698431365
transform 1 0 30912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._582__S
timestamp 1698431365
transform 1 0 29232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._583__A2
timestamp 1698431365
transform 1 0 30464 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._585__A1
timestamp 1698431365
transform -1 0 28112 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._586__A1
timestamp 1698431365
transform 1 0 30912 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._587__A1
timestamp 1698431365
transform 1 0 33712 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._590__A1
timestamp 1698431365
transform 1 0 33376 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._594__A1
timestamp 1698431365
transform 1 0 34272 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._595__B
timestamp 1698431365
transform 1 0 36400 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._599__A1
timestamp 1698431365
transform 1 0 33824 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._601__A1
timestamp 1698431365
transform 1 0 35504 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._605__A1
timestamp 1698431365
transform 1 0 35168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._607__A1
timestamp 1698431365
transform 1 0 34944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._608__B
timestamp 1698431365
transform 1 0 35504 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._612__A1
timestamp 1698431365
transform 1 0 34272 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._614__A1
timestamp 1698431365
transform 1 0 31136 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._619__A1
timestamp 1698431365
transform 1 0 30352 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._620__A1
timestamp 1698431365
transform 1 0 10864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._621__B
timestamp 1698431365
transform 1 0 12320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._622__A2
timestamp 1698431365
transform 1 0 12320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._622__B
timestamp 1698431365
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._625__A1
timestamp 1698431365
transform 1 0 9520 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._626__B
timestamp 1698431365
transform 1 0 10304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._627__A1
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._627__B
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._628__A1
timestamp 1698431365
transform 1 0 7728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._629__A1
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._630__A1
timestamp 1698431365
transform 1 0 6384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._632__A1
timestamp 1698431365
transform 1 0 7504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._633__A1
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._634__A1
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._635__A1
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._636__A1
timestamp 1698431365
transform 1 0 10528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._636__B
timestamp 1698431365
transform -1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._639__A1
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._640__A1
timestamp 1698431365
transform 1 0 6720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._642__A1
timestamp 1698431365
transform -1 0 16016 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._643__A2
timestamp 1698431365
transform 1 0 15120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._644__A1
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._645__A1
timestamp 1698431365
transform 1 0 15568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._646__A1
timestamp 1698431365
transform 1 0 17584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._646__A2
timestamp 1698431365
transform 1 0 18480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._649__A1
timestamp 1698431365
transform 1 0 11424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._650__A1
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._652__A1
timestamp 1698431365
transform 1 0 12208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._653__A1
timestamp 1698431365
transform 1 0 13664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._653__A3
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._657__A1
timestamp 1698431365
transform 1 0 8400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._658__A1
timestamp 1698431365
transform 1 0 8736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._658__A3
timestamp 1698431365
transform -1 0 8512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._661__A1
timestamp 1698431365
transform 1 0 27328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._663__A1
timestamp 1698431365
transform -1 0 26880 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._664__A1
timestamp 1698431365
transform 1 0 26768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._667__B
timestamp 1698431365
transform 1 0 24864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._668__A1
timestamp 1698431365
transform 1 0 23744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._669__A1
timestamp 1698431365
transform 1 0 17584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._670__A2
timestamp 1698431365
transform 1 0 31472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._670__B
timestamp 1698431365
transform 1 0 30912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._675__A1
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._679__A1
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._681__A1
timestamp 1698431365
transform 1 0 31024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._683__A1
timestamp 1698431365
transform 1 0 28448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._685__S
timestamp 1698431365
transform 1 0 23744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._686__A1
timestamp 1698431365
transform 1 0 22400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._689__A2
timestamp 1698431365
transform 1 0 31920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._690__A1
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._691__A1
timestamp 1698431365
transform -1 0 30800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._691__B
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._693__A1
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._695__A1
timestamp 1698431365
transform 1 0 31360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._696__A1
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._698__A1
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._699__B
timestamp 1698431365
transform 1 0 30240 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._700__A1
timestamp 1698431365
transform 1 0 23856 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._702__A2
timestamp 1698431365
transform 1 0 26768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._703__B
timestamp 1698431365
transform 1 0 27552 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._704__B2
timestamp 1698431365
transform 1 0 29680 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._705__A1
timestamp 1698431365
transform -1 0 30240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._706__A1
timestamp 1698431365
transform 1 0 29120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._706__B2
timestamp 1698431365
transform 1 0 30912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._707__A1
timestamp 1698431365
transform 1 0 30576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._709__A2
timestamp 1698431365
transform 1 0 37968 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._710__A1
timestamp 1698431365
transform 1 0 32144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._710__B2
timestamp 1698431365
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._712__A1
timestamp 1698431365
transform 1 0 30800 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._713__A1
timestamp 1698431365
transform 1 0 32480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._713__A2
timestamp 1698431365
transform -1 0 32256 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._715__A1
timestamp 1698431365
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._717__A1
timestamp 1698431365
transform 1 0 31920 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._720__A1
timestamp 1698431365
transform 1 0 15904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._721__A1
timestamp 1698431365
transform 1 0 15792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._721__A2
timestamp 1698431365
transform 1 0 16240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._722__A1
timestamp 1698431365
transform 1 0 18480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._722__A2
timestamp 1698431365
transform 1 0 16688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._723__A1
timestamp 1698431365
transform 1 0 18928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._723__A2
timestamp 1698431365
transform 1 0 16912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._723__C
timestamp 1698431365
transform 1 0 18480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._725__A1
timestamp 1698431365
transform 1 0 14672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._726__A1
timestamp 1698431365
transform 1 0 17584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._726__A2
timestamp 1698431365
transform 1 0 16688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._726__B
timestamp 1698431365
transform 1 0 16240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._727__A1
timestamp 1698431365
transform 1 0 16688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._727__A2
timestamp 1698431365
transform 1 0 18032 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._727__A3
timestamp 1698431365
transform -1 0 16912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._728__A1
timestamp 1698431365
transform 1 0 16240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._729__A1
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._730__A1
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._730__B
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._731__A1
timestamp 1698431365
transform -1 0 17472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._733__A1
timestamp 1698431365
transform 1 0 6160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._736__A1
timestamp 1698431365
transform 1 0 7504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._737__A1
timestamp 1698431365
transform 1 0 5712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._739__C
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._741__A1
timestamp 1698431365
transform 1 0 7728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._742__A1
timestamp 1698431365
transform 1 0 9632 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._742__A2
timestamp 1698431365
transform 1 0 9072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._743__A1
timestamp 1698431365
transform 1 0 7280 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._743__A2
timestamp 1698431365
transform 1 0 8288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._745__A1
timestamp 1698431365
transform 1 0 6944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._746__A1
timestamp 1698431365
transform 1 0 8176 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._747__A1
timestamp 1698431365
transform 1 0 9632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._747__A2
timestamp 1698431365
transform 1 0 9184 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._748__A1
timestamp 1698431365
transform 1 0 9632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._748__A2
timestamp 1698431365
transform 1 0 8848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._748__C
timestamp 1698431365
transform 1 0 7280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._750__A1
timestamp 1698431365
transform 1 0 8512 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._750__A2
timestamp 1698431365
transform 1 0 8960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._751__A1
timestamp 1698431365
transform 1 0 10080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._752__A1
timestamp 1698431365
transform 1 0 10528 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._752__A2
timestamp 1698431365
transform 1 0 10976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._753__A1
timestamp 1698431365
transform 1 0 10640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._753__A2
timestamp 1698431365
transform -1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._753__A3
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._754__A1
timestamp 1698431365
transform 1 0 12208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._755__A1
timestamp 1698431365
transform 1 0 7504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._755__B2
timestamp 1698431365
transform -1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._757__A1
timestamp 1698431365
transform 1 0 14000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._758__A1
timestamp 1698431365
transform 1 0 8960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._758__B2
timestamp 1698431365
transform 1 0 11200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._760__A1
timestamp 1698431365
transform 1 0 5712 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._762__A1
timestamp 1698431365
transform 1 0 8512 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._763__A1
timestamp 1698431365
transform 1 0 5152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._764__A1
timestamp 1698431365
transform 1 0 8064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._765__A1
timestamp 1698431365
transform 1 0 6944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._766__A1
timestamp 1698431365
transform 1 0 6496 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._767__A1
timestamp 1698431365
transform 1 0 8176 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._769__S
timestamp 1698431365
transform 1 0 6496 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._770__A1
timestamp 1698431365
transform 1 0 6944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._771__A1
timestamp 1698431365
transform -1 0 7840 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._771__A2
timestamp 1698431365
transform 1 0 8736 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._772__A1
timestamp 1698431365
transform 1 0 6384 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._773__A1
timestamp 1698431365
transform 1 0 16688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._773__A2
timestamp 1698431365
transform 1 0 17136 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._774__A2
timestamp 1698431365
transform 1 0 18032 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._775__A1
timestamp 1698431365
transform 1 0 18256 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._776__A1
timestamp 1698431365
transform 1 0 20272 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._778__A2
timestamp 1698431365
transform 1 0 18704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._778__A3
timestamp 1698431365
transform 1 0 17584 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._779__A2
timestamp 1698431365
transform 1 0 17136 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._779__A3
timestamp 1698431365
transform 1 0 17808 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._779__A4
timestamp 1698431365
transform 1 0 17584 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._780__B
timestamp 1698431365
transform 1 0 19376 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._782__S
timestamp 1698431365
transform 1 0 21392 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._784__A1
timestamp 1698431365
transform 1 0 19264 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._785__A1
timestamp 1698431365
transform 1 0 19040 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._788__A1
timestamp 1698431365
transform 1 0 5936 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._789__A1
timestamp 1698431365
transform 1 0 7280 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._790__B
timestamp 1698431365
transform 1 0 6496 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._793__A1
timestamp 1698431365
transform 1 0 5824 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._796__A1
timestamp 1698431365
transform 1 0 6720 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._798__A2
timestamp 1698431365
transform 1 0 23632 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._799__A1
timestamp 1698431365
transform -1 0 22624 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._800__A1
timestamp 1698431365
transform 1 0 21952 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._801__A1
timestamp 1698431365
transform 1 0 20496 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._801__A2
timestamp 1698431365
transform 1 0 20048 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._802__A1
timestamp 1698431365
transform 1 0 12880 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._803__A1
timestamp 1698431365
transform 1 0 15456 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._806__A3
timestamp 1698431365
transform 1 0 13888 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._808__A4
timestamp 1698431365
transform 1 0 14448 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._809__C
timestamp 1698431365
transform 1 0 13440 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._810__A1
timestamp 1698431365
transform 1 0 15008 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._812__A1
timestamp 1698431365
transform 1 0 18816 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._815__CLK
timestamp 1698431365
transform -1 0 31584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._815__SETN
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._816__CLK
timestamp 1698431365
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._816__RN
timestamp 1698431365
transform 1 0 28224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._817__CLK
timestamp 1698431365
transform 1 0 29680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._817__RN
timestamp 1698431365
transform 1 0 29680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._818__CLK
timestamp 1698431365
transform 1 0 30912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._818__RN
timestamp 1698431365
transform 1 0 31360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._819__CLK
timestamp 1698431365
transform 1 0 28560 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._819__RN
timestamp 1698431365
transform 1 0 28112 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._820__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._820__RN
timestamp 1698431365
transform 1 0 33824 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._821__CLK
timestamp 1698431365
transform 1 0 30016 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._821__RN
timestamp 1698431365
transform 1 0 34272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._822__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._822__RN
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._823__CLK
timestamp 1698431365
transform 1 0 34048 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._823__RN
timestamp 1698431365
transform 1 0 33600 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._824__CLK
timestamp 1698431365
transform 1 0 33712 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._824__RN
timestamp 1698431365
transform 1 0 34384 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._825__CLK
timestamp 1698431365
transform 1 0 34160 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._825__RN
timestamp 1698431365
transform 1 0 34384 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._826__CLK
timestamp 1698431365
transform 1 0 33376 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._826__RN
timestamp 1698431365
transform 1 0 33600 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._827__RN
timestamp 1698431365
transform 1 0 33712 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._828__RN
timestamp 1698431365
transform 1 0 33712 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._829__RN
timestamp 1698431365
transform 1 0 32480 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._830__RN
timestamp 1698431365
transform -1 0 31920 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._831__RN
timestamp 1698431365
transform 1 0 29792 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._832__RN
timestamp 1698431365
transform 1 0 28560 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._833__RN
timestamp 1698431365
transform -1 0 33040 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._834__CLK
timestamp 1698431365
transform 1 0 10080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._834__RN
timestamp 1698431365
transform 1 0 14560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._835__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._835__RN
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._836__CLK
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._836__RN
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._837__CLK
timestamp 1698431365
transform 1 0 9520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._837__RN
timestamp 1698431365
transform 1 0 9968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._838__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._838__RN
timestamp 1698431365
transform 1 0 17920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._839__CLK
timestamp 1698431365
transform 1 0 17584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._839__RN
timestamp 1698431365
transform 1 0 18032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._840__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._840__RN
timestamp 1698431365
transform 1 0 14560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._841__CLK
timestamp 1698431365
transform 1 0 13664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._841__RN
timestamp 1698431365
transform 1 0 14112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._842__CLK
timestamp 1698431365
transform 1 0 30016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._842__RN
timestamp 1698431365
transform 1 0 29568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._843__CLK
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._843__RN
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._844__CLK
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._844__RN
timestamp 1698431365
transform 1 0 22400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._845__CLK
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._845__RN
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._846__CLK
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._846__RN
timestamp 1698431365
transform 1 0 31584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._847__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._847__RN
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._848__CLK
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._848__RN
timestamp 1698431365
transform -1 0 28000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._849__CLK
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._849__RN
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._850__CLK
timestamp 1698431365
transform 1 0 30128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._850__RN
timestamp 1698431365
transform 1 0 31808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._851__CLK
timestamp 1698431365
transform 1 0 31024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._851__RN
timestamp 1698431365
transform 1 0 30576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._852__CLK
timestamp 1698431365
transform 1 0 26208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._852__RN
timestamp 1698431365
transform 1 0 29904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._853__CLK
timestamp 1698431365
transform 1 0 29904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._853__SETN
timestamp 1698431365
transform 1 0 30128 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._854__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._854__RN
timestamp 1698431365
transform 1 0 34272 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._855__CLK
timestamp 1698431365
transform 1 0 30016 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._855__RN
timestamp 1698431365
transform 1 0 30912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._856__CLK
timestamp 1698431365
transform 1 0 31136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._856__RN
timestamp 1698431365
transform 1 0 30688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._857__CLK
timestamp 1698431365
transform 1 0 22176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._857__SETN
timestamp 1698431365
transform 1 0 21728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._858__CLK
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._858__RN
timestamp 1698431365
transform 1 0 21392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._859__CLK
timestamp 1698431365
transform 1 0 19264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._859__RN
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._860__CLK
timestamp 1698431365
transform 1 0 11536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._860__RN
timestamp 1698431365
transform 1 0 11984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._861__CLK
timestamp 1698431365
transform 1 0 10864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._861__RN
timestamp 1698431365
transform 1 0 11312 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._862__CLK
timestamp 1698431365
transform -1 0 11088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._862__RN
timestamp 1698431365
transform 1 0 10304 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._863__CLK
timestamp 1698431365
transform 1 0 11312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._863__RN
timestamp 1698431365
transform 1 0 11760 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._864__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._864__RN
timestamp 1698431365
transform 1 0 15904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._865__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._865__RN
timestamp 1698431365
transform 1 0 14896 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._866__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._866__RN
timestamp 1698431365
transform 1 0 10080 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._867__CLK
timestamp 1698431365
transform 1 0 9744 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._867__RN
timestamp 1698431365
transform 1 0 9632 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._868__CLK
timestamp 1698431365
transform 1 0 7392 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._868__RN
timestamp 1698431365
transform 1 0 6832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._869__CLK
timestamp 1698431365
transform 1 0 9408 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._869__RN
timestamp 1698431365
transform 1 0 9856 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._870__RN
timestamp 1698431365
transform 1 0 27552 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._871__CLK
timestamp 1698431365
transform 1 0 23408 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._871__RN
timestamp 1698431365
transform 1 0 22288 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._872__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._872__RN
timestamp 1698431365
transform 1 0 16912 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._873__CLK
timestamp 1698431365
transform 1 0 9408 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._873__RN
timestamp 1698431365
transform 1 0 9184 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._874__CLK
timestamp 1698431365
transform 1 0 6272 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._874__RN
timestamp 1698431365
transform 1 0 6720 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._875__CLK
timestamp 1698431365
transform 1 0 6944 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._875__RN
timestamp 1698431365
transform 1 0 7392 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._876__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._876__RN
timestamp 1698431365
transform 1 0 25312 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._877__CLK
timestamp 1698431365
transform 1 0 14336 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._877__RN
timestamp 1698431365
transform 1 0 19936 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._878__CLK
timestamp 1698431365
transform 1 0 12208 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._878__RN
timestamp 1698431365
transform 1 0 17472 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._879__CLK
timestamp 1698431365
transform 1 0 15904 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._879__RN
timestamp 1698431365
transform 1 0 21392 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_core._880__RN
timestamp 1698431365
transform 1 0 29344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0604__I
timestamp 1698431365
transform -1 0 2352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0616__I
timestamp 1698431365
transform 1 0 18032 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0619__I
timestamp 1698431365
transform 1 0 19264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0621__I
timestamp 1698431365
transform 1 0 18704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0641__I
timestamp 1698431365
transform -1 0 19376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0669__A1
timestamp 1698431365
transform 1 0 23072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0670__A1
timestamp 1698431365
transform 1 0 24304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0673__A1
timestamp 1698431365
transform -1 0 18480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0673__A2
timestamp 1698431365
transform -1 0 15568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0674__B2
timestamp 1698431365
transform -1 0 16128 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0675__A1
timestamp 1698431365
transform 1 0 17472 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0681__A1
timestamp 1698431365
transform 1 0 17472 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0682__A1
timestamp 1698431365
transform 1 0 15456 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0685__A1
timestamp 1698431365
transform 1 0 17248 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0687__A1
timestamp 1698431365
transform 1 0 14672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0688__A1
timestamp 1698431365
transform 1 0 11536 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0689__A1
timestamp 1698431365
transform 1 0 11424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0690__A1
timestamp 1698431365
transform 1 0 11984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0705__A1
timestamp 1698431365
transform 1 0 16128 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0706__A1
timestamp 1698431365
transform 1 0 13664 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0706__B2
timestamp 1698431365
transform 1 0 16576 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0707__A1
timestamp 1698431365
transform 1 0 12432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0707__B2
timestamp 1698431365
transform -1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0708__A1
timestamp 1698431365
transform -1 0 11424 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0709__A2
timestamp 1698431365
transform 1 0 15680 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0714__A1
timestamp 1698431365
transform 1 0 12768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0715__A1
timestamp 1698431365
transform 1 0 12208 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0715__B2
timestamp 1698431365
transform 1 0 14448 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0718__A2
timestamp 1698431365
transform 1 0 24864 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0719__A2
timestamp 1698431365
transform -1 0 22400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0722__B2
timestamp 1698431365
transform 1 0 21392 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0723__A2
timestamp 1698431365
transform 1 0 18368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0724__A2
timestamp 1698431365
transform 1 0 19600 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0726__A4
timestamp 1698431365
transform 1 0 20048 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0729__A2
timestamp 1698431365
transform -1 0 17920 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0730__A2
timestamp 1698431365
transform 1 0 16688 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0733__A2
timestamp 1698431365
transform -1 0 17696 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0735__B
timestamp 1698431365
transform 1 0 19824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0736__A2
timestamp 1698431365
transform 1 0 15456 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0737__A2
timestamp 1698431365
transform 1 0 16800 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0738__A2
timestamp 1698431365
transform -1 0 14336 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0739__A2
timestamp 1698431365
transform 1 0 15008 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0742__B1
timestamp 1698431365
transform 1 0 19712 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0753__A2
timestamp 1698431365
transform 1 0 16800 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0755__A2
timestamp 1698431365
transform -1 0 15456 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0756__A2
timestamp 1698431365
transform 1 0 18144 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0758__A2
timestamp 1698431365
transform 1 0 17696 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0762__A3
timestamp 1698431365
transform 1 0 15120 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0763__A1
timestamp 1698431365
transform -1 0 14112 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0763__B2
timestamp 1698431365
transform 1 0 14896 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0769__A1
timestamp 1698431365
transform 1 0 3808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0770__A1
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0771__A1
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0772__A1
timestamp 1698431365
transform 1 0 8848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0773__A2
timestamp 1698431365
transform -1 0 8400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0775__I0
timestamp 1698431365
transform -1 0 15344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0775__I1
timestamp 1698431365
transform 1 0 14112 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0775__S
timestamp 1698431365
transform 1 0 13664 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0777__I0
timestamp 1698431365
transform -1 0 17024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0777__I1
timestamp 1698431365
transform -1 0 14448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0777__S
timestamp 1698431365
transform 1 0 13888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0779__I0
timestamp 1698431365
transform -1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0779__S
timestamp 1698431365
transform 1 0 11536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0792__A1
timestamp 1698431365
transform 1 0 4144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0793__A2
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0794__A1
timestamp 1698431365
transform 1 0 14112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0794__A2
timestamp 1698431365
transform 1 0 12880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0795__A1
timestamp 1698431365
transform 1 0 14560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0796__I1
timestamp 1698431365
transform -1 0 27104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0796__S
timestamp 1698431365
transform 1 0 26656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0797__S
timestamp 1698431365
transform 1 0 27328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0798__I1
timestamp 1698431365
transform 1 0 24864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0798__S
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0799__S
timestamp 1698431365
transform 1 0 25312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0800__I1
timestamp 1698431365
transform 1 0 26208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0800__S
timestamp 1698431365
transform 1 0 26208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0801__S
timestamp 1698431365
transform 1 0 26096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0802__I1
timestamp 1698431365
transform -1 0 25648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0802__S
timestamp 1698431365
transform 1 0 26880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0803__S
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0804__I0
timestamp 1698431365
transform 1 0 25200 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0804__I1
timestamp 1698431365
transform -1 0 22624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0804__S
timestamp 1698431365
transform -1 0 23072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0805__S
timestamp 1698431365
transform 1 0 22512 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0810__A1
timestamp 1698431365
transform 1 0 14000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0810__A2
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0811__A1
timestamp 1698431365
transform 1 0 15008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0812__I1
timestamp 1698431365
transform -1 0 21728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0812__S
timestamp 1698431365
transform 1 0 21952 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0813__S
timestamp 1698431365
transform 1 0 22288 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0814__I1
timestamp 1698431365
transform 1 0 18816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0814__S
timestamp 1698431365
transform 1 0 18368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0815__S
timestamp 1698431365
transform 1 0 18816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0816__I1
timestamp 1698431365
transform 1 0 18704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0816__S
timestamp 1698431365
transform 1 0 18256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0817__S
timestamp 1698431365
transform 1 0 18816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0818__I1
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0818__S
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0819__S
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0820__I1
timestamp 1698431365
transform 1 0 22176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0820__S
timestamp 1698431365
transform 1 0 21952 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0821__S
timestamp 1698431365
transform 1 0 22400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0822__I1
timestamp 1698431365
transform -1 0 18704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0822__S
timestamp 1698431365
transform 1 0 18032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0823__S
timestamp 1698431365
transform 1 0 20160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0824__S
timestamp 1698431365
transform 1 0 17136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0825__S
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0826__S
timestamp 1698431365
transform 1 0 15120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0827__S
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0828__A2
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0829__A1
timestamp 1698431365
transform 1 0 7616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0830__I1
timestamp 1698431365
transform 1 0 15008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0830__S
timestamp 1698431365
transform 1 0 13888 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0831__S
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0832__I1
timestamp 1698431365
transform 1 0 12992 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0832__S
timestamp 1698431365
transform 1 0 12544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0833__S
timestamp 1698431365
transform 1 0 14112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0834__S
timestamp 1698431365
transform 1 0 9184 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0835__S
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0836__I0
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0836__S
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0837__S
timestamp 1698431365
transform 1 0 7504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0838__S
timestamp 1698431365
transform -1 0 5376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0839__S
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0840__S
timestamp 1698431365
transform 1 0 5712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0841__S
timestamp 1698431365
transform 1 0 4704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0842__S
timestamp 1698431365
transform 1 0 5264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0843__S
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0844__B1
timestamp 1698431365
transform 1 0 3808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0846__A1
timestamp 1698431365
transform 1 0 9744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0847__A1
timestamp 1698431365
transform 1 0 10864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0847__A2
timestamp 1698431365
transform 1 0 10416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0848__A1
timestamp 1698431365
transform 1 0 10528 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0848__A2
timestamp 1698431365
transform 1 0 12544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0849__A2
timestamp 1698431365
transform 1 0 11648 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0850__I0
timestamp 1698431365
transform 1 0 8736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0850__S
timestamp 1698431365
transform -1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0851__A1
timestamp 1698431365
transform 1 0 10080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0851__A2
timestamp 1698431365
transform 1 0 13552 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0852__A2
timestamp 1698431365
transform -1 0 12544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0853__I0
timestamp 1698431365
transform 1 0 8960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0853__S
timestamp 1698431365
transform 1 0 11088 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0854__A1
timestamp 1698431365
transform 1 0 15344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0854__A2
timestamp 1698431365
transform 1 0 13104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0855__A1
timestamp 1698431365
transform -1 0 13776 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0855__A2
timestamp 1698431365
transform 1 0 12656 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0856__A2
timestamp 1698431365
transform 1 0 11200 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0857__A2
timestamp 1698431365
transform 1 0 12320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0858__A2
timestamp 1698431365
transform 1 0 20944 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0859__A1
timestamp 1698431365
transform 1 0 19824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0859__A2
timestamp 1698431365
transform 1 0 19376 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0860__A2
timestamp 1698431365
transform 1 0 20272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0861__A2
timestamp 1698431365
transform 1 0 20720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0862__A1
timestamp 1698431365
transform 1 0 11872 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0862__A2
timestamp 1698431365
transform 1 0 11424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0863__I0
timestamp 1698431365
transform 1 0 19488 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0864__A1
timestamp 1698431365
transform 1 0 16128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0886__A1
timestamp 1698431365
transform 1 0 7728 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0887__A1
timestamp 1698431365
transform 1 0 13104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0887__A2
timestamp 1698431365
transform 1 0 13552 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0888__A1
timestamp 1698431365
transform 1 0 22512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0888__A2
timestamp 1698431365
transform 1 0 22064 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0889__A2
timestamp 1698431365
transform 1 0 20272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0890__I0
timestamp 1698431365
transform 1 0 25312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0890__S
timestamp 1698431365
transform 1 0 24640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0891__A1
timestamp 1698431365
transform 1 0 21616 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0891__A2
timestamp 1698431365
transform 1 0 21392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0892__A2
timestamp 1698431365
transform -1 0 22624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0893__A1
timestamp 1698431365
transform 1 0 18928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0893__A2
timestamp 1698431365
transform 1 0 20048 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0894__A2
timestamp 1698431365
transform 1 0 18368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0895__A1
timestamp 1698431365
transform 1 0 18704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0895__A2
timestamp 1698431365
transform 1 0 16352 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0896__A2
timestamp 1698431365
transform 1 0 15904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0897__A2
timestamp 1698431365
transform 1 0 14000 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0898__A2
timestamp 1698431365
transform 1 0 14448 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0899__A2
timestamp 1698431365
transform 1 0 24192 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0900__A1
timestamp 1698431365
transform 1 0 21616 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0900__A2
timestamp 1698431365
transform 1 0 22064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0901__A2
timestamp 1698431365
transform 1 0 25312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0902__A2
timestamp 1698431365
transform 1 0 21616 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0903__A1
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0903__A2
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0904__I0
timestamp 1698431365
transform 1 0 19040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0905__A1
timestamp 1698431365
transform 1 0 16128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0927__A1
timestamp 1698431365
transform 1 0 7952 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0927__A2
timestamp 1698431365
transform -1 0 8624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0928__A1
timestamp 1698431365
transform 1 0 26320 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0928__A2
timestamp 1698431365
transform 1 0 26656 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0929__A2
timestamp 1698431365
transform 1 0 23744 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0930__A1
timestamp 1698431365
transform 1 0 25872 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0930__A2
timestamp 1698431365
transform 1 0 24976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0931__A2
timestamp 1698431365
transform 1 0 24640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0932__I0
timestamp 1698431365
transform 1 0 11200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0932__S
timestamp 1698431365
transform 1 0 11648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0933__I0
timestamp 1698431365
transform 1 0 27440 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0933__S
timestamp 1698431365
transform 1 0 26992 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0934__I0
timestamp 1698431365
transform -1 0 24304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0934__S
timestamp 1698431365
transform 1 0 24528 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0937__A2
timestamp 1698431365
transform 1 0 26544 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0938__A1
timestamp 1698431365
transform -1 0 23856 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0938__A2
timestamp 1698431365
transform 1 0 24080 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0939__A2
timestamp 1698431365
transform 1 0 25984 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0940__A2
timestamp 1698431365
transform 1 0 23856 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0945__A1
timestamp 1698431365
transform 1 0 8176 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0945__A2
timestamp 1698431365
transform 1 0 6384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0946__A1
timestamp 1698431365
transform 1 0 7280 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0947__I0
timestamp 1698431365
transform -1 0 3584 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0947__I1
timestamp 1698431365
transform -1 0 3136 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0947__S
timestamp 1698431365
transform 1 0 5712 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0948__S
timestamp 1698431365
transform 1 0 4032 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0949__A1
timestamp 1698431365
transform 1 0 20160 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0949__A2
timestamp 1698431365
transform 1 0 18480 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0950__A2
timestamp 1698431365
transform 1 0 19600 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0951__S
timestamp 1698431365
transform 1 0 21952 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0952__A1
timestamp 1698431365
transform -1 0 19600 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0952__A2
timestamp 1698431365
transform -1 0 20272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0953__A2
timestamp 1698431365
transform -1 0 19152 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0954__S
timestamp 1698431365
transform 1 0 21840 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0955__A1
timestamp 1698431365
transform 1 0 22176 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0955__A2
timestamp 1698431365
transform -1 0 21616 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0956__A2
timestamp 1698431365
transform 1 0 20496 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0957__S
timestamp 1698431365
transform 1 0 21392 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0958__I1
timestamp 1698431365
transform 1 0 6160 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0958__S
timestamp 1698431365
transform 1 0 7056 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0959__S
timestamp 1698431365
transform 1 0 4368 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0960__I0
timestamp 1698431365
transform 1 0 6608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0960__S
timestamp 1698431365
transform 1 0 5488 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0961__S
timestamp 1698431365
transform 1 0 4704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0962__S
timestamp 1698431365
transform 1 0 6160 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0963__S
timestamp 1698431365
transform 1 0 4928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0965__A1
timestamp 1698431365
transform 1 0 4032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0965__A2
timestamp 1698431365
transform -1 0 4704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0966__A1
timestamp 1698431365
transform 1 0 7504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0967__I0
timestamp 1698431365
transform -1 0 6608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0967__I1
timestamp 1698431365
transform -1 0 5376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0967__S
timestamp 1698431365
transform 1 0 6832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0969__I0
timestamp 1698431365
transform 1 0 7168 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0969__I1
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0969__S
timestamp 1698431365
transform 1 0 7392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0971__I0
timestamp 1698431365
transform -1 0 8064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0971__I1
timestamp 1698431365
transform -1 0 6384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0971__S
timestamp 1698431365
transform 1 0 7392 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0973__I0
timestamp 1698431365
transform 1 0 8288 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0973__I1
timestamp 1698431365
transform 1 0 6496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0973__S
timestamp 1698431365
transform 1 0 8624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0975__I1
timestamp 1698431365
transform 1 0 4144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0975__S
timestamp 1698431365
transform 1 0 7952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0977__I1
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0977__S
timestamp 1698431365
transform 1 0 7056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0985__A1
timestamp 1698431365
transform 1 0 10752 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0985__A2
timestamp 1698431365
transform -1 0 2688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0986__A1
timestamp 1698431365
transform 1 0 10640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0986__A2
timestamp 1698431365
transform 1 0 11760 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0987__A2
timestamp 1698431365
transform 1 0 9520 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0988__I0
timestamp 1698431365
transform 1 0 5712 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0988__S
timestamp 1698431365
transform 1 0 6160 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0989__I0
timestamp 1698431365
transform 1 0 10192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0989__S
timestamp 1698431365
transform 1 0 9744 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0990__A1
timestamp 1698431365
transform 1 0 10304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0990__A2
timestamp 1698431365
transform 1 0 9856 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0991__A2
timestamp 1698431365
transform 1 0 10752 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0992__A1
timestamp 1698431365
transform 1 0 10864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0992__A2
timestamp 1698431365
transform 1 0 10416 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0993__A2
timestamp 1698431365
transform 1 0 11200 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0994__I0
timestamp 1698431365
transform 1 0 11200 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0994__S
timestamp 1698431365
transform 1 0 10304 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0995__A2
timestamp 1698431365
transform 1 0 8960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0996__A2
timestamp 1698431365
transform 1 0 7392 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0997__A2
timestamp 1698431365
transform 1 0 6160 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0998__A2
timestamp 1698431365
transform 1 0 5712 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0999__A1
timestamp 1698431365
transform 1 0 9408 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._0999__A2
timestamp 1698431365
transform -1 0 9184 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1000__I0
timestamp 1698431365
transform 1 0 9856 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1000__S
timestamp 1698431365
transform 1 0 12432 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1001__I0
timestamp 1698431365
transform -1 0 7392 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1001__S
timestamp 1698431365
transform 1 0 9296 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1002__I0
timestamp 1698431365
transform -1 0 5936 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1002__S
timestamp 1698431365
transform 1 0 7616 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1003__A1
timestamp 1698431365
transform 1 0 9632 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1003__A2
timestamp 1698431365
transform 1 0 10752 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1004__A2
timestamp 1698431365
transform 1 0 10864 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1005__A1
timestamp 1698431365
transform -1 0 8288 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1005__A2
timestamp 1698431365
transform 1 0 9184 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1006__A2
timestamp 1698431365
transform 1 0 7840 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1007__A1
timestamp 1698431365
transform 1 0 7504 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1007__A2
timestamp 1698431365
transform 1 0 8288 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1008__A2
timestamp 1698431365
transform 1 0 10528 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1009__A2
timestamp 1698431365
transform 1 0 7952 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1010__A2
timestamp 1698431365
transform 1 0 8624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1013__A1
timestamp 1698431365
transform 1 0 9968 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1013__A2
timestamp 1698431365
transform -1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1014__I0
timestamp 1698431365
transform 1 0 20944 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1014__S
timestamp 1698431365
transform -1 0 20720 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1015__A1
timestamp 1698431365
transform 1 0 15680 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1015__A2
timestamp 1698431365
transform 1 0 15232 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1016__A2
timestamp 1698431365
transform 1 0 14896 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1017__A1
timestamp 1698431365
transform 1 0 18480 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1017__A2
timestamp 1698431365
transform 1 0 16128 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1018__A2
timestamp 1698431365
transform 1 0 16800 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1019__I0
timestamp 1698431365
transform 1 0 20720 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1019__S
timestamp 1698431365
transform 1 0 20272 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1020__I0
timestamp 1698431365
transform 1 0 10640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1020__S
timestamp 1698431365
transform 1 0 10192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1021__A1
timestamp 1698431365
transform 1 0 12208 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1021__A2
timestamp 1698431365
transform 1 0 11760 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1022__A2
timestamp 1698431365
transform 1 0 13328 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1023__A2
timestamp 1698431365
transform -1 0 8624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1024__A2
timestamp 1698431365
transform 1 0 10528 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1027__A1
timestamp 1698431365
transform 1 0 11872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1027__A2
timestamp 1698431365
transform 1 0 11648 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1028__A1
timestamp 1698431365
transform -1 0 13776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1029__A2
timestamp 1698431365
transform 1 0 20384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1030__A1
timestamp 1698431365
transform 1 0 20944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1030__A2
timestamp 1698431365
transform 1 0 19712 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1031__A2
timestamp 1698431365
transform 1 0 27216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1032__A1
timestamp 1698431365
transform 1 0 25424 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1033__I0
timestamp 1698431365
transform 1 0 28560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1033__I1
timestamp 1698431365
transform 1 0 26432 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1033__S
timestamp 1698431365
transform 1 0 26208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1034__S
timestamp 1698431365
transform 1 0 27104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1035__I0
timestamp 1698431365
transform -1 0 29456 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1035__I1
timestamp 1698431365
transform -1 0 24752 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1035__S
timestamp 1698431365
transform -1 0 25200 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1036__S
timestamp 1698431365
transform -1 0 27104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1037__I0
timestamp 1698431365
transform -1 0 27664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1037__I1
timestamp 1698431365
transform 1 0 25312 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1037__S
timestamp 1698431365
transform 1 0 25312 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1038__S
timestamp 1698431365
transform 1 0 26992 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1039__I1
timestamp 1698431365
transform -1 0 21616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1039__S
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1040__S
timestamp 1698431365
transform 1 0 22176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1041__A1
timestamp 1698431365
transform -1 0 14000 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1041__A2
timestamp 1698431365
transform 1 0 13328 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1042__A2
timestamp 1698431365
transform 1 0 19040 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1043__S
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1046__A1
timestamp 1698431365
transform -1 0 4704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1046__A2
timestamp 1698431365
transform -1 0 4704 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1047__A1
timestamp 1698431365
transform 1 0 8064 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1048__I1
timestamp 1698431365
transform 1 0 20496 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1048__S
timestamp 1698431365
transform 1 0 20272 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1049__S
timestamp 1698431365
transform 1 0 20720 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1050__A2
timestamp 1698431365
transform 1 0 12544 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1051__A1
timestamp 1698431365
transform 1 0 13552 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1051__A2
timestamp 1698431365
transform -1 0 12656 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1052__A2
timestamp 1698431365
transform 1 0 16128 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1053__A1
timestamp 1698431365
transform 1 0 14784 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1054__A1
timestamp 1698431365
transform -1 0 13776 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1054__A2
timestamp 1698431365
transform -1 0 13104 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1055__A2
timestamp 1698431365
transform 1 0 11760 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1056__S
timestamp 1698431365
transform -1 0 13664 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1057__I1
timestamp 1698431365
transform 1 0 18256 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1057__S
timestamp 1698431365
transform -1 0 18256 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1058__S
timestamp 1698431365
transform 1 0 18592 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1059__A1
timestamp 1698431365
transform 1 0 6384 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1059__A2
timestamp 1698431365
transform 1 0 6720 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1060__A2
timestamp 1698431365
transform 1 0 5152 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1061__S
timestamp 1698431365
transform 1 0 4816 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1062__I1
timestamp 1698431365
transform -1 0 4256 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1062__S
timestamp 1698431365
transform 1 0 7056 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1063__S
timestamp 1698431365
transform 1 0 4704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1064__S
timestamp 1698431365
transform 1 0 5264 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1065__S
timestamp 1698431365
transform 1 0 6608 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1067__A1
timestamp 1698431365
transform -1 0 2688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1067__A2
timestamp 1698431365
transform -1 0 3696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1067__B
timestamp 1698431365
transform -1 0 2240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1068__A2
timestamp 1698431365
transform 1 0 4256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1069__A1
timestamp 1698431365
transform -1 0 2688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1071__A1
timestamp 1698431365
transform 1 0 2912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1071__A2
timestamp 1698431365
transform -1 0 3584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1205__CLK
timestamp 1698431365
transform 1 0 11984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1205__RN
timestamp 1698431365
transform 1 0 16240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1206__CLK
timestamp 1698431365
transform 1 0 15232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1206__RN
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1207__CLK
timestamp 1698431365
transform -1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1207__RN
timestamp 1698431365
transform 1 0 14000 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1213__CLK
timestamp 1698431365
transform 1 0 30240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1213__RN
timestamp 1698431365
transform 1 0 29792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1214__CLK
timestamp 1698431365
transform 1 0 28224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1214__RN
timestamp 1698431365
transform 1 0 27776 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1215__CLK
timestamp 1698431365
transform 1 0 29792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1215__RN
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1216__CLK
timestamp 1698431365
transform 1 0 30912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1216__RN
timestamp 1698431365
transform 1 0 26656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1217__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1217__RN
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1221__CLK
timestamp 1698431365
transform 1 0 26432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1221__RN
timestamp 1698431365
transform 1 0 25984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1222__CLK
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1222__RN
timestamp 1698431365
transform -1 0 22064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1223__CLK
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1223__RN
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1224__CLK
timestamp 1698431365
transform 1 0 24192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1224__RN
timestamp 1698431365
transform 1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1225__CLK
timestamp 1698431365
transform 1 0 26544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1225__RN
timestamp 1698431365
transform 1 0 26096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1226__CLK
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1226__RN
timestamp 1698431365
transform -1 0 23744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1227__CLK
timestamp 1698431365
transform 1 0 15568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1227__RN
timestamp 1698431365
transform 1 0 20272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1228__CLK
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1228__RN
timestamp 1698431365
transform 1 0 19376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1229__CLK
timestamp 1698431365
transform 1 0 17360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1229__RN
timestamp 1698431365
transform 1 0 17808 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1230__CLK
timestamp 1698431365
transform 1 0 17360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1230__RN
timestamp 1698431365
transform 1 0 17808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1231__CLK
timestamp 1698431365
transform 1 0 8064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1231__RN
timestamp 1698431365
transform -1 0 11648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1232__CLK
timestamp 1698431365
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1232__RN
timestamp 1698431365
transform 1 0 9968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1233__CLK
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1233__RN
timestamp 1698431365
transform 1 0 6160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1234__CLK
timestamp 1698431365
transform 1 0 5712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1234__RN
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1235__CLK
timestamp 1698431365
transform 1 0 5712 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1235__RN
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1236__CLK
timestamp 1698431365
transform 1 0 5712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1236__RN
timestamp 1698431365
transform 1 0 6160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1237__CLK
timestamp 1698431365
transform 1 0 13888 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1237__RN
timestamp 1698431365
transform 1 0 13552 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1238__CLK
timestamp 1698431365
transform 1 0 11648 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1238__RN
timestamp 1698431365
transform 1 0 9632 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1239__CLK
timestamp 1698431365
transform 1 0 12992 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1239__RN
timestamp 1698431365
transform 1 0 12768 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1240__CLK
timestamp 1698431365
transform 1 0 11872 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1240__RN
timestamp 1698431365
transform 1 0 12320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1241__CLK
timestamp 1698431365
transform 1 0 12880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1241__RN
timestamp 1698431365
transform 1 0 15792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1242__CLK
timestamp 1698431365
transform 1 0 14560 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1242__RN
timestamp 1698431365
transform 1 0 13888 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1243__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1243__RN
timestamp 1698431365
transform 1 0 23744 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1244__CLK
timestamp 1698431365
transform 1 0 24080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1244__RN
timestamp 1698431365
transform 1 0 23632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1245__CLK
timestamp 1698431365
transform 1 0 22848 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1245__RN
timestamp 1698431365
transform 1 0 22400 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1246__CLK
timestamp 1698431365
transform 1 0 19152 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1246__RN
timestamp 1698431365
transform 1 0 19600 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1261__CLK
timestamp 1698431365
transform 1 0 26544 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1261__RN
timestamp 1698431365
transform 1 0 26096 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1262__CLK
timestamp 1698431365
transform 1 0 28112 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1262__RN
timestamp 1698431365
transform 1 0 27664 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1263__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1263__RN
timestamp 1698431365
transform 1 0 25312 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1264__CLK
timestamp 1698431365
transform 1 0 22512 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1264__RN
timestamp 1698431365
transform 1 0 22064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1265__CLK
timestamp 1698431365
transform 1 0 20160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1265__RN
timestamp 1698431365
transform 1 0 19936 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1266__CLK
timestamp 1698431365
transform 1 0 15904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1266__RN
timestamp 1698431365
transform -1 0 15456 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1267__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1267__RN
timestamp 1698431365
transform 1 0 25760 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1268__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1268__RN
timestamp 1698431365
transform 1 0 25312 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1269__CLK
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1269__RN
timestamp 1698431365
transform 1 0 23184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1270__CLK
timestamp 1698431365
transform 1 0 19040 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1270__RN
timestamp 1698431365
transform 1 0 18816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1285__RN
timestamp 1698431365
transform 1 0 29120 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1286__CLK
timestamp 1698431365
transform 1 0 29232 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1286__RN
timestamp 1698431365
transform 1 0 28336 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1287__CLK
timestamp 1698431365
transform 1 0 15008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1287__SETN
timestamp 1698431365
transform 1 0 14784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1288__CLK
timestamp 1698431365
transform 1 0 25760 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1288__RN
timestamp 1698431365
transform -1 0 30016 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1289__CLK
timestamp 1698431365
transform 1 0 29232 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1289__RN
timestamp 1698431365
transform 1 0 29568 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1291__CLK
timestamp 1698431365
transform -1 0 29904 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1291__RN
timestamp 1698431365
transform 1 0 29232 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1292__CLK
timestamp 1698431365
transform 1 0 29232 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1292__RN
timestamp 1698431365
transform -1 0 28448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1294__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1294__RN
timestamp 1698431365
transform -1 0 6272 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1295__CLK
timestamp 1698431365
transform -1 0 25648 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1295__RN
timestamp 1698431365
transform 1 0 24528 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1296__CLK
timestamp 1698431365
transform 1 0 24304 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1296__RN
timestamp 1698431365
transform 1 0 23856 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1297__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1297__RN
timestamp 1698431365
transform 1 0 25648 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1298__CLK
timestamp 1698431365
transform 1 0 5712 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1298__RN
timestamp 1698431365
transform 1 0 5712 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1299__CLK
timestamp 1698431365
transform 1 0 5712 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1299__RN
timestamp 1698431365
transform 1 0 6160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1300__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1300__RN
timestamp 1698431365
transform 1 0 5712 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1302__CLK
timestamp 1698431365
transform -1 0 7056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1302__RN
timestamp 1698431365
transform 1 0 5712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1303__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1303__RN
timestamp 1698431365
transform 1 0 6048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1304__CLK
timestamp 1698431365
transform 1 0 5712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1304__RN
timestamp 1698431365
transform 1 0 5712 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1305__CLK
timestamp 1698431365
transform 1 0 8400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1305__RN
timestamp 1698431365
transform 1 0 8848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1306__CLK
timestamp 1698431365
transform 1 0 5824 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1306__RN
timestamp 1698431365
transform 1 0 6272 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1307__CLK
timestamp 1698431365
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1307__RN
timestamp 1698431365
transform 1 0 4592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1311__CLK
timestamp 1698431365
transform 1 0 14000 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1311__RN
timestamp 1698431365
transform 1 0 13216 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1312__CLK
timestamp 1698431365
transform 1 0 6160 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1312__RN
timestamp 1698431365
transform 1 0 5712 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1313__CLK
timestamp 1698431365
transform 1 0 13440 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1313__RN
timestamp 1698431365
transform 1 0 13888 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1314__CLK
timestamp 1698431365
transform 1 0 16688 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1314__RN
timestamp 1698431365
transform 1 0 14448 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1315__CLK
timestamp 1698431365
transform -1 0 11536 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1315__RN
timestamp 1698431365
transform 1 0 16016 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1316__CLK
timestamp 1698431365
transform 1 0 14784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1316__RN
timestamp 1698431365
transform 1 0 15232 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1317__CLK
timestamp 1698431365
transform -1 0 11200 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1317__RN
timestamp 1698431365
transform 1 0 9968 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1318__CLK
timestamp 1698431365
transform 1 0 7168 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1318__RN
timestamp 1698431365
transform 1 0 7616 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1319__CLK
timestamp 1698431365
transform -1 0 9072 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1319__RN
timestamp 1698431365
transform 1 0 13888 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1320__CLK
timestamp 1698431365
transform 1 0 8848 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1320__RN
timestamp 1698431365
transform 1 0 8400 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1321__CLK
timestamp 1698431365
transform 1 0 7616 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1321__RN
timestamp 1698431365
transform 1 0 7392 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1322__CLK
timestamp 1698431365
transform -1 0 8624 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1322__RN
timestamp 1698431365
transform -1 0 13776 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1323__CLK
timestamp 1698431365
transform 1 0 10304 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1323__RN
timestamp 1698431365
transform 1 0 10752 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1324__CLK
timestamp 1698431365
transform 1 0 11984 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1324__RN
timestamp 1698431365
transform 1 0 11312 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1325__CLK
timestamp 1698431365
transform -1 0 9632 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1325__RN
timestamp 1698431365
transform 1 0 9856 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1327__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1327__RN
timestamp 1698431365
transform 1 0 24304 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1328__CLK
timestamp 1698431365
transform 1 0 15568 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1328__RN
timestamp 1698431365
transform 1 0 19824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1329__CLK
timestamp 1698431365
transform 1 0 15344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1329__RN
timestamp 1698431365
transform 1 0 20496 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1330__CLK
timestamp 1698431365
transform 1 0 25648 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1330__RN
timestamp 1698431365
transform 1 0 25200 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1331__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1331__RN
timestamp 1698431365
transform 1 0 14448 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1332__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1332__RN
timestamp 1698431365
transform 1 0 15904 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1333__CLK
timestamp 1698431365
transform 1 0 11200 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1333__RN
timestamp 1698431365
transform 1 0 10976 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1335__CLK
timestamp 1698431365
transform 1 0 29680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1335__RN
timestamp 1698431365
transform 1 0 29232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1336__CLK
timestamp 1698431365
transform 1 0 31136 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1336__RN
timestamp 1698431365
transform -1 0 27216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1337__CLK
timestamp 1698431365
transform 1 0 30352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1337__RN
timestamp 1698431365
transform 1 0 26320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1338__CLK
timestamp 1698431365
transform 1 0 31136 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1338__RN
timestamp 1698431365
transform 1 0 26432 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1339__CLK
timestamp 1698431365
transform 1 0 26096 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1339__RN
timestamp 1698431365
transform 1 0 25648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1340__CLK
timestamp 1698431365
transform 1 0 24976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1340__RN
timestamp 1698431365
transform 1 0 24528 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1343__CLK
timestamp 1698431365
transform -1 0 24640 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1343__RN
timestamp 1698431365
transform 1 0 23968 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1344__CLK
timestamp 1698431365
transform 1 0 14112 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1344__RN
timestamp 1698431365
transform 1 0 18144 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1345__CLK
timestamp 1698431365
transform -1 0 16128 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1345__RN
timestamp 1698431365
transform 1 0 16352 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1346__CLK
timestamp 1698431365
transform -1 0 17024 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1346__RN
timestamp 1698431365
transform 1 0 21280 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1347__CLK
timestamp 1698431365
transform 1 0 7168 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1347__RN
timestamp 1698431365
transform 1 0 5040 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1348__CLK
timestamp 1698431365
transform 1 0 5040 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1348__RN
timestamp 1698431365
transform 1 0 5376 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1349__CLK
timestamp 1698431365
transform 1 0 5712 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1349__RN
timestamp 1698431365
transform 1 0 6160 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1351__CLK
timestamp 1698431365
transform 1 0 4704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1351__RN
timestamp 1698431365
transform -1 0 2352 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1352__CLK
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1352__RN
timestamp 1698431365
transform -1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1353__CLK
timestamp 1698431365
transform -1 0 6048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_reg._1353__RN
timestamp 1698431365
transform -1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_sync_rclk._1__CLK
timestamp 1698431365
transform -1 0 26432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_rtc.u_sync_rclk._2__CLK
timestamp 1698431365
transform 1 0 29568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_wire1_I
timestamp 1698431365
transform 1 0 12880 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_mclk open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24528 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_rtc_clk
timestamp 1698431365
transform 1 0 19152 0 -1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_mclk
timestamp 1698431365
transform -1 0 20608 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_mclk
timestamp 1698431365
transform 1 0 22400 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_rtc_clk open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7952 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_rtc_clk
timestamp 1698431365
transform 1 0 11424 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_rtc_clk
timestamp 1698431365
transform -1 0 9184 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_rtc_clk
timestamp 1698431365
transform 1 0 9520 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_rtc_clk
timestamp 1698431365
transform 1 0 21840 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_rtc_clk
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_rtc_clk
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_rtc_clk
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_rtc_clk
timestamp 1698431365
transform 1 0 7056 0 1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_rtc_clk
timestamp 1698431365
transform 1 0 9856 0 1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_rtc_clk
timestamp 1698431365
transform 1 0 7840 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_rtc_clk
timestamp 1698431365
transform 1 0 11760 0 -1 78400
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_rtc_clk
timestamp 1698431365
transform 1 0 23632 0 1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_rtc_clk
timestamp 1698431365
transform 1 0 26880 0 -1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_rtc_clk
timestamp 1698431365
transform 1 0 24416 0 1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_rtc_clk
timestamp 1698431365
transform 1 0 27664 0 -1 72128
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_12  fanout2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8288 0 -1 25088
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout3
timestamp 1698431365
transform 1 0 5824 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout4 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout5
timestamp 1698431365
transform -1 0 8848 0 1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout6
timestamp 1698431365
transform 1 0 19264 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout7
timestamp 1698431365
transform -1 0 28000 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout8
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout9
timestamp 1698431365
transform 1 0 24976 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout10
timestamp 1698431365
transform 1 0 23744 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout11 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29792 0 -1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout12
timestamp 1698431365
transform 1 0 14448 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout13
timestamp 1698431365
transform -1 0 24080 0 1 72128
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout14
timestamp 1698431365
transform 1 0 27328 0 -1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout15
timestamp 1698431365
transform -1 0 28448 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout16
timestamp 1698431365
transform 1 0 25648 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout17
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout18
timestamp 1698431365
transform -1 0 6272 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout19
timestamp 1698431365
transform -1 0 5264 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout20
timestamp 1698431365
transform 1 0 5376 0 -1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout21
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_36 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_42 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_46 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_54
timestamp 1698431365
transform 1 0 7392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_58
timestamp 1698431365
transform 1 0 7840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_60 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_63
timestamp 1698431365
transform 1 0 8400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_133
timestamp 1698431365
transform 1 0 16240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_160
timestamp 1698431365
transform 1 0 19264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_162
timestamp 1698431365
transform 1 0 19488 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_188 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_324
timestamp 1698431365
transform 1 0 37632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698431365
transform 1 0 38080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_330
timestamp 1698431365
transform 1 0 38304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_38
timestamp 1698431365
transform 1 0 5600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_40
timestamp 1698431365
transform 1 0 5824 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_51
timestamp 1698431365
transform 1 0 7056 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_56
timestamp 1698431365
transform 1 0 7616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_58
timestamp 1698431365
transform 1 0 7840 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_231
timestamp 1698431365
transform 1 0 27216 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_263
timestamp 1698431365
transform 1 0 30800 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_330
timestamp 1698431365
transform 1 0 38304 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_46
timestamp 1698431365
transform 1 0 6496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_48
timestamp 1698431365
transform 1 0 6720 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_83
timestamp 1698431365
transform 1 0 10640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_87
timestamp 1698431365
transform 1 0 11088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_91
timestamp 1698431365
transform 1 0 11536 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_99
timestamp 1698431365
transform 1 0 12432 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_103
timestamp 1698431365
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_111
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_115
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_119
timestamp 1698431365
transform 1 0 14672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_121
timestamp 1698431365
transform 1 0 14896 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_172
timestamp 1698431365
transform 1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_183
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_238
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_329
timestamp 1698431365
transform 1 0 38192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_22
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_24
timestamp 1698431365
transform 1 0 4032 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_59
timestamp 1698431365
transform 1 0 7952 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_147
timestamp 1698431365
transform 1 0 17808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_207
timestamp 1698431365
transform 1 0 24528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_246
timestamp 1698431365
transform 1 0 28896 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_278
timestamp 1698431365
transform 1 0 32480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_314
timestamp 1698431365
transform 1 0 36512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_330
timestamp 1698431365
transform 1 0 38304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_6
timestamp 1698431365
transform 1 0 2016 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_53
timestamp 1698431365
transform 1 0 7280 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_61
timestamp 1698431365
transform 1 0 8176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_109
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_126
timestamp 1698431365
transform 1 0 15456 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_134
timestamp 1698431365
transform 1 0 16352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_217
timestamp 1698431365
transform 1 0 25648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_221
timestamp 1698431365
transform 1 0 26096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_225
timestamp 1698431365
transform 1 0 26544 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_242
timestamp 1698431365
transform 1 0 28448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_325
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_329
timestamp 1698431365
transform 1 0 38192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_36
timestamp 1698431365
transform 1 0 5376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_40
timestamp 1698431365
transform 1 0 5824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_51
timestamp 1698431365
transform 1 0 7056 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_67
timestamp 1698431365
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_76
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_80
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_84
timestamp 1698431365
transform 1 0 10752 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_86
timestamp 1698431365
transform 1 0 10976 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_121
timestamp 1698431365
transform 1 0 14896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_125
timestamp 1698431365
transform 1 0 15344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_129
timestamp 1698431365
transform 1 0 15792 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_133
timestamp 1698431365
transform 1 0 16240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_135
timestamp 1698431365
transform 1 0 16464 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_182
timestamp 1698431365
transform 1 0 21728 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_198
timestamp 1698431365
transform 1 0 23520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_237
timestamp 1698431365
transform 1 0 27888 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_269
timestamp 1698431365
transform 1 0 31472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_330
timestamp 1698431365
transform 1 0 38304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_39
timestamp 1698431365
transform 1 0 5712 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_42
timestamp 1698431365
transform 1 0 6048 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_58
timestamp 1698431365
transform 1 0 7840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_61
timestamp 1698431365
transform 1 0 8176 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_93
timestamp 1698431365
transform 1 0 11760 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_185
timestamp 1698431365
transform 1 0 22064 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_220
timestamp 1698431365
transform 1 0 25984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_224
timestamp 1698431365
transform 1 0 26432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_228
timestamp 1698431365
transform 1 0 26880 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_154
timestamp 1698431365
transform 1 0 18592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_160
timestamp 1698431365
transform 1 0 19264 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_196
timestamp 1698431365
transform 1 0 23296 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_204
timestamp 1698431365
transform 1 0 24192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_208
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_250
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_254
timestamp 1698431365
transform 1 0 29792 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_270
timestamp 1698431365
transform 1 0 31584 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_314
timestamp 1698431365
transform 1 0 36512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_330
timestamp 1698431365
transform 1 0 38304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_41
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_72
timestamp 1698431365
transform 1 0 9408 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_209
timestamp 1698431365
transform 1 0 24752 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_225
timestamp 1698431365
transform 1 0 26544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_227
timestamp 1698431365
transform 1 0 26768 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_76
timestamp 1698431365
transform 1 0 9856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_116
timestamp 1698431365
transform 1 0 14336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_120
timestamp 1698431365
transform 1 0 14784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_127
timestamp 1698431365
transform 1 0 15568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_131
timestamp 1698431365
transform 1 0 16016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_196
timestamp 1698431365
transform 1 0 23296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_200
timestamp 1698431365
transform 1 0 23744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_204
timestamp 1698431365
transform 1 0 24192 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_208
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_330
timestamp 1698431365
transform 1 0 38304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_10
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_14
timestamp 1698431365
transform 1 0 2912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_47
timestamp 1698431365
transform 1 0 6608 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_57
timestamp 1698431365
transform 1 0 7728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_93
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_97
timestamp 1698431365
transform 1 0 12208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_141
timestamp 1698431365
transform 1 0 17136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_145
timestamp 1698431365
transform 1 0 17584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_149
timestamp 1698431365
transform 1 0 18032 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_165
timestamp 1698431365
transform 1 0 19824 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_219
timestamp 1698431365
transform 1 0 25872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_223
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_227
timestamp 1698431365
transform 1 0 26768 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_329
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_37
timestamp 1698431365
transform 1 0 5488 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_41
timestamp 1698431365
transform 1 0 5936 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_62
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_76
timestamp 1698431365
transform 1 0 9856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_83
timestamp 1698431365
transform 1 0 10640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_87
timestamp 1698431365
transform 1 0 11088 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_103
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_186
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_190
timestamp 1698431365
transform 1 0 22624 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_238
timestamp 1698431365
transform 1 0 28000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_242
timestamp 1698431365
transform 1 0 28448 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_274
timestamp 1698431365
transform 1 0 32032 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_330
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_10
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_29
timestamp 1698431365
transform 1 0 4592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_33
timestamp 1698431365
transform 1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_41
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_45
timestamp 1698431365
transform 1 0 6384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_47
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_58
timestamp 1698431365
transform 1 0 7840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_60
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_71
timestamp 1698431365
transform 1 0 9296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_75
timestamp 1698431365
transform 1 0 9744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_79
timestamp 1698431365
transform 1 0 10192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_82
timestamp 1698431365
transform 1 0 10528 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_92
timestamp 1698431365
transform 1 0 11648 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_100
timestamp 1698431365
transform 1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_131
timestamp 1698431365
transform 1 0 16016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_167
timestamp 1698431365
transform 1 0 20048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_209
timestamp 1698431365
transform 1 0 24752 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_213
timestamp 1698431365
transform 1 0 25200 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_215
timestamp 1698431365
transform 1 0 25424 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_329
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_36
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_52
timestamp 1698431365
transform 1 0 7168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_56
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_63
timestamp 1698431365
transform 1 0 8400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_92
timestamp 1698431365
transform 1 0 11648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_96
timestamp 1698431365
transform 1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_100
timestamp 1698431365
transform 1 0 12544 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698431365
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698431365
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_123
timestamp 1698431365
transform 1 0 15120 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_133
timestamp 1698431365
transform 1 0 16240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_157
timestamp 1698431365
transform 1 0 18928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_165
timestamp 1698431365
transform 1 0 19824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_167
timestamp 1698431365
transform 1 0 20048 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_185
timestamp 1698431365
transform 1 0 22064 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_201
timestamp 1698431365
transform 1 0 23856 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_230
timestamp 1698431365
transform 1 0 27104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_234
timestamp 1698431365
transform 1 0 27552 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_266
timestamp 1698431365
transform 1 0 31136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_330
timestamp 1698431365
transform 1 0 38304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_41
timestamp 1698431365
transform 1 0 5936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_59
timestamp 1698431365
transform 1 0 7952 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_72
timestamp 1698431365
transform 1 0 9408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_84
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_92
timestamp 1698431365
transform 1 0 11648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_96
timestamp 1698431365
transform 1 0 12096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_100
timestamp 1698431365
transform 1 0 12544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_119
timestamp 1698431365
transform 1 0 14672 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_125
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_141
timestamp 1698431365
transform 1 0 17136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_147
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_151
timestamp 1698431365
transform 1 0 18256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_183
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_186
timestamp 1698431365
transform 1 0 22176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_190
timestamp 1698431365
transform 1 0 22624 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_198
timestamp 1698431365
transform 1 0 23520 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_200
timestamp 1698431365
transform 1 0 23744 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_235
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_329
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_36
timestamp 1698431365
transform 1 0 5376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_43
timestamp 1698431365
transform 1 0 6160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_47
timestamp 1698431365
transform 1 0 6608 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698431365
transform 1 0 10752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_88
timestamp 1698431365
transform 1 0 11200 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_109
timestamp 1698431365
transform 1 0 13552 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_111
timestamp 1698431365
transform 1 0 13776 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_114
timestamp 1698431365
transform 1 0 14112 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_118
timestamp 1698431365
transform 1 0 14560 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_134
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_152
timestamp 1698431365
transform 1 0 18368 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_187
timestamp 1698431365
transform 1 0 22288 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698431365
transform 1 0 24080 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698431365
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_250
timestamp 1698431365
transform 1 0 29344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_254
timestamp 1698431365
transform 1 0 29792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_258
timestamp 1698431365
transform 1 0 30240 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698431365
transform 1 0 32032 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_6
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_10
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_12
timestamp 1698431365
transform 1 0 2688 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_85
timestamp 1698431365
transform 1 0 10864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_89
timestamp 1698431365
transform 1 0 11312 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_116
timestamp 1698431365
transform 1 0 14336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_120
timestamp 1698431365
transform 1 0 14784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_124
timestamp 1698431365
transform 1 0 15232 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_140
timestamp 1698431365
transform 1 0 17024 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_143
timestamp 1698431365
transform 1 0 17360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_147
timestamp 1698431365
transform 1 0 17808 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_163
timestamp 1698431365
transform 1 0 19600 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_179
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_184
timestamp 1698431365
transform 1 0 21952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_188
timestamp 1698431365
transform 1 0 22400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_192
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_251
timestamp 1698431365
transform 1 0 29456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_267
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_299
timestamp 1698431365
transform 1 0 34832 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_33
timestamp 1698431365
transform 1 0 5040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_37
timestamp 1698431365
transform 1 0 5488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_41
timestamp 1698431365
transform 1 0 5936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_45
timestamp 1698431365
transform 1 0 6384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_47
timestamp 1698431365
transform 1 0 6608 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_131
timestamp 1698431365
transform 1 0 16016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_133
timestamp 1698431365
transform 1 0 16240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_147
timestamp 1698431365
transform 1 0 17808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_151
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_155
timestamp 1698431365
transform 1 0 18704 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_159
timestamp 1698431365
transform 1 0 19152 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_172
timestamp 1698431365
transform 1 0 20608 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_180
timestamp 1698431365
transform 1 0 21504 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_184
timestamp 1698431365
transform 1 0 21952 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_192
timestamp 1698431365
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_225
timestamp 1698431365
transform 1 0 26544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_229
timestamp 1698431365
transform 1 0 26992 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_261
timestamp 1698431365
transform 1 0 30576 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_330
timestamp 1698431365
transform 1 0 38304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_71
timestamp 1698431365
transform 1 0 9296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_75
timestamp 1698431365
transform 1 0 9744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_79
timestamp 1698431365
transform 1 0 10192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_88
timestamp 1698431365
transform 1 0 11200 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_158
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_208
timestamp 1698431365
transform 1 0 24640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_212
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_228
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_329
timestamp 1698431365
transform 1 0 38192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_50
timestamp 1698431365
transform 1 0 6944 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_92
timestamp 1698431365
transform 1 0 11648 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_99
timestamp 1698431365
transform 1 0 12432 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_197
timestamp 1698431365
transform 1 0 23408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_224
timestamp 1698431365
transform 1 0 26432 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_228
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_234
timestamp 1698431365
transform 1 0 27552 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_238
timestamp 1698431365
transform 1 0 28000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_255
timestamp 1698431365
transform 1 0 29904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_259
timestamp 1698431365
transform 1 0 30352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_263
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_330
timestamp 1698431365
transform 1 0 38304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_24
timestamp 1698431365
transform 1 0 4032 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698431365
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_113
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_124
timestamp 1698431365
transform 1 0 15232 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_140
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_143
timestamp 1698431365
transform 1 0 17360 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_151
timestamp 1698431365
transform 1 0 18256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_193
timestamp 1698431365
transform 1 0 22960 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_201
timestamp 1698431365
transform 1 0 23856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_203
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_206
timestamp 1698431365
transform 1 0 24416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_283
timestamp 1698431365
transform 1 0 33040 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_329
timestamp 1698431365
transform 1 0 38192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_28
timestamp 1698431365
transform 1 0 4480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_36
timestamp 1698431365
transform 1 0 5376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_38
timestamp 1698431365
transform 1 0 5600 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_41
timestamp 1698431365
transform 1 0 5936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_45
timestamp 1698431365
transform 1 0 6384 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_61
timestamp 1698431365
transform 1 0 8176 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_74
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_85
timestamp 1698431365
transform 1 0 10864 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_89
timestamp 1698431365
transform 1 0 11312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_103
timestamp 1698431365
transform 1 0 12880 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_107
timestamp 1698431365
transform 1 0 13328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_109
timestamp 1698431365
transform 1 0 13552 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_118
timestamp 1698431365
transform 1 0 14560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_122
timestamp 1698431365
transform 1 0 15008 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_158
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_190
timestamp 1698431365
transform 1 0 22624 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_194
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_267
timestamp 1698431365
transform 1 0 31248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_271
timestamp 1698431365
transform 1 0 31696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698431365
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_330
timestamp 1698431365
transform 1 0 38304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_6
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_18
timestamp 1698431365
transform 1 0 3360 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_46
timestamp 1698431365
transform 1 0 6496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_50
timestamp 1698431365
transform 1 0 6944 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_58
timestamp 1698431365
transform 1 0 7840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_64
timestamp 1698431365
transform 1 0 8512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_99
timestamp 1698431365
transform 1 0 12432 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_112
timestamp 1698431365
transform 1 0 13888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_116
timestamp 1698431365
transform 1 0 14336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_120
timestamp 1698431365
transform 1 0 14784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_122
timestamp 1698431365
transform 1 0 15008 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_125
timestamp 1698431365
transform 1 0 15344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_129
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_161
timestamp 1698431365
transform 1 0 19376 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_196
timestamp 1698431365
transform 1 0 23296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_198
timestamp 1698431365
transform 1 0 23520 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_204
timestamp 1698431365
transform 1 0 24192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_252
timestamp 1698431365
transform 1 0 29568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_294
timestamp 1698431365
transform 1 0 34272 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_310
timestamp 1698431365
transform 1 0 36064 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_37
timestamp 1698431365
transform 1 0 5488 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_53
timestamp 1698431365
transform 1 0 7280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_57
timestamp 1698431365
transform 1 0 7728 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_61
timestamp 1698431365
transform 1 0 8176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_108
timestamp 1698431365
transform 1 0 13440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_112
timestamp 1698431365
transform 1 0 13888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_116
timestamp 1698431365
transform 1 0 14336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_146
timestamp 1698431365
transform 1 0 17696 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_162
timestamp 1698431365
transform 1 0 19488 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_170
timestamp 1698431365
transform 1 0 20384 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_174
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_270
timestamp 1698431365
transform 1 0 31584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698431365
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_71
timestamp 1698431365
transform 1 0 9296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_75
timestamp 1698431365
transform 1 0 9744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_79
timestamp 1698431365
transform 1 0 10192 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_83
timestamp 1698431365
transform 1 0 10640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_85
timestamp 1698431365
transform 1 0 10864 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_122
timestamp 1698431365
transform 1 0 15008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_124
timestamp 1698431365
transform 1 0 15232 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_159
timestamp 1698431365
transform 1 0 19152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_163
timestamp 1698431365
transform 1 0 19600 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_167
timestamp 1698431365
transform 1 0 20048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_192
timestamp 1698431365
transform 1 0 22848 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_253
timestamp 1698431365
transform 1 0 29680 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_262
timestamp 1698431365
transform 1 0 30688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_266
timestamp 1698431365
transform 1 0 31136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_270
timestamp 1698431365
transform 1 0 31584 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_302
timestamp 1698431365
transform 1 0 35168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_310
timestamp 1698431365
transform 1 0 36064 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_30
timestamp 1698431365
transform 1 0 4704 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_84
timestamp 1698431365
transform 1 0 10752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_119
timestamp 1698431365
transform 1 0 14672 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698431365
transform 1 0 17920 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_216
timestamp 1698431365
transform 1 0 25536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_218
timestamp 1698431365
transform 1 0 25760 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_231
timestamp 1698431365
transform 1 0 27216 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_233
timestamp 1698431365
transform 1 0 27440 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_268
timestamp 1698431365
transform 1 0 31360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_272
timestamp 1698431365
transform 1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_330
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_30
timestamp 1698431365
transform 1 0 4704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_39
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_95
timestamp 1698431365
transform 1 0 11984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_99
timestamp 1698431365
transform 1 0 12432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_103
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_141
timestamp 1698431365
transform 1 0 17136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_145
timestamp 1698431365
transform 1 0 17584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_149
timestamp 1698431365
transform 1 0 18032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_153
timestamp 1698431365
transform 1 0 18480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_155
timestamp 1698431365
transform 1 0 18704 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_195
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_240
timestamp 1698431365
transform 1 0 28224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_267
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_271
timestamp 1698431365
transform 1 0 31696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_275
timestamp 1698431365
transform 1 0 32144 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_307
timestamp 1698431365
transform 1 0 35728 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_6
timestamp 1698431365
transform 1 0 2016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_18
timestamp 1698431365
transform 1 0 3360 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_62
timestamp 1698431365
transform 1 0 8288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_87
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_89
timestamp 1698431365
transform 1 0 11312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_92
timestamp 1698431365
transform 1 0 11648 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_102
timestamp 1698431365
transform 1 0 12768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_121
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_150
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_153
timestamp 1698431365
transform 1 0 18480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_172
timestamp 1698431365
transform 1 0 20608 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_240
timestamp 1698431365
transform 1 0 28224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_262
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_266
timestamp 1698431365
transform 1 0 31136 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_270
timestamp 1698431365
transform 1 0 31584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_330
timestamp 1698431365
transform 1 0 38304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_22
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_24
timestamp 1698431365
transform 1 0 4032 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_27
timestamp 1698431365
transform 1 0 4368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_51
timestamp 1698431365
transform 1 0 7056 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_55
timestamp 1698431365
transform 1 0 7504 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_58
timestamp 1698431365
transform 1 0 7840 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_62
timestamp 1698431365
transform 1 0 8288 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_87
timestamp 1698431365
transform 1 0 11088 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_111
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_120
timestamp 1698431365
transform 1 0 14784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_124
timestamp 1698431365
transform 1 0 15232 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_156
timestamp 1698431365
transform 1 0 18816 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_181
timestamp 1698431365
transform 1 0 21616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698431365
transform 1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_199
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_234
timestamp 1698431365
transform 1 0 27552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_259
timestamp 1698431365
transform 1 0 30352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_300
timestamp 1698431365
transform 1 0 34944 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698431365
transform 1 0 35840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698431365
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_329
timestamp 1698431365
transform 1 0 38192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_20
timestamp 1698431365
transform 1 0 3584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_24
timestamp 1698431365
transform 1 0 4032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_54
timestamp 1698431365
transform 1 0 7392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_56
timestamp 1698431365
transform 1 0 7616 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_59
timestamp 1698431365
transform 1 0 7952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_63
timestamp 1698431365
transform 1 0 8400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_148
timestamp 1698431365
transform 1 0 17920 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_198
timestamp 1698431365
transform 1 0 23520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_202
timestamp 1698431365
transform 1 0 23968 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_227
timestamp 1698431365
transform 1 0 26768 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_243
timestamp 1698431365
transform 1 0 28560 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_247
timestamp 1698431365
transform 1 0 29008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_251
timestamp 1698431365
transform 1 0 29456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_270
timestamp 1698431365
transform 1 0 31584 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_330
timestamp 1698431365
transform 1 0 38304 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_8
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_12
timestamp 1698431365
transform 1 0 2688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_16
timestamp 1698431365
transform 1 0 3136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_56
timestamp 1698431365
transform 1 0 7616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_58
timestamp 1698431365
transform 1 0 7840 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_68
timestamp 1698431365
transform 1 0 8960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_70
timestamp 1698431365
transform 1 0 9184 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_73
timestamp 1698431365
transform 1 0 9520 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_77
timestamp 1698431365
transform 1 0 9968 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_93
timestamp 1698431365
transform 1 0 11760 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698431365
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_115
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_121
timestamp 1698431365
transform 1 0 14896 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_125
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_133
timestamp 1698431365
transform 1 0 16240 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_137
timestamp 1698431365
transform 1 0 16688 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_140
timestamp 1698431365
transform 1 0 17024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_144
timestamp 1698431365
transform 1 0 17472 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_152
timestamp 1698431365
transform 1 0 18368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698431365
transform 1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_183
timestamp 1698431365
transform 1 0 21840 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_218
timestamp 1698431365
transform 1 0 25760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_222
timestamp 1698431365
transform 1 0 26208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_226
timestamp 1698431365
transform 1 0 26656 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_293
timestamp 1698431365
transform 1 0 34160 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_309
timestamp 1698431365
transform 1 0 35952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_329
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_81
timestamp 1698431365
transform 1 0 10416 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_89
timestamp 1698431365
transform 1 0 11312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_108
timestamp 1698431365
transform 1 0 13440 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_119
timestamp 1698431365
transform 1 0 14672 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_123
timestamp 1698431365
transform 1 0 15120 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_131
timestamp 1698431365
transform 1 0 16016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_133
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_154
timestamp 1698431365
transform 1 0 18592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698431365
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_216
timestamp 1698431365
transform 1 0 25536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_252
timestamp 1698431365
transform 1 0 29568 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_272
timestamp 1698431365
transform 1 0 31808 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_6
timestamp 1698431365
transform 1 0 2016 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_21
timestamp 1698431365
transform 1 0 3696 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_158
timestamp 1698431365
transform 1 0 19040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_162
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_179
timestamp 1698431365
transform 1 0 21392 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_182
timestamp 1698431365
transform 1 0 21728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_186
timestamp 1698431365
transform 1 0 22176 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_203
timestamp 1698431365
transform 1 0 24080 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_237
timestamp 1698431365
transform 1 0 27888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_42
timestamp 1698431365
transform 1 0 6048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_82
timestamp 1698431365
transform 1 0 10528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_86
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_138
timestamp 1698431365
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_176
timestamp 1698431365
transform 1 0 21056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_180
timestamp 1698431365
transform 1 0 21504 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_184
timestamp 1698431365
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_186
timestamp 1698431365
transform 1 0 22176 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_204
timestamp 1698431365
transform 1 0 24192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_224
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_262
timestamp 1698431365
transform 1 0 30688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_266
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_272
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_292
timestamp 1698431365
transform 1 0 34048 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_324
timestamp 1698431365
transform 1 0 37632 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_328
timestamp 1698431365
transform 1 0 38080 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_330
timestamp 1698431365
transform 1 0 38304 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_8
timestamp 1698431365
transform 1 0 2240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_18
timestamp 1698431365
transform 1 0 3360 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_33
timestamp 1698431365
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_49
timestamp 1698431365
transform 1 0 6832 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_102
timestamp 1698431365
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_181
timestamp 1698431365
transform 1 0 21616 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_213
timestamp 1698431365
transform 1 0 25200 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_238
timestamp 1698431365
transform 1 0 28000 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_262
timestamp 1698431365
transform 1 0 30688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_266
timestamp 1698431365
transform 1 0 31136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_270
timestamp 1698431365
transform 1 0 31584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_329
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_8
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_76
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_92
timestamp 1698431365
transform 1 0 11648 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_100
timestamp 1698431365
transform 1 0 12544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_104
timestamp 1698431365
transform 1 0 12992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_106
timestamp 1698431365
transform 1 0 13216 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_109
timestamp 1698431365
transform 1 0 13552 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_113
timestamp 1698431365
transform 1 0 14000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_117
timestamp 1698431365
transform 1 0 14448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_121
timestamp 1698431365
transform 1 0 14896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_130
timestamp 1698431365
transform 1 0 15904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_132
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_135
timestamp 1698431365
transform 1 0 16464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_153
timestamp 1698431365
transform 1 0 18480 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_185
timestamp 1698431365
transform 1 0 22064 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_201
timestamp 1698431365
transform 1 0 23856 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_248
timestamp 1698431365
transform 1 0 29120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_252
timestamp 1698431365
transform 1 0 29568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_256
timestamp 1698431365
transform 1 0 30016 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_272
timestamp 1698431365
transform 1 0 31808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_318
timestamp 1698431365
transform 1 0 36960 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_326
timestamp 1698431365
transform 1 0 37856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_330
timestamp 1698431365
transform 1 0 38304 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_12
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_16
timestamp 1698431365
transform 1 0 3136 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_18
timestamp 1698431365
transform 1 0 3360 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_51
timestamp 1698431365
transform 1 0 7056 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_55
timestamp 1698431365
transform 1 0 7504 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_65
timestamp 1698431365
transform 1 0 8624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_99
timestamp 1698431365
transform 1 0 12432 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_109
timestamp 1698431365
transform 1 0 13552 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_112
timestamp 1698431365
transform 1 0 13888 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_131
timestamp 1698431365
transform 1 0 16016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_135
timestamp 1698431365
transform 1 0 16464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_157
timestamp 1698431365
transform 1 0 18928 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_206
timestamp 1698431365
transform 1 0 24416 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_214
timestamp 1698431365
transform 1 0 25312 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_217
timestamp 1698431365
transform 1 0 25648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_226
timestamp 1698431365
transform 1 0 26656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_253
timestamp 1698431365
transform 1 0 29680 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_275
timestamp 1698431365
transform 1 0 32144 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_309
timestamp 1698431365
transform 1 0 35952 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_329
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_18
timestamp 1698431365
transform 1 0 3360 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_26
timestamp 1698431365
transform 1 0 4256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_32
timestamp 1698431365
transform 1 0 4928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_36
timestamp 1698431365
transform 1 0 5376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_40
timestamp 1698431365
transform 1 0 5824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_42
timestamp 1698431365
transform 1 0 6048 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_50
timestamp 1698431365
transform 1 0 6944 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_54
timestamp 1698431365
transform 1 0 7392 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_57
timestamp 1698431365
transform 1 0 7728 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_61
timestamp 1698431365
transform 1 0 8176 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_92
timestamp 1698431365
transform 1 0 11648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_94
timestamp 1698431365
transform 1 0 11872 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_131
timestamp 1698431365
transform 1 0 16016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_135
timestamp 1698431365
transform 1 0 16464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_144
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_147
timestamp 1698431365
transform 1 0 17808 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_151
timestamp 1698431365
transform 1 0 18256 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_167
timestamp 1698431365
transform 1 0 20048 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_175
timestamp 1698431365
transform 1 0 20944 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_216
timestamp 1698431365
transform 1 0 25536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_239
timestamp 1698431365
transform 1 0 28112 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_255
timestamp 1698431365
transform 1 0 29904 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_270
timestamp 1698431365
transform 1 0 31584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_326
timestamp 1698431365
transform 1 0 37856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_330
timestamp 1698431365
transform 1 0 38304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_18
timestamp 1698431365
transform 1 0 3360 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_22
timestamp 1698431365
transform 1 0 3808 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_24
timestamp 1698431365
transform 1 0 4032 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_27
timestamp 1698431365
transform 1 0 4368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_31
timestamp 1698431365
transform 1 0 4816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_52
timestamp 1698431365
transform 1 0 7168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_54
timestamp 1698431365
transform 1 0 7392 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_89
timestamp 1698431365
transform 1 0 11312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_93
timestamp 1698431365
transform 1 0 11760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_97
timestamp 1698431365
transform 1 0 12208 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_122
timestamp 1698431365
transform 1 0 15008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_137
timestamp 1698431365
transform 1 0 16688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_151
timestamp 1698431365
transform 1 0 18256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_155
timestamp 1698431365
transform 1 0 18704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_159
timestamp 1698431365
transform 1 0 19152 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_187
timestamp 1698431365
transform 1 0 22288 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_190
timestamp 1698431365
transform 1 0 22624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_194
timestamp 1698431365
transform 1 0 23072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_211
timestamp 1698431365
transform 1 0 24976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_215
timestamp 1698431365
transform 1 0 25424 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_219
timestamp 1698431365
transform 1 0 25872 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_221
timestamp 1698431365
transform 1 0 26096 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_224
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_240
timestamp 1698431365
transform 1 0 28224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_253
timestamp 1698431365
transform 1 0 29680 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_256
timestamp 1698431365
transform 1 0 30016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_260
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_274
timestamp 1698431365
transform 1 0 32032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_278
timestamp 1698431365
transform 1 0 32480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_282
timestamp 1698431365
transform 1 0 32928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_284
timestamp 1698431365
transform 1 0 33152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_296
timestamp 1698431365
transform 1 0 34496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_329
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_56
timestamp 1698431365
transform 1 0 7616 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_84
timestamp 1698431365
transform 1 0 10752 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_90
timestamp 1698431365
transform 1 0 11424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_94
timestamp 1698431365
transform 1 0 11872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_98
timestamp 1698431365
transform 1 0 12320 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_102
timestamp 1698431365
transform 1 0 12768 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_105
timestamp 1698431365
transform 1 0 13104 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_121
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_131
timestamp 1698431365
transform 1 0 16016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_180
timestamp 1698431365
transform 1 0 21504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_184
timestamp 1698431365
transform 1 0 21952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_188
timestamp 1698431365
transform 1 0 22400 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_204
timestamp 1698431365
transform 1 0 24192 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_216
timestamp 1698431365
transform 1 0 25536 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_254
timestamp 1698431365
transform 1 0 29792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_273
timestamp 1698431365
transform 1 0 31920 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_320
timestamp 1698431365
transform 1 0 37184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_324
timestamp 1698431365
transform 1 0 37632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_328
timestamp 1698431365
transform 1 0 38080 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_330
timestamp 1698431365
transform 1 0 38304 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_4
timestamp 1698431365
transform 1 0 1792 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_46
timestamp 1698431365
transform 1 0 6496 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_89
timestamp 1698431365
transform 1 0 11312 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_112
timestamp 1698431365
transform 1 0 13888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_116
timestamp 1698431365
transform 1 0 14336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_120
timestamp 1698431365
transform 1 0 14784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_124
timestamp 1698431365
transform 1 0 15232 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_132
timestamp 1698431365
transform 1 0 16128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_136
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_151
timestamp 1698431365
transform 1 0 18256 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_155
timestamp 1698431365
transform 1 0 18704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_157
timestamp 1698431365
transform 1 0 18928 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_189
timestamp 1698431365
transform 1 0 22512 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_191
timestamp 1698431365
transform 1 0 22736 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_226
timestamp 1698431365
transform 1 0 26656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_230
timestamp 1698431365
transform 1 0 27104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_234
timestamp 1698431365
transform 1 0 27552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_238
timestamp 1698431365
transform 1 0 28000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_242
timestamp 1698431365
transform 1 0 28448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_253
timestamp 1698431365
transform 1 0 29680 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_256
timestamp 1698431365
transform 1 0 30016 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_272
timestamp 1698431365
transform 1 0 31808 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_295
timestamp 1698431365
transform 1 0 34384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_328
timestamp 1698431365
transform 1 0 38080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_330
timestamp 1698431365
transform 1 0 38304 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_38
timestamp 1698431365
transform 1 0 5600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_42
timestamp 1698431365
transform 1 0 6048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_46
timestamp 1698431365
transform 1 0 6496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_50
timestamp 1698431365
transform 1 0 6944 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_53
timestamp 1698431365
transform 1 0 7280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_55
timestamp 1698431365
transform 1 0 7504 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_82
timestamp 1698431365
transform 1 0 10528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_158
timestamp 1698431365
transform 1 0 19040 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_193
timestamp 1698431365
transform 1 0 22960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_197
timestamp 1698431365
transform 1 0 23408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_201
timestamp 1698431365
transform 1 0 23856 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_204
timestamp 1698431365
transform 1 0 24192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_227
timestamp 1698431365
transform 1 0 26768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_244
timestamp 1698431365
transform 1 0 28672 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_260
timestamp 1698431365
transform 1 0 30464 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_268
timestamp 1698431365
transform 1 0 31360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_270
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_305
timestamp 1698431365
transform 1 0 35504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_18
timestamp 1698431365
transform 1 0 3360 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_22
timestamp 1698431365
transform 1 0 3808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_26
timestamp 1698431365
transform 1 0 4256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_57
timestamp 1698431365
transform 1 0 7728 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_61
timestamp 1698431365
transform 1 0 8176 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_83
timestamp 1698431365
transform 1 0 10640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_87
timestamp 1698431365
transform 1 0 11088 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_91
timestamp 1698431365
transform 1 0 11536 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_93
timestamp 1698431365
transform 1 0 11760 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_96
timestamp 1698431365
transform 1 0 12096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_98
timestamp 1698431365
transform 1 0 12320 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_117
timestamp 1698431365
transform 1 0 14448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_119
timestamp 1698431365
transform 1 0 14672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_122
timestamp 1698431365
transform 1 0 15008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_154
timestamp 1698431365
transform 1 0 18592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_158
timestamp 1698431365
transform 1 0 19040 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_203
timestamp 1698431365
transform 1 0 24080 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_255
timestamp 1698431365
transform 1 0 29904 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_261
timestamp 1698431365
transform 1 0 30576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_281
timestamp 1698431365
transform 1 0 32816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_297
timestamp 1698431365
transform 1 0 34608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_299
timestamp 1698431365
transform 1 0 34832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_18
timestamp 1698431365
transform 1 0 3360 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_50
timestamp 1698431365
transform 1 0 6944 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_58
timestamp 1698431365
transform 1 0 7840 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_62
timestamp 1698431365
transform 1 0 8288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_64
timestamp 1698431365
transform 1 0 8512 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_85
timestamp 1698431365
transform 1 0 10864 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_89
timestamp 1698431365
transform 1 0 11312 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_92
timestamp 1698431365
transform 1 0 11648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_126
timestamp 1698431365
transform 1 0 15456 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_130
timestamp 1698431365
transform 1 0 15904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_150
timestamp 1698431365
transform 1 0 18144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_186
timestamp 1698431365
transform 1 0 22176 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_190
timestamp 1698431365
transform 1 0 22624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_194
timestamp 1698431365
transform 1 0 23072 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_202
timestamp 1698431365
transform 1 0 23968 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_205
timestamp 1698431365
transform 1 0 24304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_207
timestamp 1698431365
transform 1 0 24528 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_227
timestamp 1698431365
transform 1 0 26768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_61
timestamp 1698431365
transform 1 0 8176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_65
timestamp 1698431365
transform 1 0 8624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_78
timestamp 1698431365
transform 1 0 10080 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_86
timestamp 1698431365
transform 1 0 10976 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_90
timestamp 1698431365
transform 1 0 11424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_94
timestamp 1698431365
transform 1 0 11872 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_102
timestamp 1698431365
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_119
timestamp 1698431365
transform 1 0 14672 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_121
timestamp 1698431365
transform 1 0 14896 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_156
timestamp 1698431365
transform 1 0 18816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_209
timestamp 1698431365
transform 1 0 24752 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_212
timestamp 1698431365
transform 1 0 25088 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_220
timestamp 1698431365
transform 1 0 25984 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_224
timestamp 1698431365
transform 1 0 26432 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_228
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_238
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_242
timestamp 1698431365
transform 1 0 28448 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_263
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_329
timestamp 1698431365
transform 1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_18
timestamp 1698431365
transform 1 0 3360 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_26
timestamp 1698431365
transform 1 0 4256 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_61
timestamp 1698431365
transform 1 0 8176 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_67
timestamp 1698431365
transform 1 0 8848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_124
timestamp 1698431365
transform 1 0 15232 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_128
timestamp 1698431365
transform 1 0 15680 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_154
timestamp 1698431365
transform 1 0 18592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_160
timestamp 1698431365
transform 1 0 19264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_164
timestamp 1698431365
transform 1 0 19712 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_180
timestamp 1698431365
transform 1 0 21504 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_205
timestamp 1698431365
transform 1 0 24304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_209
timestamp 1698431365
transform 1 0 24752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_244
timestamp 1698431365
transform 1 0 28672 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_260
timestamp 1698431365
transform 1 0 30464 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_268
timestamp 1698431365
transform 1 0 31360 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_272
timestamp 1698431365
transform 1 0 31808 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_274
timestamp 1698431365
transform 1 0 32032 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_6
timestamp 1698431365
transform 1 0 2016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_8
timestamp 1698431365
transform 1 0 2240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_41
timestamp 1698431365
transform 1 0 5936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_45
timestamp 1698431365
transform 1 0 6384 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_63
timestamp 1698431365
transform 1 0 8400 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_67
timestamp 1698431365
transform 1 0 8848 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_79
timestamp 1698431365
transform 1 0 10192 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_83
timestamp 1698431365
transform 1 0 10640 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_86
timestamp 1698431365
transform 1 0 10976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_90
timestamp 1698431365
transform 1 0 11424 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_98
timestamp 1698431365
transform 1 0 12320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_102
timestamp 1698431365
transform 1 0 12768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698431365
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_119
timestamp 1698431365
transform 1 0 14672 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_157
timestamp 1698431365
transform 1 0 18928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_161
timestamp 1698431365
transform 1 0 19376 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_165
timestamp 1698431365
transform 1 0 19824 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_173
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_215
timestamp 1698431365
transform 1 0 25424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_219
timestamp 1698431365
transform 1 0 25872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_223
timestamp 1698431365
transform 1 0 26320 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_239
timestamp 1698431365
transform 1 0 28112 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_243
timestamp 1698431365
transform 1 0 28560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_267
timestamp 1698431365
transform 1 0 31248 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_36
timestamp 1698431365
transform 1 0 5376 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_52
timestamp 1698431365
transform 1 0 7168 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_56
timestamp 1698431365
transform 1 0 7616 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_60
timestamp 1698431365
transform 1 0 8064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_64
timestamp 1698431365
transform 1 0 8512 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_68
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_84
timestamp 1698431365
transform 1 0 10752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_124
timestamp 1698431365
transform 1 0 15232 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_128
timestamp 1698431365
transform 1 0 15680 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_132
timestamp 1698431365
transform 1 0 16128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_174
timestamp 1698431365
transform 1 0 20832 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_182
timestamp 1698431365
transform 1 0 21728 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_203
timestamp 1698431365
transform 1 0 24080 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1698431365
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_218
timestamp 1698431365
transform 1 0 25760 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_259
timestamp 1698431365
transform 1 0 30352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_263
timestamp 1698431365
transform 1 0 30800 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_20
timestamp 1698431365
transform 1 0 3584 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_28
timestamp 1698431365
transform 1 0 4480 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_32
timestamp 1698431365
transform 1 0 4928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_41
timestamp 1698431365
transform 1 0 5936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_45
timestamp 1698431365
transform 1 0 6384 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_53
timestamp 1698431365
transform 1 0 7280 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_79
timestamp 1698431365
transform 1 0 10192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_103
timestamp 1698431365
transform 1 0 12880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_139
timestamp 1698431365
transform 1 0 16912 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_147
timestamp 1698431365
transform 1 0 17808 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_153
timestamp 1698431365
transform 1 0 18480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_157
timestamp 1698431365
transform 1 0 18928 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_196
timestamp 1698431365
transform 1 0 23296 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_200
timestamp 1698431365
transform 1 0 23744 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_251
timestamp 1698431365
transform 1 0 29456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_255
timestamp 1698431365
transform 1 0 29904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_257
timestamp 1698431365
transform 1 0 30128 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_330
timestamp 1698431365
transform 1 0 38304 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_34
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_50
timestamp 1698431365
transform 1 0 6944 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_54
timestamp 1698431365
transform 1 0 7392 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_62
timestamp 1698431365
transform 1 0 8288 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_109
timestamp 1698431365
transform 1 0 13552 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_113
timestamp 1698431365
transform 1 0 14000 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_129
timestamp 1698431365
transform 1 0 15792 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_137
timestamp 1698431365
transform 1 0 16688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_144
timestamp 1698431365
transform 1 0 17472 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_149
timestamp 1698431365
transform 1 0 18032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_151
timestamp 1698431365
transform 1 0 18256 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_154
timestamp 1698431365
transform 1 0 18592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_160
timestamp 1698431365
transform 1 0 19264 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_164
timestamp 1698431365
transform 1 0 19712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_168
timestamp 1698431365
transform 1 0 20160 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_207
timestamp 1698431365
transform 1 0 24528 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_263
timestamp 1698431365
transform 1 0 30800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_330
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_18
timestamp 1698431365
transform 1 0 3360 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_26
timestamp 1698431365
transform 1 0 4256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_30
timestamp 1698431365
transform 1 0 4704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_32
timestamp 1698431365
transform 1 0 4928 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_52
timestamp 1698431365
transform 1 0 7168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_56
timestamp 1698431365
transform 1 0 7616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_60
timestamp 1698431365
transform 1 0 8064 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_75
timestamp 1698431365
transform 1 0 9744 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_85
timestamp 1698431365
transform 1 0 10864 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_98
timestamp 1698431365
transform 1 0 12320 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_102
timestamp 1698431365
transform 1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_111
timestamp 1698431365
transform 1 0 13776 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_115
timestamp 1698431365
transform 1 0 14224 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_123
timestamp 1698431365
transform 1 0 15120 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_127
timestamp 1698431365
transform 1 0 15568 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_129
timestamp 1698431365
transform 1 0 15792 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_166
timestamp 1698431365
transform 1 0 19936 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_170
timestamp 1698431365
transform 1 0 20384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_192
timestamp 1698431365
transform 1 0 22848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_200
timestamp 1698431365
transform 1 0 23744 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_204
timestamp 1698431365
transform 1 0 24192 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_206
timestamp 1698431365
transform 1 0 24416 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_209
timestamp 1698431365
transform 1 0 24752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_213
timestamp 1698431365
transform 1 0 25200 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_221
timestamp 1698431365
transform 1 0 26096 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_232
timestamp 1698431365
transform 1 0 27328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_236
timestamp 1698431365
transform 1 0 27776 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_322
timestamp 1698431365
transform 1 0 37408 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_329
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_36
timestamp 1698431365
transform 1 0 5376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_40
timestamp 1698431365
transform 1 0 5824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_44
timestamp 1698431365
transform 1 0 6272 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_48
timestamp 1698431365
transform 1 0 6720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_52
timestamp 1698431365
transform 1 0 7168 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_60
timestamp 1698431365
transform 1 0 8064 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_76
timestamp 1698431365
transform 1 0 9856 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_79
timestamp 1698431365
transform 1 0 10192 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_104
timestamp 1698431365
transform 1 0 12992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_106
timestamp 1698431365
transform 1 0 13216 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_109
timestamp 1698431365
transform 1 0 13552 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_118
timestamp 1698431365
transform 1 0 14560 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_122
timestamp 1698431365
transform 1 0 15008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_124
timestamp 1698431365
transform 1 0 15232 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_127
timestamp 1698431365
transform 1 0 15568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_168
timestamp 1698431365
transform 1 0 20160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_172
timestamp 1698431365
transform 1 0 20608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_174
timestamp 1698431365
transform 1 0 20832 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_177
timestamp 1698431365
transform 1 0 21168 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_181
timestamp 1698431365
transform 1 0 21616 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_197
timestamp 1698431365
transform 1 0 23408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_205
timestamp 1698431365
transform 1 0 24304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_220
timestamp 1698431365
transform 1 0 25984 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_224
timestamp 1698431365
transform 1 0 26432 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_226
timestamp 1698431365
transform 1 0 26656 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_229
timestamp 1698431365
transform 1 0 26992 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_245
timestamp 1698431365
transform 1 0 28784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_247
timestamp 1698431365
transform 1 0 29008 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_262
timestamp 1698431365
transform 1 0 30688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_266
timestamp 1698431365
transform 1 0 31136 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_278
timestamp 1698431365
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_286
timestamp 1698431365
transform 1 0 33376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_288
timestamp 1698431365
transform 1 0 33600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_291
timestamp 1698431365
transform 1 0 33936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_295
timestamp 1698431365
transform 1 0 34384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_299
timestamp 1698431365
transform 1 0 34832 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_303
timestamp 1698431365
transform 1 0 35280 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_318
timestamp 1698431365
transform 1 0 36960 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_326
timestamp 1698431365
transform 1 0 37856 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_330
timestamp 1698431365
transform 1 0 38304 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_18
timestamp 1698431365
transform 1 0 3360 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_41
timestamp 1698431365
transform 1 0 5936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_43
timestamp 1698431365
transform 1 0 6160 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_50
timestamp 1698431365
transform 1 0 6944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_58
timestamp 1698431365
transform 1 0 7840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_68
timestamp 1698431365
transform 1 0 8960 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_72
timestamp 1698431365
transform 1 0 9408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_76
timestamp 1698431365
transform 1 0 9856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_80
timestamp 1698431365
transform 1 0 10304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_84
timestamp 1698431365
transform 1 0 10752 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_93
timestamp 1698431365
transform 1 0 11760 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_99
timestamp 1698431365
transform 1 0 12432 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_141
timestamp 1698431365
transform 1 0 17136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_160
timestamp 1698431365
transform 1 0 19264 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_172
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_193
timestamp 1698431365
transform 1 0 22960 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_197
timestamp 1698431365
transform 1 0 23408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_201
timestamp 1698431365
transform 1 0 23856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_205
timestamp 1698431365
transform 1 0 24304 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_237
timestamp 1698431365
transform 1 0 27888 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_279
timestamp 1698431365
transform 1 0 32592 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_287
timestamp 1698431365
transform 1 0 33488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_291
timestamp 1698431365
transform 1 0 33936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_327
timestamp 1698431365
transform 1 0 37968 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_20
timestamp 1698431365
transform 1 0 3584 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_28
timestamp 1698431365
transform 1 0 4480 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_32
timestamp 1698431365
transform 1 0 4928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_51
timestamp 1698431365
transform 1 0 7056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_65
timestamp 1698431365
transform 1 0 8624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_69
timestamp 1698431365
transform 1 0 9072 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_80
timestamp 1698431365
transform 1 0 10304 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_83
timestamp 1698431365
transform 1 0 10640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_87
timestamp 1698431365
transform 1 0 11088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_91
timestamp 1698431365
transform 1 0 11536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_95
timestamp 1698431365
transform 1 0 11984 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_99
timestamp 1698431365
transform 1 0 12432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_103
timestamp 1698431365
transform 1 0 12880 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_107
timestamp 1698431365
transform 1 0 13328 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_125
timestamp 1698431365
transform 1 0 15344 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_129
timestamp 1698431365
transform 1 0 15792 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_132
timestamp 1698431365
transform 1 0 16128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_156
timestamp 1698431365
transform 1 0 18816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_158
timestamp 1698431365
transform 1 0 19040 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_199
timestamp 1698431365
transform 1 0 23632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_203
timestamp 1698431365
transform 1 0 24080 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_207
timestamp 1698431365
transform 1 0 24528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_214
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_225
timestamp 1698431365
transform 1 0 26544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_229
timestamp 1698431365
transform 1 0 26992 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_239
timestamp 1698431365
transform 1 0 28112 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_257
timestamp 1698431365
transform 1 0 30128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_259
timestamp 1698431365
transform 1 0 30352 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_268
timestamp 1698431365
transform 1 0 31360 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_327
timestamp 1698431365
transform 1 0 37968 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_41
timestamp 1698431365
transform 1 0 5936 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_47
timestamp 1698431365
transform 1 0 6608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_87
timestamp 1698431365
transform 1 0 11088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_123
timestamp 1698431365
transform 1 0 15120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_127
timestamp 1698431365
transform 1 0 15568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_129
timestamp 1698431365
transform 1 0 15792 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_153
timestamp 1698431365
transform 1 0 18480 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_157
timestamp 1698431365
transform 1 0 18928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_159
timestamp 1698431365
transform 1 0 19152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_162
timestamp 1698431365
transform 1 0 19488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_166
timestamp 1698431365
transform 1 0 19936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_168
timestamp 1698431365
transform 1 0 20160 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_210
timestamp 1698431365
transform 1 0 24864 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_251
timestamp 1698431365
transform 1 0 29456 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_312
timestamp 1698431365
transform 1 0 36288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_314
timestamp 1698431365
transform 1 0 36512 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_321
timestamp 1698431365
transform 1 0 37296 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_325
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_329
timestamp 1698431365
transform 1 0 38192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_43
timestamp 1698431365
transform 1 0 6160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_47
timestamp 1698431365
transform 1 0 6608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_51
timestamp 1698431365
transform 1 0 7056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_55
timestamp 1698431365
transform 1 0 7504 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_59
timestamp 1698431365
transform 1 0 7952 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_63
timestamp 1698431365
transform 1 0 8400 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_67
timestamp 1698431365
transform 1 0 8848 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_76
timestamp 1698431365
transform 1 0 9856 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_95
timestamp 1698431365
transform 1 0 11984 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_103
timestamp 1698431365
transform 1 0 12880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_107
timestamp 1698431365
transform 1 0 13328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_111
timestamp 1698431365
transform 1 0 13776 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_115
timestamp 1698431365
transform 1 0 14224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_119
timestamp 1698431365
transform 1 0 14672 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_123
timestamp 1698431365
transform 1 0 15120 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_126
timestamp 1698431365
transform 1 0 15456 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_134
timestamp 1698431365
transform 1 0 16352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_138
timestamp 1698431365
transform 1 0 16800 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_146
timestamp 1698431365
transform 1 0 17696 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_154
timestamp 1698431365
transform 1 0 18592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_156
timestamp 1698431365
transform 1 0 18816 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_209
timestamp 1698431365
transform 1 0 24752 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_216
timestamp 1698431365
transform 1 0 25536 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_227
timestamp 1698431365
transform 1 0 26768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_231
timestamp 1698431365
transform 1 0 27216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_250
timestamp 1698431365
transform 1 0 29344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_254
timestamp 1698431365
transform 1 0 29792 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_256
timestamp 1698431365
transform 1 0 30016 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_259
timestamp 1698431365
transform 1 0 30352 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_272
timestamp 1698431365
transform 1 0 31808 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_278
timestamp 1698431365
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_286
timestamp 1698431365
transform 1 0 33376 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_290
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_317
timestamp 1698431365
transform 1 0 36848 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_321
timestamp 1698431365
transform 1 0 37296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_325
timestamp 1698431365
transform 1 0 37744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_329
timestamp 1698431365
transform 1 0 38192 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_8
timestamp 1698431365
transform 1 0 2240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_26
timestamp 1698431365
transform 1 0 4256 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_58
timestamp 1698431365
transform 1 0 7840 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_62
timestamp 1698431365
transform 1 0 8288 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_66
timestamp 1698431365
transform 1 0 8736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_70
timestamp 1698431365
transform 1 0 9184 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_90
timestamp 1698431365
transform 1 0 11424 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_100
timestamp 1698431365
transform 1 0 12544 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_104
timestamp 1698431365
transform 1 0 12992 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_115
timestamp 1698431365
transform 1 0 14224 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_143
timestamp 1698431365
transform 1 0 17360 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_147
timestamp 1698431365
transform 1 0 17808 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_163
timestamp 1698431365
transform 1 0 19600 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_238
timestamp 1698431365
transform 1 0 28000 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_242
timestamp 1698431365
transform 1 0 28448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_244
timestamp 1698431365
transform 1 0 28672 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_251
timestamp 1698431365
transform 1 0 29456 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_255
timestamp 1698431365
transform 1 0 29904 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_273
timestamp 1698431365
transform 1 0 31920 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_277
timestamp 1698431365
transform 1 0 32368 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_321
timestamp 1698431365
transform 1 0 37296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_325
timestamp 1698431365
transform 1 0 37744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_329
timestamp 1698431365
transform 1 0 38192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_20
timestamp 1698431365
transform 1 0 3584 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_30
timestamp 1698431365
transform 1 0 4704 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_34
timestamp 1698431365
transform 1 0 5152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_52
timestamp 1698431365
transform 1 0 7168 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_61
timestamp 1698431365
transform 1 0 8176 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_63
timestamp 1698431365
transform 1 0 8400 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_83
timestamp 1698431365
transform 1 0 10640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_87
timestamp 1698431365
transform 1 0 11088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_89
timestamp 1698431365
transform 1 0 11312 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_124
timestamp 1698431365
transform 1 0 15232 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_128
timestamp 1698431365
transform 1 0 15680 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_132
timestamp 1698431365
transform 1 0 16128 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_139
timestamp 1698431365
transform 1 0 16912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_160
timestamp 1698431365
transform 1 0 19264 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_168
timestamp 1698431365
transform 1 0 20160 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_172
timestamp 1698431365
transform 1 0 20608 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_207
timestamp 1698431365
transform 1 0 24528 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_209
timestamp 1698431365
transform 1 0 24752 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_216
timestamp 1698431365
transform 1 0 25536 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_220
timestamp 1698431365
transform 1 0 25984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_224
timestamp 1698431365
transform 1 0 26432 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_228
timestamp 1698431365
transform 1 0 26880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_264
timestamp 1698431365
transform 1 0 30912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_268
timestamp 1698431365
transform 1 0 31360 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_286
timestamp 1698431365
transform 1 0 33376 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_323
timestamp 1698431365
transform 1 0 37520 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_41
timestamp 1698431365
transform 1 0 5936 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_45
timestamp 1698431365
transform 1 0 6384 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_83
timestamp 1698431365
transform 1 0 10640 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_87
timestamp 1698431365
transform 1 0 11088 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_98
timestamp 1698431365
transform 1 0 12320 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_161
timestamp 1698431365
transform 1 0 19376 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_165
timestamp 1698431365
transform 1 0 19824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_169
timestamp 1698431365
transform 1 0 20272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_173
timestamp 1698431365
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_185
timestamp 1698431365
transform 1 0 22064 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_241
timestamp 1698431365
transform 1 0 28336 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_263
timestamp 1698431365
transform 1 0 30800 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_292
timestamp 1698431365
transform 1 0 34048 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_296
timestamp 1698431365
transform 1 0 34496 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_312
timestamp 1698431365
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_325
timestamp 1698431365
transform 1 0 37744 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_329
timestamp 1698431365
transform 1 0 38192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_20
timestamp 1698431365
transform 1 0 3584 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_36
timestamp 1698431365
transform 1 0 5376 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_39
timestamp 1698431365
transform 1 0 5712 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_47
timestamp 1698431365
transform 1 0 6608 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_51
timestamp 1698431365
transform 1 0 7056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_60
timestamp 1698431365
transform 1 0 8064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_62
timestamp 1698431365
transform 1 0 8288 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_69
timestamp 1698431365
transform 1 0 9072 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_76
timestamp 1698431365
transform 1 0 9856 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_116
timestamp 1698431365
transform 1 0 14336 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_120
timestamp 1698431365
transform 1 0 14784 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_138
timestamp 1698431365
transform 1 0 16800 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_146
timestamp 1698431365
transform 1 0 17696 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_165
timestamp 1698431365
transform 1 0 19824 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_181
timestamp 1698431365
transform 1 0 21616 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_208
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_220
timestamp 1698431365
transform 1 0 25984 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_226
timestamp 1698431365
transform 1 0 26656 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_247
timestamp 1698431365
transform 1 0 29008 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_263
timestamp 1698431365
transform 1 0 30800 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_271
timestamp 1698431365
transform 1 0 31696 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_273
timestamp 1698431365
transform 1 0 31920 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_286
timestamp 1698431365
transform 1 0 33376 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_318
timestamp 1698431365
transform 1 0 36960 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_326
timestamp 1698431365
transform 1 0 37856 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_330
timestamp 1698431365
transform 1 0 38304 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_18
timestamp 1698431365
transform 1 0 3360 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_41
timestamp 1698431365
transform 1 0 5936 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_45
timestamp 1698431365
transform 1 0 6384 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_49
timestamp 1698431365
transform 1 0 6832 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_57
timestamp 1698431365
transform 1 0 7728 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_61
timestamp 1698431365
transform 1 0 8176 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_64
timestamp 1698431365
transform 1 0 8512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_68
timestamp 1698431365
transform 1 0 8960 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_71
timestamp 1698431365
transform 1 0 9296 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_103
timestamp 1698431365
transform 1 0 12880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_111
timestamp 1698431365
transform 1 0 13776 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_126
timestamp 1698431365
transform 1 0 15456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_140
timestamp 1698431365
transform 1 0 17024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_144
timestamp 1698431365
transform 1 0 17472 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_163
timestamp 1698431365
transform 1 0 19600 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_167
timestamp 1698431365
transform 1 0 20048 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_193
timestamp 1698431365
transform 1 0 22960 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_208
timestamp 1698431365
transform 1 0 24640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_212
timestamp 1698431365
transform 1 0 25088 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698431365
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_255
timestamp 1698431365
transform 1 0 29904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_259
timestamp 1698431365
transform 1 0 30352 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_261
timestamp 1698431365
transform 1 0 30576 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_264
timestamp 1698431365
transform 1 0 30912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_268
timestamp 1698431365
transform 1 0 31360 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_306
timestamp 1698431365
transform 1 0 35616 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698431365
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_325
timestamp 1698431365
transform 1 0 37744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_329
timestamp 1698431365
transform 1 0 38192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_62
timestamp 1698431365
transform 1 0 8288 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_76
timestamp 1698431365
transform 1 0 9856 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_94
timestamp 1698431365
transform 1 0 11872 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_110
timestamp 1698431365
transform 1 0 13664 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_158
timestamp 1698431365
transform 1 0 19040 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_162
timestamp 1698431365
transform 1 0 19488 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_198
timestamp 1698431365
transform 1 0 23520 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_202
timestamp 1698431365
transform 1 0 23968 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_216
timestamp 1698431365
transform 1 0 25536 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_220
timestamp 1698431365
transform 1 0 25984 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_228
timestamp 1698431365
transform 1 0 26880 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_246
timestamp 1698431365
transform 1 0 28896 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_262
timestamp 1698431365
transform 1 0 30688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_266
timestamp 1698431365
transform 1 0 31136 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_279
timestamp 1698431365
transform 1 0 32592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_286
timestamp 1698431365
transform 1 0 33376 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_318
timestamp 1698431365
transform 1 0 36960 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_326
timestamp 1698431365
transform 1 0 37856 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_330
timestamp 1698431365
transform 1 0 38304 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_10
timestamp 1698431365
transform 1 0 2464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_14
timestamp 1698431365
transform 1 0 2912 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_73
timestamp 1698431365
transform 1 0 9520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_77
timestamp 1698431365
transform 1 0 9968 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_81
timestamp 1698431365
transform 1 0 10416 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_98
timestamp 1698431365
transform 1 0 12320 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_102
timestamp 1698431365
transform 1 0 12768 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_104
timestamp 1698431365
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_111
timestamp 1698431365
transform 1 0 13776 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_143
timestamp 1698431365
transform 1 0 17360 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_159
timestamp 1698431365
transform 1 0 19152 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_163
timestamp 1698431365
transform 1 0 19600 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_231
timestamp 1698431365
transform 1 0 27216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_235
timestamp 1698431365
transform 1 0 27664 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_243
timestamp 1698431365
transform 1 0 28560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_255
timestamp 1698431365
transform 1 0 29904 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_302
timestamp 1698431365
transform 1 0 35168 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_310
timestamp 1698431365
transform 1 0 36064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698431365
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_325
timestamp 1698431365
transform 1 0 37744 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_329
timestamp 1698431365
transform 1 0 38192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_8
timestamp 1698431365
transform 1 0 2240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_26
timestamp 1698431365
transform 1 0 4256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_32
timestamp 1698431365
transform 1 0 4928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_44
timestamp 1698431365
transform 1 0 6272 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_48
timestamp 1698431365
transform 1 0 6720 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_64
timestamp 1698431365
transform 1 0 8512 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_68
timestamp 1698431365
transform 1 0 8960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_110
timestamp 1698431365
transform 1 0 13664 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_114
timestamp 1698431365
transform 1 0 14112 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_118
timestamp 1698431365
transform 1 0 14560 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_121
timestamp 1698431365
transform 1 0 14896 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_137
timestamp 1698431365
transform 1 0 16688 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1698431365
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_150
timestamp 1698431365
transform 1 0 18144 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_154
timestamp 1698431365
transform 1 0 18592 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_156
timestamp 1698431365
transform 1 0 18816 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_159
timestamp 1698431365
transform 1 0 19152 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_177
timestamp 1698431365
transform 1 0 21168 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_183
timestamp 1698431365
transform 1 0 21840 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_187
timestamp 1698431365
transform 1 0 22288 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_202
timestamp 1698431365
transform 1 0 23968 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_216
timestamp 1698431365
transform 1 0 25536 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_220
timestamp 1698431365
transform 1 0 25984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_222
timestamp 1698431365
transform 1 0 26208 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_259
timestamp 1698431365
transform 1 0 30352 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_261
timestamp 1698431365
transform 1 0 30576 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_267
timestamp 1698431365
transform 1 0 31248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_277
timestamp 1698431365
transform 1 0 32368 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_279
timestamp 1698431365
transform 1 0 32592 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_314
timestamp 1698431365
transform 1 0 36512 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_330
timestamp 1698431365
transform 1 0 38304 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_20
timestamp 1698431365
transform 1 0 3584 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_28
timestamp 1698431365
transform 1 0 4480 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698431365
transform 1 0 4928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_41
timestamp 1698431365
transform 1 0 5936 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_49
timestamp 1698431365
transform 1 0 6832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_52
timestamp 1698431365
transform 1 0 7168 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_56
timestamp 1698431365
transform 1 0 7616 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_92
timestamp 1698431365
transform 1 0 11648 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_130
timestamp 1698431365
transform 1 0 15904 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_138
timestamp 1698431365
transform 1 0 16800 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_142
timestamp 1698431365
transform 1 0 17248 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_157
timestamp 1698431365
transform 1 0 18928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_165
timestamp 1698431365
transform 1 0 19824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_169
timestamp 1698431365
transform 1 0 20272 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_173
timestamp 1698431365
transform 1 0 20720 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_193
timestamp 1698431365
transform 1 0 22960 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_201
timestamp 1698431365
transform 1 0 23856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_205
timestamp 1698431365
transform 1 0 24304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_209
timestamp 1698431365
transform 1 0 24752 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_213
timestamp 1698431365
transform 1 0 25200 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_251
timestamp 1698431365
transform 1 0 29456 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_261
timestamp 1698431365
transform 1 0 30576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_265
timestamp 1698431365
transform 1 0 31024 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_271
timestamp 1698431365
transform 1 0 31696 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_275
timestamp 1698431365
transform 1 0 32144 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_307
timestamp 1698431365
transform 1 0 35728 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_325
timestamp 1698431365
transform 1 0 37744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_329
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_36
timestamp 1698431365
transform 1 0 5376 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_40
timestamp 1698431365
transform 1 0 5824 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_58
timestamp 1698431365
transform 1 0 7840 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_62
timestamp 1698431365
transform 1 0 8288 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_87
timestamp 1698431365
transform 1 0 11088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_89
timestamp 1698431365
transform 1 0 11312 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_92
timestamp 1698431365
transform 1 0 11648 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_96
timestamp 1698431365
transform 1 0 12096 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_100
timestamp 1698431365
transform 1 0 12544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_102
timestamp 1698431365
transform 1 0 12768 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_113
timestamp 1698431365
transform 1 0 14000 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_130
timestamp 1698431365
transform 1 0 15904 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_138
timestamp 1698431365
transform 1 0 16800 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_146
timestamp 1698431365
transform 1 0 17696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_148
timestamp 1698431365
transform 1 0 17920 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_183
timestamp 1698431365
transform 1 0 21840 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_187
timestamp 1698431365
transform 1 0 22288 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_191
timestamp 1698431365
transform 1 0 22736 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_207
timestamp 1698431365
transform 1 0 24528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1698431365
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_220
timestamp 1698431365
transform 1 0 25984 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_226
timestamp 1698431365
transform 1 0 26656 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_264
timestamp 1698431365
transform 1 0 30912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_268
timestamp 1698431365
transform 1 0 31360 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_286
timestamp 1698431365
transform 1 0 33376 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_290
timestamp 1698431365
transform 1 0 33824 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_294
timestamp 1698431365
transform 1 0 34272 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_330
timestamp 1698431365
transform 1 0 38304 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_41
timestamp 1698431365
transform 1 0 5936 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_45
timestamp 1698431365
transform 1 0 6384 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_55
timestamp 1698431365
transform 1 0 7504 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_82
timestamp 1698431365
transform 1 0 10528 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_86
timestamp 1698431365
transform 1 0 10976 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_89
timestamp 1698431365
transform 1 0 11312 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_93
timestamp 1698431365
transform 1 0 11760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_97
timestamp 1698431365
transform 1 0 12208 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_109
timestamp 1698431365
transform 1 0 13552 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_120
timestamp 1698431365
transform 1 0 14784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_124
timestamp 1698431365
transform 1 0 15232 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_140
timestamp 1698431365
transform 1 0 17024 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_148
timestamp 1698431365
transform 1 0 17920 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_162
timestamp 1698431365
transform 1 0 19488 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_170
timestamp 1698431365
transform 1 0 20384 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_174
timestamp 1698431365
transform 1 0 20832 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_183
timestamp 1698431365
transform 1 0 21840 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_187
timestamp 1698431365
transform 1 0 22288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_191
timestamp 1698431365
transform 1 0 22736 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_223
timestamp 1698431365
transform 1 0 26320 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_239
timestamp 1698431365
transform 1 0 28112 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_243
timestamp 1698431365
transform 1 0 28560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_279
timestamp 1698431365
transform 1 0 32592 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_295
timestamp 1698431365
transform 1 0 34384 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_303
timestamp 1698431365
transform 1 0 35280 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_309
timestamp 1698431365
transform 1 0 35952 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_325
timestamp 1698431365
transform 1 0 37744 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_329
timestamp 1698431365
transform 1 0 38192 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_6
timestamp 1698431365
transform 1 0 2016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_8
timestamp 1698431365
transform 1 0 2240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_53
timestamp 1698431365
transform 1 0 7280 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_64
timestamp 1698431365
transform 1 0 8512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_68
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_76
timestamp 1698431365
transform 1 0 9856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_80
timestamp 1698431365
transform 1 0 10304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_108
timestamp 1698431365
transform 1 0 13440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_112
timestamp 1698431365
transform 1 0 13888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_154
timestamp 1698431365
transform 1 0 18592 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_159
timestamp 1698431365
transform 1 0 19152 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_167
timestamp 1698431365
transform 1 0 20048 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_175
timestamp 1698431365
transform 1 0 20944 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_181
timestamp 1698431365
transform 1 0 21616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_195
timestamp 1698431365
transform 1 0 23184 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_203
timestamp 1698431365
transform 1 0 24080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_207
timestamp 1698431365
transform 1 0 24528 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_216
timestamp 1698431365
transform 1 0 25536 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_220
timestamp 1698431365
transform 1 0 25984 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_252
timestamp 1698431365
transform 1 0 29568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_268
timestamp 1698431365
transform 1 0 31360 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_272
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_276
timestamp 1698431365
transform 1 0 32256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_325
timestamp 1698431365
transform 1 0 37744 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_329
timestamp 1698431365
transform 1 0 38192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_10
timestamp 1698431365
transform 1 0 2464 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_14
timestamp 1698431365
transform 1 0 2912 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_30
timestamp 1698431365
transform 1 0 4704 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_52
timestamp 1698431365
transform 1 0 7168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_104
timestamp 1698431365
transform 1 0 12992 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_111
timestamp 1698431365
transform 1 0 13776 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_136
timestamp 1698431365
transform 1 0 16576 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_219
timestamp 1698431365
transform 1 0 25872 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_223
timestamp 1698431365
transform 1 0 26320 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_227
timestamp 1698431365
transform 1 0 26768 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_231
timestamp 1698431365
transform 1 0 27216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_235
timestamp 1698431365
transform 1 0 27664 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_241
timestamp 1698431365
transform 1 0 28336 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_283
timestamp 1698431365
transform 1 0 33040 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_287
timestamp 1698431365
transform 1 0 33488 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_289
timestamp 1698431365
transform 1 0 33712 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_292
timestamp 1698431365
transform 1 0 34048 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_304
timestamp 1698431365
transform 1 0 35392 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_306
timestamp 1698431365
transform 1 0 35616 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_327
timestamp 1698431365
transform 1 0 37968 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_2
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_26
timestamp 1698431365
transform 1 0 4256 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_42
timestamp 1698431365
transform 1 0 6048 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_56
timestamp 1698431365
transform 1 0 7616 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_66
timestamp 1698431365
transform 1 0 8736 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_87
timestamp 1698431365
transform 1 0 11088 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_89
timestamp 1698431365
transform 1 0 11312 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_136
timestamp 1698431365
transform 1 0 16576 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_148
timestamp 1698431365
transform 1 0 17920 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_175
timestamp 1698431365
transform 1 0 20944 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_242
timestamp 1698431365
transform 1 0 28448 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_250
timestamp 1698431365
transform 1 0 29344 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_256
timestamp 1698431365
transform 1 0 30016 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_268
timestamp 1698431365
transform 1 0 31360 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_276
timestamp 1698431365
transform 1 0 32256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_286
timestamp 1698431365
transform 1 0 33376 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_288
timestamp 1698431365
transform 1 0 33600 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_2
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_26
timestamp 1698431365
transform 1 0 4256 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_45
timestamp 1698431365
transform 1 0 6384 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_49
timestamp 1698431365
transform 1 0 6832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_51
timestamp 1698431365
transform 1 0 7056 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_59
timestamp 1698431365
transform 1 0 7952 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_63
timestamp 1698431365
transform 1 0 8400 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_65
timestamp 1698431365
transform 1 0 8624 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_102
timestamp 1698431365
transform 1 0 12768 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_104
timestamp 1698431365
transform 1 0 12992 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_111
timestamp 1698431365
transform 1 0 13776 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_113
timestamp 1698431365
transform 1 0 14000 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_126
timestamp 1698431365
transform 1 0 15456 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_130
timestamp 1698431365
transform 1 0 15904 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_134
timestamp 1698431365
transform 1 0 16352 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_138
timestamp 1698431365
transform 1 0 16800 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_186
timestamp 1698431365
transform 1 0 22176 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_190
timestamp 1698431365
transform 1 0 22624 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_198
timestamp 1698431365
transform 1 0 23520 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_233
timestamp 1698431365
transform 1 0 27440 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_237
timestamp 1698431365
transform 1 0 27888 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_241
timestamp 1698431365
transform 1 0 28336 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_251
timestamp 1698431365
transform 1 0 29456 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_262
timestamp 1698431365
transform 1 0 30688 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_266
timestamp 1698431365
transform 1 0 31136 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_278
timestamp 1698431365
transform 1 0 32480 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_282
timestamp 1698431365
transform 1 0 32928 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_290
timestamp 1698431365
transform 1 0 33824 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_294
timestamp 1698431365
transform 1 0 34272 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_297
timestamp 1698431365
transform 1 0 34608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_307
timestamp 1698431365
transform 1 0 35728 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_325
timestamp 1698431365
transform 1 0 37744 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_329
timestamp 1698431365
transform 1 0 38192 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_66
timestamp 1698431365
transform 1 0 8736 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_90
timestamp 1698431365
transform 1 0 11424 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_94
timestamp 1698431365
transform 1 0 11872 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_100
timestamp 1698431365
transform 1 0 12544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_106
timestamp 1698431365
transform 1 0 13216 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_135
timestamp 1698431365
transform 1 0 16464 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_139
timestamp 1698431365
transform 1 0 16912 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_146
timestamp 1698431365
transform 1 0 17696 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_148
timestamp 1698431365
transform 1 0 17920 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_151
timestamp 1698431365
transform 1 0 18256 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_159
timestamp 1698431365
transform 1 0 19152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_184
timestamp 1698431365
transform 1 0 21952 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_188
timestamp 1698431365
transform 1 0 22400 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_204
timestamp 1698431365
transform 1 0 24192 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_208
timestamp 1698431365
transform 1 0 24640 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_216
timestamp 1698431365
transform 1 0 25536 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_278
timestamp 1698431365
transform 1 0 32480 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_288
timestamp 1698431365
transform 1 0 33600 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_320
timestamp 1698431365
transform 1 0 37184 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_328
timestamp 1698431365
transform 1 0 38080 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_330
timestamp 1698431365
transform 1 0 38304 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_6
timestamp 1698431365
transform 1 0 2016 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_22
timestamp 1698431365
transform 1 0 3808 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_30
timestamp 1698431365
transform 1 0 4704 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_41
timestamp 1698431365
transform 1 0 5936 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_45
timestamp 1698431365
transform 1 0 6384 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_49
timestamp 1698431365
transform 1 0 6832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_53
timestamp 1698431365
transform 1 0 7280 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_85
timestamp 1698431365
transform 1 0 10864 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_101
timestamp 1698431365
transform 1 0 12656 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_104
timestamp 1698431365
transform 1 0 12992 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_139
timestamp 1698431365
transform 1 0 16912 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_155
timestamp 1698431365
transform 1 0 18704 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_165
timestamp 1698431365
transform 1 0 19824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_169
timestamp 1698431365
transform 1 0 20272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_173
timestamp 1698431365
transform 1 0 20720 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_181
timestamp 1698431365
transform 1 0 21616 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_225
timestamp 1698431365
transform 1 0 26544 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_233
timestamp 1698431365
transform 1 0 27440 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_249
timestamp 1698431365
transform 1 0 29232 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_292
timestamp 1698431365
transform 1 0 34048 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_296
timestamp 1698431365
transform 1 0 34496 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_304
timestamp 1698431365
transform 1 0 35392 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_308
timestamp 1698431365
transform 1 0 35840 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_325
timestamp 1698431365
transform 1 0 37744 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_329
timestamp 1698431365
transform 1 0 38192 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_62
timestamp 1698431365
transform 1 0 8288 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_66
timestamp 1698431365
transform 1 0 8736 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_76
timestamp 1698431365
transform 1 0 9856 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_80
timestamp 1698431365
transform 1 0 10304 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_96
timestamp 1698431365
transform 1 0 12096 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_104
timestamp 1698431365
transform 1 0 12992 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_106
timestamp 1698431365
transform 1 0 13216 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_113
timestamp 1698431365
transform 1 0 14000 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_137
timestamp 1698431365
transform 1 0 16688 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_139
timestamp 1698431365
transform 1 0 16912 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_174
timestamp 1698431365
transform 1 0 20832 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_177
timestamp 1698431365
transform 1 0 21168 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_181
timestamp 1698431365
transform 1 0 21616 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_197
timestamp 1698431365
transform 1 0 23408 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_205
timestamp 1698431365
transform 1 0 24304 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_209
timestamp 1698431365
transform 1 0 24752 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_216
timestamp 1698431365
transform 1 0 25536 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_224
timestamp 1698431365
transform 1 0 26432 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_279
timestamp 1698431365
transform 1 0 32592 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_287
timestamp 1698431365
transform 1 0 33488 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_291
timestamp 1698431365
transform 1 0 33936 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_295
timestamp 1698431365
transform 1 0 34384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_6
timestamp 1698431365
transform 1 0 2016 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_14
timestamp 1698431365
transform 1 0 2912 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_18
timestamp 1698431365
transform 1 0 3360 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1698431365
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_72
timestamp 1698431365
transform 1 0 9408 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_78
timestamp 1698431365
transform 1 0 10080 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_82
timestamp 1698431365
transform 1 0 10528 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_100
timestamp 1698431365
transform 1 0 12544 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_134
timestamp 1698431365
transform 1 0 16352 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_138
timestamp 1698431365
transform 1 0 16800 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_192
timestamp 1698431365
transform 1 0 22848 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_200
timestamp 1698431365
transform 1 0 23744 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_202
timestamp 1698431365
transform 1 0 23968 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_205
timestamp 1698431365
transform 1 0 24304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_209
timestamp 1698431365
transform 1 0 24752 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_226
timestamp 1698431365
transform 1 0 26656 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_234
timestamp 1698431365
transform 1 0 27552 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_238
timestamp 1698431365
transform 1 0 28000 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_240
timestamp 1698431365
transform 1 0 28224 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_249
timestamp 1698431365
transform 1 0 29232 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_284
timestamp 1698431365
transform 1 0 33152 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_288
timestamp 1698431365
transform 1 0 33600 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_292
timestamp 1698431365
transform 1 0 34048 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_294
timestamp 1698431365
transform 1 0 34272 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_297
timestamp 1698431365
transform 1 0 34608 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_325
timestamp 1698431365
transform 1 0 37744 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_329
timestamp 1698431365
transform 1 0 38192 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_6
timestamp 1698431365
transform 1 0 2016 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_22
timestamp 1698431365
transform 1 0 3808 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_26
timestamp 1698431365
transform 1 0 4256 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_74
timestamp 1698431365
transform 1 0 9632 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_135
timestamp 1698431365
transform 1 0 16464 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_139
timestamp 1698431365
transform 1 0 16912 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_158
timestamp 1698431365
transform 1 0 19040 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_172
timestamp 1698431365
transform 1 0 20608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_174
timestamp 1698431365
transform 1 0 20832 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_209
timestamp 1698431365
transform 1 0 24752 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_246
timestamp 1698431365
transform 1 0 28896 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_250
timestamp 1698431365
transform 1 0 29344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_254
timestamp 1698431365
transform 1 0 29792 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_258
timestamp 1698431365
transform 1 0 30240 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_267
timestamp 1698431365
transform 1 0 31248 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_275
timestamp 1698431365
transform 1 0 32144 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_279
timestamp 1698431365
transform 1 0 32592 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_288
timestamp 1698431365
transform 1 0 33600 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_324
timestamp 1698431365
transform 1 0 37632 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_328
timestamp 1698431365
transform 1 0 38080 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_330
timestamp 1698431365
transform 1 0 38304 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_6
timestamp 1698431365
transform 1 0 2016 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_14
timestamp 1698431365
transform 1 0 2912 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_18
timestamp 1698431365
transform 1 0 3360 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_41
timestamp 1698431365
transform 1 0 5936 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_45
timestamp 1698431365
transform 1 0 6384 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_70
timestamp 1698431365
transform 1 0 9184 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_72
timestamp 1698431365
transform 1 0 9408 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_75
timestamp 1698431365
transform 1 0 9744 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_102
timestamp 1698431365
transform 1 0 12768 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_104
timestamp 1698431365
transform 1 0 12992 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_111
timestamp 1698431365
transform 1 0 13776 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_115
timestamp 1698431365
transform 1 0 14224 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_119
timestamp 1698431365
transform 1 0 14672 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_144
timestamp 1698431365
transform 1 0 17472 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_152
timestamp 1698431365
transform 1 0 18368 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_156
timestamp 1698431365
transform 1 0 18816 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_193
timestamp 1698431365
transform 1 0 22960 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_197
timestamp 1698431365
transform 1 0 23408 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_201
timestamp 1698431365
transform 1 0 23856 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_205
timestamp 1698431365
transform 1 0 24304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_215
timestamp 1698431365
transform 1 0 25424 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_219
timestamp 1698431365
transform 1 0 25872 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_223
timestamp 1698431365
transform 1 0 26320 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_232
timestamp 1698431365
transform 1 0 27328 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_240
timestamp 1698431365
transform 1 0 28224 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_242
timestamp 1698431365
transform 1 0 28448 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_251
timestamp 1698431365
transform 1 0 29456 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_253
timestamp 1698431365
transform 1 0 29680 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_274
timestamp 1698431365
transform 1 0 32032 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_282
timestamp 1698431365
transform 1 0 32928 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_286
timestamp 1698431365
transform 1 0 33376 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_290
timestamp 1698431365
transform 1 0 33824 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_294
timestamp 1698431365
transform 1 0 34272 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_296
timestamp 1698431365
transform 1 0 34496 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_311
timestamp 1698431365
transform 1 0 36176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_325
timestamp 1698431365
transform 1 0 37744 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_329
timestamp 1698431365
transform 1 0 38192 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_37
timestamp 1698431365
transform 1 0 5488 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_41
timestamp 1698431365
transform 1 0 5936 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_45
timestamp 1698431365
transform 1 0 6384 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_61
timestamp 1698431365
transform 1 0 8176 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_65
timestamp 1698431365
transform 1 0 8624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_67
timestamp 1698431365
transform 1 0 8848 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_106
timestamp 1698431365
transform 1 0 13216 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_108
timestamp 1698431365
transform 1 0 13440 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_135
timestamp 1698431365
transform 1 0 16464 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_139
timestamp 1698431365
transform 1 0 16912 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_168
timestamp 1698431365
transform 1 0 20160 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_172
timestamp 1698431365
transform 1 0 20608 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_204
timestamp 1698431365
transform 1 0 24192 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_208
timestamp 1698431365
transform 1 0 24640 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_265
timestamp 1698431365
transform 1 0 31024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_269
timestamp 1698431365
transform 1 0 31472 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_273
timestamp 1698431365
transform 1 0 31920 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_277
timestamp 1698431365
transform 1 0 32368 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_279
timestamp 1698431365
transform 1 0 32592 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_282
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_314
timestamp 1698431365
transform 1 0 36512 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_330
timestamp 1698431365
transform 1 0 38304 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_6
timestamp 1698431365
transform 1 0 2016 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_18
timestamp 1698431365
transform 1 0 3360 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_24
timestamp 1698431365
transform 1 0 4032 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_32
timestamp 1698431365
transform 1 0 4928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_37
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_41
timestamp 1698431365
transform 1 0 5936 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_49
timestamp 1698431365
transform 1 0 6832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_91
timestamp 1698431365
transform 1 0 11536 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_95
timestamp 1698431365
transform 1 0 11984 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_135
timestamp 1698431365
transform 1 0 16464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_139
timestamp 1698431365
transform 1 0 16912 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_143
timestamp 1698431365
transform 1 0 17360 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_164
timestamp 1698431365
transform 1 0 19712 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_168
timestamp 1698431365
transform 1 0 20160 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_171
timestamp 1698431365
transform 1 0 20496 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_177
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_241
timestamp 1698431365
transform 1 0 28336 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_247
timestamp 1698431365
transform 1 0 29008 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_251
timestamp 1698431365
transform 1 0 29456 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_255
timestamp 1698431365
transform 1 0 29904 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_287
timestamp 1698431365
transform 1 0 33488 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_295
timestamp 1698431365
transform 1 0 34384 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_299
timestamp 1698431365
transform 1 0 34832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_301
timestamp 1698431365
transform 1 0 35056 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_312
timestamp 1698431365
transform 1 0 36288 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_314
timestamp 1698431365
transform 1 0 36512 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_325
timestamp 1698431365
transform 1 0 37744 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_329
timestamp 1698431365
transform 1 0 38192 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_36
timestamp 1698431365
transform 1 0 5376 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_40
timestamp 1698431365
transform 1 0 5824 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_44
timestamp 1698431365
transform 1 0 6272 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_52
timestamp 1698431365
transform 1 0 7168 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_56
timestamp 1698431365
transform 1 0 7616 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_60
timestamp 1698431365
transform 1 0 8064 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_68
timestamp 1698431365
transform 1 0 8960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_76
timestamp 1698431365
transform 1 0 9856 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_79
timestamp 1698431365
transform 1 0 10192 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_85
timestamp 1698431365
transform 1 0 10864 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_101
timestamp 1698431365
transform 1 0 12656 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_104
timestamp 1698431365
transform 1 0 12992 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_115
timestamp 1698431365
transform 1 0 14224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_119
timestamp 1698431365
transform 1 0 14672 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_135
timestamp 1698431365
transform 1 0 16464 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_139
timestamp 1698431365
transform 1 0 16912 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_142
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_146
timestamp 1698431365
transform 1 0 17696 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_149
timestamp 1698431365
transform 1 0 18032 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_153
timestamp 1698431365
transform 1 0 18480 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_182
timestamp 1698431365
transform 1 0 21728 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_186
timestamp 1698431365
transform 1 0 22176 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_202
timestamp 1698431365
transform 1 0 23968 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_248
timestamp 1698431365
transform 1 0 29120 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_252
timestamp 1698431365
transform 1 0 29568 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_260
timestamp 1698431365
transform 1 0 30464 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_262
timestamp 1698431365
transform 1 0 30688 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_274
timestamp 1698431365
transform 1 0 32032 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_278
timestamp 1698431365
transform 1 0 32480 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_282
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_286
timestamp 1698431365
transform 1 0 33376 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_288
timestamp 1698431365
transform 1 0 33600 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_325
timestamp 1698431365
transform 1 0 37744 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_329
timestamp 1698431365
transform 1 0 38192 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_10
timestamp 1698431365
transform 1 0 2464 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_18
timestamp 1698431365
transform 1 0 3360 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_22
timestamp 1698431365
transform 1 0 3808 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_41
timestamp 1698431365
transform 1 0 5936 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_58
timestamp 1698431365
transform 1 0 7840 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_68
timestamp 1698431365
transform 1 0 8960 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_72
timestamp 1698431365
transform 1 0 9408 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_74
timestamp 1698431365
transform 1 0 9632 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_77
timestamp 1698431365
transform 1 0 9968 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_96
timestamp 1698431365
transform 1 0 12096 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_104
timestamp 1698431365
transform 1 0 12992 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_123
timestamp 1698431365
transform 1 0 15120 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_127
timestamp 1698431365
transform 1 0 15568 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_135
timestamp 1698431365
transform 1 0 16464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_139
timestamp 1698431365
transform 1 0 16912 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_143
timestamp 1698431365
transform 1 0 17360 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_147
timestamp 1698431365
transform 1 0 17808 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_151
timestamp 1698431365
transform 1 0 18256 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_168
timestamp 1698431365
transform 1 0 20160 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_192
timestamp 1698431365
transform 1 0 22848 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_200
timestamp 1698431365
transform 1 0 23744 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_204
timestamp 1698431365
transform 1 0 24192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_206
timestamp 1698431365
transform 1 0 24416 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_209
timestamp 1698431365
transform 1 0 24752 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_213
timestamp 1698431365
transform 1 0 25200 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_217
timestamp 1698431365
transform 1 0 25648 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_221
timestamp 1698431365
transform 1 0 26096 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_225
timestamp 1698431365
transform 1 0 26544 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_241
timestamp 1698431365
transform 1 0 28336 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_281
timestamp 1698431365
transform 1 0 32816 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_297
timestamp 1698431365
transform 1 0 34608 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_305
timestamp 1698431365
transform 1 0 35504 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_325
timestamp 1698431365
transform 1 0 37744 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_329
timestamp 1698431365
transform 1 0 38192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_10
timestamp 1698431365
transform 1 0 2464 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_14
timestamp 1698431365
transform 1 0 2912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_31
timestamp 1698431365
transform 1 0 4816 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_33
timestamp 1698431365
transform 1 0 5040 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_106
timestamp 1698431365
transform 1 0 13216 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_110
timestamp 1698431365
transform 1 0 13664 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_114
timestamp 1698431365
transform 1 0 14112 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_118
timestamp 1698431365
transform 1 0 14560 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_120
timestamp 1698431365
transform 1 0 14784 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_166
timestamp 1698431365
transform 1 0 19936 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_170
timestamp 1698431365
transform 1 0 20384 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_172
timestamp 1698431365
transform 1 0 20608 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_207
timestamp 1698431365
transform 1 0 24528 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_209
timestamp 1698431365
transform 1 0 24752 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_224
timestamp 1698431365
transform 1 0 26432 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_228
timestamp 1698431365
transform 1 0 26880 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_278
timestamp 1698431365
transform 1 0 32480 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_287
timestamp 1698431365
transform 1 0 33488 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_325
timestamp 1698431365
transform 1 0 37744 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_329
timestamp 1698431365
transform 1 0 38192 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_6
timestamp 1698431365
transform 1 0 2016 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_16
timestamp 1698431365
transform 1 0 3136 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_48
timestamp 1698431365
transform 1 0 6720 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_52
timestamp 1698431365
transform 1 0 7168 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_64
timestamp 1698431365
transform 1 0 8512 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_68
timestamp 1698431365
transform 1 0 8960 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_74
timestamp 1698431365
transform 1 0 9632 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_78
timestamp 1698431365
transform 1 0 10080 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_86
timestamp 1698431365
transform 1 0 10976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_90
timestamp 1698431365
transform 1 0 11424 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_98
timestamp 1698431365
transform 1 0 12320 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_102
timestamp 1698431365
transform 1 0 12768 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_104
timestamp 1698431365
transform 1 0 12992 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_111
timestamp 1698431365
transform 1 0 13776 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_160
timestamp 1698431365
transform 1 0 19264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_162
timestamp 1698431365
transform 1 0 19488 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_173
timestamp 1698431365
transform 1 0 20720 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_232
timestamp 1698431365
transform 1 0 27328 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_236
timestamp 1698431365
transform 1 0 27776 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_244
timestamp 1698431365
transform 1 0 28672 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_247
timestamp 1698431365
transform 1 0 29008 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_279
timestamp 1698431365
transform 1 0 32592 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_283
timestamp 1698431365
transform 1 0 33040 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_299
timestamp 1698431365
transform 1 0 34832 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_310
timestamp 1698431365
transform 1 0 36064 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_314
timestamp 1698431365
transform 1 0 36512 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_323
timestamp 1698431365
transform 1 0 37520 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_6
timestamp 1698431365
transform 1 0 2016 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_14
timestamp 1698431365
transform 1 0 2912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_50
timestamp 1698431365
transform 1 0 6944 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_54
timestamp 1698431365
transform 1 0 7392 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_58
timestamp 1698431365
transform 1 0 7840 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_66
timestamp 1698431365
transform 1 0 8736 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_72
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_76
timestamp 1698431365
transform 1 0 9856 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_79
timestamp 1698431365
transform 1 0 10192 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_83
timestamp 1698431365
transform 1 0 10640 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_87
timestamp 1698431365
transform 1 0 11088 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_139
timestamp 1698431365
transform 1 0 16912 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_142
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_169
timestamp 1698431365
transform 1 0 20272 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_175
timestamp 1698431365
transform 1 0 20944 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_191
timestamp 1698431365
transform 1 0 22736 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_199
timestamp 1698431365
transform 1 0 23632 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_246
timestamp 1698431365
transform 1 0 28896 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_250
timestamp 1698431365
transform 1 0 29344 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_258
timestamp 1698431365
transform 1 0 30240 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_261
timestamp 1698431365
transform 1 0 30576 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_269
timestamp 1698431365
transform 1 0 31472 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_277
timestamp 1698431365
transform 1 0 32368 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_279
timestamp 1698431365
transform 1 0 32592 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_282
timestamp 1698431365
transform 1 0 32928 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_298
timestamp 1698431365
transform 1 0 34720 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_302
timestamp 1698431365
transform 1 0 35168 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_312
timestamp 1698431365
transform 1 0 36288 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_328
timestamp 1698431365
transform 1 0 38080 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_330
timestamp 1698431365
transform 1 0 38304 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1698431365
transform 1 0 5152 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_41
timestamp 1698431365
transform 1 0 5936 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_45
timestamp 1698431365
transform 1 0 6384 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_47
timestamp 1698431365
transform 1 0 6608 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_84
timestamp 1698431365
transform 1 0 10752 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_115
timestamp 1698431365
transform 1 0 14224 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_117
timestamp 1698431365
transform 1 0 14448 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_124
timestamp 1698431365
transform 1 0 15232 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_162
timestamp 1698431365
transform 1 0 19488 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_166
timestamp 1698431365
transform 1 0 19936 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_174
timestamp 1698431365
transform 1 0 20832 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_193
timestamp 1698431365
transform 1 0 22960 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_239
timestamp 1698431365
transform 1 0 28112 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_243
timestamp 1698431365
transform 1 0 28560 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_247
timestamp 1698431365
transform 1 0 29008 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_251
timestamp 1698431365
transform 1 0 29456 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_253
timestamp 1698431365
transform 1 0 29680 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_290
timestamp 1698431365
transform 1 0 33824 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_314
timestamp 1698431365
transform 1 0 36512 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_317
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_325
timestamp 1698431365
transform 1 0 37744 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_329
timestamp 1698431365
transform 1 0 38192 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_6
timestamp 1698431365
transform 1 0 2016 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_38
timestamp 1698431365
transform 1 0 5600 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_64
timestamp 1698431365
transform 1 0 8512 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_77
timestamp 1698431365
transform 1 0 9968 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_79
timestamp 1698431365
transform 1 0 10192 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_118
timestamp 1698431365
transform 1 0 14560 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_122
timestamp 1698431365
transform 1 0 15008 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_159
timestamp 1698431365
transform 1 0 19152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_163
timestamp 1698431365
transform 1 0 19600 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_195
timestamp 1698431365
transform 1 0 23184 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_203
timestamp 1698431365
transform 1 0 24080 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_207
timestamp 1698431365
transform 1 0 24528 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_220
timestamp 1698431365
transform 1 0 25984 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_226
timestamp 1698431365
transform 1 0 26656 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_258
timestamp 1698431365
transform 1 0 30240 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_276
timestamp 1698431365
transform 1 0 32256 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_288
timestamp 1698431365
transform 1 0 33600 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_6
timestamp 1698431365
transform 1 0 2016 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_18
timestamp 1698431365
transform 1 0 3360 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_37
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_69
timestamp 1698431365
transform 1 0 9072 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_85
timestamp 1698431365
transform 1 0 10864 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_88
timestamp 1698431365
transform 1 0 11200 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_104
timestamp 1698431365
transform 1 0 12992 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_115
timestamp 1698431365
transform 1 0 14224 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_119
timestamp 1698431365
transform 1 0 14672 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_122
timestamp 1698431365
transform 1 0 15008 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_126
timestamp 1698431365
transform 1 0 15456 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_130
timestamp 1698431365
transform 1 0 15904 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_133
timestamp 1698431365
transform 1 0 16240 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_149
timestamp 1698431365
transform 1 0 18032 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_172
timestamp 1698431365
transform 1 0 20608 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_174
timestamp 1698431365
transform 1 0 20832 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_181
timestamp 1698431365
transform 1 0 21616 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_185
timestamp 1698431365
transform 1 0 22064 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_189
timestamp 1698431365
transform 1 0 22512 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_197
timestamp 1698431365
transform 1 0 23408 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_201
timestamp 1698431365
transform 1 0 23856 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_203
timestamp 1698431365
transform 1 0 24080 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_232
timestamp 1698431365
transform 1 0 27328 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_240
timestamp 1698431365
transform 1 0 28224 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_244
timestamp 1698431365
transform 1 0 28672 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_247
timestamp 1698431365
transform 1 0 29008 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_263
timestamp 1698431365
transform 1 0 30800 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_317
timestamp 1698431365
transform 1 0 36848 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_325
timestamp 1698431365
transform 1 0 37744 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_329
timestamp 1698431365
transform 1 0 38192 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_34
timestamp 1698431365
transform 1 0 5152 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_37
timestamp 1698431365
transform 1 0 5488 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_69
timestamp 1698431365
transform 1 0 9072 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1698431365
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_195
timestamp 1698431365
transform 1 0 23184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_87_199
timestamp 1698431365
transform 1 0 23632 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_207
timestamp 1698431365
transform 1 0 24528 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_209
timestamp 1698431365
transform 1 0 24752 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_228
timestamp 1698431365
transform 1 0 26880 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_232
timestamp 1698431365
transform 1 0 27328 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_261
timestamp 1698431365
transform 1 0 30576 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_277
timestamp 1698431365
transform 1 0 32368 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_279
timestamp 1698431365
transform 1 0 32592 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_282
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_298
timestamp 1698431365
transform 1 0 34720 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_303
timestamp 1698431365
transform 1 0 35280 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_315
timestamp 1698431365
transform 1 0 36624 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_6
timestamp 1698431365
transform 1 0 2016 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_14
timestamp 1698431365
transform 1 0 2912 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_18
timestamp 1698431365
transform 1 0 3360 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_39
timestamp 1698431365
transform 1 0 5712 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_44
timestamp 1698431365
transform 1 0 6272 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_52
timestamp 1698431365
transform 1 0 7168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_54
timestamp 1698431365
transform 1 0 7392 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_63
timestamp 1698431365
transform 1 0 8400 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_67
timestamp 1698431365
transform 1 0 8848 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_71
timestamp 1698431365
transform 1 0 9296 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_74
timestamp 1698431365
transform 1 0 9632 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_78
timestamp 1698431365
transform 1 0 10080 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_94
timestamp 1698431365
transform 1 0 11872 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_102
timestamp 1698431365
transform 1 0 12768 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_104
timestamp 1698431365
transform 1 0 12992 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_171
timestamp 1698431365
transform 1 0 20496 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_203
timestamp 1698431365
transform 1 0 24080 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_207
timestamp 1698431365
transform 1 0 24528 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_239
timestamp 1698431365
transform 1 0 28112 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_243
timestamp 1698431365
transform 1 0 28560 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_247
timestamp 1698431365
transform 1 0 29008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_311
timestamp 1698431365
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_325
timestamp 1698431365
transform 1 0 37744 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_329
timestamp 1698431365
transform 1 0 38192 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_80
timestamp 1698431365
transform 1 0 10304 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_84
timestamp 1698431365
transform 1 0 10752 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_88
timestamp 1698431365
transform 1 0 11200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_124
timestamp 1698431365
transform 1 0 15232 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_128
timestamp 1698431365
transform 1 0 15680 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_132
timestamp 1698431365
transform 1 0 16128 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_158
timestamp 1698431365
transform 1 0 19040 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_162
timestamp 1698431365
transform 1 0 19488 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_164
timestamp 1698431365
transform 1 0 19712 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_199
timestamp 1698431365
transform 1 0 23632 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_203
timestamp 1698431365
transform 1 0 24080 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_207
timestamp 1698431365
transform 1 0 24528 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_209
timestamp 1698431365
transform 1 0 24752 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_276
timestamp 1698431365
transform 1 0 32256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_282
timestamp 1698431365
transform 1 0 32928 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_314
timestamp 1698431365
transform 1 0 36512 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_330
timestamp 1698431365
transform 1 0 38304 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_10
timestamp 1698431365
transform 1 0 2464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_14
timestamp 1698431365
transform 1 0 2912 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_16
timestamp 1698431365
transform 1 0 3136 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_32
timestamp 1698431365
transform 1 0 4928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1698431365
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_41
timestamp 1698431365
transform 1 0 5936 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_45
timestamp 1698431365
transform 1 0 6384 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_49
timestamp 1698431365
transform 1 0 6832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_51
timestamp 1698431365
transform 1 0 7056 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_86
timestamp 1698431365
transform 1 0 10976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_90
timestamp 1698431365
transform 1 0 11424 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_92
timestamp 1698431365
transform 1 0 11648 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_95
timestamp 1698431365
transform 1 0 11984 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_123
timestamp 1698431365
transform 1 0 15120 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_163
timestamp 1698431365
transform 1 0 19600 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_167
timestamp 1698431365
transform 1 0 20048 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_241
timestamp 1698431365
transform 1 0 28336 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_247
timestamp 1698431365
transform 1 0 29008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_311
timestamp 1698431365
transform 1 0 36176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_325
timestamp 1698431365
transform 1 0 37744 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_329
timestamp 1698431365
transform 1 0 38192 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_2
timestamp 1698431365
transform 1 0 1568 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_10
timestamp 1698431365
transform 1 0 2464 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_48
timestamp 1698431365
transform 1 0 6720 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_52
timestamp 1698431365
transform 1 0 7168 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_56
timestamp 1698431365
transform 1 0 7616 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_58
timestamp 1698431365
transform 1 0 7840 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_61
timestamp 1698431365
transform 1 0 8176 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_74
timestamp 1698431365
transform 1 0 9632 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_80
timestamp 1698431365
transform 1 0 10304 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_94
timestamp 1698431365
transform 1 0 11872 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_96
timestamp 1698431365
transform 1 0 12096 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_105
timestamp 1698431365
transform 1 0 13104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_109
timestamp 1698431365
transform 1 0 13552 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_113
timestamp 1698431365
transform 1 0 14000 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_118
timestamp 1698431365
transform 1 0 14560 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_122
timestamp 1698431365
transform 1 0 15008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_126
timestamp 1698431365
transform 1 0 15456 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_130
timestamp 1698431365
transform 1 0 15904 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_142
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_144
timestamp 1698431365
transform 1 0 17472 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_151
timestamp 1698431365
transform 1 0 18256 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_155
timestamp 1698431365
transform 1 0 18704 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_187
timestamp 1698431365
transform 1 0 22288 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_203
timestamp 1698431365
transform 1 0 24080 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_207
timestamp 1698431365
transform 1 0 24528 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_209
timestamp 1698431365
transform 1 0 24752 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_212
timestamp 1698431365
transform 1 0 25088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698431365
transform 1 0 32256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_282
timestamp 1698431365
transform 1 0 32928 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_314
timestamp 1698431365
transform 1 0 36512 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_330
timestamp 1698431365
transform 1 0 38304 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_6
timestamp 1698431365
transform 1 0 2016 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_22
timestamp 1698431365
transform 1 0 3808 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_24
timestamp 1698431365
transform 1 0 4032 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_29
timestamp 1698431365
transform 1 0 4592 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_33
timestamp 1698431365
transform 1 0 5040 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_46
timestamp 1698431365
transform 1 0 6496 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_50
timestamp 1698431365
transform 1 0 6944 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_88
timestamp 1698431365
transform 1 0 11200 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_115
timestamp 1698431365
transform 1 0 14224 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_119
timestamp 1698431365
transform 1 0 14672 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_123
timestamp 1698431365
transform 1 0 15120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_169
timestamp 1698431365
transform 1 0 20272 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_173
timestamp 1698431365
transform 1 0 20720 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_177
timestamp 1698431365
transform 1 0 21168 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_241
timestamp 1698431365
transform 1 0 28336 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_247
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_311
timestamp 1698431365
transform 1 0 36176 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_317
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_325
timestamp 1698431365
transform 1 0 37744 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_329
timestamp 1698431365
transform 1 0 38192 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_6
timestamp 1698431365
transform 1 0 2016 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_22
timestamp 1698431365
transform 1 0 3808 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_32
timestamp 1698431365
transform 1 0 4928 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_38
timestamp 1698431365
transform 1 0 5600 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_48
timestamp 1698431365
transform 1 0 6720 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_64
timestamp 1698431365
transform 1 0 8512 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_68
timestamp 1698431365
transform 1 0 8960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_72
timestamp 1698431365
transform 1 0 9408 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_74
timestamp 1698431365
transform 1 0 9632 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_77
timestamp 1698431365
transform 1 0 9968 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_81
timestamp 1698431365
transform 1 0 10416 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_132
timestamp 1698431365
transform 1 0 16128 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_136
timestamp 1698431365
transform 1 0 16576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_158
timestamp 1698431365
transform 1 0 19040 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_166
timestamp 1698431365
transform 1 0 19936 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_168
timestamp 1698431365
transform 1 0 20160 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_171
timestamp 1698431365
transform 1 0 20496 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_190
timestamp 1698431365
transform 1 0 22624 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_206
timestamp 1698431365
transform 1 0 24416 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_212
timestamp 1698431365
transform 1 0 25088 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_276
timestamp 1698431365
transform 1 0 32256 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_282
timestamp 1698431365
transform 1 0 32928 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_314
timestamp 1698431365
transform 1 0 36512 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_330
timestamp 1698431365
transform 1 0 38304 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_6
timestamp 1698431365
transform 1 0 2016 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_14
timestamp 1698431365
transform 1 0 2912 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_30
timestamp 1698431365
transform 1 0 4704 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_32
timestamp 1698431365
transform 1 0 4928 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_37
timestamp 1698431365
transform 1 0 5488 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_51
timestamp 1698431365
transform 1 0 7056 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_94
timestamp 1698431365
transform 1 0 11872 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_102
timestamp 1698431365
transform 1 0 12768 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_104
timestamp 1698431365
transform 1 0 12992 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_107
timestamp 1698431365
transform 1 0 13328 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_94_131
timestamp 1698431365
transform 1 0 16016 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_163
timestamp 1698431365
transform 1 0 19600 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_171
timestamp 1698431365
transform 1 0 20496 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_211
timestamp 1698431365
transform 1 0 24976 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_215
timestamp 1698431365
transform 1 0 25424 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_94_219
timestamp 1698431365
transform 1 0 25872 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_235
timestamp 1698431365
transform 1 0 27664 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_243
timestamp 1698431365
transform 1 0 28560 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_247
timestamp 1698431365
transform 1 0 29008 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_311
timestamp 1698431365
transform 1 0 36176 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_317
timestamp 1698431365
transform 1 0 36848 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_325
timestamp 1698431365
transform 1 0 37744 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_329
timestamp 1698431365
transform 1 0 38192 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_60
timestamp 1698431365
transform 1 0 8064 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_80
timestamp 1698431365
transform 1 0 10304 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_84
timestamp 1698431365
transform 1 0 10752 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_88
timestamp 1698431365
transform 1 0 11200 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_91
timestamp 1698431365
transform 1 0 11536 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_119
timestamp 1698431365
transform 1 0 14672 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_131
timestamp 1698431365
transform 1 0 16016 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_135
timestamp 1698431365
transform 1 0 16464 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_139
timestamp 1698431365
transform 1 0 16912 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_95_142
timestamp 1698431365
transform 1 0 17248 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95_158
timestamp 1698431365
transform 1 0 19040 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_166
timestamp 1698431365
transform 1 0 19936 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_168
timestamp 1698431365
transform 1 0 20160 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_203
timestamp 1698431365
transform 1 0 24080 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_207
timestamp 1698431365
transform 1 0 24528 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_209
timestamp 1698431365
transform 1 0 24752 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_212
timestamp 1698431365
transform 1 0 25088 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_216
timestamp 1698431365
transform 1 0 25536 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_95_282
timestamp 1698431365
transform 1 0 32928 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_95_314
timestamp 1698431365
transform 1 0 36512 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_330
timestamp 1698431365
transform 1 0 38304 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_6
timestamp 1698431365
transform 1 0 2016 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_14
timestamp 1698431365
transform 1 0 2912 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_20
timestamp 1698431365
transform 1 0 3584 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_49
timestamp 1698431365
transform 1 0 6832 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_53
timestamp 1698431365
transform 1 0 7280 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_93
timestamp 1698431365
transform 1 0 11760 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_97
timestamp 1698431365
transform 1 0 12208 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_107
timestamp 1698431365
transform 1 0 13328 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_96_137
timestamp 1698431365
transform 1 0 16688 0 1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_153
timestamp 1698431365
transform 1 0 18480 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_161
timestamp 1698431365
transform 1 0 19376 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_96_198
timestamp 1698431365
transform 1 0 23520 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_230
timestamp 1698431365
transform 1 0 27104 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_238
timestamp 1698431365
transform 1 0 28000 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_242
timestamp 1698431365
transform 1 0 28448 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_244
timestamp 1698431365
transform 1 0 28672 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_247
timestamp 1698431365
transform 1 0 29008 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_311
timestamp 1698431365
transform 1 0 36176 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_317
timestamp 1698431365
transform 1 0 36848 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_325
timestamp 1698431365
transform 1 0 37744 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_329
timestamp 1698431365
transform 1 0 38192 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_38
timestamp 1698431365
transform 1 0 5600 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_42
timestamp 1698431365
transform 1 0 6048 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_46
timestamp 1698431365
transform 1 0 6496 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_50
timestamp 1698431365
transform 1 0 6944 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_52
timestamp 1698431365
transform 1 0 7168 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_67
timestamp 1698431365
transform 1 0 8848 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_69
timestamp 1698431365
transform 1 0 9072 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_97_72
timestamp 1698431365
transform 1 0 9408 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_80
timestamp 1698431365
transform 1 0 10304 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_84
timestamp 1698431365
transform 1 0 10752 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_142
timestamp 1698431365
transform 1 0 17248 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_97_146
timestamp 1698431365
transform 1 0 17696 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_97_162
timestamp 1698431365
transform 1 0 19488 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_170
timestamp 1698431365
transform 1 0 20384 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_173
timestamp 1698431365
transform 1 0 20720 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_177
timestamp 1698431365
transform 1 0 21168 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_179
timestamp 1698431365
transform 1 0 21392 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_97_192
timestamp 1698431365
transform 1 0 22848 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_208
timestamp 1698431365
transform 1 0 24640 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_212
timestamp 1698431365
transform 1 0 25088 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_276
timestamp 1698431365
transform 1 0 32256 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_282
timestamp 1698431365
transform 1 0 32928 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_97_314
timestamp 1698431365
transform 1 0 36512 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_330
timestamp 1698431365
transform 1 0 38304 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_98_6
timestamp 1698431365
transform 1 0 2016 0 1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_98_22
timestamp 1698431365
transform 1 0 3808 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_30
timestamp 1698431365
transform 1 0 4704 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_34
timestamp 1698431365
transform 1 0 5152 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_37
timestamp 1698431365
transform 1 0 5488 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_39
timestamp 1698431365
transform 1 0 5712 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_51
timestamp 1698431365
transform 1 0 7056 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_55
timestamp 1698431365
transform 1 0 7504 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_57
timestamp 1698431365
transform 1 0 7728 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_68
timestamp 1698431365
transform 1 0 8960 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_82
timestamp 1698431365
transform 1 0 10528 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_86
timestamp 1698431365
transform 1 0 10976 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_96
timestamp 1698431365
transform 1 0 12096 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_100
timestamp 1698431365
transform 1 0 12544 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_102
timestamp 1698431365
transform 1 0 12768 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_107
timestamp 1698431365
transform 1 0 13328 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_109
timestamp 1698431365
transform 1 0 13552 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_125
timestamp 1698431365
transform 1 0 15344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_127
timestamp 1698431365
transform 1 0 15568 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_164
timestamp 1698431365
transform 1 0 19712 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_168
timestamp 1698431365
transform 1 0 20160 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_172
timestamp 1698431365
transform 1 0 20608 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_174
timestamp 1698431365
transform 1 0 20832 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_98_177
timestamp 1698431365
transform 1 0 21168 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_241
timestamp 1698431365
transform 1 0 28336 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_98_247
timestamp 1698431365
transform 1 0 29008 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_311
timestamp 1698431365
transform 1 0 36176 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_98_317
timestamp 1698431365
transform 1 0 36848 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_325
timestamp 1698431365
transform 1 0 37744 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_329
timestamp 1698431365
transform 1 0 38192 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_99_6
timestamp 1698431365
transform 1 0 2016 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_99_22
timestamp 1698431365
transform 1 0 3808 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_30
timestamp 1698431365
transform 1 0 4704 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_90
timestamp 1698431365
transform 1 0 11424 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_103
timestamp 1698431365
transform 1 0 12880 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_107
timestamp 1698431365
transform 1 0 13328 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_110
timestamp 1698431365
transform 1 0 13664 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_114
timestamp 1698431365
transform 1 0 14112 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_128
timestamp 1698431365
transform 1 0 15680 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_165
timestamp 1698431365
transform 1 0 19824 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_169
timestamp 1698431365
transform 1 0 20272 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_99_173
timestamp 1698431365
transform 1 0 20720 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_181
timestamp 1698431365
transform 1 0 21616 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_183
timestamp 1698431365
transform 1 0 21840 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_197
timestamp 1698431365
transform 1 0 23408 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_99_201
timestamp 1698431365
transform 1 0 23856 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_209
timestamp 1698431365
transform 1 0 24752 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_212
timestamp 1698431365
transform 1 0 25088 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_276
timestamp 1698431365
transform 1 0 32256 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_99_282
timestamp 1698431365
transform 1 0 32928 0 -1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_99_314
timestamp 1698431365
transform 1 0 36512 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_330
timestamp 1698431365
transform 1 0 38304 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_100_6
timestamp 1698431365
transform 1 0 2016 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_22
timestamp 1698431365
transform 1 0 3808 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_34
timestamp 1698431365
transform 1 0 5152 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_37
timestamp 1698431365
transform 1 0 5488 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_43
timestamp 1698431365
transform 1 0 6160 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_100_47
timestamp 1698431365
transform 1 0 6608 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_100_63
timestamp 1698431365
transform 1 0 8400 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_71
timestamp 1698431365
transform 1 0 9296 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_74
timestamp 1698431365
transform 1 0 9632 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_100
timestamp 1698431365
transform 1 0 12544 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_104
timestamp 1698431365
transform 1 0 12992 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_107
timestamp 1698431365
transform 1 0 13328 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_113
timestamp 1698431365
transform 1 0 14000 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_128
timestamp 1698431365
transform 1 0 15680 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_177
timestamp 1698431365
transform 1 0 21168 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_181
timestamp 1698431365
transform 1 0 21616 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_183
timestamp 1698431365
transform 1 0 21840 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_100_194
timestamp 1698431365
transform 1 0 23072 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_100_226
timestamp 1698431365
transform 1 0 26656 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_242
timestamp 1698431365
transform 1 0 28448 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_244
timestamp 1698431365
transform 1 0 28672 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_100_247
timestamp 1698431365
transform 1 0 29008 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_311
timestamp 1698431365
transform 1 0 36176 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_100_317
timestamp 1698431365
transform 1 0 36848 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_325
timestamp 1698431365
transform 1 0 37744 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_329
timestamp 1698431365
transform 1 0 38192 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_46
timestamp 1698431365
transform 1 0 6496 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_50
timestamp 1698431365
transform 1 0 6944 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_54
timestamp 1698431365
transform 1 0 7392 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_58
timestamp 1698431365
transform 1 0 7840 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_66
timestamp 1698431365
transform 1 0 8736 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_72
timestamp 1698431365
transform 1 0 9408 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_80
timestamp 1698431365
transform 1 0 10304 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_92
timestamp 1698431365
transform 1 0 11648 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_112
timestamp 1698431365
transform 1 0 13888 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_119
timestamp 1698431365
transform 1 0 14672 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_123
timestamp 1698431365
transform 1 0 15120 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_125
timestamp 1698431365
transform 1 0 15344 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_128
timestamp 1698431365
transform 1 0 15680 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_139
timestamp 1698431365
transform 1 0 16912 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_154
timestamp 1698431365
transform 1 0 18592 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_101_158
timestamp 1698431365
transform 1 0 19040 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_212
timestamp 1698431365
transform 1 0 25088 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_216
timestamp 1698431365
transform 1 0 25536 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_101_220
timestamp 1698431365
transform 1 0 25984 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_101_252
timestamp 1698431365
transform 1 0 29568 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_268
timestamp 1698431365
transform 1 0 31360 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_276
timestamp 1698431365
transform 1 0 32256 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_101_282
timestamp 1698431365
transform 1 0 32928 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_101_314
timestamp 1698431365
transform 1 0 36512 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_330
timestamp 1698431365
transform 1 0 38304 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_102_6
timestamp 1698431365
transform 1 0 2016 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_14
timestamp 1698431365
transform 1 0 2912 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_31
timestamp 1698431365
transform 1 0 4816 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_37
timestamp 1698431365
transform 1 0 5488 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_54
timestamp 1698431365
transform 1 0 7392 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_58
timestamp 1698431365
transform 1 0 7840 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_68
timestamp 1698431365
transform 1 0 8960 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_102_72
timestamp 1698431365
transform 1 0 9408 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_88
timestamp 1698431365
transform 1 0 11200 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_163
timestamp 1698431365
transform 1 0 19600 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_167
timestamp 1698431365
transform 1 0 20048 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_171
timestamp 1698431365
transform 1 0 20496 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_102_177
timestamp 1698431365
transform 1 0 21168 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_185
timestamp 1698431365
transform 1 0 22064 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_187
timestamp 1698431365
transform 1 0 22288 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_102_195
timestamp 1698431365
transform 1 0 23184 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_102_227
timestamp 1698431365
transform 1 0 26768 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_243
timestamp 1698431365
transform 1 0 28560 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_102_247
timestamp 1698431365
transform 1 0 29008 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_311
timestamp 1698431365
transform 1 0 36176 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_102_317
timestamp 1698431365
transform 1 0 36848 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_325
timestamp 1698431365
transform 1 0 37744 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_329
timestamp 1698431365
transform 1 0 38192 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_103_6
timestamp 1698431365
transform 1 0 2016 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_14
timestamp 1698431365
transform 1 0 2912 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_18
timestamp 1698431365
transform 1 0 3360 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_54
timestamp 1698431365
transform 1 0 7392 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_68
timestamp 1698431365
transform 1 0 8960 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_72
timestamp 1698431365
transform 1 0 9408 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_103_77
timestamp 1698431365
transform 1 0 9968 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_95
timestamp 1698431365
transform 1 0 11984 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_112
timestamp 1698431365
transform 1 0 13888 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_114
timestamp 1698431365
transform 1 0 14112 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_120
timestamp 1698431365
transform 1 0 14784 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_103_124
timestamp 1698431365
transform 1 0 15232 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_142
timestamp 1698431365
transform 1 0 17248 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_146
timestamp 1698431365
transform 1 0 17696 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_150
timestamp 1698431365
transform 1 0 18144 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_168
timestamp 1698431365
transform 1 0 20160 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_170
timestamp 1698431365
transform 1 0 20384 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_103_188
timestamp 1698431365
transform 1 0 22400 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_204
timestamp 1698431365
transform 1 0 24192 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_208
timestamp 1698431365
transform 1 0 24640 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_212
timestamp 1698431365
transform 1 0 25088 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_276
timestamp 1698431365
transform 1 0 32256 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_103_282
timestamp 1698431365
transform 1 0 32928 0 -1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_103_314
timestamp 1698431365
transform 1 0 36512 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_330
timestamp 1698431365
transform 1 0 38304 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_104_2
timestamp 1698431365
transform 1 0 1568 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104_18
timestamp 1698431365
transform 1 0 3360 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_26
timestamp 1698431365
transform 1 0 4256 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_30
timestamp 1698431365
transform 1 0 4704 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_33
timestamp 1698431365
transform 1 0 5040 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_37
timestamp 1698431365
transform 1 0 5488 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_41
timestamp 1698431365
transform 1 0 5936 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_43
timestamp 1698431365
transform 1 0 6160 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_78
timestamp 1698431365
transform 1 0 10080 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_82
timestamp 1698431365
transform 1 0 10528 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104_86
timestamp 1698431365
transform 1 0 10976 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_94
timestamp 1698431365
transform 1 0 11872 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_98
timestamp 1698431365
transform 1 0 12320 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_101
timestamp 1698431365
transform 1 0 12656 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_107
timestamp 1698431365
transform 1 0 13328 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_104_119
timestamp 1698431365
transform 1 0 14672 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104_135
timestamp 1698431365
transform 1 0 16464 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_143
timestamp 1698431365
transform 1 0 17360 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_147
timestamp 1698431365
transform 1 0 17808 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_104_151
timestamp 1698431365
transform 1 0 18256 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_167
timestamp 1698431365
transform 1 0 20048 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_171
timestamp 1698431365
transform 1 0 20496 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104_192
timestamp 1698431365
transform 1 0 22848 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_104_224
timestamp 1698431365
transform 1 0 26432 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_240
timestamp 1698431365
transform 1 0 28224 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_244
timestamp 1698431365
transform 1 0 28672 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_104_247
timestamp 1698431365
transform 1 0 29008 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_311
timestamp 1698431365
transform 1 0 36176 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104_317
timestamp 1698431365
transform 1 0 36848 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_325
timestamp 1698431365
transform 1 0 37744 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_329
timestamp 1698431365
transform 1 0 38192 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_105_6
timestamp 1698431365
transform 1 0 2016 0 -1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_105_38
timestamp 1698431365
transform 1 0 5600 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_56
timestamp 1698431365
transform 1 0 7616 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_64
timestamp 1698431365
transform 1 0 8512 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_68
timestamp 1698431365
transform 1 0 8960 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_72
timestamp 1698431365
transform 1 0 9408 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_82
timestamp 1698431365
transform 1 0 10528 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_105_86
timestamp 1698431365
transform 1 0 10976 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_102
timestamp 1698431365
transform 1 0 12768 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_106
timestamp 1698431365
transform 1 0 13216 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_108
timestamp 1698431365
transform 1 0 13440 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_111
timestamp 1698431365
transform 1 0 13776 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_113
timestamp 1698431365
transform 1 0 14000 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_116
timestamp 1698431365
transform 1 0 14336 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_130
timestamp 1698431365
transform 1 0 15904 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_142
timestamp 1698431365
transform 1 0 17248 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_152
timestamp 1698431365
transform 1 0 18368 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_156
timestamp 1698431365
transform 1 0 18816 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_164
timestamp 1698431365
transform 1 0 19712 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_200
timestamp 1698431365
transform 1 0 23744 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_204
timestamp 1698431365
transform 1 0 24192 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_208
timestamp 1698431365
transform 1 0 24640 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_212
timestamp 1698431365
transform 1 0 25088 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_276
timestamp 1698431365
transform 1 0 32256 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_105_282
timestamp 1698431365
transform 1 0 32928 0 -1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_105_314
timestamp 1698431365
transform 1 0 36512 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_330
timestamp 1698431365
transform 1 0 38304 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_106_6
timestamp 1698431365
transform 1 0 2016 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_106_22
timestamp 1698431365
transform 1 0 3808 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_30
timestamp 1698431365
transform 1 0 4704 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_34
timestamp 1698431365
transform 1 0 5152 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_106_37
timestamp 1698431365
transform 1 0 5488 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_45
timestamp 1698431365
transform 1 0 6384 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_49
timestamp 1698431365
transform 1 0 6832 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_51
timestamp 1698431365
transform 1 0 7056 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_69
timestamp 1698431365
transform 1 0 9072 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_73
timestamp 1698431365
transform 1 0 9520 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_83
timestamp 1698431365
transform 1 0 10640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_87
timestamp 1698431365
transform 1 0 11088 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_91
timestamp 1698431365
transform 1 0 11536 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_97
timestamp 1698431365
transform 1 0 12208 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_101
timestamp 1698431365
transform 1 0 12656 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_115
timestamp 1698431365
transform 1 0 14224 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_106_165
timestamp 1698431365
transform 1 0 19824 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_173
timestamp 1698431365
transform 1 0 20720 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_177
timestamp 1698431365
transform 1 0 21168 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_241
timestamp 1698431365
transform 1 0 28336 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_247
timestamp 1698431365
transform 1 0 29008 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_311
timestamp 1698431365
transform 1 0 36176 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_106_317
timestamp 1698431365
transform 1 0 36848 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_325
timestamp 1698431365
transform 1 0 37744 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_329
timestamp 1698431365
transform 1 0 38192 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107_2
timestamp 1698431365
transform 1 0 1568 0 -1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_34
timestamp 1698431365
transform 1 0 5152 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_72
timestamp 1698431365
transform 1 0 9408 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_93
timestamp 1698431365
transform 1 0 11760 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_128
timestamp 1698431365
transform 1 0 15680 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_132
timestamp 1698431365
transform 1 0 16128 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_136
timestamp 1698431365
transform 1 0 16576 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_176
timestamp 1698431365
transform 1 0 21056 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_107_180
timestamp 1698431365
transform 1 0 21504 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107_196
timestamp 1698431365
transform 1 0 23296 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_204
timestamp 1698431365
transform 1 0 24192 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_208
timestamp 1698431365
transform 1 0 24640 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_212
timestamp 1698431365
transform 1 0 25088 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_276
timestamp 1698431365
transform 1 0 32256 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107_282
timestamp 1698431365
transform 1 0 32928 0 -1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_107_314
timestamp 1698431365
transform 1 0 36512 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_330
timestamp 1698431365
transform 1 0 38304 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_108_6
timestamp 1698431365
transform 1 0 2016 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_108_22
timestamp 1698431365
transform 1 0 3808 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_30
timestamp 1698431365
transform 1 0 4704 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_34
timestamp 1698431365
transform 1 0 5152 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_108_37
timestamp 1698431365
transform 1 0 5488 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_108_53
timestamp 1698431365
transform 1 0 7280 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_61
timestamp 1698431365
transform 1 0 8176 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_65
timestamp 1698431365
transform 1 0 8624 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_103
timestamp 1698431365
transform 1 0 12880 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_108_122
timestamp 1698431365
transform 1 0 15008 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_108_154
timestamp 1698431365
transform 1 0 18592 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_170
timestamp 1698431365
transform 1 0 20384 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_174
timestamp 1698431365
transform 1 0 20832 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_108_177
timestamp 1698431365
transform 1 0 21168 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_241
timestamp 1698431365
transform 1 0 28336 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_108_247
timestamp 1698431365
transform 1 0 29008 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_311
timestamp 1698431365
transform 1 0 36176 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_108_317
timestamp 1698431365
transform 1 0 36848 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_325
timestamp 1698431365
transform 1 0 37744 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_329
timestamp 1698431365
transform 1 0 38192 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_109_6
timestamp 1698431365
transform 1 0 2016 0 -1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_109_38
timestamp 1698431365
transform 1 0 5600 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_109_54
timestamp 1698431365
transform 1 0 7392 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_62
timestamp 1698431365
transform 1 0 8288 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_65
timestamp 1698431365
transform 1 0 8624 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_69
timestamp 1698431365
transform 1 0 9072 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_106
timestamp 1698431365
transform 1 0 13216 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_110
timestamp 1698431365
transform 1 0 13664 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_109_114
timestamp 1698431365
transform 1 0 14112 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_109_130
timestamp 1698431365
transform 1 0 15904 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_138
timestamp 1698431365
transform 1 0 16800 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_142
timestamp 1698431365
transform 1 0 17248 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_206
timestamp 1698431365
transform 1 0 24416 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_212
timestamp 1698431365
transform 1 0 25088 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_276
timestamp 1698431365
transform 1 0 32256 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_109_282
timestamp 1698431365
transform 1 0 32928 0 -1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_109_314
timestamp 1698431365
transform 1 0 36512 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_330
timestamp 1698431365
transform 1 0 38304 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_110_6
timestamp 1698431365
transform 1 0 2016 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_110_22
timestamp 1698431365
transform 1 0 3808 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_30
timestamp 1698431365
transform 1 0 4704 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_34
timestamp 1698431365
transform 1 0 5152 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_37
timestamp 1698431365
transform 1 0 5488 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_101
timestamp 1698431365
transform 1 0 12656 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_107
timestamp 1698431365
transform 1 0 13328 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_111
timestamp 1698431365
transform 1 0 13776 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_177
timestamp 1698431365
transform 1 0 21168 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_241
timestamp 1698431365
transform 1 0 28336 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_247
timestamp 1698431365
transform 1 0 29008 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_311
timestamp 1698431365
transform 1 0 36176 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_110_317
timestamp 1698431365
transform 1 0 36848 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_325
timestamp 1698431365
transform 1 0 37744 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_329
timestamp 1698431365
transform 1 0 38192 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_2
timestamp 1698431365
transform 1 0 1568 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_66
timestamp 1698431365
transform 1 0 8736 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_72
timestamp 1698431365
transform 1 0 9408 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_136
timestamp 1698431365
transform 1 0 16576 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_142
timestamp 1698431365
transform 1 0 17248 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_206
timestamp 1698431365
transform 1 0 24416 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_212
timestamp 1698431365
transform 1 0 25088 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_276
timestamp 1698431365
transform 1 0 32256 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_111_282
timestamp 1698431365
transform 1 0 32928 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_111_314
timestamp 1698431365
transform 1 0 36512 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_330
timestamp 1698431365
transform 1 0 38304 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_112_6
timestamp 1698431365
transform 1 0 2016 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_112_22
timestamp 1698431365
transform 1 0 3808 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_30
timestamp 1698431365
transform 1 0 4704 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_34
timestamp 1698431365
transform 1 0 5152 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_37
timestamp 1698431365
transform 1 0 5488 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_101
timestamp 1698431365
transform 1 0 12656 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_107
timestamp 1698431365
transform 1 0 13328 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_171
timestamp 1698431365
transform 1 0 20496 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_177
timestamp 1698431365
transform 1 0 21168 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_241
timestamp 1698431365
transform 1 0 28336 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_247
timestamp 1698431365
transform 1 0 29008 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_311
timestamp 1698431365
transform 1 0 36176 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_112_317
timestamp 1698431365
transform 1 0 36848 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_325
timestamp 1698431365
transform 1 0 37744 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_329
timestamp 1698431365
transform 1 0 38192 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_6
timestamp 1698431365
transform 1 0 2016 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_72
timestamp 1698431365
transform 1 0 9408 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_136
timestamp 1698431365
transform 1 0 16576 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_142
timestamp 1698431365
transform 1 0 17248 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_206
timestamp 1698431365
transform 1 0 24416 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_212
timestamp 1698431365
transform 1 0 25088 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_276
timestamp 1698431365
transform 1 0 32256 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_113_282
timestamp 1698431365
transform 1 0 32928 0 -1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_113_314
timestamp 1698431365
transform 1 0 36512 0 -1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_330
timestamp 1698431365
transform 1 0 38304 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_114_2
timestamp 1698431365
transform 1 0 1568 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_34
timestamp 1698431365
transform 1 0 5152 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_37
timestamp 1698431365
transform 1 0 5488 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_101
timestamp 1698431365
transform 1 0 12656 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_107
timestamp 1698431365
transform 1 0 13328 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_171
timestamp 1698431365
transform 1 0 20496 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_177
timestamp 1698431365
transform 1 0 21168 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_241
timestamp 1698431365
transform 1 0 28336 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_247
timestamp 1698431365
transform 1 0 29008 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_311
timestamp 1698431365
transform 1 0 36176 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_114_317
timestamp 1698431365
transform 1 0 36848 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_325
timestamp 1698431365
transform 1 0 37744 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_329
timestamp 1698431365
transform 1 0 38192 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_6
timestamp 1698431365
transform 1 0 2016 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_72
timestamp 1698431365
transform 1 0 9408 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_136
timestamp 1698431365
transform 1 0 16576 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_142
timestamp 1698431365
transform 1 0 17248 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_206
timestamp 1698431365
transform 1 0 24416 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_212
timestamp 1698431365
transform 1 0 25088 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_276
timestamp 1698431365
transform 1 0 32256 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_115_282
timestamp 1698431365
transform 1 0 32928 0 -1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_115_314
timestamp 1698431365
transform 1 0 36512 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_330
timestamp 1698431365
transform 1 0 38304 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_116_6
timestamp 1698431365
transform 1 0 2016 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_22
timestamp 1698431365
transform 1 0 3808 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_30
timestamp 1698431365
transform 1 0 4704 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_34
timestamp 1698431365
transform 1 0 5152 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_37
timestamp 1698431365
transform 1 0 5488 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_101
timestamp 1698431365
transform 1 0 12656 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_107
timestamp 1698431365
transform 1 0 13328 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_171
timestamp 1698431365
transform 1 0 20496 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_177
timestamp 1698431365
transform 1 0 21168 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_241
timestamp 1698431365
transform 1 0 28336 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_247
timestamp 1698431365
transform 1 0 29008 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_311
timestamp 1698431365
transform 1 0 36176 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_317
timestamp 1698431365
transform 1 0 36848 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_325
timestamp 1698431365
transform 1 0 37744 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_329
timestamp 1698431365
transform 1 0 38192 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_2
timestamp 1698431365
transform 1 0 1568 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_66
timestamp 1698431365
transform 1 0 8736 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_72
timestamp 1698431365
transform 1 0 9408 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_136
timestamp 1698431365
transform 1 0 16576 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_142
timestamp 1698431365
transform 1 0 17248 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_206
timestamp 1698431365
transform 1 0 24416 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_212
timestamp 1698431365
transform 1 0 25088 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_276
timestamp 1698431365
transform 1 0 32256 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_117_282
timestamp 1698431365
transform 1 0 32928 0 -1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_117_314
timestamp 1698431365
transform 1 0 36512 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_330
timestamp 1698431365
transform 1 0 38304 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_118_6
timestamp 1698431365
transform 1 0 2016 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_22
timestamp 1698431365
transform 1 0 3808 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_30
timestamp 1698431365
transform 1 0 4704 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_36
timestamp 1698431365
transform 1 0 5376 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_70
timestamp 1698431365
transform 1 0 9184 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_104
timestamp 1698431365
transform 1 0 12992 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_138
timestamp 1698431365
transform 1 0 16800 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_172
timestamp 1698431365
transform 1 0 20608 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_206
timestamp 1698431365
transform 1 0 24416 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_240
timestamp 1698431365
transform 1 0 28224 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_248
timestamp 1698431365
transform 1 0 29120 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_252
timestamp 1698431365
transform 1 0 29568 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_261
timestamp 1698431365
transform 1 0 30576 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_269
timestamp 1698431365
transform 1 0 31472 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_271
timestamp 1698431365
transform 1 0 31696 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_274
timestamp 1698431365
transform 1 0 32032 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_118_308
timestamp 1698431365
transform 1 0 35840 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_324
timestamp 1698431365
transform 1 0 37632 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_328
timestamp 1698431365
transform 1 0 38080 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_330
timestamp 1698431365
transform 1 0 38304 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  hold1 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28672 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold3
timestamp 1698431365
transform -1 0 18592 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold4
timestamp 1698431365
transform -1 0 28448 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold5
timestamp 1698431365
transform 1 0 13664 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold6
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  hold7 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output1
timestamp 1698431365
transform -1 0 30576 0 1 95648
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_24 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2016 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_25
timestamp 1698431365
transform -1 0 2016 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_26
timestamp 1698431365
transform -1 0 2016 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_27
timestamp 1698431365
transform -1 0 2016 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_28
timestamp 1698431365
transform -1 0 2016 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_29
timestamp 1698431365
transform -1 0 2016 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_30
timestamp 1698431365
transform -1 0 2016 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_31
timestamp 1698431365
transform -1 0 2016 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_32
timestamp 1698431365
transform -1 0 2016 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_33
timestamp 1698431365
transform -1 0 2016 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_34
timestamp 1698431365
transform -1 0 2016 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_35
timestamp 1698431365
transform -1 0 2016 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_36
timestamp 1698431365
transform -1 0 2016 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_37
timestamp 1698431365
transform -1 0 2016 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_38
timestamp 1698431365
transform -1 0 2016 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_39
timestamp 1698431365
transform -1 0 2016 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_40
timestamp 1698431365
transform -1 0 2016 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_41
timestamp 1698431365
transform -1 0 2016 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_42
timestamp 1698431365
transform -1 0 2016 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_43
timestamp 1698431365
transform -1 0 2464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_44
timestamp 1698431365
transform -1 0 2016 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_45
timestamp 1698431365
transform -1 0 2016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_46
timestamp 1698431365
transform -1 0 2016 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_47
timestamp 1698431365
transform -1 0 2016 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_48
timestamp 1698431365
transform -1 0 2016 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_49
timestamp 1698431365
transform -1 0 2016 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_50
timestamp 1698431365
transform -1 0 2464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_51
timestamp 1698431365
transform -1 0 2016 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_52
timestamp 1698431365
transform -1 0 2016 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_53
timestamp 1698431365
transform -1 0 2016 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_54
timestamp 1698431365
transform -1 0 2016 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_55
timestamp 1698431365
transform -1 0 2016 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  peri_top_56
timestamp 1698431365
transform -1 0 2016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_119 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_120
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_121
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_122
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_123
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_124
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_125
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_126
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_127
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_128
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_129
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_130
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_131
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_132
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_133
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_134
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_135
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_136
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_137
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_138
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_139
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_140
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_141
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_142
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_143
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_144
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_145
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_146
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_147
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_148
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_149
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_150
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_151
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_152
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_153
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_154
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_155
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_156
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_157
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_158
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_159
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_160
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_161
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_162
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 38640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_163
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_164
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 38640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_165
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 38640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_166
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 38640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_167
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 38640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_168
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 38640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_169
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 38640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_170
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 38640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_171
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 38640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_172
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 38640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_173
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 38640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_174
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 38640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_175
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 38640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_176
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 38640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_177
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 38640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_178
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 38640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_179
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 38640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_180
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 38640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_181
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 38640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_182
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 38640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_183
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 38640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_184
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 38640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_185
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 38640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_186
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 38640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_187
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 38640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_188
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 38640 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_189
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 38640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_190
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 38640 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_191
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 38640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_192
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 38640 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_193
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 38640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_194
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 38640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_195
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 38640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_196
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 38640 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_197
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 38640 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_198
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 38640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_199
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 38640 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_200
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 38640 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_201
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 38640 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_202
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 38640 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_203
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 38640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_204
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 38640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_205
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 38640 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_206
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 38640 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_207
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 38640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_208
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 38640 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_209
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 38640 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_210
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 38640 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_211
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 38640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_212
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 38640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Left_213
timestamp 1698431365
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Right_94
timestamp 1698431365
transform -1 0 38640 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Left_214
timestamp 1698431365
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Right_95
timestamp 1698431365
transform -1 0 38640 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Left_215
timestamp 1698431365
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Right_96
timestamp 1698431365
transform -1 0 38640 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Left_216
timestamp 1698431365
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Right_97
timestamp 1698431365
transform -1 0 38640 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Left_217
timestamp 1698431365
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Right_98
timestamp 1698431365
transform -1 0 38640 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Left_218
timestamp 1698431365
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Right_99
timestamp 1698431365
transform -1 0 38640 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Left_219
timestamp 1698431365
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Right_100
timestamp 1698431365
transform -1 0 38640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Left_220
timestamp 1698431365
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Right_101
timestamp 1698431365
transform -1 0 38640 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Left_221
timestamp 1698431365
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Right_102
timestamp 1698431365
transform -1 0 38640 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Left_222
timestamp 1698431365
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Right_103
timestamp 1698431365
transform -1 0 38640 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Left_223
timestamp 1698431365
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Right_104
timestamp 1698431365
transform -1 0 38640 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Left_224
timestamp 1698431365
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Right_105
timestamp 1698431365
transform -1 0 38640 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Left_225
timestamp 1698431365
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Right_106
timestamp 1698431365
transform -1 0 38640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Left_226
timestamp 1698431365
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Right_107
timestamp 1698431365
transform -1 0 38640 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Left_227
timestamp 1698431365
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Right_108
timestamp 1698431365
transform -1 0 38640 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Left_228
timestamp 1698431365
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Right_109
timestamp 1698431365
transform -1 0 38640 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Left_229
timestamp 1698431365
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Right_110
timestamp 1698431365
transform -1 0 38640 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Left_230
timestamp 1698431365
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Right_111
timestamp 1698431365
transform -1 0 38640 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Left_231
timestamp 1698431365
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Right_112
timestamp 1698431365
transform -1 0 38640 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Left_232
timestamp 1698431365
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Right_113
timestamp 1698431365
transform -1 0 38640 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Left_233
timestamp 1698431365
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Right_114
timestamp 1698431365
transform -1 0 38640 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Left_234
timestamp 1698431365
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Right_115
timestamp 1698431365
transform -1 0 38640 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Left_235
timestamp 1698431365
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Right_116
timestamp 1698431365
transform -1 0 38640 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Left_236
timestamp 1698431365
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Right_117
timestamp 1698431365
transform -1 0 38640 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Left_237
timestamp 1698431365
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Right_118
timestamp 1698431365
transform -1 0 38640 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_238 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_239
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_240
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_241
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_242
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_243
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_244
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_245
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_246
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_247
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_248
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_249
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_250
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_251
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_252
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_253
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_254
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_255
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_256
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_257
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_258
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_259
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_260
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_261
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_262
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_263
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_264
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_265
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_266
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_267
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_268
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_269
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_270
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_271
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_272
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_273
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_274
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_275
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_276
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_277
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_278
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_279
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_280
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_281
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_282
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_283
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_284
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_285
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_286
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_287
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_288
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_289
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_290
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_291
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_292
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_293
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_294
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_295
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_296
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_297
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_298
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_299
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_300
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_301
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_302
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_303
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_304
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_305
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_306
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_307
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_308
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_309
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_310
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_311
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_312
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_313
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_314
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_315
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_316
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_317
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_318
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_319
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_320
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_321
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_322
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_323
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_324
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_325
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_326
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_327
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_328
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_329
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_330
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_331
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_332
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_333
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_334
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_335
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_336
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_337
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_338
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_339
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_340
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_341
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_342
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_343
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_344
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_345
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_346
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_347
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_348
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_349
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_350
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_351
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_352
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_353
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_354
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_355
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_356
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_357
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_358
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_359
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_360
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_361
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_362
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_363
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_364
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_365
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_366
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_367
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_368
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_369
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_370
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_371
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_372
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_373
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_374
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_375
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_376
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_377
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_378
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_379
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_380
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_381
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_382
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_383
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_384
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_385
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_386
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_387
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_388
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_389
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_390
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_391
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_392
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_393
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_394
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_395
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_396
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_397
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_398
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_399
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_400
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_401
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_402
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_403
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_404
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_405
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_406
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_407
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_408
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_409
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_410
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_411
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_412
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_416
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_417
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_422
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_427
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_428
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_429
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_431
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_432
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_433
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_434
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_435
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_436
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_437
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_438
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_439
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_440
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_441
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_442
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_443
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_444
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_445
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_446
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_447
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_448
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_449
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_450
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_451
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_452
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_453
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_454
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_455
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_456
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_457
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_458
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_459
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_460
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_461
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_462
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_463
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_464
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_465
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_466
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_467
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_468
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_469
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_470
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_471
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_472
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_473
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_474
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_475
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_476
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_477
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_478
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_479
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_480
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_481
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_482
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_483
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_484
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_485
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_486
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_487
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_488
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_489
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_490
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_491
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_492
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_493
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_494
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_495
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_496
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_497
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_498
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_499
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_500
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_501
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_502
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_503
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_504
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_505
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_506
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_507
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_508
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_509
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_510
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_511
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_512
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_513
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_514
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_515
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_516
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_517
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_518
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_519
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_520
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_521
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_522
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_523
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_524
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_525
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_526
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_527
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_528
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_529
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_530
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_531
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_532
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_533
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_534
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_535
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_536
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_537
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_538
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_539
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_540
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_541
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_542
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_543
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_544
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_545
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_546
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_547
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_548
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_549
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_550
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_551
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_552
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_553
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_554
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_555
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_556
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_557
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_558
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_559
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_560
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_561
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_562
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_563
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_564
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_565
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_566
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_567
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_568
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_569
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_570
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_571
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_572
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_573
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_574
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_575
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_576
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_577
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_578
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_579
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_580
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_581
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_582
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_583
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_584
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_585
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_586
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_587
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_588
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_589
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_590
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_591
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_592
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_593
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_594
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_595
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_596
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_597
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_598
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_599
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_600
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_601
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_602
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_603
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_604
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_605
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_606
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_607
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_608
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_609
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_610
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_611
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_612
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_613
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_614
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_615
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_616
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_617
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_618
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_619
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_620
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_621
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_622
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_623
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_624
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_625
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_626
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_627
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_628
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_629
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_630
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_631
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_632
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_633
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_634
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_635
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_636
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_637
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_638
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_639
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_640
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_641
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_642
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_643
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_644
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_645
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_646
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_647
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_648
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_649
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_650
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_651
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_652
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_653
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_654
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_655
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_656
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_657
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_658
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_659
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_660
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_661
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_662
timestamp 1698431365
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_663
timestamp 1698431365
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_664
timestamp 1698431365
transform 1 0 32704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_665
timestamp 1698431365
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_666
timestamp 1698431365
transform 1 0 13104 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_667
timestamp 1698431365
transform 1 0 20944 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_668
timestamp 1698431365
transform 1 0 28784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_669
timestamp 1698431365
transform 1 0 36624 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_670
timestamp 1698431365
transform 1 0 9184 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_671
timestamp 1698431365
transform 1 0 17024 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_672
timestamp 1698431365
transform 1 0 24864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_673
timestamp 1698431365
transform 1 0 32704 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_674
timestamp 1698431365
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_675
timestamp 1698431365
transform 1 0 13104 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_676
timestamp 1698431365
transform 1 0 20944 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_677
timestamp 1698431365
transform 1 0 28784 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_678
timestamp 1698431365
transform 1 0 36624 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_679
timestamp 1698431365
transform 1 0 9184 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_680
timestamp 1698431365
transform 1 0 17024 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_681
timestamp 1698431365
transform 1 0 24864 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_682
timestamp 1698431365
transform 1 0 32704 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_683
timestamp 1698431365
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_684
timestamp 1698431365
transform 1 0 13104 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_685
timestamp 1698431365
transform 1 0 20944 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_686
timestamp 1698431365
transform 1 0 28784 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_687
timestamp 1698431365
transform 1 0 36624 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_688
timestamp 1698431365
transform 1 0 9184 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_689
timestamp 1698431365
transform 1 0 17024 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_690
timestamp 1698431365
transform 1 0 24864 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_691
timestamp 1698431365
transform 1 0 32704 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_692
timestamp 1698431365
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_693
timestamp 1698431365
transform 1 0 13104 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_694
timestamp 1698431365
transform 1 0 20944 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_695
timestamp 1698431365
transform 1 0 28784 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_696
timestamp 1698431365
transform 1 0 36624 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_697
timestamp 1698431365
transform 1 0 9184 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_698
timestamp 1698431365
transform 1 0 17024 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_699
timestamp 1698431365
transform 1 0 24864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_700
timestamp 1698431365
transform 1 0 32704 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_701
timestamp 1698431365
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_702
timestamp 1698431365
transform 1 0 13104 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_703
timestamp 1698431365
transform 1 0 20944 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_704
timestamp 1698431365
transform 1 0 28784 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_705
timestamp 1698431365
transform 1 0 36624 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_706
timestamp 1698431365
transform 1 0 9184 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_707
timestamp 1698431365
transform 1 0 17024 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_708
timestamp 1698431365
transform 1 0 24864 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_709
timestamp 1698431365
transform 1 0 32704 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_710
timestamp 1698431365
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_711
timestamp 1698431365
transform 1 0 13104 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_712
timestamp 1698431365
transform 1 0 20944 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_713
timestamp 1698431365
transform 1 0 28784 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_714
timestamp 1698431365
transform 1 0 36624 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_715
timestamp 1698431365
transform 1 0 9184 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_716
timestamp 1698431365
transform 1 0 17024 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_717
timestamp 1698431365
transform 1 0 24864 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_718
timestamp 1698431365
transform 1 0 32704 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_719
timestamp 1698431365
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_720
timestamp 1698431365
transform 1 0 13104 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_721
timestamp 1698431365
transform 1 0 20944 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_722
timestamp 1698431365
transform 1 0 28784 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_723
timestamp 1698431365
transform 1 0 36624 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_724
timestamp 1698431365
transform 1 0 9184 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_725
timestamp 1698431365
transform 1 0 17024 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_726
timestamp 1698431365
transform 1 0 24864 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_727
timestamp 1698431365
transform 1 0 32704 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_728
timestamp 1698431365
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_729
timestamp 1698431365
transform 1 0 13104 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_730
timestamp 1698431365
transform 1 0 20944 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_731
timestamp 1698431365
transform 1 0 28784 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_732
timestamp 1698431365
transform 1 0 36624 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_733
timestamp 1698431365
transform 1 0 9184 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_734
timestamp 1698431365
transform 1 0 17024 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_735
timestamp 1698431365
transform 1 0 24864 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_736
timestamp 1698431365
transform 1 0 32704 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_737
timestamp 1698431365
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_738
timestamp 1698431365
transform 1 0 13104 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_739
timestamp 1698431365
transform 1 0 20944 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_740
timestamp 1698431365
transform 1 0 28784 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_741
timestamp 1698431365
transform 1 0 36624 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_742
timestamp 1698431365
transform 1 0 9184 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_743
timestamp 1698431365
transform 1 0 17024 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_744
timestamp 1698431365
transform 1 0 24864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_745
timestamp 1698431365
transform 1 0 32704 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_746
timestamp 1698431365
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_747
timestamp 1698431365
transform 1 0 13104 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_748
timestamp 1698431365
transform 1 0 20944 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_749
timestamp 1698431365
transform 1 0 28784 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_750
timestamp 1698431365
transform 1 0 36624 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_751
timestamp 1698431365
transform 1 0 9184 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_752
timestamp 1698431365
transform 1 0 17024 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_753
timestamp 1698431365
transform 1 0 24864 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_754
timestamp 1698431365
transform 1 0 32704 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_755
timestamp 1698431365
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_756
timestamp 1698431365
transform 1 0 13104 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_757
timestamp 1698431365
transform 1 0 20944 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_758
timestamp 1698431365
transform 1 0 28784 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_759
timestamp 1698431365
transform 1 0 36624 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_760
timestamp 1698431365
transform 1 0 9184 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_761
timestamp 1698431365
transform 1 0 17024 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_762
timestamp 1698431365
transform 1 0 24864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_763
timestamp 1698431365
transform 1 0 32704 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_764
timestamp 1698431365
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_765
timestamp 1698431365
transform 1 0 13104 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_766
timestamp 1698431365
transform 1 0 20944 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_767
timestamp 1698431365
transform 1 0 28784 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_768
timestamp 1698431365
transform 1 0 36624 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_769
timestamp 1698431365
transform 1 0 9184 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_770
timestamp 1698431365
transform 1 0 17024 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_771
timestamp 1698431365
transform 1 0 24864 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_772
timestamp 1698431365
transform 1 0 32704 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_773
timestamp 1698431365
transform 1 0 5152 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_774
timestamp 1698431365
transform 1 0 8960 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_775
timestamp 1698431365
transform 1 0 12768 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_776
timestamp 1698431365
transform 1 0 16576 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_777
timestamp 1698431365
transform 1 0 20384 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_778
timestamp 1698431365
transform 1 0 24192 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_779
timestamp 1698431365
transform 1 0 28000 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_780
timestamp 1698431365
transform 1 0 31808 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_781
timestamp 1698431365
transform 1 0 35616 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  u_rst_sync._1__59 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rst_sync._1_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21056 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rst_sync._2_
timestamp 1698431365
transform 1 0 21056 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_rst_sync.u_buf.genblk1.u_mux_22
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rst_sync.u_buf.genblk1.u_mux open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27216 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_async_reg_bus._092_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_async_reg_bus._093_
timestamp 1698431365
transform -1 0 21616 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_async_reg_bus._094_
timestamp 1698431365
transform -1 0 20048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_async_reg_bus._095_
timestamp 1698431365
transform -1 0 7616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_async_reg_bus._096_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20496 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_async_reg_bus._097_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_async_reg_bus._098_
timestamp 1698431365
transform -1 0 17024 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_async_reg_bus._099_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_rtc.u_async_reg_bus._099__23
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_async_reg_bus._100_
timestamp 1698431365
transform -1 0 17808 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_async_reg_bus._101_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_async_reg_bus._102_
timestamp 1698431365
transform 1 0 6160 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_async_reg_bus._103_
timestamp 1698431365
transform 1 0 6384 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_async_reg_bus._104_
timestamp 1698431365
transform -1 0 6048 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_async_reg_bus._105_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_async_reg_bus._106_
timestamp 1698431365
transform -1 0 3808 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_async_reg_bus._107_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6048 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_async_reg_bus._108_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_async_reg_bus._109_
timestamp 1698431365
transform 1 0 7392 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_async_reg_bus._110_
timestamp 1698431365
transform -1 0 8288 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_async_reg_bus._111_
timestamp 1698431365
transform 1 0 8288 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_async_reg_bus._112_
timestamp 1698431365
transform 1 0 8400 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_async_reg_bus._113_
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_async_reg_bus._181_
timestamp 1698431365
transform -1 0 18256 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_async_reg_bus._182_
timestamp 1698431365
transform -1 0 19264 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_async_reg_bus._183_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._184_
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._185_
timestamp 1698431365
transform 1 0 9296 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._186_
timestamp 1698431365
transform -1 0 14896 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._187_
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._188_
timestamp 1698431365
transform 1 0 13216 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._189_
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._190_
timestamp 1698431365
transform 1 0 4144 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._191_
timestamp 1698431365
transform -1 0 10640 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._192_
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._226_
timestamp 1698431365
transform 1 0 17024 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_async_reg_bus._227_
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  u_rtc.u_async_reg_bus._231_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._232_
timestamp 1698431365
transform 1 0 2016 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  u_rtc.u_async_reg_bus._233_
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_rtc.u_async_reg_bus._234_
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  u_rtc.u_async_reg_bus._235_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._236_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._237_
timestamp 1698431365
transform 1 0 2688 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  u_rtc.u_async_reg_bus._238_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 58016
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  u_rtc.u_async_reg_bus._239_
timestamp 1698431365
transform 1 0 2688 0 -1 58016
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._240_
timestamp 1698431365
transform 1 0 2576 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._241_
timestamp 1698431365
transform 1 0 2688 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._242_
timestamp 1698431365
transform 1 0 2688 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._243_
timestamp 1698431365
transform 1 0 2688 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._244_
timestamp 1698431365
transform 1 0 2688 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._245_
timestamp 1698431365
transform 1 0 2688 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._246_
timestamp 1698431365
transform 1 0 2688 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._247_
timestamp 1698431365
transform 1 0 2688 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._248_
timestamp 1698431365
transform 1 0 2688 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._249_
timestamp 1698431365
transform 1 0 2688 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_rtc.u_async_reg_bus._250_
timestamp 1698431365
transform 1 0 2688 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._251_
timestamp 1698431365
transform 1 0 3584 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._252_
timestamp 1698431365
transform 1 0 3584 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._253_
timestamp 1698431365
transform 1 0 2688 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  u_rtc.u_async_reg_bus._254_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  u_rtc.u_async_reg_bus._255_
timestamp 1698431365
transform 1 0 2576 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  u_rtc.u_async_reg_bus._256_
timestamp 1698431365
transform 1 0 2688 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  u_rtc.u_async_reg_bus._257_
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  u_rtc.u_async_reg_bus._258_
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  u_rtc.u_async_reg_bus._259_
timestamp 1698431365
transform 1 0 2688 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._260_
timestamp 1698431365
transform 1 0 3360 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._261_
timestamp 1698431365
transform 1 0 1792 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._262_
timestamp 1698431365
transform 1 0 2688 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._263_
timestamp 1698431365
transform 1 0 2688 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._264_
timestamp 1698431365
transform 1 0 2352 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._265_
timestamp 1698431365
transform 1 0 2016 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._266_
timestamp 1698431365
transform 1 0 2688 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._267_
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._268_
timestamp 1698431365
transform 1 0 2688 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._269_
timestamp 1698431365
transform 1 0 2016 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_rtc.u_async_reg_bus._270_
timestamp 1698431365
transform 1 0 2688 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._400_
timestamp 1698431365
transform -1 0 7504 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._401_
timestamp 1698431365
transform -1 0 18368 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._402_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._403_
timestamp 1698431365
transform 1 0 7280 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._404_
timestamp 1698431365
transform 1 0 7616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_4  u_rtc.u_core._405_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30128 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._406_
timestamp 1698431365
transform -1 0 37296 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._407_
timestamp 1698431365
transform -1 0 32480 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._408_
timestamp 1698431365
transform -1 0 34384 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._409_
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  u_rtc.u_core._410_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31696 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_rtc.u_core._411_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32032 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  u_rtc.u_core._412_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._413_
timestamp 1698431365
transform 1 0 29904 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  u_rtc.u_core._414_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._415_
timestamp 1698431365
transform 1 0 33936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  u_rtc.u_core._416_
timestamp 1698431365
transform -1 0 24192 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  u_rtc.u_core._417_
timestamp 1698431365
transform 1 0 24192 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._418_
timestamp 1698431365
transform -1 0 24864 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._419_
timestamp 1698431365
transform -1 0 23520 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._420_
timestamp 1698431365
transform -1 0 23408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._421_
timestamp 1698431365
transform -1 0 21952 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._422_
timestamp 1698431365
transform 1 0 19152 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._423_
timestamp 1698431365
transform 1 0 13888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._424_
timestamp 1698431365
transform 1 0 13440 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._425_
timestamp 1698431365
transform -1 0 8400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._426_
timestamp 1698431365
transform -1 0 9856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._427_
timestamp 1698431365
transform 1 0 24304 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._428_
timestamp 1698431365
transform 1 0 25200 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._429_
timestamp 1698431365
transform 1 0 29904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._430_
timestamp 1698431365
transform -1 0 32480 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._431_
timestamp 1698431365
transform 1 0 28336 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_4  u_rtc.u_core._432_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31024 0 -1 64288
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._433_
timestamp 1698431365
transform 1 0 13440 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_rtc.u_core._434_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._435_
timestamp 1698431365
transform -1 0 8960 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._436_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8848 0 -1 79968
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_rtc.u_core._437_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11872 0 1 76832
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._438_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  u_rtc.u_core._439_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._440_
timestamp 1698431365
transform -1 0 10864 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  u_rtc.u_core._441_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 1 62720
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._442_
timestamp 1698431365
transform -1 0 9408 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._443_
timestamp 1698431365
transform 1 0 7392 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._444_
timestamp 1698431365
transform 1 0 7840 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  u_rtc.u_core._445_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  u_rtc.u_core._446_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._447_
timestamp 1698431365
transform -1 0 9184 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._448_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10752 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._449_
timestamp 1698431365
transform -1 0 9184 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  u_rtc.u_core._450_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10192 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._451_
timestamp 1698431365
transform 1 0 8848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._452_
timestamp 1698431365
transform 1 0 8400 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_rtc.u_core._453_
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._454_
timestamp 1698431365
transform 1 0 8624 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._455_
timestamp 1698431365
transform 1 0 9520 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  u_rtc.u_core._456_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9856 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._457_
timestamp 1698431365
transform -1 0 10752 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_core._458_
timestamp 1698431365
transform -1 0 29344 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._459_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  u_rtc.u_core._460_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35952 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_rtc.u_core._461_
timestamp 1698431365
transform -1 0 32368 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  u_rtc.u_core._462_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_rtc.u_core._463_
timestamp 1698431365
transform 1 0 32368 0 1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_core._464_
timestamp 1698431365
transform 1 0 34160 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  u_rtc.u_core._465_
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_core._466_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30912 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_rtc.u_core._467_
timestamp 1698431365
transform -1 0 37520 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._468_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  u_rtc.u_core._469_
timestamp 1698431365
transform 1 0 33824 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  u_rtc.u_core._470_
timestamp 1698431365
transform -1 0 31808 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._471_
timestamp 1698431365
transform 1 0 32704 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  u_rtc.u_core._472_
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._473_
timestamp 1698431365
transform -1 0 36288 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._474_
timestamp 1698431365
transform -1 0 36848 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_core._475_
timestamp 1698431365
transform -1 0 37968 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  u_rtc.u_core._476_
timestamp 1698431365
transform -1 0 36960 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._477_
timestamp 1698431365
transform -1 0 38416 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._478_
timestamp 1698431365
transform -1 0 38192 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  u_rtc.u_core._479_
timestamp 1698431365
transform 1 0 33936 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._480_
timestamp 1698431365
transform 1 0 32256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  u_rtc.u_core._481_
timestamp 1698431365
transform 1 0 33488 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._482_
timestamp 1698431365
transform 1 0 32032 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._483_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33824 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._484_
timestamp 1698431365
transform -1 0 33040 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  u_rtc.u_core._485_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34720 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._486_
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  u_rtc.u_core._487_
timestamp 1698431365
transform -1 0 37968 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._488_
timestamp 1698431365
transform 1 0 37520 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._489_
timestamp 1698431365
transform -1 0 34496 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._490_
timestamp 1698431365
transform -1 0 32704 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  u_rtc.u_core._491_
timestamp 1698431365
transform -1 0 34608 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._492_
timestamp 1698431365
transform 1 0 31024 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_rtc.u_core._493_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35504 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_rtc.u_core._494_
timestamp 1698431365
transform 1 0 33376 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._495_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_rtc.u_core._496_
timestamp 1698431365
transform 1 0 32480 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._497_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36736 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._498_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_core._499_
timestamp 1698431365
transform 1 0 35504 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  u_rtc.u_core._500_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35504 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._501_
timestamp 1698431365
transform -1 0 38080 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._502_
timestamp 1698431365
transform 1 0 36848 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._503_
timestamp 1698431365
transform -1 0 35504 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._504_
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  u_rtc.u_core._505_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38192 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._506_
timestamp 1698431365
transform -1 0 36512 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  u_rtc.u_core._507_
timestamp 1698431365
transform -1 0 36848 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._508_
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._509_
timestamp 1698431365
transform -1 0 38304 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._510_
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  u_rtc.u_core._511_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36624 0 1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  u_rtc.u_core._512_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._513_
timestamp 1698431365
transform -1 0 12432 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._514_
timestamp 1698431365
transform -1 0 14560 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  u_rtc.u_core._515_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15456 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._516_
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_rtc.u_core._517_
timestamp 1698431365
transform -1 0 22960 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  u_rtc.u_core._518_
timestamp 1698431365
transform -1 0 16912 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  u_rtc.u_core._519_
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  u_rtc.u_core._520_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._521_
timestamp 1698431365
transform -1 0 35056 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._522_
timestamp 1698431365
transform 1 0 34384 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_core._523_
timestamp 1698431365
transform -1 0 36624 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._524_
timestamp 1698431365
transform -1 0 37856 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._525_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  u_rtc.u_core._526_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34944 0 -1 42336
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  u_rtc.u_core._527_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34608 0 1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_rtc.u_core._528_
timestamp 1698431365
transform -1 0 34944 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._529_
timestamp 1698431365
transform 1 0 31584 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  u_rtc.u_core._530_
timestamp 1698431365
transform -1 0 31920 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._531_
timestamp 1698431365
transform -1 0 31248 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  u_rtc.u_core._532_
timestamp 1698431365
transform -1 0 36624 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._533_
timestamp 1698431365
transform 1 0 32144 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  u_rtc.u_core._534_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34384 0 -1 39200
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._535_
timestamp 1698431365
transform 1 0 37856 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  u_rtc.u_core._536_
timestamp 1698431365
transform -1 0 38416 0 -1 40768
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._537_
timestamp 1698431365
transform 1 0 30464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  u_rtc.u_core._538_
timestamp 1698431365
transform 1 0 31248 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  u_rtc.u_core._539_
timestamp 1698431365
transform -1 0 34384 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_rtc.u_core._540_
timestamp 1698431365
transform 1 0 31920 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  u_rtc.u_core._541_
timestamp 1698431365
transform -1 0 30688 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._542_
timestamp 1698431365
transform -1 0 29792 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._543_
timestamp 1698431365
transform 1 0 22960 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  u_rtc.u_core._544_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_rtc.u_core._545_
timestamp 1698431365
transform 1 0 28000 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._546_
timestamp 1698431365
transform -1 0 27552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._547_
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  u_rtc.u_core._548_
timestamp 1698431365
transform -1 0 24640 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_rtc.u_core._549_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_rtc.u_core._550_
timestamp 1698431365
transform 1 0 10976 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_core._551_
timestamp 1698431365
transform -1 0 11424 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  u_rtc.u_core._552_
timestamp 1698431365
transform -1 0 13104 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._554_
timestamp 1698431365
transform 1 0 30912 0 1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  u_rtc.u_core._555_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30912 0 1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._556_
timestamp 1698431365
transform -1 0 32032 0 1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._557_
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._558_
timestamp 1698431365
transform 1 0 34832 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_core._559_
timestamp 1698431365
transform -1 0 37968 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._560_
timestamp 1698431365
transform -1 0 37744 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._561_
timestamp 1698431365
transform -1 0 37744 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._562_
timestamp 1698431365
transform -1 0 37744 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._563_
timestamp 1698431365
transform -1 0 37744 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_core._564_
timestamp 1698431365
transform -1 0 36512 0 1 68992
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._565_
timestamp 1698431365
transform -1 0 32816 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._566_
timestamp 1698431365
transform -1 0 33488 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  u_rtc.u_core._567_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32032 0 -1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._568_
timestamp 1698431365
transform 1 0 30016 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._569_
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._570_
timestamp 1698431365
transform -1 0 32032 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._571_
timestamp 1698431365
transform -1 0 30800 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._572_
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._573_
timestamp 1698431365
transform -1 0 32144 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._574_
timestamp 1698431365
transform -1 0 30576 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._575_
timestamp 1698431365
transform -1 0 28224 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._576_
timestamp 1698431365
transform -1 0 29904 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._577_
timestamp 1698431365
transform 1 0 30800 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._578_
timestamp 1698431365
transform -1 0 30800 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._579_
timestamp 1698431365
transform -1 0 32144 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_core._580_
timestamp 1698431365
transform -1 0 31808 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._581_
timestamp 1698431365
transform -1 0 30128 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_core._582_
timestamp 1698431365
transform -1 0 31584 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._583_
timestamp 1698431365
transform -1 0 31360 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._584_
timestamp 1698431365
transform -1 0 31248 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._585_
timestamp 1698431365
transform -1 0 28784 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._586_
timestamp 1698431365
transform -1 0 30688 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._587_
timestamp 1698431365
transform 1 0 30352 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._588_
timestamp 1698431365
transform -1 0 33488 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._589_
timestamp 1698431365
transform -1 0 30240 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._590_
timestamp 1698431365
transform 1 0 31696 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._591_
timestamp 1698431365
transform 1 0 29792 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  u_rtc.u_core._592_
timestamp 1698431365
transform -1 0 32480 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._593_
timestamp 1698431365
transform 1 0 33936 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._594_
timestamp 1698431365
transform 1 0 34496 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._595_
timestamp 1698431365
transform -1 0 37744 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._596_
timestamp 1698431365
transform 1 0 36848 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._597_
timestamp 1698431365
transform -1 0 35952 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._598_
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._599_
timestamp 1698431365
transform -1 0 36624 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._600_
timestamp 1698431365
transform -1 0 36624 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._601_
timestamp 1698431365
transform -1 0 36624 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._602_
timestamp 1698431365
transform -1 0 36176 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._603_
timestamp 1698431365
transform -1 0 35280 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._604_
timestamp 1698431365
transform 1 0 35952 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._605_
timestamp 1698431365
transform -1 0 36288 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._606_
timestamp 1698431365
transform 1 0 36848 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._607_
timestamp 1698431365
transform -1 0 36064 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._608_
timestamp 1698431365
transform 1 0 35728 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._609_
timestamp 1698431365
transform 1 0 35392 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._610_
timestamp 1698431365
transform -1 0 35280 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._611_
timestamp 1698431365
transform 1 0 37520 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._612_
timestamp 1698431365
transform -1 0 35392 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._613_
timestamp 1698431365
transform -1 0 33600 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._614_
timestamp 1698431365
transform -1 0 32256 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  u_rtc.u_core._615_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32592 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._616_
timestamp 1698431365
transform -1 0 31472 0 -1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._617_
timestamp 1698431365
transform 1 0 29232 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._618_
timestamp 1698431365
transform -1 0 31696 0 1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._619_
timestamp 1698431365
transform -1 0 30352 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._620_
timestamp 1698431365
transform 1 0 10080 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._621_
timestamp 1698431365
transform 1 0 10752 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._622_
timestamp 1698431365
transform -1 0 12544 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._623_
timestamp 1698431365
transform -1 0 11648 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._624_
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  u_rtc.u_core._625_
timestamp 1698431365
transform -1 0 9408 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._626_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._627_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._628_
timestamp 1698431365
transform 1 0 6608 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._629_
timestamp 1698431365
transform 1 0 8064 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._630_
timestamp 1698431365
transform 1 0 5600 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  u_rtc.u_core._631_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6720 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._632_
timestamp 1698431365
transform 1 0 6720 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._633_
timestamp 1698431365
transform -1 0 7168 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_core._634_
timestamp 1698431365
transform 1 0 6720 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  u_rtc.u_core._635_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._636_
timestamp 1698431365
transform 1 0 9632 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._637_
timestamp 1698431365
transform -1 0 9296 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._638_
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._639_
timestamp 1698431365
transform 1 0 8064 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._640_
timestamp 1698431365
transform 1 0 5936 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  u_rtc.u_core._641_
timestamp 1698431365
transform -1 0 8064 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._642_
timestamp 1698431365
transform 1 0 15008 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._643_
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._644_
timestamp 1698431365
transform -1 0 16016 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._645_
timestamp 1698431365
transform -1 0 15344 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._646_
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._647_
timestamp 1698431365
transform -1 0 12880 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._648_
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._649_
timestamp 1698431365
transform -1 0 11200 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._650_
timestamp 1698431365
transform 1 0 12544 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._651_
timestamp 1698431365
transform 1 0 14112 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._652_
timestamp 1698431365
transform 1 0 11424 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._653_
timestamp 1698431365
transform -1 0 12880 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._654_
timestamp 1698431365
transform -1 0 12320 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._655_
timestamp 1698431365
transform 1 0 11088 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._656_
timestamp 1698431365
transform -1 0 12096 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._657_
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._658_
timestamp 1698431365
transform 1 0 8960 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._659_
timestamp 1698431365
transform 1 0 9744 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._660_
timestamp 1698431365
transform -1 0 10864 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._661_
timestamp 1698431365
transform 1 0 26544 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._662_
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_rtc.u_core._663_
timestamp 1698431365
transform -1 0 26656 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._664_
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._665_
timestamp 1698431365
transform 1 0 25648 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._666_
timestamp 1698431365
transform -1 0 24528 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._667_
timestamp 1698431365
transform -1 0 25984 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._668_
timestamp 1698431365
transform -1 0 24976 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._669_
timestamp 1698431365
transform 1 0 18704 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  u_rtc.u_core._670_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 20384
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._671_
timestamp 1698431365
transform 1 0 22064 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._672_
timestamp 1698431365
transform -1 0 22512 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._673_
timestamp 1698431365
transform -1 0 21504 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  u_rtc.u_core._674_
timestamp 1698431365
transform 1 0 19264 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._675_
timestamp 1698431365
transform 1 0 18480 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._676_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._677_
timestamp 1698431365
transform 1 0 20048 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  u_rtc.u_core._678_
timestamp 1698431365
transform 1 0 18704 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._679_
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._680_
timestamp 1698431365
transform 1 0 25872 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._681_
timestamp 1698431365
transform -1 0 29904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._682_
timestamp 1698431365
transform -1 0 29680 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._683_
timestamp 1698431365
transform 1 0 26320 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._684_
timestamp 1698431365
transform -1 0 25312 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_core._685_
timestamp 1698431365
transform -1 0 23520 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._686_
timestamp 1698431365
transform 1 0 22624 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._687_
timestamp 1698431365
transform -1 0 28224 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._688_
timestamp 1698431365
transform -1 0 24192 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._689_
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._690_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  u_rtc.u_core._691_
timestamp 1698431365
transform -1 0 29904 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._692_
timestamp 1698431365
transform 1 0 28672 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._693_
timestamp 1698431365
transform -1 0 28560 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._694_
timestamp 1698431365
transform 1 0 30016 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._695_
timestamp 1698431365
transform 1 0 29792 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._696_
timestamp 1698431365
transform 1 0 26096 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._697_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._698_
timestamp 1698431365
transform -1 0 28336 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  u_rtc.u_core._699_
timestamp 1698431365
transform 1 0 31024 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._700_
timestamp 1698431365
transform -1 0 25088 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._701_
timestamp 1698431365
transform 1 0 25088 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_core._702_
timestamp 1698431365
transform 1 0 25648 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._703_
timestamp 1698431365
transform 1 0 26432 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  u_rtc.u_core._704_
timestamp 1698431365
transform 1 0 26320 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._705_
timestamp 1698431365
transform 1 0 30240 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  u_rtc.u_core._706_
timestamp 1698431365
transform 1 0 29344 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._707_
timestamp 1698431365
transform -1 0 31808 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._708_
timestamp 1698431365
transform 1 0 30464 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._709_
timestamp 1698431365
transform -1 0 35728 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._710_
timestamp 1698431365
transform -1 0 31920 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._711_
timestamp 1698431365
transform 1 0 31472 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._712_
timestamp 1698431365
transform 1 0 30688 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._713_
timestamp 1698431365
transform 1 0 31248 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._714_
timestamp 1698431365
transform 1 0 33376 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._715_
timestamp 1698431365
transform 1 0 31248 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._716_
timestamp 1698431365
transform -1 0 32368 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._717_
timestamp 1698431365
transform 1 0 31136 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._718_
timestamp 1698431365
transform -1 0 33376 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._719_
timestamp 1698431365
transform -1 0 31136 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._720_
timestamp 1698431365
transform 1 0 16128 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._721_
timestamp 1698431365
transform 1 0 16464 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._722_
timestamp 1698431365
transform 1 0 17472 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._723_
timestamp 1698431365
transform -1 0 18256 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._724_
timestamp 1698431365
transform -1 0 17472 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._725_
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._726_
timestamp 1698431365
transform -1 0 18928 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_core._727_
timestamp 1698431365
transform 1 0 16912 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._728_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._729_
timestamp 1698431365
transform 1 0 14112 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._730_
timestamp 1698431365
transform -1 0 18144 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._731_
timestamp 1698431365
transform -1 0 18144 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._732_
timestamp 1698431365
transform -1 0 16016 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._733_
timestamp 1698431365
transform 1 0 6384 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._734_
timestamp 1698431365
transform -1 0 10304 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_core._735_
timestamp 1698431365
transform -1 0 11312 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._736_
timestamp 1698431365
transform 1 0 7728 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._737_
timestamp 1698431365
transform 1 0 5936 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._738_
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._739_
timestamp 1698431365
transform -1 0 9184 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._740_
timestamp 1698431365
transform -1 0 7616 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._741_
timestamp 1698431365
transform 1 0 7280 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._742_
timestamp 1698431365
transform -1 0 9072 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._743_
timestamp 1698431365
transform -1 0 8064 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._744_
timestamp 1698431365
transform 1 0 7280 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._745_
timestamp 1698431365
transform 1 0 6272 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._746_
timestamp 1698431365
transform -1 0 9072 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._747_
timestamp 1698431365
transform -1 0 8960 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  u_rtc.u_core._748_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8624 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._749_
timestamp 1698431365
transform -1 0 7840 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._750_
timestamp 1698431365
transform -1 0 10640 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  u_rtc.u_core._751_
timestamp 1698431365
transform 1 0 9968 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._752_
timestamp 1698431365
transform 1 0 11200 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._753_
timestamp 1698431365
transform -1 0 12992 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._754_
timestamp 1698431365
transform -1 0 12208 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._755_
timestamp 1698431365
transform -1 0 8736 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._756_
timestamp 1698431365
transform 1 0 10416 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._757_
timestamp 1698431365
transform 1 0 10976 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._758_
timestamp 1698431365
transform -1 0 10192 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._759_
timestamp 1698431365
transform 1 0 11648 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._760_
timestamp 1698431365
transform 1 0 4592 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._761_
timestamp 1698431365
transform -1 0 7728 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._762_
timestamp 1698431365
transform 1 0 7056 0 -1 61152
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._763_
timestamp 1698431365
transform 1 0 4704 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_core._764_
timestamp 1698431365
transform -1 0 7840 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._765_
timestamp 1698431365
transform 1 0 6048 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._766_
timestamp 1698431365
transform -1 0 6272 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._767_
timestamp 1698431365
transform -1 0 7952 0 1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._768_
timestamp 1698431365
transform 1 0 6720 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_core._769_
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._770_
timestamp 1698431365
transform 1 0 6160 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._771_
timestamp 1698431365
transform -1 0 8512 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._772_
timestamp 1698431365
transform 1 0 6608 0 1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._773_
timestamp 1698431365
transform 1 0 17808 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  u_rtc.u_core._774_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18704 0 1 65856
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  u_rtc.u_core._775_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  u_rtc.u_core._776_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20496 0 -1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._777_
timestamp 1698431365
transform 1 0 20496 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._778_
timestamp 1698431365
transform 1 0 18928 0 1 64288
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  u_rtc.u_core._779_
timestamp 1698431365
transform 1 0 18704 0 -1 67424
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._780_
timestamp 1698431365
transform 1 0 18704 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._781_
timestamp 1698431365
transform 1 0 19600 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_core._782_
timestamp 1698431365
transform -1 0 20608 0 1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._783_
timestamp 1698431365
transform 1 0 18816 0 -1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  u_rtc.u_core._784_
timestamp 1698431365
transform 1 0 19488 0 -1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  u_rtc.u_core._785_
timestamp 1698431365
transform 1 0 19712 0 1 62720
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._786_
timestamp 1698431365
transform 1 0 19264 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_core._787_
timestamp 1698431365
transform -1 0 8512 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._788_
timestamp 1698431365
transform 1 0 5376 0 -1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._789_
timestamp 1698431365
transform 1 0 5824 0 1 79968
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_core._790_
timestamp 1698431365
transform -1 0 6496 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._791_
timestamp 1698431365
transform 1 0 6496 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._792_
timestamp 1698431365
transform -1 0 6832 0 1 78400
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._793_
timestamp 1698431365
transform -1 0 5264 0 1 78400
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._794_
timestamp 1698431365
transform -1 0 3584 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._795_
timestamp 1698431365
transform 1 0 7056 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._796_
timestamp 1698431365
transform -1 0 6496 0 1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_core._797_
timestamp 1698431365
transform -1 0 4592 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  u_rtc.u_core._798_
timestamp 1698431365
transform -1 0 23408 0 -1 81536
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._799_
timestamp 1698431365
transform -1 0 23184 0 1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_core._800_
timestamp 1698431365
transform 1 0 22176 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_core._801_
timestamp 1698431365
transform -1 0 19824 0 -1 81536
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._802_
timestamp 1698431365
transform 1 0 13664 0 1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._803_
timestamp 1698431365
transform 1 0 15904 0 1 81536
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  u_rtc.u_core._804_
timestamp 1698431365
transform -1 0 18704 0 -1 81536
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._805_
timestamp 1698431365
transform 1 0 15792 0 -1 81536
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_rtc.u_core._806_
timestamp 1698431365
transform 1 0 14224 0 1 79968
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_core._807_
timestamp 1698431365
transform 1 0 16128 0 -1 83104
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_rtc.u_core._808_
timestamp 1698431365
transform -1 0 15680 0 1 81536
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_rtc.u_core._809_
timestamp 1698431365
transform -1 0 15680 0 -1 81536
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._810_
timestamp 1698431365
transform -1 0 14784 0 -1 84672
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_core._811_
timestamp 1698431365
transform -1 0 14672 0 -1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_core._812_
timestamp 1698431365
transform 1 0 18592 0 1 83104
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_core._813_
timestamp 1698431365
transform -1 0 18592 0 -1 83104
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_core._814_
timestamp 1698431365
transform -1 0 18592 0 1 83104
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_4  u_rtc.u_core._815_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31808 0 1 29792
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._816_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 -1 37632
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._817_
timestamp 1698431365
transform 1 0 30128 0 1 26656
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_4  u_rtc.u_core._818_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30464 0 1 25088
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._819_
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._820_
timestamp 1698431365
transform 1 0 29344 0 1 61152
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._821_
timestamp 1698431365
transform 1 0 30240 0 1 59584
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._822_
timestamp 1698431365
transform 1 0 33040 0 -1 56448
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._823_
timestamp 1698431365
transform 1 0 34496 0 -1 54880
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._824_
timestamp 1698431365
transform 1 0 34608 0 -1 58016
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._825_
timestamp 1698431365
transform 1 0 34608 0 -1 61152
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._826_
timestamp 1698431365
transform 1 0 33824 0 -1 62720
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._827_
timestamp 1698431365
transform 1 0 33936 0 -1 65856
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._828_
timestamp 1698431365
transform 1 0 33936 0 -1 67424
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._829_
timestamp 1698431365
transform 1 0 33712 0 -1 70560
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._830_
timestamp 1698431365
transform 1 0 32816 0 1 70560
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._831_
timestamp 1698431365
transform 1 0 30016 0 1 68992
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._832_
timestamp 1698431365
transform 1 0 29008 0 1 65856
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._833_
timestamp 1698431365
transform 1 0 28672 0 -1 67424
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._834_
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._835_
timestamp 1698431365
transform -1 0 9184 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._836_
timestamp 1698431365
transform 1 0 7952 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._837_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._838_
timestamp 1698431365
transform -1 0 17024 0 -1 12544
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._839_
timestamp 1698431365
transform -1 0 17360 0 1 17248
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._840_
timestamp 1698431365
transform 1 0 10864 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._841_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._842_
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._843_
timestamp 1698431365
transform -1 0 27664 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._844_
timestamp 1698431365
transform 1 0 18480 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._845_
timestamp 1698431365
transform 1 0 17360 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._846_
timestamp 1698431365
transform -1 0 31360 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._847_
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._848_
timestamp 1698431365
transform -1 0 27552 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._849_
timestamp 1698431365
transform -1 0 33040 0 1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_4  u_rtc.u_core._850_
timestamp 1698431365
transform 1 0 29792 0 1 20384
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_4  u_rtc.u_core._851_
timestamp 1698431365
transform 1 0 25872 0 -1 40768
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._852_
timestamp 1698431365
transform 1 0 26768 0 -1 42336
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_4  u_rtc.u_core._853_
timestamp 1698431365
transform 1 0 30352 0 1 45472
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._854_
timestamp 1698431365
transform 1 0 33488 0 -1 48608
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._855_
timestamp 1698431365
transform 1 0 31136 0 1 51744
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._856_
timestamp 1698431365
transform 1 0 31584 0 1 50176
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_2  u_rtc.u_core._857_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._858_
timestamp 1698431365
transform -1 0 20496 0 1 29792
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._859_
timestamp 1698431365
transform -1 0 19040 0 1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._860_
timestamp 1698431365
transform -1 0 11312 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._861_
timestamp 1698431365
transform 1 0 6608 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._862_
timestamp 1698431365
transform 1 0 6608 0 1 48608
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._863_
timestamp 1698431365
transform 1 0 7056 0 1 45472
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._864_
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._865_
timestamp 1698431365
transform 1 0 11200 0 -1 39200
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._866_
timestamp 1698431365
transform 1 0 5152 0 -1 62720
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._867_
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._868_
timestamp 1698431365
transform 1 0 3472 0 -1 56448
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._869_
timestamp 1698431365
transform -1 0 9184 0 -1 67424
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._870_
timestamp 1698431365
transform -1 0 25200 0 1 67424
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._871_
timestamp 1698431365
transform -1 0 21504 0 -1 72128
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._872_
timestamp 1698431365
transform -1 0 20944 0 1 61152
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._873_
timestamp 1698431365
transform 1 0 5376 0 -1 81536
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._874_
timestamp 1698431365
transform 1 0 1568 0 -1 79968
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._875_
timestamp 1698431365
transform 1 0 2912 0 -1 75264
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._876_
timestamp 1698431365
transform -1 0 24864 0 -1 83104
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._877_
timestamp 1698431365
transform 1 0 15680 0 1 79968
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._878_
timestamp 1698431365
transform 1 0 13328 0 1 83104
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_core._879_
timestamp 1698431365
transform 1 0 16912 0 1 81536
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_core._880_
timestamp 1698431365
transform 1 0 25312 0 -1 65856
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0602_
timestamp 1698431365
transform -1 0 7392 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0603_
timestamp 1698431365
transform -1 0 5824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0604_
timestamp 1698431365
transform 1 0 2352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0605_
timestamp 1698431365
transform -1 0 18816 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0606_
timestamp 1698431365
transform -1 0 14000 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0607_
timestamp 1698431365
transform -1 0 13216 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0608_
timestamp 1698431365
transform -1 0 12208 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0609_
timestamp 1698431365
transform -1 0 9968 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_rtc.u_reg._0610_
timestamp 1698431365
transform 1 0 9408 0 -1 81536
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0611_
timestamp 1698431365
transform -1 0 11760 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0612_
timestamp 1698431365
transform 1 0 10752 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0613_
timestamp 1698431365
transform -1 0 20944 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0614_
timestamp 1698431365
transform 1 0 18928 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0615_
timestamp 1698431365
transform 1 0 19936 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0616_
timestamp 1698431365
transform 1 0 18256 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0617_
timestamp 1698431365
transform 1 0 18704 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_rtc.u_reg._0618_
timestamp 1698431365
transform -1 0 19824 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0619_
timestamp 1698431365
transform -1 0 19264 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0620_
timestamp 1698431365
transform 1 0 18144 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0621_
timestamp 1698431365
transform 1 0 17584 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0622_
timestamp 1698431365
transform -1 0 15792 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_rtc.u_reg._0623_
timestamp 1698431365
transform -1 0 16464 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0624_
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0625_
timestamp 1698431365
transform -1 0 14560 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0626_
timestamp 1698431365
transform -1 0 18592 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0627_
timestamp 1698431365
transform -1 0 19040 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0628_
timestamp 1698431365
transform -1 0 14560 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0629_
timestamp 1698431365
transform 1 0 13216 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0630_
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0631_
timestamp 1698431365
transform -1 0 17808 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0632_
timestamp 1698431365
transform -1 0 13104 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_rtc.u_reg._0633_
timestamp 1698431365
transform -1 0 13104 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0634_
timestamp 1698431365
transform -1 0 4704 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0637_
timestamp 1698431365
transform 1 0 5824 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0638_
timestamp 1698431365
transform 1 0 3584 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0639_
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_rtc.u_reg._0640_
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0641_
timestamp 1698431365
transform 1 0 19376 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0645_
timestamp 1698431365
transform -1 0 28112 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0646_
timestamp 1698431365
transform -1 0 26656 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0652_
timestamp 1698431365
transform -1 0 4816 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0667_
timestamp 1698431365
transform 1 0 2800 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_rtc.u_reg._0668_
timestamp 1698431365
transform -1 0 2688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0669_
timestamp 1698431365
transform 1 0 21728 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0670_
timestamp 1698431365
transform -1 0 23968 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0671_
timestamp 1698431365
transform 1 0 21616 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_reg._0672_
timestamp 1698431365
transform -1 0 23632 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0673_
timestamp 1698431365
transform -1 0 18256 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0674_
timestamp 1698431365
transform 1 0 16016 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0675_
timestamp 1698431365
transform 1 0 15456 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  u_rtc.u_reg._0676_
timestamp 1698431365
transform 1 0 15232 0 1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_reg._0677_
timestamp 1698431365
transform 1 0 15792 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  u_rtc.u_reg._0678_
timestamp 1698431365
transform -1 0 18480 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0679_
timestamp 1698431365
transform 1 0 14336 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  u_rtc.u_reg._0680_
timestamp 1698431365
transform 1 0 14448 0 -1 62720
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0681_
timestamp 1698431365
transform -1 0 17248 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0682_
timestamp 1698431365
transform 1 0 14000 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_reg._0683_
timestamp 1698431365
transform 1 0 13552 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_reg._0684_
timestamp 1698431365
transform 1 0 15680 0 -1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0685_
timestamp 1698431365
transform 1 0 14112 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  u_rtc.u_reg._0686_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14560 0 -1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0687_
timestamp 1698431365
transform -1 0 14672 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0688_
timestamp 1698431365
transform 1 0 12096 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0689_
timestamp 1698431365
transform 1 0 11760 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0690_
timestamp 1698431365
transform 1 0 10752 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  u_rtc.u_reg._0691_
timestamp 1698431365
transform 1 0 12880 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  u_rtc.u_reg._0692_
timestamp 1698431365
transform 1 0 14672 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0693_
timestamp 1698431365
transform 1 0 13328 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_reg._0694_
timestamp 1698431365
transform -1 0 17472 0 1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  u_rtc.u_reg._0695_
timestamp 1698431365
transform 1 0 10416 0 -1 75264
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  u_rtc.u_reg._0696_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13440 0 -1 79968
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  u_rtc.u_reg._0697_
timestamp 1698431365
transform 1 0 13440 0 1 76832
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0698_
timestamp 1698431365
transform 1 0 21504 0 -1 79968
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0699_
timestamp 1698431365
transform 1 0 19600 0 1 78400
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0700_
timestamp 1698431365
transform 1 0 22848 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  u_rtc.u_reg._0701_
timestamp 1698431365
transform -1 0 16016 0 -1 78400
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  u_rtc.u_reg._0702_
timestamp 1698431365
transform 1 0 14112 0 1 78400
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  u_rtc.u_reg._0703_
timestamp 1698431365
transform 1 0 14672 0 -1 76832
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  u_rtc.u_reg._0704_
timestamp 1698431365
transform 1 0 14448 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  u_rtc.u_reg._0705_
timestamp 1698431365
transform 1 0 14000 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  u_rtc.u_reg._0706_
timestamp 1698431365
transform -1 0 16576 0 1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  u_rtc.u_reg._0707_
timestamp 1698431365
transform -1 0 14784 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  u_rtc.u_reg._0708_
timestamp 1698431365
transform -1 0 14000 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0709_
timestamp 1698431365
transform 1 0 14112 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0710_
timestamp 1698431365
transform 1 0 13328 0 -1 59584
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_rtc.u_reg._0711_
timestamp 1698431365
transform -1 0 16464 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  u_rtc.u_reg._0712_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15232 0 1 61152
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  u_rtc.u_reg._0713_
timestamp 1698431365
transform 1 0 14448 0 -1 64288
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_reg._0714_
timestamp 1698431365
transform 1 0 13440 0 -1 65856
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0715_
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  u_rtc.u_reg._0716_
timestamp 1698431365
transform 1 0 14784 0 1 62720
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  u_rtc.u_reg._0717_
timestamp 1698431365
transform -1 0 16464 0 1 64288
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0718_
timestamp 1698431365
transform -1 0 24640 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0719_
timestamp 1698431365
transform 1 0 22400 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0720_
timestamp 1698431365
transform 1 0 22960 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  u_rtc.u_reg._0721_
timestamp 1698431365
transform 1 0 23072 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0722_
timestamp 1698431365
transform 1 0 18256 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0723_
timestamp 1698431365
transform -1 0 18368 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  u_rtc.u_reg._0724_
timestamp 1698431365
transform 1 0 16688 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_rtc.u_reg._0725_
timestamp 1698431365
transform -1 0 19264 0 1 67424
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  u_rtc.u_reg._0726_
timestamp 1698431365
transform 1 0 18144 0 1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0727_
timestamp 1698431365
transform 1 0 15792 0 -1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  u_rtc.u_reg._0728_
timestamp 1698431365
transform 1 0 18256 0 1 68992
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0729_
timestamp 1698431365
transform 1 0 17920 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0730_
timestamp 1698431365
transform 1 0 15344 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_reg._0731_
timestamp 1698431365
transform -1 0 16912 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  u_rtc.u_reg._0732_
timestamp 1698431365
transform -1 0 18704 0 -1 67424
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0733_
timestamp 1698431365
transform -1 0 19040 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  u_rtc.u_reg._0734_
timestamp 1698431365
transform 1 0 17808 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  u_rtc.u_reg._0735_
timestamp 1698431365
transform -1 0 19600 0 1 50176
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0736_
timestamp 1698431365
transform 1 0 15680 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0737_
timestamp 1698431365
transform 1 0 17024 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0738_
timestamp 1698431365
transform 1 0 14336 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0739_
timestamp 1698431365
transform 1 0 15680 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  u_rtc.u_reg._0740_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0741_
timestamp 1698431365
transform -1 0 15232 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  u_rtc.u_reg._0742_
timestamp 1698431365
transform 1 0 17360 0 -1 68992
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0743_
timestamp 1698431365
transform 1 0 10752 0 1 81536
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  u_rtc.u_reg._0744_
timestamp 1698431365
transform -1 0 10528 0 1 79968
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0745_
timestamp 1698431365
transform 1 0 9744 0 1 81536
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  u_rtc.u_reg._0746_
timestamp 1698431365
transform 1 0 10528 0 -1 83104
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  u_rtc.u_reg._0747_
timestamp 1698431365
transform -1 0 13104 0 1 83104
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  u_rtc.u_reg._0748_
timestamp 1698431365
transform -1 0 11424 0 -1 81536
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0749_
timestamp 1698431365
transform 1 0 11088 0 1 79968
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_reg._0750_
timestamp 1698431365
transform 1 0 11760 0 1 81536
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  u_rtc.u_reg._0751_
timestamp 1698431365
transform 1 0 11536 0 -1 81536
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  u_rtc.u_reg._0752_
timestamp 1698431365
transform 1 0 17472 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  u_rtc.u_reg._0753_
timestamp 1698431365
transform 1 0 18368 0 -1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  u_rtc.u_reg._0754_
timestamp 1698431365
transform -1 0 19936 0 1 58016
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0755_
timestamp 1698431365
transform 1 0 15680 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  u_rtc.u_reg._0756_
timestamp 1698431365
transform 1 0 19712 0 -1 58016
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_rtc.u_reg._0757_
timestamp 1698431365
transform 1 0 16912 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  u_rtc.u_reg._0758_
timestamp 1698431365
transform 1 0 18368 0 1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_reg._0759_
timestamp 1698431365
transform -1 0 19152 0 -1 59584
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0760_
timestamp 1698431365
transform -1 0 17024 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  u_rtc.u_reg._0761_
timestamp 1698431365
transform 1 0 16240 0 1 68992
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_reg._0762_
timestamp 1698431365
transform -1 0 16240 0 1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_rtc.u_reg._0763_
timestamp 1698431365
transform 1 0 14112 0 1 67424
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  u_rtc.u_reg._0764_
timestamp 1698431365
transform 1 0 15120 0 -1 67424
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  u_rtc.u_reg._0765_
timestamp 1698431365
transform -1 0 19152 0 -1 70560
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  u_rtc.u_reg._0766_
timestamp 1698431365
transform 1 0 25200 0 1 67424
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  u_rtc.u_reg._0767_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 1 6272
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_reg._0768_
timestamp 1698431365
transform 1 0 4368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  u_rtc.u_reg._0769_
timestamp 1698431365
transform 1 0 5712 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0770_
timestamp 1698431365
transform 1 0 4704 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0771_
timestamp 1698431365
transform 1 0 7504 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  u_rtc.u_reg._0772_
timestamp 1698431365
transform 1 0 5712 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_reg._0773_
timestamp 1698431365
transform 1 0 6720 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_rtc.u_reg._0774_
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0775_
timestamp 1698431365
transform 1 0 14336 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0776_
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0777_
timestamp 1698431365
transform 1 0 15120 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0778_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0779_
timestamp 1698431365
transform 1 0 11760 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0780_
timestamp 1698431365
transform 1 0 11088 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_reg._0791_
timestamp 1698431365
transform -1 0 6384 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_reg._0792_
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  u_rtc.u_reg._0793_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7056 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0794_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._0795_
timestamp 1698431365
transform 1 0 14784 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0796_
timestamp 1698431365
transform 1 0 27104 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0797_
timestamp 1698431365
transform 1 0 26992 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0798_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0799_
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0800_
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0801_
timestamp 1698431365
transform 1 0 26320 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0802_
timestamp 1698431365
transform 1 0 27104 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0803_
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0804_
timestamp 1698431365
transform 1 0 23296 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0805_
timestamp 1698431365
transform 1 0 22736 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0810_
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._0811_
timestamp 1698431365
transform 1 0 15008 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0812_
timestamp 1698431365
transform 1 0 22400 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0813_
timestamp 1698431365
transform 1 0 22512 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0814_
timestamp 1698431365
transform 1 0 19040 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0815_
timestamp 1698431365
transform 1 0 19040 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0816_
timestamp 1698431365
transform 1 0 18928 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0817_
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0818_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0819_
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0820_
timestamp 1698431365
transform 1 0 22400 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0821_
timestamp 1698431365
transform 1 0 22624 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0822_
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0823_
timestamp 1698431365
transform 1 0 20384 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0824_
timestamp 1698431365
transform 1 0 17360 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0825_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0826_
timestamp 1698431365
transform 1 0 15344 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0827_
timestamp 1698431365
transform 1 0 15344 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  u_rtc.u_reg._0828_
timestamp 1698431365
transform -1 0 5824 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._0829_
timestamp 1698431365
transform -1 0 7616 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0830_
timestamp 1698431365
transform 1 0 14336 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0831_
timestamp 1698431365
transform 1 0 13440 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0832_
timestamp 1698431365
transform 1 0 13216 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0833_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0834_
timestamp 1698431365
transform 1 0 9408 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0835_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0836_
timestamp 1698431365
transform 1 0 3584 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0837_
timestamp 1698431365
transform 1 0 5600 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0838_
timestamp 1698431365
transform 1 0 3472 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0839_
timestamp 1698431365
transform 1 0 2912 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0840_
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0841_
timestamp 1698431365
transform 1 0 2800 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0842_
timestamp 1698431365
transform 1 0 3584 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0843_
timestamp 1698431365
transform 1 0 3136 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  u_rtc.u_reg._0844_
timestamp 1698431365
transform -1 0 4704 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_rtc.u_reg._0845_
timestamp 1698431365
transform 1 0 6048 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  u_rtc.u_reg._0846_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._0847_
timestamp 1698431365
transform 1 0 11312 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0848_
timestamp 1698431365
transform -1 0 12320 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0849_
timestamp 1698431365
transform 1 0 10752 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0850_
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0851_
timestamp 1698431365
transform -1 0 12992 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0852_
timestamp 1698431365
transform 1 0 11424 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0853_
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0854_
timestamp 1698431365
transform -1 0 15344 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0855_
timestamp 1698431365
transform 1 0 13776 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0856_
timestamp 1698431365
transform -1 0 13104 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0857_
timestamp 1698431365
transform 1 0 11424 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0858_
timestamp 1698431365
transform -1 0 21728 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0859_
timestamp 1698431365
transform 1 0 20048 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0860_
timestamp 1698431365
transform 1 0 22064 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0861_
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  u_rtc.u_reg._0862_
timestamp 1698431365
transform 1 0 12656 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0863_
timestamp 1698431365
transform 1 0 19040 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0864_
timestamp 1698431365
transform 1 0 16352 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0865_
timestamp 1698431365
transform -1 0 18144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0884_
timestamp 1698431365
transform -1 0 5152 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_rtc.u_reg._0885_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  u_rtc.u_reg._0886_
timestamp 1698431365
transform 1 0 7952 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._0887_
timestamp 1698431365
transform -1 0 15120 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0888_
timestamp 1698431365
transform -1 0 23184 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0889_
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0890_
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0891_
timestamp 1698431365
transform -1 0 22512 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0892_
timestamp 1698431365
transform 1 0 21280 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0893_
timestamp 1698431365
transform -1 0 19824 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0894_
timestamp 1698431365
transform 1 0 18592 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0895_
timestamp 1698431365
transform -1 0 18816 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0896_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0897_
timestamp 1698431365
transform 1 0 13440 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0898_
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0899_
timestamp 1698431365
transform -1 0 23968 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0900_
timestamp 1698431365
transform 1 0 22512 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0901_
timestamp 1698431365
transform -1 0 24192 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0902_
timestamp 1698431365
transform 1 0 21840 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  u_rtc.u_reg._0903_
timestamp 1698431365
transform 1 0 13440 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0904_
timestamp 1698431365
transform -1 0 20944 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0905_
timestamp 1698431365
transform 1 0 16352 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0906_
timestamp 1698431365
transform -1 0 18144 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  u_rtc.u_reg._0925_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  u_rtc.u_reg._0927_
timestamp 1698431365
transform 1 0 8176 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0928_
timestamp 1698431365
transform -1 0 26432 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0929_
timestamp 1698431365
transform 1 0 23968 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0930_
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0931_
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0932_
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0933_
timestamp 1698431365
transform -1 0 28448 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0934_
timestamp 1698431365
transform -1 0 26656 0 1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0937_
timestamp 1698431365
transform -1 0 27328 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0938_
timestamp 1698431365
transform 1 0 24528 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0939_
timestamp 1698431365
transform -1 0 26768 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0940_
timestamp 1698431365
transform 1 0 23968 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0945_
timestamp 1698431365
transform 1 0 5600 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._0946_
timestamp 1698431365
transform -1 0 7280 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0947_
timestamp 1698431365
transform 1 0 3584 0 1 67424
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0948_
timestamp 1698431365
transform 1 0 3136 0 -1 67424
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0949_
timestamp 1698431365
transform -1 0 20944 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0950_
timestamp 1698431365
transform 1 0 19824 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0951_
timestamp 1698431365
transform 1 0 21168 0 1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0952_
timestamp 1698431365
transform -1 0 20944 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0953_
timestamp 1698431365
transform 1 0 19600 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0954_
timestamp 1698431365
transform 1 0 21504 0 -1 72128
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0955_
timestamp 1698431365
transform 1 0 21392 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0956_
timestamp 1698431365
transform 1 0 20496 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0957_
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0958_
timestamp 1698431365
transform 1 0 5376 0 -1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0959_
timestamp 1698431365
transform 1 0 3472 0 1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0960_
timestamp 1698431365
transform 1 0 3584 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0961_
timestamp 1698431365
transform 1 0 3024 0 1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0962_
timestamp 1698431365
transform 1 0 3584 0 1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0963_
timestamp 1698431365
transform 1 0 3024 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0965_
timestamp 1698431365
transform 1 0 4704 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._0966_
timestamp 1698431365
transform -1 0 7280 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0967_
timestamp 1698431365
transform 1 0 5376 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0968_
timestamp 1698431365
transform 1 0 3584 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0969_
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0970_
timestamp 1698431365
transform 1 0 3584 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0971_
timestamp 1698431365
transform 1 0 5488 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0972_
timestamp 1698431365
transform 1 0 3472 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0973_
timestamp 1698431365
transform 1 0 6720 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0974_
timestamp 1698431365
transform 1 0 5600 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0975_
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0976_
timestamp 1698431365
transform 1 0 1904 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0977_
timestamp 1698431365
transform 1 0 5376 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0978_
timestamp 1698431365
transform 1 0 3584 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  u_rtc.u_reg._0985_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0986_
timestamp 1698431365
transform -1 0 11536 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0987_
timestamp 1698431365
transform 1 0 9744 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0988_
timestamp 1698431365
transform 1 0 3584 0 1 62720
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0989_
timestamp 1698431365
transform 1 0 10416 0 1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0990_
timestamp 1698431365
transform 1 0 10976 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0991_
timestamp 1698431365
transform -1 0 12544 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._0992_
timestamp 1698431365
transform 1 0 11536 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._0993_
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._0994_
timestamp 1698431365
transform 1 0 11424 0 1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0995_
timestamp 1698431365
transform -1 0 9968 0 -1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0996_
timestamp 1698431365
transform 1 0 7616 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._0997_
timestamp 1698431365
transform -1 0 6160 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._0998_
timestamp 1698431365
transform 1 0 4256 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._0999_
timestamp 1698431365
transform -1 0 11424 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1000_
timestamp 1698431365
transform 1 0 10080 0 -1 87808
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1001_
timestamp 1698431365
transform 1 0 7392 0 1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1002_
timestamp 1698431365
transform 1 0 5712 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1003_
timestamp 1698431365
transform 1 0 9856 0 -1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1004_
timestamp 1698431365
transform 1 0 9744 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1005_
timestamp 1698431365
transform 1 0 8288 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1006_
timestamp 1698431365
transform 1 0 8064 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1007_
timestamp 1698431365
transform 1 0 8512 0 -1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1008_
timestamp 1698431365
transform -1 0 10304 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._1009_
timestamp 1698431365
transform -1 0 9184 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._1010_
timestamp 1698431365
transform 1 0 7504 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._1013_
timestamp 1698431365
transform -1 0 11984 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1014_
timestamp 1698431365
transform -1 0 22848 0 1 78400
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1015_
timestamp 1698431365
transform -1 0 17024 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1016_
timestamp 1698431365
transform 1 0 15568 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1017_
timestamp 1698431365
transform 1 0 17584 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1018_
timestamp 1698431365
transform 1 0 17248 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1019_
timestamp 1698431365
transform -1 0 22624 0 -1 76832
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1020_
timestamp 1698431365
transform 1 0 11424 0 1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1021_
timestamp 1698431365
transform 1 0 12432 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1022_
timestamp 1698431365
transform 1 0 12208 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._1023_
timestamp 1698431365
transform 1 0 9744 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._1024_
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._1027_
timestamp 1698431365
transform 1 0 12096 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._1028_
timestamp 1698431365
transform -1 0 15456 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1029_
timestamp 1698431365
transform -1 0 20608 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1030_
timestamp 1698431365
transform -1 0 22064 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1031_
timestamp 1698431365
transform 1 0 27440 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1032_
timestamp 1698431365
transform 1 0 25648 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1033_
timestamp 1698431365
transform -1 0 28336 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1034_
timestamp 1698431365
transform 1 0 27328 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1035_
timestamp 1698431365
transform -1 0 27104 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1036_
timestamp 1698431365
transform 1 0 27104 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1037_
timestamp 1698431365
transform -1 0 27216 0 1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1038_
timestamp 1698431365
transform 1 0 27216 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1039_
timestamp 1698431365
transform -1 0 23296 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1040_
timestamp 1698431365
transform 1 0 22400 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._1041_
timestamp 1698431365
transform 1 0 14000 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._1042_
timestamp 1698431365
transform -1 0 20160 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1043_
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._1046_
timestamp 1698431365
transform 1 0 4704 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_rtc.u_reg._1047_
timestamp 1698431365
transform -1 0 7168 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1048_
timestamp 1698431365
transform -1 0 22400 0 -1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1049_
timestamp 1698431365
transform 1 0 21168 0 1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1050_
timestamp 1698431365
transform 1 0 13216 0 -1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1051_
timestamp 1698431365
transform -1 0 14672 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1052_
timestamp 1698431365
transform -1 0 17024 0 -1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1053_
timestamp 1698431365
transform 1 0 15008 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._1054_
timestamp 1698431365
transform -1 0 13888 0 -1 84672
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._1055_
timestamp 1698431365
transform 1 0 12432 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1056_
timestamp 1698431365
transform 1 0 13328 0 1 87808
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1057_
timestamp 1698431365
transform 1 0 18480 0 -1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1058_
timestamp 1698431365
transform 1 0 18144 0 1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_rtc.u_reg._1059_
timestamp 1698431365
transform -1 0 6496 0 -1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_rtc.u_reg._1060_
timestamp 1698431365
transform 1 0 4256 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1061_
timestamp 1698431365
transform 1 0 3136 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1062_
timestamp 1698431365
transform 1 0 5376 0 -1 78400
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1063_
timestamp 1698431365
transform 1 0 3024 0 1 76832
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1064_
timestamp 1698431365
transform 1 0 3584 0 1 72128
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_reg._1065_
timestamp 1698431365
transform 1 0 3248 0 1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1067_
timestamp 1698431365
transform 1 0 3472 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1068_
timestamp 1698431365
transform -1 0 6048 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_rtc.u_reg._1069_
timestamp 1698431365
transform -1 0 4368 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1070_
timestamp 1698431365
transform -1 0 3696 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_rtc.u_reg._1071_
timestamp 1698431365
transform -1 0 4704 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_rtc.u_reg._1072_
timestamp 1698431365
transform 1 0 4368 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1205_
timestamp 1698431365
transform 1 0 12208 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1206_
timestamp 1698431365
transform 1 0 11312 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1207_
timestamp 1698431365
transform 1 0 9296 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1213_
timestamp 1698431365
transform 1 0 25984 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1214_
timestamp 1698431365
transform 1 0 22848 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1215_
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1216_
timestamp 1698431365
transform 1 0 26880 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1217_
timestamp 1698431365
transform 1 0 21056 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1221_
timestamp 1698431365
transform 1 0 21952 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1222_
timestamp 1698431365
transform 1 0 18032 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1223_
timestamp 1698431365
transform 1 0 18032 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1224_
timestamp 1698431365
transform 1 0 21056 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1225_
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1226_
timestamp 1698431365
transform 1 0 19488 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1227_
timestamp 1698431365
transform 1 0 16240 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1228_
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1229_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1230_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1231_
timestamp 1698431365
transform 1 0 7616 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1232_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1233_
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1234_
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1235_
timestamp 1698431365
transform 1 0 1680 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1236_
timestamp 1698431365
transform 1 0 1680 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1237_
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1238_
timestamp 1698431365
transform 1 0 7616 0 1 56448
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1239_
timestamp 1698431365
transform 1 0 8960 0 1 58016
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1240_
timestamp 1698431365
transform 1 0 7840 0 1 53312
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1241_
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1242_
timestamp 1698431365
transform 1 0 10528 0 -1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1243_
timestamp 1698431365
transform 1 0 19712 0 -1 51744
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1244_
timestamp 1698431365
transform 1 0 19824 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1245_
timestamp 1698431365
transform 1 0 18368 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1246_
timestamp 1698431365
transform -1 0 18928 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1261_
timestamp 1698431365
transform -1 0 25872 0 1 56448
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1262_
timestamp 1698431365
transform -1 0 27440 0 1 58016
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1263_
timestamp 1698431365
transform 1 0 21056 0 -1 58016
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1264_
timestamp 1698431365
transform 1 0 18032 0 -1 54880
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1265_
timestamp 1698431365
transform 1 0 16128 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1266_
timestamp 1698431365
transform 1 0 11424 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1267_
timestamp 1698431365
transform 1 0 21728 0 1 51744
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1268_
timestamp 1698431365
transform 1 0 20720 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1269_
timestamp 1698431365
transform 1 0 19152 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1270_
timestamp 1698431365
transform 1 0 15008 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1285_
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1286_
timestamp 1698431365
transform 1 0 23856 0 1 68992
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  u_rtc.u_reg._1287_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14784 0 -1 36064
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1288_
timestamp 1698431365
transform 1 0 25984 0 -1 59584
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1289_
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1291_
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1292_
timestamp 1698431365
transform 1 0 24192 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1294_
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1295_
timestamp 1698431365
transform 1 0 20720 0 -1 67424
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1296_
timestamp 1698431365
transform -1 0 23632 0 -1 73696
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1297_
timestamp 1698431365
transform 1 0 20944 0 -1 62720
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1298_
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1299_
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1300_
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1302_
timestamp 1698431365
transform 1 0 1792 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1303_
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1304_
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1305_
timestamp 1698431365
transform 1 0 4368 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1306_
timestamp 1698431365
transform 1 0 1792 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1307_
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1311_
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1312_
timestamp 1698431365
transform 1 0 1680 0 -1 64288
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1313_
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1314_
timestamp 1698431365
transform 1 0 10640 0 -1 62720
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1315_
timestamp 1698431365
transform 1 0 12208 0 -1 68992
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_reg._1316_
timestamp 1698431365
transform 1 0 10528 0 -1 70560
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_reg._1317_
timestamp 1698431365
transform 1 0 6720 0 1 68992
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1318_
timestamp 1698431365
transform 1 0 3136 0 -1 68992
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1319_
timestamp 1698431365
transform 1 0 9072 0 1 87808
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1320_
timestamp 1698431365
transform 1 0 5376 0 -1 87808
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1321_
timestamp 1698431365
transform 1 0 3584 0 -1 84672
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1322_
timestamp 1698431365
transform 1 0 9408 0 -1 89376
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1323_
timestamp 1698431365
transform 1 0 6272 0 1 84672
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1324_
timestamp 1698431365
transform 1 0 7504 0 1 78400
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1325_
timestamp 1698431365
transform 1 0 5376 0 -1 73696
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1327_
timestamp 1698431365
transform -1 0 24080 0 -1 78400
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1328_
timestamp 1698431365
transform 1 0 15792 0 1 73696
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1329_
timestamp 1698431365
transform 1 0 16464 0 1 75264
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1330_
timestamp 1698431365
transform -1 0 24976 0 1 76832
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1331_
timestamp 1698431365
transform 1 0 10864 0 -1 76832
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1332_
timestamp 1698431365
transform 1 0 11424 0 -1 73696
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1333_
timestamp 1698431365
transform 1 0 7168 0 1 73696
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1335_
timestamp 1698431365
transform 1 0 24976 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1336_
timestamp 1698431365
transform 1 0 27104 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1337_
timestamp 1698431365
transform 1 0 26544 0 -1 53312
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1338_
timestamp 1698431365
transform 1 0 27104 0 -1 54880
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1339_
timestamp 1698431365
transform 1 0 21616 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1340_
timestamp 1698431365
transform 1 0 20720 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1343_
timestamp 1698431365
transform 1 0 19936 0 -1 86240
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1344_
timestamp 1698431365
transform 1 0 14336 0 1 86240
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1345_
timestamp 1698431365
transform 1 0 11872 0 -1 87808
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1346_
timestamp 1698431365
transform 1 0 17248 0 -1 87808
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1347_
timestamp 1698431365
transform 1 0 1568 0 -1 83104
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1348_
timestamp 1698431365
transform 1 0 1568 0 -1 78400
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1349_
timestamp 1698431365
transform 1 0 1568 0 -1 73696
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1351_
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_reg._1352_
timestamp 1698431365
transform -1 0 5376 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_rtc.u_reg._1353_
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  u_rtc.u_sync_rclk._1__60
timestamp 1698431365
transform -1 0 23296 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_sync_rclk._1_
timestamp 1698431365
transform 1 0 22176 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_sync_rclk._2_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_rtc.u_sync_rclk.u_buf.genblk1.u_mux_57
timestamp 1698431365
transform -1 0 29344 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_sync_rclk.u_buf.genblk1.u_mux
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_sync_sclk._1_
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  u_rtc.u_sync_sclk._1__61
timestamp 1698431365
transform 1 0 21952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_rtc.u_sync_sclk._2_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_rtc.u_sync_sclk.u_buf.genblk1.u_mux_58
timestamp 1698431365
transform -1 0 27888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_rtc.u_sync_sclk.u_buf.genblk1.u_mux
timestamp 1698431365
transform 1 0 25760 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  wire1
timestamp 1698431365
transform 1 0 13328 0 1 86240
box -86 -86 982 870
<< labels >>
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 mclk
port 0 nsew signal input
flabel metal3 s 0 95200 800 95312 0 FreeSans 448 0 0 0 reg_ack
port 1 nsew signal tristate
flabel metal3 s 0 17920 800 18032 0 FreeSans 448 0 0 0 reg_addr[0]
port 2 nsew signal input
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 reg_addr[10]
port 3 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 reg_addr[1]
port 4 nsew signal input
flabel metal3 s 0 15680 800 15792 0 FreeSans 448 0 0 0 reg_addr[2]
port 5 nsew signal input
flabel metal3 s 0 14560 800 14672 0 FreeSans 448 0 0 0 reg_addr[3]
port 6 nsew signal input
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 reg_addr[4]
port 7 nsew signal input
flabel metal3 s 0 12320 800 12432 0 FreeSans 448 0 0 0 reg_addr[5]
port 8 nsew signal input
flabel metal3 s 0 11200 800 11312 0 FreeSans 448 0 0 0 reg_addr[6]
port 9 nsew signal input
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 reg_addr[7]
port 10 nsew signal input
flabel metal3 s 0 8960 800 9072 0 FreeSans 448 0 0 0 reg_addr[8]
port 11 nsew signal input
flabel metal3 s 0 7840 800 7952 0 FreeSans 448 0 0 0 reg_addr[9]
port 12 nsew signal input
flabel metal3 s 0 22400 800 22512 0 FreeSans 448 0 0 0 reg_be[0]
port 13 nsew signal input
flabel metal3 s 0 21280 800 21392 0 FreeSans 448 0 0 0 reg_be[1]
port 14 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 reg_be[2]
port 15 nsew signal input
flabel metal3 s 0 19040 800 19152 0 FreeSans 448 0 0 0 reg_be[3]
port 16 nsew signal input
flabel metal3 s 0 4480 800 4592 0 FreeSans 448 0 0 0 reg_cs
port 17 nsew signal input
flabel metal3 s 0 94080 800 94192 0 FreeSans 448 0 0 0 reg_rdata[0]
port 18 nsew signal tristate
flabel metal3 s 0 82880 800 82992 0 FreeSans 448 0 0 0 reg_rdata[10]
port 19 nsew signal tristate
flabel metal3 s 0 81760 800 81872 0 FreeSans 448 0 0 0 reg_rdata[11]
port 20 nsew signal tristate
flabel metal3 s 0 80640 800 80752 0 FreeSans 448 0 0 0 reg_rdata[12]
port 21 nsew signal tristate
flabel metal3 s 0 79520 800 79632 0 FreeSans 448 0 0 0 reg_rdata[13]
port 22 nsew signal tristate
flabel metal3 s 0 78400 800 78512 0 FreeSans 448 0 0 0 reg_rdata[14]
port 23 nsew signal tristate
flabel metal3 s 0 77280 800 77392 0 FreeSans 448 0 0 0 reg_rdata[15]
port 24 nsew signal tristate
flabel metal3 s 0 76160 800 76272 0 FreeSans 448 0 0 0 reg_rdata[16]
port 25 nsew signal tristate
flabel metal3 s 0 75040 800 75152 0 FreeSans 448 0 0 0 reg_rdata[17]
port 26 nsew signal tristate
flabel metal3 s 0 73920 800 74032 0 FreeSans 448 0 0 0 reg_rdata[18]
port 27 nsew signal tristate
flabel metal3 s 0 72800 800 72912 0 FreeSans 448 0 0 0 reg_rdata[19]
port 28 nsew signal tristate
flabel metal3 s 0 92960 800 93072 0 FreeSans 448 0 0 0 reg_rdata[1]
port 29 nsew signal tristate
flabel metal3 s 0 71680 800 71792 0 FreeSans 448 0 0 0 reg_rdata[20]
port 30 nsew signal tristate
flabel metal3 s 0 70560 800 70672 0 FreeSans 448 0 0 0 reg_rdata[21]
port 31 nsew signal tristate
flabel metal3 s 0 69440 800 69552 0 FreeSans 448 0 0 0 reg_rdata[22]
port 32 nsew signal tristate
flabel metal3 s 0 68320 800 68432 0 FreeSans 448 0 0 0 reg_rdata[23]
port 33 nsew signal tristate
flabel metal3 s 0 67200 800 67312 0 FreeSans 448 0 0 0 reg_rdata[24]
port 34 nsew signal tristate
flabel metal3 s 0 66080 800 66192 0 FreeSans 448 0 0 0 reg_rdata[25]
port 35 nsew signal tristate
flabel metal3 s 0 64960 800 65072 0 FreeSans 448 0 0 0 reg_rdata[26]
port 36 nsew signal tristate
flabel metal3 s 0 63840 800 63952 0 FreeSans 448 0 0 0 reg_rdata[27]
port 37 nsew signal tristate
flabel metal3 s 0 62720 800 62832 0 FreeSans 448 0 0 0 reg_rdata[28]
port 38 nsew signal tristate
flabel metal3 s 0 61600 800 61712 0 FreeSans 448 0 0 0 reg_rdata[29]
port 39 nsew signal tristate
flabel metal3 s 0 91840 800 91952 0 FreeSans 448 0 0 0 reg_rdata[2]
port 40 nsew signal tristate
flabel metal3 s 0 60480 800 60592 0 FreeSans 448 0 0 0 reg_rdata[30]
port 41 nsew signal tristate
flabel metal3 s 0 59360 800 59472 0 FreeSans 448 0 0 0 reg_rdata[31]
port 42 nsew signal tristate
flabel metal3 s 0 90720 800 90832 0 FreeSans 448 0 0 0 reg_rdata[3]
port 43 nsew signal tristate
flabel metal3 s 0 89600 800 89712 0 FreeSans 448 0 0 0 reg_rdata[4]
port 44 nsew signal tristate
flabel metal3 s 0 88480 800 88592 0 FreeSans 448 0 0 0 reg_rdata[5]
port 45 nsew signal tristate
flabel metal3 s 0 87360 800 87472 0 FreeSans 448 0 0 0 reg_rdata[6]
port 46 nsew signal tristate
flabel metal3 s 0 86240 800 86352 0 FreeSans 448 0 0 0 reg_rdata[7]
port 47 nsew signal tristate
flabel metal3 s 0 85120 800 85232 0 FreeSans 448 0 0 0 reg_rdata[8]
port 48 nsew signal tristate
flabel metal3 s 0 84000 800 84112 0 FreeSans 448 0 0 0 reg_rdata[9]
port 49 nsew signal tristate
flabel metal3 s 0 58240 800 58352 0 FreeSans 448 0 0 0 reg_wdata[0]
port 50 nsew signal input
flabel metal3 s 0 47040 800 47152 0 FreeSans 448 0 0 0 reg_wdata[10]
port 51 nsew signal input
flabel metal3 s 0 45920 800 46032 0 FreeSans 448 0 0 0 reg_wdata[11]
port 52 nsew signal input
flabel metal3 s 0 44800 800 44912 0 FreeSans 448 0 0 0 reg_wdata[12]
port 53 nsew signal input
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 reg_wdata[13]
port 54 nsew signal input
flabel metal3 s 0 42560 800 42672 0 FreeSans 448 0 0 0 reg_wdata[14]
port 55 nsew signal input
flabel metal3 s 0 41440 800 41552 0 FreeSans 448 0 0 0 reg_wdata[15]
port 56 nsew signal input
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 reg_wdata[16]
port 57 nsew signal input
flabel metal3 s 0 39200 800 39312 0 FreeSans 448 0 0 0 reg_wdata[17]
port 58 nsew signal input
flabel metal3 s 0 38080 800 38192 0 FreeSans 448 0 0 0 reg_wdata[18]
port 59 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 reg_wdata[19]
port 60 nsew signal input
flabel metal3 s 0 57120 800 57232 0 FreeSans 448 0 0 0 reg_wdata[1]
port 61 nsew signal input
flabel metal3 s 0 35840 800 35952 0 FreeSans 448 0 0 0 reg_wdata[20]
port 62 nsew signal input
flabel metal3 s 0 34720 800 34832 0 FreeSans 448 0 0 0 reg_wdata[21]
port 63 nsew signal input
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 reg_wdata[22]
port 64 nsew signal input
flabel metal3 s 0 32480 800 32592 0 FreeSans 448 0 0 0 reg_wdata[23]
port 65 nsew signal input
flabel metal3 s 0 31360 800 31472 0 FreeSans 448 0 0 0 reg_wdata[24]
port 66 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 reg_wdata[25]
port 67 nsew signal input
flabel metal3 s 0 29120 800 29232 0 FreeSans 448 0 0 0 reg_wdata[26]
port 68 nsew signal input
flabel metal3 s 0 28000 800 28112 0 FreeSans 448 0 0 0 reg_wdata[27]
port 69 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 reg_wdata[28]
port 70 nsew signal input
flabel metal3 s 0 25760 800 25872 0 FreeSans 448 0 0 0 reg_wdata[29]
port 71 nsew signal input
flabel metal3 s 0 56000 800 56112 0 FreeSans 448 0 0 0 reg_wdata[2]
port 72 nsew signal input
flabel metal3 s 0 24640 800 24752 0 FreeSans 448 0 0 0 reg_wdata[30]
port 73 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 reg_wdata[31]
port 74 nsew signal input
flabel metal3 s 0 54880 800 54992 0 FreeSans 448 0 0 0 reg_wdata[3]
port 75 nsew signal input
flabel metal3 s 0 53760 800 53872 0 FreeSans 448 0 0 0 reg_wdata[4]
port 76 nsew signal input
flabel metal3 s 0 52640 800 52752 0 FreeSans 448 0 0 0 reg_wdata[5]
port 77 nsew signal input
flabel metal3 s 0 51520 800 51632 0 FreeSans 448 0 0 0 reg_wdata[6]
port 78 nsew signal input
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 reg_wdata[7]
port 79 nsew signal input
flabel metal3 s 0 49280 800 49392 0 FreeSans 448 0 0 0 reg_wdata[8]
port 80 nsew signal input
flabel metal3 s 0 48160 800 48272 0 FreeSans 448 0 0 0 reg_wdata[9]
port 81 nsew signal input
flabel metal3 s 0 5600 800 5712 0 FreeSans 448 0 0 0 reg_wr
port 82 nsew signal input
flabel metal2 s 9856 99200 9968 100000 0 FreeSans 448 90 0 0 rtc_clk
port 83 nsew signal input
flabel metal2 s 29792 99200 29904 100000 0 FreeSans 448 90 0 0 rtc_intr
port 84 nsew signal tristate
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 s_reset_n
port 85 nsew signal input
flabel metal4 s 3988 3076 5228 96492 0 FreeSans 5120 90 0 0 vdd
port 86 nsew power bidirectional
flabel metal4 s 23988 3076 25228 96492 0 FreeSans 5120 90 0 0 vdd
port 86 nsew power bidirectional
flabel metal4 s 13988 3076 15228 96492 0 FreeSans 5120 90 0 0 vss
port 87 nsew ground bidirectional
flabel metal4 s 33988 3076 35228 96492 0 FreeSans 5120 90 0 0 vss
port 87 nsew ground bidirectional
rlabel metal1 19992 96432 19992 96432 0 vdd
rlabel metal1 19992 95648 19992 95648 0 vss
rlabel metal2 22344 5432 22344 5432 0 clknet_0_mclk
rlabel metal2 22008 23184 22008 23184 0 clknet_0_rtc_clk
rlabel metal2 16856 5432 16856 5432 0 clknet_1_0__leaf_mclk
rlabel metal2 25368 5544 25368 5544 0 clknet_1_1__leaf_mclk
rlabel metal2 1848 4312 1848 4312 0 clknet_4_0_0_rtc_clk
rlabel metal2 3192 74536 3192 74536 0 clknet_4_10_0_rtc_clk
rlabel metal2 15456 73192 15456 73192 0 clknet_4_11_0_rtc_clk
rlabel metal2 25816 47824 25816 47824 0 clknet_4_12_0_rtc_clk
rlabel metal2 25368 63112 25368 63112 0 clknet_4_13_0_rtc_clk
rlabel metal3 22344 85848 22344 85848 0 clknet_4_14_0_rtc_clk
rlabel metal2 25256 67816 25256 67816 0 clknet_4_15_0_rtc_clk
rlabel metal3 16632 16856 16632 16856 0 clknet_4_1_0_rtc_clk
rlabel metal2 1848 41944 1848 41944 0 clknet_4_2_0_rtc_clk
rlabel metal2 15512 39648 15512 39648 0 clknet_4_3_0_rtc_clk
rlabel metal3 20552 15288 20552 15288 0 clknet_4_4_0_rtc_clk
rlabel metal2 28392 11648 28392 11648 0 clknet_4_5_0_rtc_clk
rlabel metal2 21784 39648 21784 39648 0 clknet_4_6_0_rtc_clk
rlabel metal2 26264 43848 26264 43848 0 clknet_4_7_0_rtc_clk
rlabel metal2 1848 53368 1848 53368 0 clknet_4_8_0_rtc_clk
rlabel metal2 16688 62552 16688 62552 0 clknet_4_9_0_rtc_clk
rlabel metal2 29848 3598 29848 3598 0 mclk
rlabel metal2 30240 96040 30240 96040 0 net1
rlabel metal3 24248 66024 24248 66024 0 net10
rlabel metal2 25704 62664 25704 62664 0 net11
rlabel metal2 15400 47040 15400 47040 0 net12
rlabel metal2 17752 85736 17752 85736 0 net13
rlabel metal3 24696 85736 24696 85736 0 net14
rlabel metal2 27384 12656 27384 12656 0 net15
rlabel metal3 24752 26152 24752 26152 0 net16
rlabel metal2 15176 21448 15176 21448 0 net17
rlabel metal3 24192 40936 24192 40936 0 net18
rlabel metal3 25088 24808 25088 24808 0 net19
rlabel metal2 15736 16128 15736 16128 0 net2
rlabel metal2 20776 62888 20776 62888 0 net20
rlabel metal2 21560 66304 21560 66304 0 net21
rlabel metal2 24696 7392 24696 7392 0 net22
rlabel metal3 18088 7672 18088 7672 0 net23
rlabel metal3 1246 95256 1246 95256 0 net24
rlabel metal3 1246 94136 1246 94136 0 net25
rlabel metal3 1246 93016 1246 93016 0 net26
rlabel metal3 1246 91896 1246 91896 0 net27
rlabel metal3 1246 90776 1246 90776 0 net28
rlabel metal3 1246 89656 1246 89656 0 net29
rlabel metal2 26264 48664 26264 48664 0 net3
rlabel metal3 1246 88536 1246 88536 0 net30
rlabel metal3 1246 87416 1246 87416 0 net31
rlabel metal3 1246 86296 1246 86296 0 net32
rlabel metal3 1246 85176 1246 85176 0 net33
rlabel metal3 1246 84056 1246 84056 0 net34
rlabel metal3 1246 82936 1246 82936 0 net35
rlabel metal3 1246 81816 1246 81816 0 net36
rlabel metal3 1246 80696 1246 80696 0 net37
rlabel metal3 1246 79576 1246 79576 0 net38
rlabel metal3 1246 78456 1246 78456 0 net39
rlabel metal2 15792 31752 15792 31752 0 net4
rlabel metal2 1736 77224 1736 77224 0 net40
rlabel metal3 1246 76216 1246 76216 0 net41
rlabel metal3 1246 75096 1246 75096 0 net42
rlabel metal2 2184 73920 2184 73920 0 net43
rlabel metal3 1246 72856 1246 72856 0 net44
rlabel metal3 1246 71736 1246 71736 0 net45
rlabel metal3 1246 70616 1246 70616 0 net46
rlabel metal3 1246 69496 1246 69496 0 net47
rlabel metal3 1246 68376 1246 68376 0 net48
rlabel metal3 1246 67256 1246 67256 0 net49
rlabel metal2 20776 65632 20776 65632 0 net5
rlabel metal3 1470 66136 1470 66136 0 net50
rlabel metal3 1246 65016 1246 65016 0 net51
rlabel metal3 1246 63896 1246 63896 0 net52
rlabel metal3 1246 62776 1246 62776 0 net53
rlabel metal3 1246 61656 1246 61656 0 net54
rlabel metal3 1246 60536 1246 60536 0 net55
rlabel metal3 1246 59416 1246 59416 0 net56
rlabel metal3 28672 9128 28672 9128 0 net57
rlabel metal2 27608 7504 27608 7504 0 net58
rlabel metal2 20440 4200 20440 4200 0 net59
rlabel metal2 21392 17416 21392 17416 0 net6
rlabel metal2 22904 8512 22904 8512 0 net60
rlabel metal2 22232 5992 22232 5992 0 net61
rlabel metal2 19320 46760 19320 46760 0 net62
rlabel metal3 21056 4424 21056 4424 0 net63
rlabel metal2 25816 9464 25816 9464 0 net64
rlabel metal2 13944 3976 13944 3976 0 net65
rlabel metal2 26320 6776 26320 6776 0 net66
rlabel metal3 14672 6776 14672 6776 0 net67
rlabel metal2 21784 3976 21784 3976 0 net68
rlabel metal3 17472 3416 17472 3416 0 net69
rlabel metal3 28224 14280 28224 14280 0 net7
rlabel metal2 19656 39760 19656 39760 0 net8
rlabel metal2 21224 26600 21224 26600 0 net9
rlabel metal2 2632 16744 2632 16744 0 reg_addr[2]
rlabel metal2 1792 15848 1792 15848 0 reg_addr[3]
rlabel metal3 2296 24584 2296 24584 0 reg_addr[4]
rlabel metal2 1904 23688 1904 23688 0 reg_be[0]
rlabel metal2 1848 21728 1848 21728 0 reg_be[1]
rlabel metal2 2520 20384 2520 20384 0 reg_be[2]
rlabel metal2 2520 19544 2520 19544 0 reg_be[3]
rlabel metal3 1638 58296 1638 58296 0 reg_wdata[0]
rlabel metal2 2184 47152 2184 47152 0 reg_wdata[10]
rlabel metal3 1638 45976 1638 45976 0 reg_wdata[11]
rlabel metal2 2520 44912 2520 44912 0 reg_wdata[12]
rlabel metal3 1624 43792 1624 43792 0 reg_wdata[13]
rlabel metal3 2142 42616 2142 42616 0 reg_wdata[14]
rlabel metal2 2632 42000 2632 42000 0 reg_wdata[15]
rlabel metal2 2632 40656 2632 40656 0 reg_wdata[16]
rlabel metal2 2520 39312 2520 39312 0 reg_wdata[17]
rlabel metal2 2856 38752 2856 38752 0 reg_wdata[18]
rlabel metal2 2520 37072 2520 37072 0 reg_wdata[19]
rlabel metal2 2632 57344 2632 57344 0 reg_wdata[1]
rlabel metal2 2464 33208 2464 33208 0 reg_wdata[20]
rlabel metal2 2632 35504 2632 35504 0 reg_wdata[21]
rlabel metal2 2688 18984 2688 18984 0 reg_wdata[22]
rlabel metal2 1960 22064 1960 22064 0 reg_wdata[23]
rlabel metal2 2184 31304 2184 31304 0 reg_wdata[24]
rlabel metal2 2856 30296 2856 30296 0 reg_wdata[25]
rlabel metal2 2520 28672 2520 28672 0 reg_wdata[26]
rlabel metal2 2184 24416 2184 24416 0 reg_wdata[27]
rlabel metal2 2968 16912 2968 16912 0 reg_wdata[28]
rlabel metal3 1246 25816 1246 25816 0 reg_wdata[29]
rlabel metal3 1582 56056 1582 56056 0 reg_wdata[2]
rlabel metal3 1862 24696 1862 24696 0 reg_wdata[30]
rlabel metal2 2184 22960 2184 22960 0 reg_wdata[31]
rlabel metal2 2632 54992 2632 54992 0 reg_wdata[3]
rlabel metal2 2520 53760 2520 53760 0 reg_wdata[4]
rlabel metal2 2072 52752 2072 52752 0 reg_wdata[5]
rlabel metal3 1358 51576 1358 51576 0 reg_wdata[6]
rlabel metal3 1470 50456 1470 50456 0 reg_wdata[7]
rlabel metal2 2520 49504 2520 49504 0 reg_wdata[8]
rlabel metal3 1638 48216 1638 48216 0 reg_wdata[9]
rlabel metal2 2072 5712 2072 5712 0 reg_wr
rlabel metal2 12936 90440 12936 90440 0 rtc_clk
rlabel metal2 30072 96656 30072 96656 0 rtc_intr
rlabel metal2 25480 3864 25480 3864 0 s_reset_n
rlabel metal3 25368 4424 25368 4424 0 u_rst_sync.in_data_2s
rlabel metal2 20888 3584 20888 3584 0 u_rst_sync.in_data_s
rlabel metal2 28168 6944 28168 6944 0 u_rst_sync.srst_n
rlabel metal3 29400 45752 29400 45752 0 u_rtc.cfg_date\[0\]
rlabel metal3 29792 31080 29792 31080 0 u_rtc.cfg_date\[10\]
rlabel metal2 30464 26376 30464 26376 0 u_rtc.cfg_date\[11\]
rlabel metal3 25536 32312 25536 32312 0 u_rtc.cfg_date\[12\]
rlabel metal2 25704 27552 25704 27552 0 u_rtc.cfg_date\[16\]
rlabel metal3 21112 26488 21112 26488 0 u_rtc.cfg_date\[17\]
rlabel metal2 21784 23576 21784 23576 0 u_rtc.cfg_date\[18\]
rlabel metal2 23016 21000 23016 21000 0 u_rtc.cfg_date\[19\]
rlabel metal3 29792 48440 29792 48440 0 u_rtc.cfg_date\[1\]
rlabel metal2 25816 12376 25816 12376 0 u_rtc.cfg_date\[20\]
rlabel metal3 23128 12936 23128 12936 0 u_rtc.cfg_date\[21\]
rlabel metal2 18648 13496 18648 13496 0 u_rtc.cfg_date\[22\]
rlabel metal2 18648 21112 18648 21112 0 u_rtc.cfg_date\[23\]
rlabel metal2 15176 10752 15176 10752 0 u_rtc.cfg_date\[24\]
rlabel metal2 17080 22960 17080 22960 0 u_rtc.cfg_date\[25\]
rlabel metal2 11368 24472 11368 24472 0 u_rtc.cfg_date\[26\]
rlabel metal2 8792 21896 8792 21896 0 u_rtc.cfg_date\[27\]
rlabel metal2 5320 11480 5320 11480 0 u_rtc.cfg_date\[28\]
rlabel metal2 5320 15736 5320 15736 0 u_rtc.cfg_date\[29\]
rlabel metal2 30296 53368 30296 53368 0 u_rtc.cfg_date\[2\]
rlabel metal2 5432 11648 5432 11648 0 u_rtc.cfg_date\[30\]
rlabel metal2 5432 21056 5432 21056 0 u_rtc.cfg_date\[31\]
rlabel metal2 31304 53368 31304 53368 0 u_rtc.cfg_date\[3\]
rlabel metal2 24360 40600 24360 40600 0 u_rtc.cfg_date\[4\]
rlabel metal3 23520 41944 23520 41944 0 u_rtc.cfg_date\[5\]
rlabel metal3 29064 34328 29064 34328 0 u_rtc.cfg_date\[8\]
rlabel metal2 26488 36400 26488 36400 0 u_rtc.cfg_date\[9\]
rlabel metal2 27944 46928 27944 46928 0 u_rtc.cfg_fast_date
rlabel metal3 27944 63896 27944 63896 0 u_rtc.cfg_fast_time
rlabel metal3 11704 35448 11704 35448 0 u_rtc.cfg_hmode
rlabel metal2 1624 28280 1624 28280 0 u_rtc.cfg_rtc_capture
rlabel metal2 30800 62552 30800 62552 0 u_rtc.cfg_rtc_halt
rlabel metal2 26040 61936 26040 61936 0 u_rtc.cfg_rtc_reset
rlabel metal2 5320 30632 5320 30632 0 u_rtc.cfg_rtc_update
rlabel metal3 23128 85736 23128 85736 0 u_rtc.cfg_time\[0\]
rlabel metal2 19880 71960 19880 71960 0 u_rtc.cfg_time\[10\]
rlabel metal3 21448 62440 21448 62440 0 u_rtc.cfg_time\[11\]
rlabel metal2 4872 62664 4872 62664 0 u_rtc.cfg_time\[12\]
rlabel metal2 4872 51800 4872 51800 0 u_rtc.cfg_time\[13\]
rlabel metal3 5544 56728 5544 56728 0 u_rtc.cfg_time\[14\]
rlabel metal3 6496 46872 6496 46872 0 u_rtc.cfg_time\[16\]
rlabel metal3 5712 44184 5712 44184 0 u_rtc.cfg_time\[17\]
rlabel metal2 5320 40768 5320 40768 0 u_rtc.cfg_time\[18\]
rlabel metal3 8792 39032 8792 39032 0 u_rtc.cfg_time\[19\]
rlabel metal2 18088 86184 18088 86184 0 u_rtc.cfg_time\[1\]
rlabel metal2 3304 34496 3304 34496 0 u_rtc.cfg_time\[20\]
rlabel metal3 5544 34776 5544 34776 0 u_rtc.cfg_time\[21\]
rlabel metal2 16016 32760 16016 32760 0 u_rtc.cfg_time\[24\]
rlabel metal2 15400 30296 15400 30296 0 u_rtc.cfg_time\[25\]
rlabel metal2 13048 29512 13048 29512 0 u_rtc.cfg_time\[26\]
rlabel metal2 15624 85848 15624 85848 0 u_rtc.cfg_time\[2\]
rlabel metal2 19432 86968 19432 86968 0 u_rtc.cfg_time\[3\]
rlabel metal2 5320 83160 5320 83160 0 u_rtc.cfg_time\[4\]
rlabel metal2 5320 78288 5320 78288 0 u_rtc.cfg_time\[5\]
rlabel metal2 5488 75656 5488 75656 0 u_rtc.cfg_time\[6\]
rlabel via2 5432 67144 5432 67144 0 u_rtc.cfg_time\[8\]
rlabel metal2 22568 66472 22568 66472 0 u_rtc.cfg_time\[9\]
rlabel metal2 16520 21616 16520 21616 0 u_rtc.date_c\[0\]
rlabel metal3 15316 16968 15316 16968 0 u_rtc.date_c\[1\]
rlabel metal2 12096 20104 12096 20104 0 u_rtc.date_c\[2\]
rlabel metal2 10360 23072 10360 23072 0 u_rtc.date_c\[3\]
rlabel metal2 19320 45584 19320 45584 0 u_rtc.date_d\[0\]
rlabel metal2 17752 48888 17752 48888 0 u_rtc.date_d\[1\]
rlabel metal3 25256 50680 25256 50680 0 u_rtc.date_d\[2\]
rlabel metal2 23464 45528 23464 45528 0 u_rtc.date_d\[3\]
rlabel metal3 33320 38920 33320 38920 0 u_rtc.date_m\[0\]
rlabel metal2 26488 37464 26488 37464 0 u_rtc.date_m\[1\]
rlabel metal2 30408 31472 30408 31472 0 u_rtc.date_m\[2\]
rlabel metal2 33040 29400 33040 29400 0 u_rtc.date_m\[3\]
rlabel metal3 5880 20552 5880 20552 0 u_rtc.date_tc\[0\]
rlabel metal2 6328 15596 6328 15596 0 u_rtc.date_tc\[1\]
rlabel metal2 5880 16352 5880 16352 0 u_rtc.date_tc\[2\]
rlabel metal2 7112 16800 7112 16800 0 u_rtc.date_tc\[3\]
rlabel metal2 22960 38696 22960 38696 0 u_rtc.date_td\[0\]
rlabel metal2 26824 43344 26824 43344 0 u_rtc.date_td\[1\]
rlabel metal2 26376 19656 26376 19656 0 u_rtc.date_tm
rlabel metal3 23128 19992 23128 19992 0 u_rtc.date_ty\[0\]
rlabel metal3 24416 16856 24416 16856 0 u_rtc.date_ty\[1\]
rlabel metal3 21392 15176 21392 15176 0 u_rtc.date_ty\[2\]
rlabel metal3 21896 18200 21896 18200 0 u_rtc.date_ty\[3\]
rlabel metal2 24024 22456 24024 22456 0 u_rtc.date_y\[0\]
rlabel metal2 24696 21952 24696 21952 0 u_rtc.date_y\[1\]
rlabel metal3 22064 25704 22064 25704 0 u_rtc.date_y\[2\]
rlabel metal2 20440 21672 20440 21672 0 u_rtc.date_y\[3\]
rlabel metal2 8680 17248 8680 17248 0 u_rtc.inc_date_c
rlabel metal2 31752 42952 31752 42952 0 u_rtc.inc_date_d
rlabel metal2 30296 40152 30296 40152 0 u_rtc.inc_date_m
rlabel metal2 26600 42784 26600 42784 0 u_rtc.inc_date_td
rlabel metal2 28504 19880 28504 19880 0 u_rtc.inc_date_tm
rlabel metal3 25928 15960 25928 15960 0 u_rtc.inc_date_ty
rlabel metal2 26712 23744 26712 23744 0 u_rtc.inc_date_y
rlabel metal3 17304 34664 17304 34664 0 u_rtc.inc_time_dow
rlabel metal3 9464 48104 9464 48104 0 u_rtc.inc_time_h
rlabel metal2 8456 68040 8456 68040 0 u_rtc.inc_time_m
rlabel metal2 30296 64344 30296 64344 0 u_rtc.inc_time_s
rlabel metal2 10360 42448 10360 42448 0 u_rtc.inc_time_th
rlabel metal2 19992 65128 19992 65128 0 u_rtc.inc_time_tm
rlabel metal2 8512 80248 8512 80248 0 u_rtc.inc_time_ts
rlabel metal2 27272 8372 27272 8372 0 u_rtc.rst_rn
rlabel metal2 20664 7616 20664 7616 0 u_rtc.rst_sn
rlabel metal2 2408 6664 2408 6664 0 u_rtc.rtc_reg_ack
rlabel metal2 3136 17416 3136 17416 0 u_rtc.rtc_reg_addr\[2\]
rlabel metal3 3976 26264 3976 26264 0 u_rtc.rtc_reg_addr\[3\]
rlabel metal2 3192 25872 3192 25872 0 u_rtc.rtc_reg_addr\[4\]
rlabel metal3 3136 27048 3136 27048 0 u_rtc.rtc_reg_be\[0\]
rlabel metal2 7840 25704 7840 25704 0 u_rtc.rtc_reg_be\[1\]
rlabel metal2 4088 35840 4088 35840 0 u_rtc.rtc_reg_be\[2\]
rlabel metal2 5432 23016 5432 23016 0 u_rtc.rtc_reg_be\[3\]
rlabel metal3 3080 6384 3080 6384 0 u_rtc.rtc_reg_cs
rlabel metal3 15848 87584 15848 87584 0 u_rtc.rtc_reg_wdata\[0\]
rlabel metal2 25480 33992 25480 33992 0 u_rtc.rtc_reg_wdata\[10\]
rlabel metal2 21392 44072 21392 44072 0 u_rtc.rtc_reg_wdata\[11\]
rlabel metal2 3304 45080 3304 45080 0 u_rtc.rtc_reg_wdata\[12\]
rlabel metal3 4760 48888 4760 48888 0 u_rtc.rtc_reg_wdata\[13\]
rlabel metal2 4088 53536 4088 53536 0 u_rtc.rtc_reg_wdata\[14\]
rlabel metal2 3192 42672 3192 42672 0 u_rtc.rtc_reg_wdata\[15\]
rlabel metal2 19824 38920 19824 38920 0 u_rtc.rtc_reg_wdata\[16\]
rlabel metal2 3304 39256 3304 39256 0 u_rtc.rtc_reg_wdata\[17\]
rlabel metal2 19544 24808 19544 24808 0 u_rtc.rtc_reg_wdata\[18\]
rlabel metal3 21336 22456 21336 22456 0 u_rtc.rtc_reg_wdata\[19\]
rlabel metal2 3696 46312 3696 46312 0 u_rtc.rtc_reg_wdata\[1\]
rlabel metal2 22232 15680 22232 15680 0 u_rtc.rtc_reg_wdata\[20\]
rlabel metal2 3192 35840 3192 35840 0 u_rtc.rtc_reg_wdata\[21\]
rlabel metal2 3864 18368 3864 18368 0 u_rtc.rtc_reg_wdata\[22\]
rlabel metal2 2296 23184 2296 23184 0 u_rtc.rtc_reg_wdata\[23\]
rlabel metal2 14000 31528 14000 31528 0 u_rtc.rtc_reg_wdata\[24\]
rlabel metal2 3192 30408 3192 30408 0 u_rtc.rtc_reg_wdata\[25\]
rlabel metal2 2856 28560 2856 28560 0 u_rtc.rtc_reg_wdata\[26\]
rlabel metal2 2520 23128 2520 23128 0 u_rtc.rtc_reg_wdata\[27\]
rlabel metal2 3192 15848 3192 15848 0 u_rtc.rtc_reg_wdata\[28\]
rlabel metal2 3304 17192 3304 17192 0 u_rtc.rtc_reg_wdata\[29\]
rlabel metal2 24696 53760 24696 53760 0 u_rtc.rtc_reg_wdata\[2\]
rlabel metal2 3304 18424 3304 18424 0 u_rtc.rtc_reg_wdata\[30\]
rlabel metal2 2520 22288 2520 22288 0 u_rtc.rtc_reg_wdata\[31\]
rlabel metal2 3304 55328 3304 55328 0 u_rtc.rtc_reg_wdata\[3\]
rlabel metal3 22120 41272 22120 41272 0 u_rtc.rtc_reg_wdata\[4\]
rlabel metal2 3304 53032 3304 53032 0 u_rtc.rtc_reg_wdata\[5\]
rlabel metal2 3192 71680 3192 71680 0 u_rtc.rtc_reg_wdata\[6\]
rlabel metal3 3472 64568 3472 64568 0 u_rtc.rtc_reg_wdata\[7\]
rlabel metal2 3248 49672 3248 49672 0 u_rtc.rtc_reg_wdata\[8\]
rlabel metal2 3304 48328 3304 48328 0 u_rtc.rtc_reg_wdata\[9\]
rlabel metal2 3248 5992 3248 5992 0 u_rtc.rtc_reg_wr
rlabel metal2 18032 48104 18032 48104 0 u_rtc.time_dow\[0\]
rlabel metal2 16744 47320 16744 47320 0 u_rtc.time_dow\[1\]
rlabel metal2 15792 49224 15792 49224 0 u_rtc.time_dow\[2\]
rlabel metal2 12600 43176 12600 43176 0 u_rtc.time_h\[0\]
rlabel metal2 17416 56784 17416 56784 0 u_rtc.time_h\[1\]
rlabel metal2 15960 55552 15960 55552 0 u_rtc.time_h\[2\]
rlabel metal2 15456 55048 15456 55048 0 u_rtc.time_h\[3\]
rlabel metal2 7896 65968 7896 65968 0 u_rtc.time_m\[0\]
rlabel metal2 19208 68376 19208 68376 0 u_rtc.time_m\[1\]
rlabel metal2 17752 57344 17752 57344 0 u_rtc.time_m\[2\]
rlabel metal2 18200 62832 18200 62832 0 u_rtc.time_m\[3\]
rlabel metal2 22568 80976 22568 80976 0 u_rtc.time_s\[0\]
rlabel metal2 16912 82936 16912 82936 0 u_rtc.time_s\[1\]
rlabel metal2 16296 83048 16296 83048 0 u_rtc.time_s\[2\]
rlabel metal2 15288 79688 15288 79688 0 u_rtc.time_s\[3\]
rlabel metal2 7560 33264 7560 33264 0 u_rtc.time_th\[0\]
rlabel metal2 8792 35560 8792 35560 0 u_rtc.time_th\[1\]
rlabel metal2 7168 63112 7168 63112 0 u_rtc.time_tm\[0\]
rlabel metal2 15456 49784 15456 49784 0 u_rtc.time_tm\[1\]
rlabel metal2 18200 53984 18200 53984 0 u_rtc.time_tm\[2\]
rlabel metal3 7784 80136 7784 80136 0 u_rtc.time_ts\[0\]
rlabel metal2 10360 80640 10360 80640 0 u_rtc.time_ts\[1\]
rlabel metal2 6720 74648 6720 74648 0 u_rtc.time_ts\[2\]
rlabel metal3 16856 5880 16856 5880 0 u_rtc.u_async_reg_bus._000_
rlabel metal2 2184 6720 2184 6720 0 u_rtc.u_async_reg_bus._001_
rlabel metal2 6328 6832 6328 6832 0 u_rtc.u_async_reg_bus._002_
rlabel metal2 9856 5096 9856 5096 0 u_rtc.u_async_reg_bus._003_
rlabel metal2 9128 5208 9128 5208 0 u_rtc.u_async_reg_bus._004_
rlabel metal2 17752 7448 17752 7448 0 u_rtc.u_async_reg_bus._038_
rlabel metal2 18368 7448 18368 7448 0 u_rtc.u_async_reg_bus._039_
rlabel metal2 19768 7840 19768 7840 0 u_rtc.u_async_reg_bus._040_
rlabel metal2 20328 7504 20328 7504 0 u_rtc.u_async_reg_bus._041_
rlabel metal2 19768 4760 19768 4760 0 u_rtc.u_async_reg_bus._042_
rlabel metal3 7224 6552 7224 6552 0 u_rtc.u_async_reg_bus._043_
rlabel metal3 19376 8120 19376 8120 0 u_rtc.u_async_reg_bus._044_
rlabel metal2 18312 6328 18312 6328 0 u_rtc.u_async_reg_bus._045_
rlabel metal2 17528 6272 17528 6272 0 u_rtc.u_async_reg_bus._046_
rlabel metal2 17640 8288 17640 8288 0 u_rtc.u_async_reg_bus._047_
rlabel metal2 8792 6048 8792 6048 0 u_rtc.u_async_reg_bus._048_
rlabel metal2 6440 4816 6440 4816 0 u_rtc.u_async_reg_bus._049_
rlabel metal2 5712 6664 5712 6664 0 u_rtc.u_async_reg_bus._050_
rlabel metal2 5768 6944 5768 6944 0 u_rtc.u_async_reg_bus._051_
rlabel metal2 5992 5488 5992 5488 0 u_rtc.u_async_reg_bus._052_
rlabel metal2 8960 6104 8960 6104 0 u_rtc.u_async_reg_bus._053_
rlabel metal3 8344 6888 8344 6888 0 u_rtc.u_async_reg_bus._054_
rlabel metal2 8456 6776 8456 6776 0 u_rtc.u_async_reg_bus._055_
rlabel metal2 8736 4424 8736 4424 0 u_rtc.u_async_reg_bus._056_
rlabel metal2 18424 8624 18424 8624 0 u_rtc.u_async_reg_bus._091_
rlabel metal2 16744 6608 16744 6608 0 u_rtc.u_async_reg_bus.in_flag
rlabel metal3 13496 6552 13496 6552 0 u_rtc.u_async_reg_bus.in_flag_s
rlabel metal2 8568 5824 8568 5824 0 u_rtc.u_async_reg_bus.in_flag_ss
rlabel metal2 20776 6272 20776 6272 0 u_rtc.u_async_reg_bus.in_state\[0\]
rlabel metal2 21224 7952 21224 7952 0 u_rtc.u_async_reg_bus.in_state\[1\]
rlabel metal2 10136 4984 10136 4984 0 u_rtc.u_async_reg_bus.out_flag
rlabel metal2 17976 3752 17976 3752 0 u_rtc.u_async_reg_bus.out_flag_s
rlabel metal2 16968 4032 16968 4032 0 u_rtc.u_async_reg_bus.out_flag_ss
rlabel metal2 7896 6720 7896 6720 0 u_rtc.u_async_reg_bus.out_state\[0\]
rlabel metal2 6664 6888 6664 6888 0 u_rtc.u_async_reg_bus.out_state\[1\]
rlabel metal3 28448 65464 28448 65464 0 u_rtc.u_core._000_
rlabel metal2 32536 30520 32536 30520 0 u_rtc.u_core._001_
rlabel metal2 29624 36904 29624 36904 0 u_rtc.u_core._002_
rlabel metal2 30744 28728 30744 28728 0 u_rtc.u_core._003_
rlabel metal2 31192 25760 31192 25760 0 u_rtc.u_core._004_
rlabel metal2 29736 57064 29736 57064 0 u_rtc.u_core._005_
rlabel metal2 29904 60088 29904 60088 0 u_rtc.u_core._006_
rlabel metal2 31752 59696 31752 59696 0 u_rtc.u_core._007_
rlabel metal2 33768 56448 33768 56448 0 u_rtc.u_core._008_
rlabel metal2 35280 54488 35280 54488 0 u_rtc.u_core._009_
rlabel metal2 35336 57344 35336 57344 0 u_rtc.u_core._010_
rlabel metal2 35504 60760 35504 60760 0 u_rtc.u_core._011_
rlabel metal2 34440 62384 34440 62384 0 u_rtc.u_core._012_
rlabel metal2 34664 65184 34664 65184 0 u_rtc.u_core._013_
rlabel metal2 34552 67144 34552 67144 0 u_rtc.u_core._014_
rlabel metal2 34440 70280 34440 70280 0 u_rtc.u_core._015_
rlabel metal2 33544 70280 33544 70280 0 u_rtc.u_core._016_
rlabel metal2 30744 69552 30744 69552 0 u_rtc.u_core._017_
rlabel metal2 29624 66920 29624 66920 0 u_rtc.u_core._018_
rlabel metal2 29288 67480 29288 67480 0 u_rtc.u_core._019_
rlabel metal2 11032 11648 11032 11648 0 u_rtc.u_core._020_
rlabel metal2 8232 15512 8232 15512 0 u_rtc.u_core._021_
rlabel metal2 8680 12208 8680 12208 0 u_rtc.u_core._022_
rlabel metal2 6104 17192 6104 17192 0 u_rtc.u_core._023_
rlabel metal2 16016 12152 16016 12152 0 u_rtc.u_core._024_
rlabel metal2 16632 17976 16632 17976 0 u_rtc.u_core._025_
rlabel metal2 11592 22792 11592 22792 0 u_rtc.u_core._026_
rlabel metal2 10136 20720 10136 20720 0 u_rtc.u_core._027_
rlabel metal2 25928 14616 25928 14616 0 u_rtc.u_core._028_
rlabel metal2 26936 14784 26936 14784 0 u_rtc.u_core._029_
rlabel metal2 19208 16016 19208 16016 0 u_rtc.u_core._030_
rlabel metal2 18088 18704 18088 18704 0 u_rtc.u_core._031_
rlabel metal2 30632 23240 30632 23240 0 u_rtc.u_core._032_
rlabel metal2 23240 26544 23240 26544 0 u_rtc.u_core._033_
rlabel metal2 26152 25200 26152 25200 0 u_rtc.u_core._034_
rlabel metal3 31304 19768 31304 19768 0 u_rtc.u_core._035_
rlabel metal3 29960 20776 29960 20776 0 u_rtc.u_core._036_
rlabel metal2 26488 40656 26488 40656 0 u_rtc.u_core._037_
rlabel metal2 27272 41608 27272 41608 0 u_rtc.u_core._038_
rlabel metal2 31192 45584 31192 45584 0 u_rtc.u_core._039_
rlabel metal2 32536 48328 32536 48328 0 u_rtc.u_core._040_
rlabel metal2 31976 52136 31976 52136 0 u_rtc.u_core._041_
rlabel metal2 32200 51240 32200 51240 0 u_rtc.u_core._042_
rlabel metal2 17864 33992 17864 33992 0 u_rtc.u_core._043_
rlabel metal2 17752 30520 17752 30520 0 u_rtc.u_core._044_
rlabel metal2 15512 28336 15512 28336 0 u_rtc.u_core._045_
rlabel metal2 8288 33992 8288 33992 0 u_rtc.u_core._046_
rlabel metal2 7112 34552 7112 34552 0 u_rtc.u_core._047_
rlabel metal2 7448 48440 7448 48440 0 u_rtc.u_core._048_
rlabel metal2 7560 45136 7560 45136 0 u_rtc.u_core._049_
rlabel metal2 11760 40376 11760 40376 0 u_rtc.u_core._050_
rlabel metal2 11928 40096 11928 40096 0 u_rtc.u_core._051_
rlabel metal2 5824 61544 5824 61544 0 u_rtc.u_core._052_
rlabel metal2 6104 52472 6104 52472 0 u_rtc.u_core._053_
rlabel metal2 4200 56168 4200 56168 0 u_rtc.u_core._054_
rlabel metal2 8456 66808 8456 66808 0 u_rtc.u_core._055_
rlabel metal2 24472 67928 24472 67928 0 u_rtc.u_core._056_
rlabel metal2 20328 71456 20328 71456 0 u_rtc.u_core._057_
rlabel metal3 19880 62328 19880 62328 0 u_rtc.u_core._058_
rlabel metal2 6104 80864 6104 80864 0 u_rtc.u_core._059_
rlabel metal2 3304 79296 3304 79296 0 u_rtc.u_core._060_
rlabel metal2 3640 75152 3640 75152 0 u_rtc.u_core._061_
rlabel metal2 22456 82264 22456 82264 0 u_rtc.u_core._062_
rlabel metal2 16296 80696 16296 80696 0 u_rtc.u_core._063_
rlabel metal3 14000 82712 14000 82712 0 u_rtc.u_core._064_
rlabel metal2 17528 82600 17528 82600 0 u_rtc.u_core._065_
rlabel metal2 7112 58128 7112 58128 0 u_rtc.u_core._066_
rlabel metal2 18088 63560 18088 63560 0 u_rtc.u_core._067_
rlabel metal2 7952 77784 7952 77784 0 u_rtc.u_core._068_
rlabel metal2 8344 79072 8344 79072 0 u_rtc.u_core._069_
rlabel metal3 9184 36344 9184 36344 0 u_rtc.u_core._070_
rlabel metal2 25816 16184 25816 16184 0 u_rtc.u_core._071_
rlabel metal2 35448 45416 35448 45416 0 u_rtc.u_core._072_
rlabel metal3 34272 46872 34272 46872 0 u_rtc.u_core._073_
rlabel metal2 33992 46872 33992 46872 0 u_rtc.u_core._074_
rlabel metal2 33208 47656 33208 47656 0 u_rtc.u_core._075_
rlabel metal2 31976 35504 31976 35504 0 u_rtc.u_core._076_
rlabel metal2 34888 35560 34888 35560 0 u_rtc.u_core._077_
rlabel metal2 35784 31696 35784 31696 0 u_rtc.u_core._078_
rlabel metal2 30184 27328 30184 27328 0 u_rtc.u_core._079_
rlabel metal2 27832 20104 27832 20104 0 u_rtc.u_core._080_
rlabel metal2 34216 39984 34216 39984 0 u_rtc.u_core._081_
rlabel metal2 25480 22400 25480 22400 0 u_rtc.u_core._082_
rlabel metal2 29680 22456 29680 22456 0 u_rtc.u_core._083_
rlabel metal3 23912 20776 23912 20776 0 u_rtc.u_core._084_
rlabel metal2 22120 18032 22120 18032 0 u_rtc.u_core._085_
rlabel metal2 23128 18032 23128 18032 0 u_rtc.u_core._086_
rlabel metal2 21672 16576 21672 16576 0 u_rtc.u_core._087_
rlabel metal3 21000 17640 21000 17640 0 u_rtc.u_core._088_
rlabel metal3 13216 15848 13216 15848 0 u_rtc.u_core._089_
rlabel metal2 14504 19040 14504 19040 0 u_rtc.u_core._090_
rlabel metal2 7784 15204 7784 15204 0 u_rtc.u_core._091_
rlabel metal3 8288 16856 8288 16856 0 u_rtc.u_core._092_
rlabel metal3 24192 13160 24192 13160 0 u_rtc.u_core._093_
rlabel metal2 27160 41440 27160 41440 0 u_rtc.u_core._094_
rlabel metal3 30576 46088 30576 46088 0 u_rtc.u_core._095_
rlabel metal2 32200 58688 32200 58688 0 u_rtc.u_core._096_
rlabel metal2 29792 59864 29792 59864 0 u_rtc.u_core._097_
rlabel metal2 13944 79352 13944 79352 0 u_rtc.u_core._098_
rlabel metal2 13832 79856 13832 79856 0 u_rtc.u_core._099_
rlabel metal2 6552 79128 6552 79128 0 u_rtc.u_core._100_
rlabel metal2 18760 67760 18760 67760 0 u_rtc.u_core._101_
rlabel metal2 17304 64400 17304 64400 0 u_rtc.u_core._102_
rlabel metal2 8008 56392 8008 56392 0 u_rtc.u_core._103_
rlabel metal3 8288 54488 8288 54488 0 u_rtc.u_core._104_
rlabel metal2 8344 56784 8344 56784 0 u_rtc.u_core._105_
rlabel metal3 10024 41944 10024 41944 0 u_rtc.u_core._106_
rlabel metal2 9128 41048 9128 41048 0 u_rtc.u_core._107_
rlabel metal3 9240 39592 9240 39592 0 u_rtc.u_core._108_
rlabel metal2 9464 40824 9464 40824 0 u_rtc.u_core._109_
rlabel metal2 8736 42168 8736 42168 0 u_rtc.u_core._110_
rlabel metal2 9576 41608 9576 41608 0 u_rtc.u_core._111_
rlabel metal2 9016 42840 9016 42840 0 u_rtc.u_core._112_
rlabel metal3 9184 42504 9184 42504 0 u_rtc.u_core._113_
rlabel metal2 9128 37688 9128 37688 0 u_rtc.u_core._114_
rlabel metal2 10248 37520 10248 37520 0 u_rtc.u_core._115_
rlabel metal2 10360 34104 10360 34104 0 u_rtc.u_core._116_
rlabel metal2 33880 31416 33880 31416 0 u_rtc.u_core._117_
rlabel metal2 34776 41496 34776 41496 0 u_rtc.u_core._118_
rlabel metal2 32256 39704 32256 39704 0 u_rtc.u_core._119_
rlabel metal2 32592 39032 32592 39032 0 u_rtc.u_core._120_
rlabel metal2 34328 42784 34328 42784 0 u_rtc.u_core._121_
rlabel metal3 34552 41944 34552 41944 0 u_rtc.u_core._122_
rlabel metal2 33544 38752 33544 38752 0 u_rtc.u_core._123_
rlabel metal3 32928 40152 32928 40152 0 u_rtc.u_core._124_
rlabel metal3 36568 38920 36568 38920 0 u_rtc.u_core._125_
rlabel metal3 35784 39032 35784 39032 0 u_rtc.u_core._126_
rlabel metal2 33656 34608 33656 34608 0 u_rtc.u_core._127_
rlabel metal2 34328 35504 34328 35504 0 u_rtc.u_core._128_
rlabel metal3 34552 40936 34552 40936 0 u_rtc.u_core._129_
rlabel metal2 36232 35616 36232 35616 0 u_rtc.u_core._130_
rlabel metal3 35448 45192 35448 45192 0 u_rtc.u_core._131_
rlabel metal2 36960 45192 36960 45192 0 u_rtc.u_core._132_
rlabel metal2 35784 41496 35784 41496 0 u_rtc.u_core._133_
rlabel metal2 36568 41188 36568 41188 0 u_rtc.u_core._134_
rlabel metal2 36456 35952 36456 35952 0 u_rtc.u_core._135_
rlabel metal2 36120 41832 36120 41832 0 u_rtc.u_core._136_
rlabel metal3 36176 34776 36176 34776 0 u_rtc.u_core._137_
rlabel metal2 32536 35224 32536 35224 0 u_rtc.u_core._138_
rlabel metal2 33992 33488 33992 33488 0 u_rtc.u_core._139_
rlabel metal3 33320 31080 33320 31080 0 u_rtc.u_core._140_
rlabel metal2 32984 32032 32984 32032 0 u_rtc.u_core._141_
rlabel metal3 33824 33320 33824 33320 0 u_rtc.u_core._142_
rlabel metal2 35672 34832 35672 34832 0 u_rtc.u_core._143_
rlabel metal2 37912 36064 37912 36064 0 u_rtc.u_core._144_
rlabel metal2 37800 43400 37800 43400 0 u_rtc.u_core._145_
rlabel metal2 37688 36456 37688 36456 0 u_rtc.u_core._146_
rlabel metal2 37128 41272 37128 41272 0 u_rtc.u_core._147_
rlabel metal2 32200 37184 32200 37184 0 u_rtc.u_core._148_
rlabel metal2 37352 37632 37352 37632 0 u_rtc.u_core._149_
rlabel metal3 34552 36344 34552 36344 0 u_rtc.u_core._150_
rlabel metal2 35000 33824 35000 33824 0 u_rtc.u_core._151_
rlabel metal2 37240 32872 37240 32872 0 u_rtc.u_core._152_
rlabel metal2 36400 34776 36400 34776 0 u_rtc.u_core._153_
rlabel metal2 33712 47208 33712 47208 0 u_rtc.u_core._154_
rlabel metal2 36120 33320 36120 33320 0 u_rtc.u_core._155_
rlabel metal2 33432 34496 33432 34496 0 u_rtc.u_core._156_
rlabel metal2 35784 34496 35784 34496 0 u_rtc.u_core._157_
rlabel metal2 36288 35000 36288 35000 0 u_rtc.u_core._158_
rlabel metal3 36232 34664 36232 34664 0 u_rtc.u_core._159_
rlabel metal2 37296 35896 37296 35896 0 u_rtc.u_core._160_
rlabel metal2 35168 35000 35168 35000 0 u_rtc.u_core._161_
rlabel metal2 36680 35784 36680 35784 0 u_rtc.u_core._162_
rlabel metal3 36792 39144 36792 39144 0 u_rtc.u_core._163_
rlabel metal3 35560 38696 35560 38696 0 u_rtc.u_core._164_
rlabel metal2 36176 35896 36176 35896 0 u_rtc.u_core._165_
rlabel metal2 38192 39816 38192 39816 0 u_rtc.u_core._166_
rlabel metal2 37576 40656 37576 40656 0 u_rtc.u_core._167_
rlabel metal2 37072 39704 37072 39704 0 u_rtc.u_core._168_
rlabel metal2 35504 41272 35504 41272 0 u_rtc.u_core._169_
rlabel metal2 37128 42112 37128 42112 0 u_rtc.u_core._170_
rlabel metal2 11928 17920 11928 17920 0 u_rtc.u_core._171_
rlabel metal2 15736 19208 15736 19208 0 u_rtc.u_core._172_
rlabel metal2 15400 18536 15400 18536 0 u_rtc.u_core._173_
rlabel metal2 21448 18928 21448 18928 0 u_rtc.u_core._174_
rlabel metal3 18984 18424 18984 18424 0 u_rtc.u_core._175_
rlabel metal2 16632 19264 16632 19264 0 u_rtc.u_core._176_
rlabel metal2 24248 20384 24248 20384 0 u_rtc.u_core._177_
rlabel metal3 31024 22568 31024 22568 0 u_rtc.u_core._178_
rlabel metal2 36008 44688 36008 44688 0 u_rtc.u_core._179_
rlabel metal2 35056 44184 35056 44184 0 u_rtc.u_core._180_
rlabel metal2 36288 42728 36288 42728 0 u_rtc.u_core._181_
rlabel metal2 35112 40488 35112 40488 0 u_rtc.u_core._182_
rlabel metal2 37352 42224 37352 42224 0 u_rtc.u_core._183_
rlabel metal2 33208 42448 33208 42448 0 u_rtc.u_core._184_
rlabel metal2 33656 41832 33656 41832 0 u_rtc.u_core._185_
rlabel metal2 31752 41384 31752 41384 0 u_rtc.u_core._186_
rlabel metal2 32312 42224 32312 42224 0 u_rtc.u_core._187_
rlabel metal2 31248 42728 31248 42728 0 u_rtc.u_core._188_
rlabel metal2 35224 38920 35224 38920 0 u_rtc.u_core._189_
rlabel metal3 33712 38808 33712 38808 0 u_rtc.u_core._190_
rlabel metal2 36008 39536 36008 39536 0 u_rtc.u_core._191_
rlabel metal2 38024 39984 38024 39984 0 u_rtc.u_core._192_
rlabel metal2 32424 41944 32424 41944 0 u_rtc.u_core._193_
rlabel metal3 31416 41160 31416 41160 0 u_rtc.u_core._194_
rlabel metal2 32816 34776 32816 34776 0 u_rtc.u_core._195_
rlabel metal2 27160 18928 27160 18928 0 u_rtc.u_core._196_
rlabel metal2 26376 21672 26376 21672 0 u_rtc.u_core._197_
rlabel metal2 25368 20888 25368 20888 0 u_rtc.u_core._198_
rlabel metal2 28280 21056 28280 21056 0 u_rtc.u_core._199_
rlabel metal2 23352 17416 23352 17416 0 u_rtc.u_core._200_
rlabel metal2 23688 18032 23688 18032 0 u_rtc.u_core._201_
rlabel metal2 18536 17136 18536 17136 0 u_rtc.u_core._202_
rlabel metal3 9464 16968 9464 16968 0 u_rtc.u_core._203_
rlabel metal2 11144 17528 11144 17528 0 u_rtc.u_core._204_
rlabel metal2 31528 66808 31528 66808 0 u_rtc.u_core._205_
rlabel metal2 30016 67592 30016 67592 0 u_rtc.u_core._206_
rlabel metal2 31304 58968 31304 58968 0 u_rtc.u_core._207_
rlabel metal3 33768 57624 33768 57624 0 u_rtc.u_core._208_
rlabel metal2 36904 58352 36904 58352 0 u_rtc.u_core._209_
rlabel metal3 36904 59976 36904 59976 0 u_rtc.u_core._210_
rlabel metal2 36008 62524 36008 62524 0 u_rtc.u_core._211_
rlabel metal2 37352 64960 37352 64960 0 u_rtc.u_core._212_
rlabel metal2 37352 66528 37352 66528 0 u_rtc.u_core._213_
rlabel metal2 35672 67088 35672 67088 0 u_rtc.u_core._214_
rlabel metal2 33432 70392 33432 70392 0 u_rtc.u_core._215_
rlabel metal2 32200 67480 32200 67480 0 u_rtc.u_core._216_
rlabel metal2 31416 67368 31416 67368 0 u_rtc.u_core._217_
rlabel metal2 31192 33376 31192 33376 0 u_rtc.u_core._218_
rlabel metal2 31864 33656 31864 33656 0 u_rtc.u_core._219_
rlabel metal2 28616 41328 28616 41328 0 u_rtc.u_core._220_
rlabel metal3 27160 41160 27160 41160 0 u_rtc.u_core._221_
rlabel metal2 30408 36848 30408 36848 0 u_rtc.u_core._222_
rlabel metal2 29904 36232 29904 36232 0 u_rtc.u_core._223_
rlabel metal2 29064 36568 29064 36568 0 u_rtc.u_core._224_
rlabel metal2 31080 32032 31080 32032 0 u_rtc.u_core._225_
rlabel metal2 29960 29064 29960 29064 0 u_rtc.u_core._226_
rlabel metal2 31080 30968 31080 30968 0 u_rtc.u_core._227_
rlabel metal2 30968 26544 30968 26544 0 u_rtc.u_core._228_
rlabel metal2 29960 60928 29960 60928 0 u_rtc.u_core._229_
rlabel metal3 30408 59864 30408 59864 0 u_rtc.u_core._230_
rlabel metal3 29232 58408 29232 58408 0 u_rtc.u_core._231_
rlabel metal3 32424 60760 32424 60760 0 u_rtc.u_core._232_
rlabel metal2 29624 60200 29624 60200 0 u_rtc.u_core._233_
rlabel metal2 31976 59920 31976 59920 0 u_rtc.u_core._234_
rlabel metal2 32312 59640 32312 59640 0 u_rtc.u_core._235_
rlabel metal2 34664 57120 34664 57120 0 u_rtc.u_core._236_
rlabel metal2 37464 55776 37464 55776 0 u_rtc.u_core._237_
rlabel metal2 35784 55664 35784 55664 0 u_rtc.u_core._238_
rlabel metal2 36456 57512 36456 57512 0 u_rtc.u_core._239_
rlabel metal2 36344 60816 36344 60816 0 u_rtc.u_core._240_
rlabel metal3 35504 63000 35504 63000 0 u_rtc.u_core._241_
rlabel metal2 36176 64680 36176 64680 0 u_rtc.u_core._242_
rlabel metal3 36512 67816 36512 67816 0 u_rtc.u_core._243_
rlabel metal2 35952 68824 35952 68824 0 u_rtc.u_core._244_
rlabel metal2 35672 69664 35672 69664 0 u_rtc.u_core._245_
rlabel metal2 35224 69720 35224 69720 0 u_rtc.u_core._246_
rlabel metal2 32088 70224 32088 70224 0 u_rtc.u_core._247_
rlabel metal2 31864 68320 31864 68320 0 u_rtc.u_core._248_
rlabel metal3 30072 67704 30072 67704 0 u_rtc.u_core._249_
rlabel metal2 30352 67704 30352 67704 0 u_rtc.u_core._250_
rlabel metal2 10584 12656 10584 12656 0 u_rtc.u_core._251_
rlabel metal2 11200 12936 11200 12936 0 u_rtc.u_core._252_
rlabel metal2 11536 12936 11536 12936 0 u_rtc.u_core._253_
rlabel metal3 7224 14504 7224 14504 0 u_rtc.u_core._254_
rlabel metal2 7168 15624 7168 15624 0 u_rtc.u_core._255_
rlabel metal2 8904 12992 8904 12992 0 u_rtc.u_core._256_
rlabel metal2 7560 16128 7560 16128 0 u_rtc.u_core._257_
rlabel metal2 8008 14616 8008 14616 0 u_rtc.u_core._258_
rlabel metal3 7896 15064 7896 15064 0 u_rtc.u_core._259_
rlabel metal3 6664 15400 6664 15400 0 u_rtc.u_core._260_
rlabel metal2 7000 11760 7000 11760 0 u_rtc.u_core._261_
rlabel metal2 7560 12208 7560 12208 0 u_rtc.u_core._262_
rlabel metal2 7560 13160 7560 13160 0 u_rtc.u_core._263_
rlabel metal2 8232 12544 8232 12544 0 u_rtc.u_core._264_
rlabel metal3 9296 12824 9296 12824 0 u_rtc.u_core._265_
rlabel metal2 7896 16184 7896 16184 0 u_rtc.u_core._266_
rlabel metal3 8064 16632 8064 16632 0 u_rtc.u_core._267_
rlabel metal2 7448 17920 7448 17920 0 u_rtc.u_core._268_
rlabel metal2 15456 10808 15456 10808 0 u_rtc.u_core._269_
rlabel metal2 15848 13048 15848 13048 0 u_rtc.u_core._270_
rlabel metal2 15064 19712 15064 19712 0 u_rtc.u_core._271_
rlabel metal2 16520 16632 16520 16632 0 u_rtc.u_core._272_
rlabel metal2 12320 20104 12320 20104 0 u_rtc.u_core._273_
rlabel metal2 12824 15624 12824 15624 0 u_rtc.u_core._274_
rlabel metal2 10472 20608 10472 20608 0 u_rtc.u_core._275_
rlabel metal3 14056 19208 14056 19208 0 u_rtc.u_core._276_
rlabel metal2 11256 23016 11256 23016 0 u_rtc.u_core._277_
rlabel metal3 11872 22232 11872 22232 0 u_rtc.u_core._278_
rlabel metal2 11592 20160 11592 20160 0 u_rtc.u_core._279_
rlabel metal2 12264 21112 12264 21112 0 u_rtc.u_core._280_
rlabel metal2 8904 20664 8904 20664 0 u_rtc.u_core._281_
rlabel metal3 10024 20104 10024 20104 0 u_rtc.u_core._282_
rlabel metal2 10752 20216 10752 20216 0 u_rtc.u_core._283_
rlabel metal3 26656 13496 26656 13496 0 u_rtc.u_core._284_
rlabel metal2 25256 15484 25256 15484 0 u_rtc.u_core._285_
rlabel metal2 26152 18200 26152 18200 0 u_rtc.u_core._286_
rlabel metal2 25872 15848 25872 15848 0 u_rtc.u_core._287_
rlabel metal2 24584 16128 24584 16128 0 u_rtc.u_core._288_
rlabel metal2 24808 16184 24808 16184 0 u_rtc.u_core._289_
rlabel metal2 19768 16044 19768 16044 0 u_rtc.u_core._290_
rlabel metal2 25480 20496 25480 20496 0 u_rtc.u_core._291_
rlabel metal2 21112 16800 21112 16800 0 u_rtc.u_core._292_
rlabel metal2 21448 16968 21448 16968 0 u_rtc.u_core._293_
rlabel metal3 20160 16632 20160 16632 0 u_rtc.u_core._294_
rlabel metal2 19208 19544 19208 19544 0 u_rtc.u_core._295_
rlabel metal2 19768 18032 19768 18032 0 u_rtc.u_core._296_
rlabel metal3 19768 19208 19768 19208 0 u_rtc.u_core._297_
rlabel metal2 26712 26096 26712 26096 0 u_rtc.u_core._298_
rlabel metal2 27048 23464 27048 23464 0 u_rtc.u_core._299_
rlabel metal2 24472 23800 24472 23800 0 u_rtc.u_core._300_
rlabel metal2 27048 24192 27048 24192 0 u_rtc.u_core._301_
rlabel metal3 23744 24024 23744 24024 0 u_rtc.u_core._302_
rlabel metal2 23128 24192 23128 24192 0 u_rtc.u_core._303_
rlabel metal3 26880 24584 26880 24584 0 u_rtc.u_core._304_
rlabel metal2 29736 20720 29736 20720 0 u_rtc.u_core._305_
rlabel metal2 26040 24304 26040 24304 0 u_rtc.u_core._306_
rlabel metal2 30688 19992 30688 19992 0 u_rtc.u_core._307_
rlabel metal3 30408 19880 30408 19880 0 u_rtc.u_core._308_
rlabel metal2 28056 19656 28056 19656 0 u_rtc.u_core._309_
rlabel metal2 29288 21000 29288 21000 0 u_rtc.u_core._310_
rlabel metal2 29176 21280 29176 21280 0 u_rtc.u_core._311_
rlabel metal2 24696 41216 24696 41216 0 u_rtc.u_core._312_
rlabel metal3 31976 48216 31976 48216 0 u_rtc.u_core._313_
rlabel metal3 24920 41048 24920 41048 0 u_rtc.u_core._314_
rlabel metal2 26656 41384 26656 41384 0 u_rtc.u_core._315_
rlabel metal2 26488 41664 26488 41664 0 u_rtc.u_core._316_
rlabel metal3 31864 47432 31864 47432 0 u_rtc.u_core._317_
rlabel metal2 30296 44352 30296 44352 0 u_rtc.u_core._318_
rlabel metal2 31080 45080 31080 45080 0 u_rtc.u_core._319_
rlabel metal3 33488 46760 33488 46760 0 u_rtc.u_core._320_
rlabel metal2 31416 47656 31416 47656 0 u_rtc.u_core._321_
rlabel metal2 31360 52920 31360 52920 0 u_rtc.u_core._322_
rlabel metal2 31696 49112 31696 49112 0 u_rtc.u_core._323_
rlabel metal3 33376 49000 33376 49000 0 u_rtc.u_core._324_
rlabel metal2 32424 52192 32424 52192 0 u_rtc.u_core._325_
rlabel metal3 30968 52136 30968 52136 0 u_rtc.u_core._326_
rlabel metal3 31640 49112 31640 49112 0 u_rtc.u_core._327_
rlabel metal2 16408 33712 16408 33712 0 u_rtc.u_core._328_
rlabel metal2 16968 34552 16968 34552 0 u_rtc.u_core._329_
rlabel metal2 17752 33488 17752 33488 0 u_rtc.u_core._330_
rlabel metal2 17304 34104 17304 34104 0 u_rtc.u_core._331_
rlabel metal3 16520 30744 16520 30744 0 u_rtc.u_core._332_
rlabel metal2 17976 31080 17976 31080 0 u_rtc.u_core._333_
rlabel metal2 18032 30744 18032 30744 0 u_rtc.u_core._334_
rlabel metal3 15176 27944 15176 27944 0 u_rtc.u_core._335_
rlabel metal2 17528 28840 17528 28840 0 u_rtc.u_core._336_
rlabel metal3 16856 27832 16856 27832 0 u_rtc.u_core._337_
rlabel metal2 7000 32760 7000 32760 0 u_rtc.u_core._338_
rlabel metal2 8456 34216 8456 34216 0 u_rtc.u_core._339_
rlabel metal2 9016 34888 9016 34888 0 u_rtc.u_core._340_
rlabel metal2 7336 34384 7336 34384 0 u_rtc.u_core._341_
rlabel metal3 9184 35784 9184 35784 0 u_rtc.u_core._342_
rlabel metal2 7448 34888 7448 34888 0 u_rtc.u_core._343_
rlabel metal2 7784 47880 7784 47880 0 u_rtc.u_core._344_
rlabel metal2 7672 49000 7672 49000 0 u_rtc.u_core._345_
rlabel metal2 7448 48272 7448 48272 0 u_rtc.u_core._346_
rlabel metal2 7336 44352 7336 44352 0 u_rtc.u_core._347_
rlabel metal2 8792 44016 8792 44016 0 u_rtc.u_core._348_
rlabel metal2 8008 44688 8008 44688 0 u_rtc.u_core._349_
rlabel metal2 7728 44520 7728 44520 0 u_rtc.u_core._350_
rlabel metal2 10696 41496 10696 41496 0 u_rtc.u_core._351_
rlabel metal2 11144 42000 11144 42000 0 u_rtc.u_core._352_
rlabel metal2 11760 43400 11760 43400 0 u_rtc.u_core._353_
rlabel metal2 12152 43288 12152 43288 0 u_rtc.u_core._354_
rlabel metal2 11368 42392 11368 42392 0 u_rtc.u_core._355_
rlabel metal3 9408 41048 9408 41048 0 u_rtc.u_core._356_
rlabel metal2 12600 42000 12600 42000 0 u_rtc.u_core._357_
rlabel metal2 9408 39704 9408 39704 0 u_rtc.u_core._358_
rlabel metal2 7224 61544 7224 61544 0 u_rtc.u_core._359_
rlabel metal2 7672 62552 7672 62552 0 u_rtc.u_core._360_
rlabel metal2 5264 52136 5264 52136 0 u_rtc.u_core._361_
rlabel metal2 6776 54432 6776 54432 0 u_rtc.u_core._362_
rlabel metal3 6216 53032 6216 53032 0 u_rtc.u_core._363_
rlabel metal2 7280 57848 7280 57848 0 u_rtc.u_core._364_
rlabel metal2 6104 57288 6104 57288 0 u_rtc.u_core._365_
rlabel metal2 6720 66472 6720 66472 0 u_rtc.u_core._366_
rlabel metal2 7560 67200 7560 67200 0 u_rtc.u_core._367_
rlabel metal3 20328 65352 20328 65352 0 u_rtc.u_core._368_
rlabel metal2 19656 65968 19656 65968 0 u_rtc.u_core._369_
rlabel metal3 20720 65240 20720 65240 0 u_rtc.u_core._370_
rlabel metal2 20944 65688 20944 65688 0 u_rtc.u_core._371_
rlabel metal2 19656 64120 19656 64120 0 u_rtc.u_core._372_
rlabel metal2 19880 67984 19880 67984 0 u_rtc.u_core._373_
rlabel metal2 19768 68768 19768 68768 0 u_rtc.u_core._374_
rlabel metal2 20104 69720 20104 69720 0 u_rtc.u_core._375_
rlabel metal2 19768 63056 19768 63056 0 u_rtc.u_core._376_
rlabel metal2 20216 62832 20216 62832 0 u_rtc.u_core._377_
rlabel metal3 20048 63000 20048 63000 0 u_rtc.u_core._378_
rlabel metal2 7896 80584 7896 80584 0 u_rtc.u_core._379_
rlabel metal2 5992 80752 5992 80752 0 u_rtc.u_core._380_
rlabel metal2 6104 77336 6104 77336 0 u_rtc.u_core._381_
rlabel metal2 7000 77616 7000 77616 0 u_rtc.u_core._382_
rlabel metal2 5376 78680 5376 78680 0 u_rtc.u_core._383_
rlabel metal3 3976 78904 3976 78904 0 u_rtc.u_core._384_
rlabel metal2 6384 75656 6384 75656 0 u_rtc.u_core._385_
rlabel metal3 5152 75768 5152 75768 0 u_rtc.u_core._386_
rlabel metal2 22288 81704 22288 81704 0 u_rtc.u_core._387_
rlabel metal2 22792 82544 22792 82544 0 u_rtc.u_core._388_
rlabel metal3 18648 83496 18648 83496 0 u_rtc.u_core._389_
rlabel metal2 16520 81312 16520 81312 0 u_rtc.u_core._390_
rlabel metal2 15960 81424 15960 81424 0 u_rtc.u_core._391_
rlabel metal3 17080 81144 17080 81144 0 u_rtc.u_core._392_
rlabel metal2 15176 80640 15176 80640 0 u_rtc.u_core._393_
rlabel metal3 17248 82712 17248 82712 0 u_rtc.u_core._394_
rlabel metal2 15064 81200 15064 81200 0 u_rtc.u_core._395_
rlabel metal3 15176 82040 15176 82040 0 u_rtc.u_core._396_
rlabel metal3 14952 82712 14952 82712 0 u_rtc.u_core._397_
rlabel metal3 18760 83384 18760 83384 0 u_rtc.u_core._398_
rlabel metal2 17416 83160 17416 83160 0 u_rtc.u_core._399_
rlabel metal2 29176 64624 29176 64624 0 u_rtc.u_core.pulse_1s
rlabel metal2 29624 46928 29624 46928 0 u_rtc.u_core.rtc_div\[0\]
rlabel metal2 36120 70560 36120 70560 0 u_rtc.u_core.rtc_div\[10\]
rlabel metal2 36344 70056 36344 70056 0 u_rtc.u_core.rtc_div\[11\]
rlabel metal2 33096 70392 33096 70392 0 u_rtc.u_core.rtc_div\[12\]
rlabel metal3 32312 66024 32312 66024 0 u_rtc.u_core.rtc_div\[13\]
rlabel metal3 31808 66808 31808 66808 0 u_rtc.u_core.rtc_div\[14\]
rlabel metal2 30632 61096 30632 61096 0 u_rtc.u_core.rtc_div\[1\]
rlabel metal2 32424 60480 32424 60480 0 u_rtc.u_core.rtc_div\[2\]
rlabel metal2 36792 56616 36792 56616 0 u_rtc.u_core.rtc_div\[3\]
rlabel metal2 37576 56896 37576 56896 0 u_rtc.u_core.rtc_div\[4\]
rlabel metal2 38360 58072 38360 58072 0 u_rtc.u_core.rtc_div\[5\]
rlabel metal2 37576 60144 37576 60144 0 u_rtc.u_core.rtc_div\[6\]
rlabel metal2 37576 62720 37576 62720 0 u_rtc.u_core.rtc_div\[7\]
rlabel metal3 37016 65464 37016 65464 0 u_rtc.u_core.rtc_div\[8\]
rlabel metal2 37688 67536 37688 67536 0 u_rtc.u_core.rtc_div\[9\]
rlabel metal2 2296 4984 2296 4984 0 u_rtc.u_reg._0000_
rlabel metal3 13272 32536 13272 32536 0 u_rtc.u_reg._0001_
rlabel metal2 13608 29120 13608 29120 0 u_rtc.u_reg._0002_
rlabel metal2 10024 29288 10024 29288 0 u_rtc.u_reg._0003_
rlabel metal2 26712 34776 26712 34776 0 u_rtc.u_reg._0009_
rlabel metal2 23576 35168 23576 35168 0 u_rtc.u_reg._0010_
rlabel metal2 26600 30688 26600 30688 0 u_rtc.u_reg._0011_
rlabel metal2 27608 29680 27608 29680 0 u_rtc.u_reg._0012_
rlabel metal3 22400 31864 22400 31864 0 u_rtc.u_reg._0013_
rlabel metal2 22736 27048 22736 27048 0 u_rtc.u_reg._0017_
rlabel metal2 19320 26544 19320 26544 0 u_rtc.u_reg._0018_
rlabel metal2 18872 23128 18872 23128 0 u_rtc.u_reg._0019_
rlabel metal2 21896 21280 21896 21280 0 u_rtc.u_reg._0020_
rlabel metal2 22848 11368 22848 11368 0 u_rtc.u_reg._0021_
rlabel metal2 20384 10584 20384 10584 0 u_rtc.u_reg._0022_
rlabel metal2 16968 13216 16968 13216 0 u_rtc.u_reg._0023_
rlabel metal2 15624 22064 15624 22064 0 u_rtc.u_reg._0024_
rlabel metal2 13888 11368 13888 11368 0 u_rtc.u_reg._0025_
rlabel metal3 13776 23688 13776 23688 0 u_rtc.u_reg._0026_
rlabel metal2 8344 24192 8344 24192 0 u_rtc.u_reg._0027_
rlabel metal2 5880 22064 5880 22064 0 u_rtc.u_reg._0028_
rlabel metal2 2296 11648 2296 11648 0 u_rtc.u_reg._0029_
rlabel metal2 2296 15568 2296 15568 0 u_rtc.u_reg._0030_
rlabel metal2 2408 11872 2408 11872 0 u_rtc.u_reg._0031_
rlabel metal2 2408 22176 2408 22176 0 u_rtc.u_reg._0032_
rlabel metal2 10136 52584 10136 52584 0 u_rtc.u_reg._0033_
rlabel metal2 8232 57008 8232 57008 0 u_rtc.u_reg._0034_
rlabel metal2 9576 57680 9576 57680 0 u_rtc.u_reg._0035_
rlabel metal2 8568 53872 8568 53872 0 u_rtc.u_reg._0036_
rlabel metal2 14056 44632 14056 44632 0 u_rtc.u_reg._0037_
rlabel metal2 11704 49448 11704 49448 0 u_rtc.u_reg._0038_
rlabel metal2 20328 51744 20328 51744 0 u_rtc.u_reg._0039_
rlabel metal2 20552 45248 20552 45248 0 u_rtc.u_reg._0040_
rlabel metal2 19096 37520 19096 37520 0 u_rtc.u_reg._0041_
rlabel metal2 17864 39312 17864 39312 0 u_rtc.u_reg._0042_
rlabel metal2 21560 56728 21560 56728 0 u_rtc.u_reg._0057_
rlabel metal2 25368 58072 25368 58072 0 u_rtc.u_reg._0058_
rlabel metal2 21672 57904 21672 57904 0 u_rtc.u_reg._0059_
rlabel metal2 18816 54488 18816 54488 0 u_rtc.u_reg._0060_
rlabel metal2 16744 42952 16744 42952 0 u_rtc.u_reg._0061_
rlabel metal3 12880 47544 12880 47544 0 u_rtc.u_reg._0062_
rlabel metal2 22456 52192 22456 52192 0 u_rtc.u_reg._0063_
rlabel metal3 21784 47544 21784 47544 0 u_rtc.u_reg._0064_
rlabel metal3 20272 35112 20272 35112 0 u_rtc.u_reg._0065_
rlabel metal3 16800 37464 16800 37464 0 u_rtc.u_reg._0066_
rlabel metal3 24976 68600 24976 68600 0 u_rtc.u_reg._0081_
rlabel metal2 24584 69496 24584 69496 0 u_rtc.u_reg._0082_
rlabel metal2 12824 35392 12824 35392 0 u_rtc.u_reg._0083_
rlabel metal2 26824 58520 26824 58520 0 u_rtc.u_reg._0084_
rlabel metal2 26376 61824 26376 61824 0 u_rtc.u_reg._0085_
rlabel metal3 25256 63224 25256 63224 0 u_rtc.u_reg._0087_
rlabel metal2 24248 46032 24248 46032 0 u_rtc.u_reg._0088_
rlabel metal2 2296 66136 2296 66136 0 u_rtc.u_reg._0090_
rlabel metal2 21448 66752 21448 66752 0 u_rtc.u_reg._0091_
rlabel metal2 21784 72632 21784 72632 0 u_rtc.u_reg._0092_
rlabel metal2 21504 61768 21504 61768 0 u_rtc.u_reg._0093_
rlabel metal2 2296 61040 2296 61040 0 u_rtc.u_reg._0094_
rlabel via1 2296 51358 2296 51358 0 u_rtc.u_reg._0095_
rlabel metal3 2800 56616 2800 56616 0 u_rtc.u_reg._0096_
rlabel metal2 3864 46368 3864 46368 0 u_rtc.u_reg._0098_
rlabel metal2 2296 43792 2296 43792 0 u_rtc.u_reg._0099_
rlabel metal2 2296 40096 2296 40096 0 u_rtc.u_reg._0100_
rlabel metal2 5096 38724 5096 38724 0 u_rtc.u_reg._0101_
rlabel metal2 2184 35392 2184 35392 0 u_rtc.u_reg._0102_
rlabel metal2 2296 34384 2296 34384 0 u_rtc.u_reg._0103_
rlabel metal2 10024 63224 10024 63224 0 u_rtc.u_reg._0107_
rlabel metal2 2408 63616 2408 63616 0 u_rtc.u_reg._0108_
rlabel metal2 10696 66752 10696 66752 0 u_rtc.u_reg._0109_
rlabel metal2 12152 61600 12152 61600 0 u_rtc.u_reg._0110_
rlabel metal2 12936 68880 12936 68880 0 u_rtc.u_reg._0111_
rlabel metal2 11704 69888 11704 69888 0 u_rtc.u_reg._0112_
rlabel metal2 7448 69552 7448 69552 0 u_rtc.u_reg._0113_
rlabel metal3 4088 66136 4088 66136 0 u_rtc.u_reg._0114_
rlabel metal2 10360 87920 10360 87920 0 u_rtc.u_reg._0115_
rlabel metal3 6888 86856 6888 86856 0 u_rtc.u_reg._0116_
rlabel metal3 4928 83720 4928 83720 0 u_rtc.u_reg._0117_
rlabel metal2 10024 87864 10024 87864 0 u_rtc.u_reg._0118_
rlabel metal3 7672 84504 7672 84504 0 u_rtc.u_reg._0119_
rlabel metal2 9912 78512 9912 78512 0 u_rtc.u_reg._0120_
rlabel metal2 7784 72968 7784 72968 0 u_rtc.u_reg._0121_
rlabel metal2 23352 78120 23352 78120 0 u_rtc.u_reg._0123_
rlabel metal2 16408 74144 16408 74144 0 u_rtc.u_reg._0124_
rlabel metal2 17360 75656 17360 75656 0 u_rtc.u_reg._0125_
rlabel metal2 22344 76944 22344 76944 0 u_rtc.u_reg._0126_
rlabel metal2 11648 75880 11648 75880 0 u_rtc.u_reg._0127_
rlabel metal2 12320 74312 12320 74312 0 u_rtc.u_reg._0128_
rlabel metal3 8792 73528 8792 73528 0 u_rtc.u_reg._0129_
rlabel metal2 25928 45528 25928 45528 0 u_rtc.u_reg._0131_
rlabel metal2 27664 48216 27664 48216 0 u_rtc.u_reg._0132_
rlabel metal2 27272 53200 27272 53200 0 u_rtc.u_reg._0133_
rlabel metal2 27496 53032 27496 53032 0 u_rtc.u_reg._0134_
rlabel metal2 22344 39872 22344 39872 0 u_rtc.u_reg._0135_
rlabel metal2 21448 42224 21448 42224 0 u_rtc.u_reg._0136_
rlabel metal2 21056 85848 21056 85848 0 u_rtc.u_reg._0139_
rlabel metal2 15400 86352 15400 86352 0 u_rtc.u_reg._0140_
rlabel metal2 12600 87696 12600 87696 0 u_rtc.u_reg._0141_
rlabel metal2 18424 87136 18424 87136 0 u_rtc.u_reg._0142_
rlabel metal2 2296 82992 2296 82992 0 u_rtc.u_reg._0143_
rlabel metal2 3304 77728 3304 77728 0 u_rtc.u_reg._0144_
rlabel metal2 2296 73640 2296 73640 0 u_rtc.u_reg._0145_
rlabel metal2 2296 29176 2296 29176 0 u_rtc.u_reg._0147_
rlabel metal2 4760 28336 4760 28336 0 u_rtc.u_reg._0148_
rlabel metal2 6664 26544 6664 26544 0 u_rtc.u_reg._0224_
rlabel metal2 6328 26264 6328 26264 0 u_rtc.u_reg._0225_
rlabel metal2 2800 6552 2800 6552 0 u_rtc.u_reg._0226_
rlabel metal2 17752 44688 17752 44688 0 u_rtc.u_reg._0227_
rlabel metal2 11480 82096 11480 82096 0 u_rtc.u_reg._0228_
rlabel metal2 12880 82936 12880 82936 0 u_rtc.u_reg._0229_
rlabel metal3 11088 86520 11088 86520 0 u_rtc.u_reg._0230_
rlabel metal2 9184 84504 9184 84504 0 u_rtc.u_reg._0231_
rlabel metal3 7280 81032 7280 81032 0 u_rtc.u_reg._0232_
rlabel metal3 10584 80472 10584 80472 0 u_rtc.u_reg._0233_
rlabel metal2 11480 79576 11480 79576 0 u_rtc.u_reg._0234_
rlabel metal3 20104 57624 20104 57624 0 u_rtc.u_reg._0235_
rlabel metal3 19768 65464 19768 65464 0 u_rtc.u_reg._0236_
rlabel metal2 20216 58352 20216 58352 0 u_rtc.u_reg._0237_
rlabel metal2 19936 58408 19936 58408 0 u_rtc.u_reg._0238_
rlabel metal3 19544 56280 19544 56280 0 u_rtc.u_reg._0239_
rlabel metal2 18648 57120 18648 57120 0 u_rtc.u_reg._0240_
rlabel metal2 18984 43456 18984 43456 0 u_rtc.u_reg._0241_
rlabel metal2 18424 39704 18424 39704 0 u_rtc.u_reg._0242_
rlabel metal2 18088 42840 18088 42840 0 u_rtc.u_reg._0243_
rlabel metal2 17808 68600 17808 68600 0 u_rtc.u_reg._0244_
rlabel metal2 15960 67480 15960 67480 0 u_rtc.u_reg._0245_
rlabel metal2 15512 44296 15512 44296 0 u_rtc.u_reg._0246_
rlabel metal2 13944 55720 13944 55720 0 u_rtc.u_reg._0247_
rlabel metal2 15344 77112 15344 77112 0 u_rtc.u_reg._0248_
rlabel metal2 17752 76608 17752 76608 0 u_rtc.u_reg._0249_
rlabel metal2 14616 77280 14616 77280 0 u_rtc.u_reg._0250_
rlabel metal2 11256 52304 11256 52304 0 u_rtc.u_reg._0251_
rlabel metal2 15400 56952 15400 56952 0 u_rtc.u_reg._0252_
rlabel metal3 17024 41384 17024 41384 0 u_rtc.u_reg._0253_
rlabel metal2 10248 62216 10248 62216 0 u_rtc.u_reg._0254_
rlabel metal2 15400 63280 15400 63280 0 u_rtc.u_reg._0255_
rlabel metal2 4088 23520 4088 23520 0 u_rtc.u_reg._0256_
rlabel metal3 8848 72520 8848 72520 0 u_rtc.u_reg._0259_
rlabel metal2 3864 65072 3864 65072 0 u_rtc.u_reg._0260_
rlabel metal3 8792 48776 8792 48776 0 u_rtc.u_reg._0261_
rlabel metal3 24360 63112 24360 63112 0 u_rtc.u_reg._0262_
rlabel metal3 20608 45640 20608 45640 0 u_rtc.u_reg._0263_
rlabel metal2 26488 68096 26488 68096 0 u_rtc.u_reg._0267_
rlabel metal2 26320 70168 26320 70168 0 u_rtc.u_reg._0268_
rlabel metal3 4928 21000 4928 21000 0 u_rtc.u_reg._0274_
rlabel metal2 2520 6104 2520 6104 0 u_rtc.u_reg._0289_
rlabel metal2 23016 48664 23016 48664 0 u_rtc.u_reg._0290_
rlabel metal2 22792 46256 22792 46256 0 u_rtc.u_reg._0291_
rlabel metal2 22792 40992 22792 40992 0 u_rtc.u_reg._0292_
rlabel metal2 18312 46368 18312 46368 0 u_rtc.u_reg._0293_
rlabel metal2 18088 45528 18088 45528 0 u_rtc.u_reg._0294_
rlabel metal2 16520 44464 16520 44464 0 u_rtc.u_reg._0295_
rlabel metal2 16688 55496 16688 55496 0 u_rtc.u_reg._0296_
rlabel metal2 15960 60872 15960 60872 0 u_rtc.u_reg._0297_
rlabel metal3 16968 45864 16968 45864 0 u_rtc.u_reg._0298_
rlabel metal2 17304 46536 17304 46536 0 u_rtc.u_reg._0299_
rlabel metal2 14840 64792 14840 64792 0 u_rtc.u_reg._0300_
rlabel metal2 15680 62104 15680 62104 0 u_rtc.u_reg._0301_
rlabel metal2 16184 51464 16184 51464 0 u_rtc.u_reg._0302_
rlabel metal2 15568 50904 15568 50904 0 u_rtc.u_reg._0303_
rlabel metal3 15064 63672 15064 63672 0 u_rtc.u_reg._0304_
rlabel metal2 15400 51688 15400 51688 0 u_rtc.u_reg._0305_
rlabel metal2 15288 50848 15288 50848 0 u_rtc.u_reg._0306_
rlabel metal2 15624 52640 15624 52640 0 u_rtc.u_reg._0307_
rlabel metal2 13496 53984 13496 53984 0 u_rtc.u_reg._0308_
rlabel metal2 13440 54488 13440 54488 0 u_rtc.u_reg._0309_
rlabel metal2 13104 53816 13104 53816 0 u_rtc.u_reg._0310_
rlabel metal2 12992 54488 12992 54488 0 u_rtc.u_reg._0311_
rlabel metal2 14672 53928 14672 53928 0 u_rtc.u_reg._0312_
rlabel metal2 15064 53872 15064 53872 0 u_rtc.u_reg._0313_
rlabel metal2 17304 63168 17304 63168 0 u_rtc.u_reg._0314_
rlabel metal2 16968 62720 16968 62720 0 u_rtc.u_reg._0315_
rlabel metal2 11984 79576 11984 79576 0 u_rtc.u_reg._0316_
rlabel metal2 12936 78792 12936 78792 0 u_rtc.u_reg._0317_
rlabel metal2 15288 76608 15288 76608 0 u_rtc.u_reg._0318_
rlabel metal2 23240 79072 23240 79072 0 u_rtc.u_reg._0319_
rlabel metal3 21896 78680 21896 78680 0 u_rtc.u_reg._0320_
rlabel metal3 19656 76552 19656 76552 0 u_rtc.u_reg._0321_
rlabel metal2 15400 78232 15400 78232 0 u_rtc.u_reg._0322_
rlabel metal2 15960 77672 15960 77672 0 u_rtc.u_reg._0323_
rlabel metal3 14280 75432 14280 75432 0 u_rtc.u_reg._0324_
rlabel metal2 15624 56000 15624 56000 0 u_rtc.u_reg._0325_
rlabel metal2 15288 57120 15288 57120 0 u_rtc.u_reg._0326_
rlabel metal2 16072 58520 16072 58520 0 u_rtc.u_reg._0327_
rlabel metal2 14056 55832 14056 55832 0 u_rtc.u_reg._0328_
rlabel metal2 12600 58520 12600 58520 0 u_rtc.u_reg._0329_
rlabel metal2 15288 58912 15288 58912 0 u_rtc.u_reg._0330_
rlabel metal2 14672 59192 14672 59192 0 u_rtc.u_reg._0331_
rlabel metal2 13832 61600 13832 61600 0 u_rtc.u_reg._0332_
rlabel metal2 15624 62664 15624 62664 0 u_rtc.u_reg._0333_
rlabel metal2 16072 64400 16072 64400 0 u_rtc.u_reg._0334_
rlabel metal2 14168 65184 14168 65184 0 u_rtc.u_reg._0335_
rlabel metal2 14952 63448 14952 63448 0 u_rtc.u_reg._0336_
rlabel metal2 15512 64008 15512 64008 0 u_rtc.u_reg._0337_
rlabel metal3 21504 64904 21504 64904 0 u_rtc.u_reg._0338_
rlabel metal2 23688 50120 23688 50120 0 u_rtc.u_reg._0339_
rlabel metal2 23576 49448 23576 49448 0 u_rtc.u_reg._0340_
rlabel metal2 24136 39368 24136 39368 0 u_rtc.u_reg._0341_
rlabel metal3 21672 50456 21672 50456 0 u_rtc.u_reg._0342_
rlabel metal2 18424 48888 18424 48888 0 u_rtc.u_reg._0343_
rlabel metal2 17640 44464 17640 44464 0 u_rtc.u_reg._0344_
rlabel metal3 18312 48888 18312 48888 0 u_rtc.u_reg._0345_
rlabel metal3 19488 49112 19488 49112 0 u_rtc.u_reg._0346_
rlabel metal2 19488 49224 19488 49224 0 u_rtc.u_reg._0347_
rlabel metal2 16968 68992 16968 68992 0 u_rtc.u_reg._0348_
rlabel metal3 19768 50680 19768 50680 0 u_rtc.u_reg._0349_
rlabel metal2 19096 49112 19096 49112 0 u_rtc.u_reg._0350_
rlabel metal2 16520 49448 16520 49448 0 u_rtc.u_reg._0351_
rlabel metal2 16184 67984 16184 67984 0 u_rtc.u_reg._0352_
rlabel metal2 17976 50092 17976 50092 0 u_rtc.u_reg._0353_
rlabel metal2 17976 51240 17976 51240 0 u_rtc.u_reg._0354_
rlabel metal2 18200 50288 18200 50288 0 u_rtc.u_reg._0355_
rlabel metal2 19152 57848 19152 57848 0 u_rtc.u_reg._0356_
rlabel metal2 16856 55496 16856 55496 0 u_rtc.u_reg._0357_
rlabel metal2 17640 56112 17640 56112 0 u_rtc.u_reg._0358_
rlabel metal2 17864 55776 17864 55776 0 u_rtc.u_reg._0359_
rlabel metal3 17472 55832 17472 55832 0 u_rtc.u_reg._0360_
rlabel metal4 18536 57456 18536 57456 0 u_rtc.u_reg._0361_
rlabel metal3 14952 67816 14952 67816 0 u_rtc.u_reg._0362_
rlabel metal2 18312 69216 18312 69216 0 u_rtc.u_reg._0363_
rlabel metal2 10976 81256 10976 81256 0 u_rtc.u_reg._0364_
rlabel metal2 9800 80808 9800 80808 0 u_rtc.u_reg._0365_
rlabel metal2 12376 81928 12376 81928 0 u_rtc.u_reg._0366_
rlabel metal2 11928 81648 11928 81648 0 u_rtc.u_reg._0367_
rlabel metal2 12152 82824 12152 82824 0 u_rtc.u_reg._0368_
rlabel metal2 10696 81200 10696 81200 0 u_rtc.u_reg._0369_
rlabel metal2 11704 80640 11704 80640 0 u_rtc.u_reg._0370_
rlabel metal2 12432 81144 12432 81144 0 u_rtc.u_reg._0371_
rlabel metal2 16408 69832 16408 69832 0 u_rtc.u_reg._0372_
rlabel metal2 18872 56952 18872 56952 0 u_rtc.u_reg._0373_
rlabel metal2 19320 58128 19320 58128 0 u_rtc.u_reg._0374_
rlabel metal2 18592 59304 18592 59304 0 u_rtc.u_reg._0375_
rlabel metal2 16856 52248 16856 52248 0 u_rtc.u_reg._0376_
rlabel metal2 20608 57848 20608 57848 0 u_rtc.u_reg._0377_
rlabel metal2 18088 57512 18088 57512 0 u_rtc.u_reg._0378_
rlabel metal2 19096 58968 19096 58968 0 u_rtc.u_reg._0379_
rlabel metal2 17248 62888 17248 62888 0 u_rtc.u_reg._0380_
rlabel metal3 17640 70168 17640 70168 0 u_rtc.u_reg._0381_
rlabel metal2 17528 69832 17528 69832 0 u_rtc.u_reg._0382_
rlabel metal2 15512 68152 15512 68152 0 u_rtc.u_reg._0383_
rlabel metal2 15400 67312 15400 67312 0 u_rtc.u_reg._0384_
rlabel metal2 17752 69552 17752 69552 0 u_rtc.u_reg._0385_
rlabel metal2 25592 68264 25592 68264 0 u_rtc.u_reg._0386_
rlabel metal3 4088 6776 4088 6776 0 u_rtc.u_reg._0387_
rlabel metal3 5600 27160 5600 27160 0 u_rtc.u_reg._0388_
rlabel metal2 6832 44632 6832 44632 0 u_rtc.u_reg._0389_
rlabel metal2 7616 30296 7616 30296 0 u_rtc.u_reg._0390_
rlabel metal2 9800 29680 9800 29680 0 u_rtc.u_reg._0391_
rlabel metal2 7392 46536 7392 46536 0 u_rtc.u_reg._0392_
rlabel metal2 7392 27272 7392 27272 0 u_rtc.u_reg._0393_
rlabel metal3 14392 28784 14392 28784 0 u_rtc.u_reg._0394_
rlabel metal2 14560 31976 14560 31976 0 u_rtc.u_reg._0395_
rlabel metal2 14728 28840 14728 28840 0 u_rtc.u_reg._0396_
rlabel metal2 12040 29064 12040 29064 0 u_rtc.u_reg._0397_
rlabel metal2 5544 25872 5544 25872 0 u_rtc.u_reg._0403_
rlabel metal2 5880 24584 5880 24584 0 u_rtc.u_reg._0404_
rlabel metal2 15400 35952 15400 35952 0 u_rtc.u_reg._0405_
rlabel metal2 13608 35448 13608 35448 0 u_rtc.u_reg._0406_
rlabel metal3 21168 35784 21168 35784 0 u_rtc.u_reg._0407_
rlabel metal2 27608 35952 27608 35952 0 u_rtc.u_reg._0408_
rlabel metal2 25648 35672 25648 35672 0 u_rtc.u_reg._0409_
rlabel metal2 26712 31360 26712 31360 0 u_rtc.u_reg._0410_
rlabel metal2 29624 30968 29624 30968 0 u_rtc.u_reg._0411_
rlabel metal2 23352 32144 23352 32144 0 u_rtc.u_reg._0412_
rlabel metal2 15176 25368 15176 25368 0 u_rtc.u_reg._0414_
rlabel metal2 16632 20832 16632 20832 0 u_rtc.u_reg._0415_
rlabel metal2 22680 29120 22680 29120 0 u_rtc.u_reg._0416_
rlabel metal2 19600 27272 19600 27272 0 u_rtc.u_reg._0417_
rlabel metal2 19656 24192 19656 24192 0 u_rtc.u_reg._0418_
rlabel metal3 21840 21000 21840 21000 0 u_rtc.u_reg._0419_
rlabel metal2 22680 14112 22680 14112 0 u_rtc.u_reg._0420_
rlabel metal2 21000 14000 21000 14000 0 u_rtc.u_reg._0421_
rlabel metal2 17752 17416 17752 17416 0 u_rtc.u_reg._0422_
rlabel metal2 15736 21560 15736 21560 0 u_rtc.u_reg._0423_
rlabel metal2 5208 23408 5208 23408 0 u_rtc.u_reg._0424_
rlabel metal2 6664 24360 6664 24360 0 u_rtc.u_reg._0425_
rlabel metal2 13944 15848 13944 15848 0 u_rtc.u_reg._0426_
rlabel metal2 13776 23576 13776 23576 0 u_rtc.u_reg._0427_
rlabel metal2 10024 24976 10024 24976 0 u_rtc.u_reg._0428_
rlabel metal2 6216 21616 6216 21616 0 u_rtc.u_reg._0429_
rlabel metal2 3528 13664 3528 13664 0 u_rtc.u_reg._0430_
rlabel metal2 3416 16520 3416 16520 0 u_rtc.u_reg._0431_
rlabel metal2 3808 11592 3808 11592 0 u_rtc.u_reg._0432_
rlabel metal3 8288 27608 8288 27608 0 u_rtc.u_reg._0433_
rlabel metal2 11480 45136 11480 45136 0 u_rtc.u_reg._0434_
rlabel metal2 20552 45976 20552 45976 0 u_rtc.u_reg._0435_
rlabel metal3 11648 52248 11648 52248 0 u_rtc.u_reg._0436_
rlabel metal3 12320 56952 12320 56952 0 u_rtc.u_reg._0437_
rlabel metal2 14504 45024 14504 45024 0 u_rtc.u_reg._0438_
rlabel metal2 12432 49000 12432 49000 0 u_rtc.u_reg._0439_
rlabel metal2 21056 52136 21056 52136 0 u_rtc.u_reg._0440_
rlabel metal2 22008 45976 22008 45976 0 u_rtc.u_reg._0441_
rlabel metal2 17976 38752 17976 38752 0 u_rtc.u_reg._0442_
rlabel metal3 17136 38808 17136 38808 0 u_rtc.u_reg._0443_
rlabel metal3 5096 27048 5096 27048 0 u_rtc.u_reg._0448_
rlabel metal2 8344 27832 8344 27832 0 u_rtc.u_reg._0449_
rlabel metal2 13720 45640 13720 45640 0 u_rtc.u_reg._0450_
rlabel metal2 15960 44912 15960 44912 0 u_rtc.u_reg._0451_
rlabel metal2 22680 55664 22680 55664 0 u_rtc.u_reg._0452_
rlabel metal2 22008 57120 22008 57120 0 u_rtc.u_reg._0453_
rlabel metal2 19320 54544 19320 54544 0 u_rtc.u_reg._0454_
rlabel metal2 17976 44968 17976 44968 0 u_rtc.u_reg._0455_
rlabel metal2 13944 47376 13944 47376 0 u_rtc.u_reg._0456_
rlabel metal2 23464 52976 23464 52976 0 u_rtc.u_reg._0457_
rlabel metal3 23128 47432 23128 47432 0 u_rtc.u_reg._0458_
rlabel metal3 18872 37240 18872 37240 0 u_rtc.u_reg._0459_
rlabel metal2 17528 37184 17528 37184 0 u_rtc.u_reg._0460_
rlabel metal3 7504 29512 7504 29512 0 u_rtc.u_reg._0465_
rlabel metal3 19544 35168 19544 35168 0 u_rtc.u_reg._0467_
rlabel metal2 26264 67256 26264 67256 0 u_rtc.u_reg._0468_
rlabel metal2 25592 67256 25592 67256 0 u_rtc.u_reg._0469_
rlabel metal2 25256 63000 25256 63000 0 u_rtc.u_reg._0471_
rlabel metal3 25536 45864 25536 45864 0 u_rtc.u_reg._0472_
rlabel metal2 6104 47096 6104 47096 0 u_rtc.u_reg._0476_
rlabel metal2 22008 65744 22008 65744 0 u_rtc.u_reg._0477_
rlabel metal2 3752 67312 3752 67312 0 u_rtc.u_reg._0478_
rlabel metal2 20664 67144 20664 67144 0 u_rtc.u_reg._0479_
rlabel metal2 21784 67032 21784 67032 0 u_rtc.u_reg._0480_
rlabel metal2 20440 58800 20440 58800 0 u_rtc.u_reg._0481_
rlabel metal3 21000 59416 21000 59416 0 u_rtc.u_reg._0482_
rlabel metal2 21336 59080 21336 59080 0 u_rtc.u_reg._0483_
rlabel metal2 20776 59976 20776 59976 0 u_rtc.u_reg._0484_
rlabel metal2 5656 61264 5656 61264 0 u_rtc.u_reg._0485_
rlabel metal2 3808 50568 3808 50568 0 u_rtc.u_reg._0486_
rlabel metal2 3864 55888 3864 55888 0 u_rtc.u_reg._0487_
rlabel metal3 5544 36344 5544 36344 0 u_rtc.u_reg._0488_
rlabel metal2 3080 35000 3080 35000 0 u_rtc.u_reg._0489_
rlabel metal3 4928 45192 4928 45192 0 u_rtc.u_reg._0490_
rlabel metal2 5768 43176 5768 43176 0 u_rtc.u_reg._0491_
rlabel metal2 3976 39816 3976 39816 0 u_rtc.u_reg._0492_
rlabel metal3 6608 39368 6608 39368 0 u_rtc.u_reg._0493_
rlabel metal2 2520 34160 2520 34160 0 u_rtc.u_reg._0494_
rlabel metal2 5656 34608 5656 34608 0 u_rtc.u_reg._0495_
rlabel metal2 9968 46872 9968 46872 0 u_rtc.u_reg._0499_
rlabel metal2 10472 62888 10472 62888 0 u_rtc.u_reg._0500_
rlabel metal2 11480 61600 11480 61600 0 u_rtc.u_reg._0501_
rlabel metal2 11816 69048 11816 69048 0 u_rtc.u_reg._0502_
rlabel metal3 8960 70168 8960 70168 0 u_rtc.u_reg._0503_
rlabel metal2 4984 66360 4984 66360 0 u_rtc.u_reg._0504_
rlabel metal3 9352 47656 9352 47656 0 u_rtc.u_reg._0505_
rlabel metal2 10360 86184 10360 86184 0 u_rtc.u_reg._0506_
rlabel metal2 8792 84000 8792 84000 0 u_rtc.u_reg._0507_
rlabel metal2 9576 77952 9576 77952 0 u_rtc.u_reg._0508_
rlabel metal3 8512 74648 8512 74648 0 u_rtc.u_reg._0509_
rlabel metal2 20664 79408 20664 79408 0 u_rtc.u_reg._0511_
rlabel metal2 16464 74760 16464 74760 0 u_rtc.u_reg._0512_
rlabel metal2 17864 75768 17864 75768 0 u_rtc.u_reg._0513_
rlabel metal2 12936 74592 12936 74592 0 u_rtc.u_reg._0514_
rlabel metal2 10248 74088 10248 74088 0 u_rtc.u_reg._0515_
rlabel metal3 13328 37352 13328 37352 0 u_rtc.u_reg._0517_
rlabel metal2 26152 45024 26152 45024 0 u_rtc.u_reg._0518_
rlabel metal2 21336 44352 21336 44352 0 u_rtc.u_reg._0519_
rlabel metal2 21784 44744 21784 44744 0 u_rtc.u_reg._0520_
rlabel metal3 27048 45080 27048 45080 0 u_rtc.u_reg._0521_
rlabel metal2 28056 49392 28056 49392 0 u_rtc.u_reg._0522_
rlabel metal2 26824 53816 26824 53816 0 u_rtc.u_reg._0523_
rlabel metal2 27832 51408 27832 51408 0 u_rtc.u_reg._0524_
rlabel metal2 23016 40656 23016 40656 0 u_rtc.u_reg._0525_
rlabel metal3 16912 43512 16912 43512 0 u_rtc.u_reg._0526_
rlabel metal2 21784 43176 21784 43176 0 u_rtc.u_reg._0527_
rlabel metal2 5264 47432 5264 47432 0 u_rtc.u_reg._0528_
rlabel metal2 15400 85792 15400 85792 0 u_rtc.u_reg._0529_
rlabel metal2 22008 84504 22008 84504 0 u_rtc.u_reg._0530_
rlabel metal2 13720 82880 13720 82880 0 u_rtc.u_reg._0531_
rlabel metal3 14784 85848 14784 85848 0 u_rtc.u_reg._0532_
rlabel metal2 16128 85960 16128 85960 0 u_rtc.u_reg._0533_
rlabel metal2 13384 84336 13384 84336 0 u_rtc.u_reg._0534_
rlabel metal2 12712 85008 12712 85008 0 u_rtc.u_reg._0535_
rlabel metal2 18760 85568 18760 85568 0 u_rtc.u_reg._0536_
rlabel metal2 4872 81984 4872 81984 0 u_rtc.u_reg._0537_
rlabel metal3 4088 82040 4088 82040 0 u_rtc.u_reg._0538_
rlabel metal2 3640 77616 3640 77616 0 u_rtc.u_reg._0539_
rlabel metal2 3864 73416 3864 73416 0 u_rtc.u_reg._0540_
rlabel metal2 3248 28616 3248 28616 0 u_rtc.u_reg._0541_
rlabel metal2 4200 27160 4200 27160 0 u_rtc.u_reg._0542_
rlabel metal2 3528 29064 3528 29064 0 u_rtc.u_reg._0543_
rlabel metal2 4200 28392 4200 28392 0 u_rtc.u_reg._0544_
rlabel metal2 22232 78512 22232 78512 0 u_rtc.u_reg.cfg_alarm1\[0\]
rlabel metal2 13496 56392 13496 56392 0 u_rtc.u_reg.cfg_alarm1\[10\]
rlabel metal3 13608 57624 13608 57624 0 u_rtc.u_reg.cfg_alarm1\[11\]
rlabel metal2 16744 45584 16744 45584 0 u_rtc.u_reg.cfg_alarm1\[12\]
rlabel metal2 14280 48944 14280 48944 0 u_rtc.u_reg.cfg_alarm1\[13\]
rlabel metal2 15176 50680 15176 50680 0 u_rtc.u_reg.cfg_alarm1\[14\]
rlabel metal2 23576 45640 23576 45640 0 u_rtc.u_reg.cfg_alarm1\[15\]
rlabel metal2 22120 37744 22120 37744 0 u_rtc.u_reg.cfg_alarm1\[16\]
rlabel metal2 17640 40824 17640 40824 0 u_rtc.u_reg.cfg_alarm1\[17\]
rlabel metal3 18984 74312 18984 74312 0 u_rtc.u_reg.cfg_alarm1\[1\]
rlabel metal2 20216 76160 20216 76160 0 u_rtc.u_reg.cfg_alarm1\[2\]
rlabel metal3 20608 77224 20608 77224 0 u_rtc.u_reg.cfg_alarm1\[3\]
rlabel metal2 15736 77728 15736 77728 0 u_rtc.u_reg.cfg_alarm1\[4\]
rlabel metal2 15288 73528 15288 73528 0 u_rtc.u_reg.cfg_alarm1\[5\]
rlabel metal2 10920 74872 10920 74872 0 u_rtc.u_reg.cfg_alarm1\[6\]
rlabel metal2 13160 53200 13160 53200 0 u_rtc.u_reg.cfg_alarm1\[8\]
rlabel metal2 13160 56560 13160 56560 0 u_rtc.u_reg.cfg_alarm1\[9\]
rlabel metal2 12824 87080 12824 87080 0 u_rtc.u_reg.cfg_alarm2\[0\]
rlabel metal2 20048 58296 20048 58296 0 u_rtc.u_reg.cfg_alarm2\[10\]
rlabel metal2 18872 55608 18872 55608 0 u_rtc.u_reg.cfg_alarm2\[11\]
rlabel metal2 18536 48272 18536 48272 0 u_rtc.u_reg.cfg_alarm2\[12\]
rlabel metal3 15624 49000 15624 49000 0 u_rtc.u_reg.cfg_alarm2\[13\]
rlabel metal2 18312 52528 18312 52528 0 u_rtc.u_reg.cfg_alarm2\[14\]
rlabel metal3 23688 48440 23688 48440 0 u_rtc.u_reg.cfg_alarm2\[15\]
rlabel metal3 23240 35896 23240 35896 0 u_rtc.u_reg.cfg_alarm2\[16\]
rlabel metal2 18144 40488 18144 40488 0 u_rtc.u_reg.cfg_alarm2\[17\]
rlabel metal2 9128 86912 9128 86912 0 u_rtc.u_reg.cfg_alarm2\[1\]
rlabel metal2 7336 83888 7336 83888 0 u_rtc.u_reg.cfg_alarm2\[2\]
rlabel metal2 12040 86800 12040 86800 0 u_rtc.u_reg.cfg_alarm2\[3\]
rlabel metal2 9800 84616 9800 84616 0 u_rtc.u_reg.cfg_alarm2\[4\]
rlabel metal2 11424 78792 11424 78792 0 u_rtc.u_reg.cfg_alarm2\[5\]
rlabel metal2 9128 73724 9128 73724 0 u_rtc.u_reg.cfg_alarm2\[6\]
rlabel metal2 22176 56616 22176 56616 0 u_rtc.u_reg.cfg_alarm2\[8\]
rlabel metal2 23688 57904 23688 57904 0 u_rtc.u_reg.cfg_alarm2\[9\]
rlabel metal3 28392 68824 28392 68824 0 u_rtc.u_reg.cfg_alrm1_ie
rlabel metal2 15624 61824 15624 61824 0 u_rtc.u_reg.cfg_alrm1_mode\[0\]
rlabel metal2 15400 61824 15400 61824 0 u_rtc.u_reg.cfg_alrm1_mode\[1\]
rlabel metal2 13160 66640 13160 66640 0 u_rtc.u_reg.cfg_alrm1_mode\[2\]
rlabel metal2 15960 62832 15960 62832 0 u_rtc.u_reg.cfg_alrm1_mode\[3\]
rlabel metal2 27608 69832 27608 69832 0 u_rtc.u_reg.cfg_alrm2_ie
rlabel metal2 16520 68992 16520 68992 0 u_rtc.u_reg.cfg_alrm2_mode\[0\]
rlabel metal2 15680 69272 15680 69272 0 u_rtc.u_reg.cfg_alrm2_mode\[1\]
rlabel metal2 16688 67032 16688 67032 0 u_rtc.u_reg.cfg_alrm2_mode\[2\]
rlabel metal2 16296 67536 16296 67536 0 u_rtc.u_reg.cfg_alrm2_mode\[3\]
rlabel metal2 28392 8260 28392 8260 0 u_rtc.u_sync_rclk.in_data_2s
rlabel metal2 25928 9016 25928 9016 0 u_rtc.u_sync_rclk.in_data_s
rlabel metal3 27944 6104 27944 6104 0 u_rtc.u_sync_sclk.in_data_2s
rlabel metal3 26712 6552 26712 6552 0 u_rtc.u_sync_sclk.in_data_s
<< properties >>
string FIXED_BBOX 0 0 40000 100000
<< end >>
