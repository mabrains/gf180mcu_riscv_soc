magic
tech gf180mcuD
magscale 1 5
timestamp 1699167808
<< obsm1 >>
rect 672 463 74872 75686
<< metal2 >>
rect 57120 76962 57176 77362
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 5376 0 5432 400
rect 5712 0 5768 400
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 50064 0 50120 400
rect 50400 0 50456 400
rect 50736 0 50792 400
rect 51072 0 51128 400
rect 51408 0 51464 400
rect 51744 0 51800 400
rect 52080 0 52136 400
rect 52416 0 52472 400
rect 52752 0 52808 400
rect 53088 0 53144 400
rect 53424 0 53480 400
rect 53760 0 53816 400
rect 54096 0 54152 400
rect 54432 0 54488 400
rect 54768 0 54824 400
rect 55104 0 55160 400
rect 55440 0 55496 400
rect 55776 0 55832 400
rect 56112 0 56168 400
rect 56448 0 56504 400
rect 56784 0 56840 400
rect 57120 0 57176 400
rect 57456 0 57512 400
rect 57792 0 57848 400
rect 58128 0 58184 400
rect 58464 0 58520 400
rect 58800 0 58856 400
rect 59136 0 59192 400
rect 59472 0 59528 400
rect 59808 0 59864 400
rect 60144 0 60200 400
rect 60480 0 60536 400
rect 60816 0 60872 400
rect 61152 0 61208 400
rect 61488 0 61544 400
rect 61824 0 61880 400
rect 62160 0 62216 400
rect 62496 0 62552 400
rect 62832 0 62888 400
rect 63168 0 63224 400
rect 63504 0 63560 400
rect 63840 0 63896 400
rect 64848 0 64904 400
rect 65184 0 65240 400
rect 65520 0 65576 400
rect 67200 0 67256 400
rect 67536 0 67592 400
rect 67872 0 67928 400
rect 68208 0 68264 400
rect 68544 0 68600 400
rect 68880 0 68936 400
rect 69216 0 69272 400
rect 69552 0 69608 400
rect 69888 0 69944 400
rect 70224 0 70280 400
rect 70560 0 70616 400
rect 70896 0 70952 400
rect 71232 0 71288 400
rect 71568 0 71624 400
rect 71904 0 71960 400
rect 72240 0 72296 400
rect 72576 0 72632 400
rect 72912 0 72968 400
rect 73248 0 73304 400
rect 73584 0 73640 400
rect 73920 0 73976 400
rect 74256 0 74312 400
rect 74592 0 74648 400
rect 74928 0 74984 400
rect 75264 0 75320 400
<< obsm2 >>
rect 854 76932 57090 76962
rect 57206 76932 75306 76962
rect 854 430 75306 76932
rect 854 9 978 430
rect 1094 9 1314 430
rect 1430 9 1650 430
rect 1766 9 1986 430
rect 2102 9 2322 430
rect 2438 9 2658 430
rect 2774 9 2994 430
rect 3110 9 3330 430
rect 3446 9 3666 430
rect 3782 9 4002 430
rect 4118 9 4338 430
rect 4454 9 4674 430
rect 4790 9 5010 430
rect 5126 9 5346 430
rect 5462 9 5682 430
rect 5798 9 6018 430
rect 6134 9 6354 430
rect 6470 9 6690 430
rect 6806 9 7026 430
rect 7142 9 7362 430
rect 7478 9 7698 430
rect 7814 9 8034 430
rect 8150 9 8370 430
rect 8486 9 8706 430
rect 8822 9 9042 430
rect 9158 9 9378 430
rect 9494 9 9714 430
rect 9830 9 10050 430
rect 10166 9 10386 430
rect 10502 9 10722 430
rect 10838 9 11058 430
rect 11174 9 11394 430
rect 11510 9 50034 430
rect 50150 9 50370 430
rect 50486 9 50706 430
rect 50822 9 51042 430
rect 51158 9 51378 430
rect 51494 9 51714 430
rect 51830 9 52050 430
rect 52166 9 52386 430
rect 52502 9 52722 430
rect 52838 9 53058 430
rect 53174 9 53394 430
rect 53510 9 53730 430
rect 53846 9 54066 430
rect 54182 9 54402 430
rect 54518 9 54738 430
rect 54854 9 55074 430
rect 55190 9 55410 430
rect 55526 9 55746 430
rect 55862 9 56082 430
rect 56198 9 56418 430
rect 56534 9 56754 430
rect 56870 9 57090 430
rect 57206 9 57426 430
rect 57542 9 57762 430
rect 57878 9 58098 430
rect 58214 9 58434 430
rect 58550 9 58770 430
rect 58886 9 59106 430
rect 59222 9 59442 430
rect 59558 9 59778 430
rect 59894 9 60114 430
rect 60230 9 60450 430
rect 60566 9 60786 430
rect 60902 9 61122 430
rect 61238 9 61458 430
rect 61574 9 61794 430
rect 61910 9 62130 430
rect 62246 9 62466 430
rect 62582 9 62802 430
rect 62918 9 63138 430
rect 63254 9 63474 430
rect 63590 9 63810 430
rect 63926 9 64818 430
rect 64934 9 65154 430
rect 65270 9 65490 430
rect 65606 9 67170 430
rect 67286 9 67506 430
rect 67622 9 67842 430
rect 67958 9 68178 430
rect 68294 9 68514 430
rect 68630 9 68850 430
rect 68966 9 69186 430
rect 69302 9 69522 430
rect 69638 9 69858 430
rect 69974 9 70194 430
rect 70310 9 70530 430
rect 70646 9 70866 430
rect 70982 9 71202 430
rect 71318 9 71538 430
rect 71654 9 71874 430
rect 71990 9 72210 430
rect 72326 9 72546 430
rect 72662 9 72882 430
rect 72998 9 73218 430
rect 73334 9 73554 430
rect 73670 9 73890 430
rect 74006 9 74226 430
rect 74342 9 74562 430
rect 74678 9 74898 430
rect 75014 9 75234 430
<< metal3 >>
rect 75170 55440 75570 55496
rect 75170 55104 75570 55160
rect 75170 54768 75570 54824
rect 75170 54432 75570 54488
rect 75170 54096 75570 54152
rect 75170 53760 75570 53816
rect 75170 53424 75570 53480
rect 75170 53088 75570 53144
rect 75170 52752 75570 52808
rect 75170 52416 75570 52472
rect 75170 52080 75570 52136
rect 75170 51744 75570 51800
rect 75170 51408 75570 51464
rect 75170 51072 75570 51128
rect 75170 50736 75570 50792
rect 75170 50400 75570 50456
rect 75170 50064 75570 50120
rect 75170 49728 75570 49784
rect 75170 49392 75570 49448
rect 75170 49056 75570 49112
rect 75170 48720 75570 48776
rect 75170 48384 75570 48440
rect 75170 48048 75570 48104
rect 75170 47712 75570 47768
rect 75170 47376 75570 47432
rect 75170 47040 75570 47096
rect 75170 46704 75570 46760
rect 75170 46368 75570 46424
rect 75170 46032 75570 46088
rect 75170 45696 75570 45752
rect 75170 45360 75570 45416
rect 75170 45024 75570 45080
rect 75170 44688 75570 44744
rect 75170 44352 75570 44408
rect 75170 44016 75570 44072
rect 75170 43680 75570 43736
rect 75170 43344 75570 43400
rect 75170 43008 75570 43064
rect 75170 42672 75570 42728
rect 75170 42336 75570 42392
rect 75170 42000 75570 42056
rect 75170 41664 75570 41720
rect 75170 41328 75570 41384
rect 75170 40992 75570 41048
rect 75170 40656 75570 40712
rect 75170 40320 75570 40376
rect 75170 39984 75570 40040
rect 75170 39648 75570 39704
rect 75170 39312 75570 39368
rect 75170 38976 75570 39032
rect 75170 38640 75570 38696
rect 75170 38304 75570 38360
rect 75170 37968 75570 38024
rect 75170 37632 75570 37688
rect 75170 37296 75570 37352
rect 75170 36960 75570 37016
rect 75170 36624 75570 36680
rect 75170 36288 75570 36344
rect 75170 35952 75570 36008
rect 75170 35616 75570 35672
rect 75170 35280 75570 35336
rect 75170 34944 75570 35000
rect 75170 34608 75570 34664
rect 75170 34272 75570 34328
rect 75170 33936 75570 33992
rect 75170 33600 75570 33656
rect 75170 33264 75570 33320
rect 75170 32928 75570 32984
rect 75170 32592 75570 32648
rect 75170 32256 75570 32312
rect 75170 31920 75570 31976
rect 75170 31584 75570 31640
rect 75170 31248 75570 31304
rect 75170 30912 75570 30968
rect 0 30576 400 30632
rect 75170 30576 75570 30632
rect 75170 30240 75570 30296
rect 75170 29904 75570 29960
rect 75170 29568 75570 29624
rect 75170 29232 75570 29288
rect 75170 28896 75570 28952
rect 75170 28560 75570 28616
rect 75170 28224 75570 28280
rect 75170 27888 75570 27944
rect 75170 27552 75570 27608
rect 75170 27216 75570 27272
rect 75170 26880 75570 26936
rect 75170 26544 75570 26600
rect 75170 26208 75570 26264
rect 75170 25872 75570 25928
rect 75170 25536 75570 25592
rect 75170 25200 75570 25256
rect 75170 24864 75570 24920
rect 75170 24528 75570 24584
rect 75170 24192 75570 24248
rect 75170 23856 75570 23912
rect 75170 23520 75570 23576
rect 75170 23184 75570 23240
rect 75170 22848 75570 22904
rect 75170 22512 75570 22568
rect 75170 22176 75570 22232
rect 75170 21840 75570 21896
rect 75170 21504 75570 21560
rect 75170 21168 75570 21224
rect 75170 20832 75570 20888
rect 75170 20496 75570 20552
rect 75170 20160 75570 20216
rect 75170 19824 75570 19880
rect 75170 19488 75570 19544
rect 75170 19152 75570 19208
rect 75170 18816 75570 18872
rect 75170 18480 75570 18536
rect 75170 18144 75570 18200
rect 75170 17808 75570 17864
rect 75170 17472 75570 17528
rect 75170 17136 75570 17192
rect 75170 16800 75570 16856
rect 75170 16464 75570 16520
rect 75170 16128 75570 16184
rect 75170 15792 75570 15848
rect 75170 15456 75570 15512
rect 75170 15120 75570 15176
rect 75170 14784 75570 14840
rect 75170 14448 75570 14504
rect 75170 14112 75570 14168
rect 75170 13776 75570 13832
rect 75170 13440 75570 13496
rect 75170 13104 75570 13160
rect 75170 12768 75570 12824
rect 75170 12432 75570 12488
rect 75170 12096 75570 12152
rect 75170 11760 75570 11816
rect 75170 11424 75570 11480
rect 75170 11088 75570 11144
rect 75170 10752 75570 10808
rect 75170 10416 75570 10472
rect 75170 10080 75570 10136
rect 75170 9744 75570 9800
rect 75170 9408 75570 9464
rect 75170 9072 75570 9128
rect 75170 8736 75570 8792
rect 75170 8400 75570 8456
rect 75170 8064 75570 8120
rect 75170 7728 75570 7784
rect 75170 7392 75570 7448
rect 75170 7056 75570 7112
rect 75170 6720 75570 6776
rect 75170 6384 75570 6440
rect 75170 6048 75570 6104
rect 75170 5712 75570 5768
rect 75170 5376 75570 5432
rect 75170 5040 75570 5096
rect 75170 4704 75570 4760
rect 75170 4368 75570 4424
rect 75170 4032 75570 4088
rect 75170 3696 75570 3752
rect 75170 3360 75570 3416
rect 75170 3024 75570 3080
rect 75170 2688 75570 2744
rect 75170 2352 75570 2408
rect 75170 2016 75570 2072
rect 75170 1680 75570 1736
rect 75170 1344 75570 1400
rect 75170 1008 75570 1064
rect 75170 672 75570 728
rect 75170 336 75570 392
rect 75170 0 75570 56
<< obsm3 >>
rect 400 55526 75311 75670
rect 400 55410 75140 55526
rect 400 55190 75311 55410
rect 400 55074 75140 55190
rect 400 54854 75311 55074
rect 400 54738 75140 54854
rect 400 54518 75311 54738
rect 400 54402 75140 54518
rect 400 54182 75311 54402
rect 400 54066 75140 54182
rect 400 53846 75311 54066
rect 400 53730 75140 53846
rect 400 53510 75311 53730
rect 400 53394 75140 53510
rect 400 53174 75311 53394
rect 400 53058 75140 53174
rect 400 52838 75311 53058
rect 400 52722 75140 52838
rect 400 52502 75311 52722
rect 400 52386 75140 52502
rect 400 52166 75311 52386
rect 400 52050 75140 52166
rect 400 51830 75311 52050
rect 400 51714 75140 51830
rect 400 51494 75311 51714
rect 400 51378 75140 51494
rect 400 51158 75311 51378
rect 400 51042 75140 51158
rect 400 50822 75311 51042
rect 400 50706 75140 50822
rect 400 50486 75311 50706
rect 400 50370 75140 50486
rect 400 50150 75311 50370
rect 400 50034 75140 50150
rect 400 49814 75311 50034
rect 400 49698 75140 49814
rect 400 49478 75311 49698
rect 400 49362 75140 49478
rect 400 49142 75311 49362
rect 400 49026 75140 49142
rect 400 48806 75311 49026
rect 400 48690 75140 48806
rect 400 48470 75311 48690
rect 400 48354 75140 48470
rect 400 48134 75311 48354
rect 400 48018 75140 48134
rect 400 47798 75311 48018
rect 400 47682 75140 47798
rect 400 47462 75311 47682
rect 400 47346 75140 47462
rect 400 47126 75311 47346
rect 400 47010 75140 47126
rect 400 46790 75311 47010
rect 400 46674 75140 46790
rect 400 46454 75311 46674
rect 400 46338 75140 46454
rect 400 46118 75311 46338
rect 400 46002 75140 46118
rect 400 45782 75311 46002
rect 400 45666 75140 45782
rect 400 45446 75311 45666
rect 400 45330 75140 45446
rect 400 45110 75311 45330
rect 400 44994 75140 45110
rect 400 44774 75311 44994
rect 400 44658 75140 44774
rect 400 44438 75311 44658
rect 400 44322 75140 44438
rect 400 44102 75311 44322
rect 400 43986 75140 44102
rect 400 43766 75311 43986
rect 400 43650 75140 43766
rect 400 43430 75311 43650
rect 400 43314 75140 43430
rect 400 43094 75311 43314
rect 400 42978 75140 43094
rect 400 42758 75311 42978
rect 400 42642 75140 42758
rect 400 42422 75311 42642
rect 400 42306 75140 42422
rect 400 42086 75311 42306
rect 400 41970 75140 42086
rect 400 41750 75311 41970
rect 400 41634 75140 41750
rect 400 41414 75311 41634
rect 400 41298 75140 41414
rect 400 41078 75311 41298
rect 400 40962 75140 41078
rect 400 40742 75311 40962
rect 400 40626 75140 40742
rect 400 40406 75311 40626
rect 400 40290 75140 40406
rect 400 40070 75311 40290
rect 400 39954 75140 40070
rect 400 39734 75311 39954
rect 400 39618 75140 39734
rect 400 39398 75311 39618
rect 400 39282 75140 39398
rect 400 39062 75311 39282
rect 400 38946 75140 39062
rect 400 38726 75311 38946
rect 400 38610 75140 38726
rect 400 38390 75311 38610
rect 400 38274 75140 38390
rect 400 38054 75311 38274
rect 400 37938 75140 38054
rect 400 37718 75311 37938
rect 400 37602 75140 37718
rect 400 37382 75311 37602
rect 400 37266 75140 37382
rect 400 37046 75311 37266
rect 400 36930 75140 37046
rect 400 36710 75311 36930
rect 400 36594 75140 36710
rect 400 36374 75311 36594
rect 400 36258 75140 36374
rect 400 36038 75311 36258
rect 400 35922 75140 36038
rect 400 35702 75311 35922
rect 400 35586 75140 35702
rect 400 35366 75311 35586
rect 400 35250 75140 35366
rect 400 35030 75311 35250
rect 400 34914 75140 35030
rect 400 34694 75311 34914
rect 400 34578 75140 34694
rect 400 34358 75311 34578
rect 400 34242 75140 34358
rect 400 34022 75311 34242
rect 400 33906 75140 34022
rect 400 33686 75311 33906
rect 400 33570 75140 33686
rect 400 33350 75311 33570
rect 400 33234 75140 33350
rect 400 33014 75311 33234
rect 400 32898 75140 33014
rect 400 32678 75311 32898
rect 400 32562 75140 32678
rect 400 32342 75311 32562
rect 400 32226 75140 32342
rect 400 32006 75311 32226
rect 400 31890 75140 32006
rect 400 31670 75311 31890
rect 400 31554 75140 31670
rect 400 31334 75311 31554
rect 400 31218 75140 31334
rect 400 30998 75311 31218
rect 400 30882 75140 30998
rect 400 30662 75311 30882
rect 430 30546 75140 30662
rect 400 30326 75311 30546
rect 400 30210 75140 30326
rect 400 29990 75311 30210
rect 400 29874 75140 29990
rect 400 29654 75311 29874
rect 400 29538 75140 29654
rect 400 29318 75311 29538
rect 400 29202 75140 29318
rect 400 28982 75311 29202
rect 400 28866 75140 28982
rect 400 28646 75311 28866
rect 400 28530 75140 28646
rect 400 28310 75311 28530
rect 400 28194 75140 28310
rect 400 27974 75311 28194
rect 400 27858 75140 27974
rect 400 27638 75311 27858
rect 400 27522 75140 27638
rect 400 27302 75311 27522
rect 400 27186 75140 27302
rect 400 26966 75311 27186
rect 400 26850 75140 26966
rect 400 26630 75311 26850
rect 400 26514 75140 26630
rect 400 26294 75311 26514
rect 400 26178 75140 26294
rect 400 25958 75311 26178
rect 400 25842 75140 25958
rect 400 25622 75311 25842
rect 400 25506 75140 25622
rect 400 25286 75311 25506
rect 400 25170 75140 25286
rect 400 24950 75311 25170
rect 400 24834 75140 24950
rect 400 24614 75311 24834
rect 400 24498 75140 24614
rect 400 24278 75311 24498
rect 400 24162 75140 24278
rect 400 23942 75311 24162
rect 400 23826 75140 23942
rect 400 23606 75311 23826
rect 400 23490 75140 23606
rect 400 23270 75311 23490
rect 400 23154 75140 23270
rect 400 22934 75311 23154
rect 400 22818 75140 22934
rect 400 22598 75311 22818
rect 400 22482 75140 22598
rect 400 22262 75311 22482
rect 400 22146 75140 22262
rect 400 21926 75311 22146
rect 400 21810 75140 21926
rect 400 21590 75311 21810
rect 400 21474 75140 21590
rect 400 21254 75311 21474
rect 400 21138 75140 21254
rect 400 20918 75311 21138
rect 400 20802 75140 20918
rect 400 20582 75311 20802
rect 400 20466 75140 20582
rect 400 20246 75311 20466
rect 400 20130 75140 20246
rect 400 19910 75311 20130
rect 400 19794 75140 19910
rect 400 19574 75311 19794
rect 400 19458 75140 19574
rect 400 19238 75311 19458
rect 400 19122 75140 19238
rect 400 18902 75311 19122
rect 400 18786 75140 18902
rect 400 18566 75311 18786
rect 400 18450 75140 18566
rect 400 18230 75311 18450
rect 400 18114 75140 18230
rect 400 17894 75311 18114
rect 400 17778 75140 17894
rect 400 17558 75311 17778
rect 400 17442 75140 17558
rect 400 17222 75311 17442
rect 400 17106 75140 17222
rect 400 16886 75311 17106
rect 400 16770 75140 16886
rect 400 16550 75311 16770
rect 400 16434 75140 16550
rect 400 16214 75311 16434
rect 400 16098 75140 16214
rect 400 15878 75311 16098
rect 400 15762 75140 15878
rect 400 15542 75311 15762
rect 400 15426 75140 15542
rect 400 15206 75311 15426
rect 400 15090 75140 15206
rect 400 14870 75311 15090
rect 400 14754 75140 14870
rect 400 14534 75311 14754
rect 400 14418 75140 14534
rect 400 14198 75311 14418
rect 400 14082 75140 14198
rect 400 13862 75311 14082
rect 400 13746 75140 13862
rect 400 13526 75311 13746
rect 400 13410 75140 13526
rect 400 13190 75311 13410
rect 400 13074 75140 13190
rect 400 12854 75311 13074
rect 400 12738 75140 12854
rect 400 12518 75311 12738
rect 400 12402 75140 12518
rect 400 12182 75311 12402
rect 400 12066 75140 12182
rect 400 11846 75311 12066
rect 400 11730 75140 11846
rect 400 11510 75311 11730
rect 400 11394 75140 11510
rect 400 11174 75311 11394
rect 400 11058 75140 11174
rect 400 10838 75311 11058
rect 400 10722 75140 10838
rect 400 10502 75311 10722
rect 400 10386 75140 10502
rect 400 10166 75311 10386
rect 400 10050 75140 10166
rect 400 9830 75311 10050
rect 400 9714 75140 9830
rect 400 9494 75311 9714
rect 400 9378 75140 9494
rect 400 9158 75311 9378
rect 400 9042 75140 9158
rect 400 8822 75311 9042
rect 400 8706 75140 8822
rect 400 8486 75311 8706
rect 400 8370 75140 8486
rect 400 8150 75311 8370
rect 400 8034 75140 8150
rect 400 7814 75311 8034
rect 400 7698 75140 7814
rect 400 7478 75311 7698
rect 400 7362 75140 7478
rect 400 7142 75311 7362
rect 400 7026 75140 7142
rect 400 6806 75311 7026
rect 400 6690 75140 6806
rect 400 6470 75311 6690
rect 400 6354 75140 6470
rect 400 6134 75311 6354
rect 400 6018 75140 6134
rect 400 5798 75311 6018
rect 400 5682 75140 5798
rect 400 5462 75311 5682
rect 400 5346 75140 5462
rect 400 5126 75311 5346
rect 400 5010 75140 5126
rect 400 4790 75311 5010
rect 400 4674 75140 4790
rect 400 4454 75311 4674
rect 400 4338 75140 4454
rect 400 4118 75311 4338
rect 400 4002 75140 4118
rect 400 3782 75311 4002
rect 400 3666 75140 3782
rect 400 3446 75311 3666
rect 400 3330 75140 3446
rect 400 3110 75311 3330
rect 400 2994 75140 3110
rect 400 2774 75311 2994
rect 400 2658 75140 2774
rect 400 2438 75311 2658
rect 400 2322 75140 2438
rect 400 2102 75311 2322
rect 400 1986 75140 2102
rect 400 1766 75311 1986
rect 400 1650 75140 1766
rect 400 1430 75311 1650
rect 400 1314 75140 1430
rect 400 1094 75311 1314
rect 400 978 75140 1094
rect 400 758 75311 978
rect 400 642 75140 758
rect 400 422 75311 642
rect 400 306 75140 422
rect 400 86 75311 306
rect 400 14 75140 86
<< metal4 >>
rect 2224 1538 2384 75686
rect 9904 1538 10064 75686
rect 17584 1538 17744 75686
rect 25264 1538 25424 75686
rect 32944 1538 33104 75686
rect 40624 1538 40784 75686
rect 48304 1538 48464 75686
rect 55984 1538 56144 75686
rect 63664 1538 63824 75686
rect 71344 1538 71504 75686
<< obsm4 >>
rect 5838 1689 9874 73463
rect 10094 1689 17554 73463
rect 17774 1689 25234 73463
rect 25454 1689 32914 73463
rect 33134 1689 40594 73463
rect 40814 1689 48274 73463
rect 48494 1689 55954 73463
rect 56174 1689 63634 73463
rect 63854 1689 71314 73463
rect 71534 1689 74522 73463
<< obsm5 >>
rect 8406 10823 74530 55507
<< labels >>
rlabel metal4 s 2224 1538 2384 75686 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 75686 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 75686 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 75686 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 75686 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 75686 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 75686 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 75686 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 75686 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 75686 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 75170 55440 75570 55496 6 clk
port 3 nsew signal input
rlabel metal3 s 75170 14784 75570 14840 6 i_dbus_ack
port 4 nsew signal input
rlabel metal3 s 75170 13104 75570 13160 6 i_dbus_rdt[0]
port 5 nsew signal input
rlabel metal3 s 75170 55104 75570 55160 6 i_dbus_rdt[10]
port 6 nsew signal input
rlabel metal3 s 75170 47376 75570 47432 6 i_dbus_rdt[11]
port 7 nsew signal input
rlabel metal3 s 75170 50400 75570 50456 6 i_dbus_rdt[12]
port 8 nsew signal input
rlabel metal3 s 75170 43680 75570 43736 6 i_dbus_rdt[13]
port 9 nsew signal input
rlabel metal3 s 75170 42672 75570 42728 6 i_dbus_rdt[14]
port 10 nsew signal input
rlabel metal3 s 75170 35280 75570 35336 6 i_dbus_rdt[15]
port 11 nsew signal input
rlabel metal3 s 75170 40320 75570 40376 6 i_dbus_rdt[16]
port 12 nsew signal input
rlabel metal3 s 75170 39648 75570 39704 6 i_dbus_rdt[17]
port 13 nsew signal input
rlabel metal3 s 75170 43008 75570 43064 6 i_dbus_rdt[18]
port 14 nsew signal input
rlabel metal3 s 75170 47712 75570 47768 6 i_dbus_rdt[19]
port 15 nsew signal input
rlabel metal3 s 75170 25872 75570 25928 6 i_dbus_rdt[1]
port 16 nsew signal input
rlabel metal3 s 75170 54768 75570 54824 6 i_dbus_rdt[20]
port 17 nsew signal input
rlabel metal3 s 75170 41664 75570 41720 6 i_dbus_rdt[21]
port 18 nsew signal input
rlabel metal3 s 75170 45360 75570 45416 6 i_dbus_rdt[22]
port 19 nsew signal input
rlabel metal3 s 75170 34272 75570 34328 6 i_dbus_rdt[23]
port 20 nsew signal input
rlabel metal3 s 75170 51072 75570 51128 6 i_dbus_rdt[24]
port 21 nsew signal input
rlabel metal3 s 75170 35616 75570 35672 6 i_dbus_rdt[25]
port 22 nsew signal input
rlabel metal3 s 75170 51408 75570 51464 6 i_dbus_rdt[26]
port 23 nsew signal input
rlabel metal3 s 75170 38304 75570 38360 6 i_dbus_rdt[27]
port 24 nsew signal input
rlabel metal3 s 75170 29568 75570 29624 6 i_dbus_rdt[28]
port 25 nsew signal input
rlabel metal3 s 75170 54432 75570 54488 6 i_dbus_rdt[29]
port 26 nsew signal input
rlabel metal3 s 75170 12096 75570 12152 6 i_dbus_rdt[2]
port 27 nsew signal input
rlabel metal3 s 75170 52416 75570 52472 6 i_dbus_rdt[30]
port 28 nsew signal input
rlabel metal3 s 75170 29232 75570 29288 6 i_dbus_rdt[31]
port 29 nsew signal input
rlabel metal3 s 75170 23856 75570 23912 6 i_dbus_rdt[3]
port 30 nsew signal input
rlabel metal3 s 75170 22848 75570 22904 6 i_dbus_rdt[4]
port 31 nsew signal input
rlabel metal3 s 75170 22512 75570 22568 6 i_dbus_rdt[5]
port 32 nsew signal input
rlabel metal3 s 75170 52080 75570 52136 6 i_dbus_rdt[6]
port 33 nsew signal input
rlabel metal3 s 75170 33600 75570 33656 6 i_dbus_rdt[7]
port 34 nsew signal input
rlabel metal3 s 75170 31248 75570 31304 6 i_dbus_rdt[8]
port 35 nsew signal input
rlabel metal3 s 75170 34608 75570 34664 6 i_dbus_rdt[9]
port 36 nsew signal input
rlabel metal2 s 0 0 56 400 6 i_ext_rd[0]
port 37 nsew signal input
rlabel metal2 s 336 0 392 400 6 i_ext_rd[10]
port 38 nsew signal input
rlabel metal2 s 672 0 728 400 6 i_ext_rd[11]
port 39 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 i_ext_rd[12]
port 40 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 i_ext_rd[13]
port 41 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 i_ext_rd[14]
port 42 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 i_ext_rd[15]
port 43 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 i_ext_rd[16]
port 44 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 i_ext_rd[17]
port 45 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 i_ext_rd[18]
port 46 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 i_ext_rd[19]
port 47 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 i_ext_rd[1]
port 48 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 i_ext_rd[20]
port 49 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 i_ext_rd[21]
port 50 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 i_ext_rd[22]
port 51 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 i_ext_rd[23]
port 52 nsew signal input
rlabel metal2 s 5376 0 5432 400 6 i_ext_rd[24]
port 53 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 i_ext_rd[25]
port 54 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 i_ext_rd[26]
port 55 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 i_ext_rd[27]
port 56 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 i_ext_rd[28]
port 57 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 i_ext_rd[29]
port 58 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 i_ext_rd[2]
port 59 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 i_ext_rd[30]
port 60 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 i_ext_rd[31]
port 61 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 i_ext_rd[3]
port 62 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 i_ext_rd[4]
port 63 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 i_ext_rd[5]
port 64 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 i_ext_rd[6]
port 65 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 i_ext_rd[7]
port 66 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 i_ext_rd[8]
port 67 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 i_ext_rd[9]
port 68 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 i_ext_ready
port 69 nsew signal input
rlabel metal3 s 75170 18144 75570 18200 6 i_ibus_ack
port 70 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 i_ibus_rdt[0]
port 71 nsew signal input
rlabel metal3 s 75170 20832 75570 20888 6 i_ibus_rdt[10]
port 72 nsew signal input
rlabel metal3 s 75170 19152 75570 19208 6 i_ibus_rdt[11]
port 73 nsew signal input
rlabel metal3 s 75170 27888 75570 27944 6 i_ibus_rdt[12]
port 74 nsew signal input
rlabel metal3 s 75170 26880 75570 26936 6 i_ibus_rdt[13]
port 75 nsew signal input
rlabel metal3 s 75170 26208 75570 26264 6 i_ibus_rdt[14]
port 76 nsew signal input
rlabel metal3 s 75170 28560 75570 28616 6 i_ibus_rdt[15]
port 77 nsew signal input
rlabel metal3 s 75170 32592 75570 32648 6 i_ibus_rdt[16]
port 78 nsew signal input
rlabel metal3 s 75170 25536 75570 25592 6 i_ibus_rdt[17]
port 79 nsew signal input
rlabel metal3 s 75170 12432 75570 12488 6 i_ibus_rdt[18]
port 80 nsew signal input
rlabel metal3 s 75170 13440 75570 13496 6 i_ibus_rdt[19]
port 81 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 i_ibus_rdt[1]
port 82 nsew signal input
rlabel metal2 s 68880 0 68936 400 6 i_ibus_rdt[20]
port 83 nsew signal input
rlabel metal3 s 75170 19488 75570 19544 6 i_ibus_rdt[21]
port 84 nsew signal input
rlabel metal2 s 74592 0 74648 400 6 i_ibus_rdt[22]
port 85 nsew signal input
rlabel metal3 s 75170 16128 75570 16184 6 i_ibus_rdt[23]
port 86 nsew signal input
rlabel metal3 s 75170 17136 75570 17192 6 i_ibus_rdt[24]
port 87 nsew signal input
rlabel metal2 s 74928 0 74984 400 6 i_ibus_rdt[25]
port 88 nsew signal input
rlabel metal2 s 67872 0 67928 400 6 i_ibus_rdt[26]
port 89 nsew signal input
rlabel metal2 s 72912 0 72968 400 6 i_ibus_rdt[27]
port 90 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 i_ibus_rdt[28]
port 91 nsew signal input
rlabel metal2 s 73920 0 73976 400 6 i_ibus_rdt[29]
port 92 nsew signal input
rlabel metal2 s 68544 0 68600 400 6 i_ibus_rdt[2]
port 93 nsew signal input
rlabel metal2 s 73248 0 73304 400 6 i_ibus_rdt[30]
port 94 nsew signal input
rlabel metal3 s 75170 16464 75570 16520 6 i_ibus_rdt[31]
port 95 nsew signal input
rlabel metal3 s 75170 28896 75570 28952 6 i_ibus_rdt[3]
port 96 nsew signal input
rlabel metal3 s 75170 21840 75570 21896 6 i_ibus_rdt[4]
port 97 nsew signal input
rlabel metal3 s 75170 18816 75570 18872 6 i_ibus_rdt[5]
port 98 nsew signal input
rlabel metal3 s 75170 23184 75570 23240 6 i_ibus_rdt[6]
port 99 nsew signal input
rlabel metal3 s 75170 20160 75570 20216 6 i_ibus_rdt[7]
port 100 nsew signal input
rlabel metal3 s 75170 19824 75570 19880 6 i_ibus_rdt[8]
port 101 nsew signal input
rlabel metal3 s 75170 21168 75570 21224 6 i_ibus_rdt[9]
port 102 nsew signal input
rlabel metal2 s 75264 0 75320 400 6 i_rst
port 103 nsew signal input
rlabel metal2 s 71232 0 71288 400 6 i_timer_irq
port 104 nsew signal input
rlabel metal3 s 0 30576 400 30632 6 o_dbus_adr[0]
port 105 nsew signal output
rlabel metal2 s 72240 0 72296 400 6 o_dbus_adr[10]
port 106 nsew signal output
rlabel metal2 s 69888 0 69944 400 6 o_dbus_adr[11]
port 107 nsew signal output
rlabel metal2 s 71904 0 71960 400 6 o_dbus_adr[12]
port 108 nsew signal output
rlabel metal2 s 69552 0 69608 400 6 o_dbus_adr[13]
port 109 nsew signal output
rlabel metal2 s 70896 0 70952 400 6 o_dbus_adr[14]
port 110 nsew signal output
rlabel metal2 s 70560 0 70616 400 6 o_dbus_adr[15]
port 111 nsew signal output
rlabel metal2 s 69216 0 69272 400 6 o_dbus_adr[16]
port 112 nsew signal output
rlabel metal2 s 71568 0 71624 400 6 o_dbus_adr[17]
port 113 nsew signal output
rlabel metal2 s 72576 0 72632 400 6 o_dbus_adr[18]
port 114 nsew signal output
rlabel metal2 s 70224 0 70280 400 6 o_dbus_adr[19]
port 115 nsew signal output
rlabel metal3 s 75170 44688 75570 44744 6 o_dbus_adr[1]
port 116 nsew signal output
rlabel metal2 s 68208 0 68264 400 6 o_dbus_adr[20]
port 117 nsew signal output
rlabel metal2 s 74256 0 74312 400 6 o_dbus_adr[21]
port 118 nsew signal output
rlabel metal2 s 52416 0 52472 400 6 o_dbus_adr[22]
port 119 nsew signal output
rlabel metal2 s 50064 0 50120 400 6 o_dbus_adr[23]
port 120 nsew signal output
rlabel metal2 s 50400 0 50456 400 6 o_dbus_adr[24]
port 121 nsew signal output
rlabel metal2 s 51744 0 51800 400 6 o_dbus_adr[25]
port 122 nsew signal output
rlabel metal2 s 67200 0 67256 400 6 o_dbus_adr[26]
port 123 nsew signal output
rlabel metal2 s 67536 0 67592 400 6 o_dbus_adr[27]
port 124 nsew signal output
rlabel metal2 s 55104 0 55160 400 6 o_dbus_adr[28]
port 125 nsew signal output
rlabel metal2 s 56784 0 56840 400 6 o_dbus_adr[29]
port 126 nsew signal output
rlabel metal3 s 75170 0 75570 56 6 o_dbus_adr[2]
port 127 nsew signal output
rlabel metal2 s 57456 0 57512 400 6 o_dbus_adr[30]
port 128 nsew signal output
rlabel metal2 s 58800 0 58856 400 6 o_dbus_adr[31]
port 129 nsew signal output
rlabel metal3 s 75170 1344 75570 1400 6 o_dbus_adr[3]
port 130 nsew signal output
rlabel metal2 s 61824 0 61880 400 6 o_dbus_adr[4]
port 131 nsew signal output
rlabel metal2 s 59808 0 59864 400 6 o_dbus_adr[5]
port 132 nsew signal output
rlabel metal2 s 61152 0 61208 400 6 o_dbus_adr[6]
port 133 nsew signal output
rlabel metal2 s 63840 0 63896 400 6 o_dbus_adr[7]
port 134 nsew signal output
rlabel metal2 s 63504 0 63560 400 6 o_dbus_adr[8]
port 135 nsew signal output
rlabel metal2 s 62160 0 62216 400 6 o_dbus_adr[9]
port 136 nsew signal output
rlabel metal3 s 75170 20496 75570 20552 6 o_dbus_cyc
port 137 nsew signal output
rlabel metal3 s 75170 13776 75570 13832 6 o_dbus_dat[0]
port 138 nsew signal output
rlabel metal3 s 75170 48048 75570 48104 6 o_dbus_dat[10]
port 139 nsew signal output
rlabel metal3 s 75170 32256 75570 32312 6 o_dbus_dat[11]
port 140 nsew signal output
rlabel metal3 s 75170 39312 75570 39368 6 o_dbus_dat[12]
port 141 nsew signal output
rlabel metal3 s 75170 35952 75570 36008 6 o_dbus_dat[13]
port 142 nsew signal output
rlabel metal3 s 75170 40992 75570 41048 6 o_dbus_dat[14]
port 143 nsew signal output
rlabel metal3 s 75170 47040 75570 47096 6 o_dbus_dat[15]
port 144 nsew signal output
rlabel metal3 s 75170 48720 75570 48776 6 o_dbus_dat[16]
port 145 nsew signal output
rlabel metal3 s 75170 38640 75570 38696 6 o_dbus_dat[17]
port 146 nsew signal output
rlabel metal3 s 75170 46704 75570 46760 6 o_dbus_dat[18]
port 147 nsew signal output
rlabel metal3 s 75170 42000 75570 42056 6 o_dbus_dat[19]
port 148 nsew signal output
rlabel metal3 s 75170 27552 75570 27608 6 o_dbus_dat[1]
port 149 nsew signal output
rlabel metal3 s 75170 36960 75570 37016 6 o_dbus_dat[20]
port 150 nsew signal output
rlabel metal3 s 75170 37968 75570 38024 6 o_dbus_dat[21]
port 151 nsew signal output
rlabel metal3 s 75170 34944 75570 35000 6 o_dbus_dat[22]
port 152 nsew signal output
rlabel metal3 s 75170 36288 75570 36344 6 o_dbus_dat[23]
port 153 nsew signal output
rlabel metal3 s 75170 43344 75570 43400 6 o_dbus_dat[24]
port 154 nsew signal output
rlabel metal3 s 75170 37632 75570 37688 6 o_dbus_dat[25]
port 155 nsew signal output
rlabel metal3 s 75170 38976 75570 39032 6 o_dbus_dat[26]
port 156 nsew signal output
rlabel metal3 s 75170 32928 75570 32984 6 o_dbus_dat[27]
port 157 nsew signal output
rlabel metal3 s 75170 53760 75570 53816 6 o_dbus_dat[28]
port 158 nsew signal output
rlabel metal3 s 75170 41328 75570 41384 6 o_dbus_dat[29]
port 159 nsew signal output
rlabel metal3 s 75170 14448 75570 14504 6 o_dbus_dat[2]
port 160 nsew signal output
rlabel metal3 s 75170 31584 75570 31640 6 o_dbus_dat[30]
port 161 nsew signal output
rlabel metal3 s 75170 30240 75570 30296 6 o_dbus_dat[31]
port 162 nsew signal output
rlabel metal3 s 75170 23520 75570 23576 6 o_dbus_dat[3]
port 163 nsew signal output
rlabel metal3 s 75170 17472 75570 17528 6 o_dbus_dat[4]
port 164 nsew signal output
rlabel metal3 s 75170 21504 75570 21560 6 o_dbus_dat[5]
port 165 nsew signal output
rlabel metal3 s 75170 22176 75570 22232 6 o_dbus_dat[6]
port 166 nsew signal output
rlabel metal3 s 75170 31920 75570 31976 6 o_dbus_dat[7]
port 167 nsew signal output
rlabel metal3 s 75170 50736 75570 50792 6 o_dbus_dat[8]
port 168 nsew signal output
rlabel metal3 s 75170 33264 75570 33320 6 o_dbus_dat[9]
port 169 nsew signal output
rlabel metal3 s 75170 14112 75570 14168 6 o_dbus_sel[0]
port 170 nsew signal output
rlabel metal3 s 75170 24528 75570 24584 6 o_dbus_sel[1]
port 171 nsew signal output
rlabel metal3 s 75170 15792 75570 15848 6 o_dbus_sel[2]
port 172 nsew signal output
rlabel metal3 s 75170 15456 75570 15512 6 o_dbus_sel[3]
port 173 nsew signal output
rlabel metal3 s 75170 18480 75570 18536 6 o_dbus_we
port 174 nsew signal output
rlabel metal3 s 75170 25200 75570 25256 6 o_ext_funct3[0]
port 175 nsew signal output
rlabel metal3 s 75170 24192 75570 24248 6 o_ext_funct3[1]
port 176 nsew signal output
rlabel metal3 s 75170 24864 75570 24920 6 o_ext_funct3[2]
port 177 nsew signal output
rlabel metal3 s 75170 11424 75570 11480 6 o_ext_rs1[0]
port 178 nsew signal output
rlabel metal2 s 60480 0 60536 400 6 o_ext_rs1[10]
port 179 nsew signal output
rlabel metal2 s 59136 0 59192 400 6 o_ext_rs1[11]
port 180 nsew signal output
rlabel metal2 s 57792 0 57848 400 6 o_ext_rs1[12]
port 181 nsew signal output
rlabel metal2 s 58464 0 58520 400 6 o_ext_rs1[13]
port 182 nsew signal output
rlabel metal2 s 57120 0 57176 400 6 o_ext_rs1[14]
port 183 nsew signal output
rlabel metal2 s 56112 0 56168 400 6 o_ext_rs1[15]
port 184 nsew signal output
rlabel metal2 s 55440 0 55496 400 6 o_ext_rs1[16]
port 185 nsew signal output
rlabel metal2 s 54432 0 54488 400 6 o_ext_rs1[17]
port 186 nsew signal output
rlabel metal2 s 52752 0 52808 400 6 o_ext_rs1[18]
port 187 nsew signal output
rlabel metal2 s 53424 0 53480 400 6 o_ext_rs1[19]
port 188 nsew signal output
rlabel metal3 s 75170 11088 75570 11144 6 o_ext_rs1[1]
port 189 nsew signal output
rlabel metal2 s 54096 0 54152 400 6 o_ext_rs1[20]
port 190 nsew signal output
rlabel metal2 s 53760 0 53816 400 6 o_ext_rs1[21]
port 191 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 o_ext_rs1[22]
port 192 nsew signal output
rlabel metal2 s 51072 0 51128 400 6 o_ext_rs1[23]
port 193 nsew signal output
rlabel metal2 s 50736 0 50792 400 6 o_ext_rs1[24]
port 194 nsew signal output
rlabel metal2 s 51408 0 51464 400 6 o_ext_rs1[25]
port 195 nsew signal output
rlabel metal2 s 53088 0 53144 400 6 o_ext_rs1[26]
port 196 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 o_ext_rs1[27]
port 197 nsew signal output
rlabel metal2 s 55776 0 55832 400 6 o_ext_rs1[28]
port 198 nsew signal output
rlabel metal2 s 56448 0 56504 400 6 o_ext_rs1[29]
port 199 nsew signal output
rlabel metal3 s 75170 672 75570 728 6 o_ext_rs1[2]
port 200 nsew signal output
rlabel metal2 s 58128 0 58184 400 6 o_ext_rs1[30]
port 201 nsew signal output
rlabel metal2 s 59472 0 59528 400 6 o_ext_rs1[31]
port 202 nsew signal output
rlabel metal3 s 75170 8064 75570 8120 6 o_ext_rs1[3]
port 203 nsew signal output
rlabel metal2 s 61488 0 61544 400 6 o_ext_rs1[4]
port 204 nsew signal output
rlabel metal2 s 60144 0 60200 400 6 o_ext_rs1[5]
port 205 nsew signal output
rlabel metal2 s 60816 0 60872 400 6 o_ext_rs1[6]
port 206 nsew signal output
rlabel metal2 s 62832 0 62888 400 6 o_ext_rs1[7]
port 207 nsew signal output
rlabel metal2 s 63168 0 63224 400 6 o_ext_rs1[8]
port 208 nsew signal output
rlabel metal2 s 62496 0 62552 400 6 o_ext_rs1[9]
port 209 nsew signal output
rlabel metal3 s 75170 12768 75570 12824 6 o_ext_rs2[0]
port 210 nsew signal output
rlabel metal3 s 75170 33936 75570 33992 6 o_ext_rs2[10]
port 211 nsew signal output
rlabel metal3 s 75170 50064 75570 50120 6 o_ext_rs2[11]
port 212 nsew signal output
rlabel metal3 s 75170 40656 75570 40712 6 o_ext_rs2[12]
port 213 nsew signal output
rlabel metal3 s 75170 36624 75570 36680 6 o_ext_rs2[13]
port 214 nsew signal output
rlabel metal3 s 75170 45024 75570 45080 6 o_ext_rs2[14]
port 215 nsew signal output
rlabel metal3 s 75170 45696 75570 45752 6 o_ext_rs2[15]
port 216 nsew signal output
rlabel metal3 s 75170 26544 75570 26600 6 o_ext_rs2[16]
port 217 nsew signal output
rlabel metal3 s 75170 46368 75570 46424 6 o_ext_rs2[17]
port 218 nsew signal output
rlabel metal3 s 75170 49392 75570 49448 6 o_ext_rs2[18]
port 219 nsew signal output
rlabel metal3 s 75170 42336 75570 42392 6 o_ext_rs2[19]
port 220 nsew signal output
rlabel metal3 s 75170 27216 75570 27272 6 o_ext_rs2[1]
port 221 nsew signal output
rlabel metal3 s 75170 39984 75570 40040 6 o_ext_rs2[20]
port 222 nsew signal output
rlabel metal3 s 75170 51744 75570 51800 6 o_ext_rs2[21]
port 223 nsew signal output
rlabel metal3 s 75170 44016 75570 44072 6 o_ext_rs2[22]
port 224 nsew signal output
rlabel metal3 s 75170 44352 75570 44408 6 o_ext_rs2[23]
port 225 nsew signal output
rlabel metal3 s 75170 49056 75570 49112 6 o_ext_rs2[24]
port 226 nsew signal output
rlabel metal3 s 75170 46032 75570 46088 6 o_ext_rs2[25]
port 227 nsew signal output
rlabel metal3 s 75170 53088 75570 53144 6 o_ext_rs2[26]
port 228 nsew signal output
rlabel metal3 s 75170 54096 75570 54152 6 o_ext_rs2[27]
port 229 nsew signal output
rlabel metal3 s 75170 52752 75570 52808 6 o_ext_rs2[28]
port 230 nsew signal output
rlabel metal3 s 75170 28224 75570 28280 6 o_ext_rs2[29]
port 231 nsew signal output
rlabel metal3 s 75170 49728 75570 49784 6 o_ext_rs2[2]
port 232 nsew signal output
rlabel metal3 s 75170 37296 75570 37352 6 o_ext_rs2[30]
port 233 nsew signal output
rlabel metal3 s 75170 53424 75570 53480 6 o_ext_rs2[31]
port 234 nsew signal output
rlabel metal3 s 75170 15120 75570 15176 6 o_ext_rs2[3]
port 235 nsew signal output
rlabel metal3 s 75170 16800 75570 16856 6 o_ext_rs2[4]
port 236 nsew signal output
rlabel metal3 s 75170 17808 75570 17864 6 o_ext_rs2[5]
port 237 nsew signal output
rlabel metal3 s 75170 30576 75570 30632 6 o_ext_rs2[6]
port 238 nsew signal output
rlabel metal3 s 75170 48384 75570 48440 6 o_ext_rs2[7]
port 239 nsew signal output
rlabel metal3 s 75170 29904 75570 29960 6 o_ext_rs2[8]
port 240 nsew signal output
rlabel metal3 s 75170 30912 75570 30968 6 o_ext_rs2[9]
port 241 nsew signal output
rlabel metal3 s 75170 9408 75570 9464 6 o_ibus_adr[0]
port 242 nsew signal output
rlabel metal3 s 75170 2352 75570 2408 6 o_ibus_adr[10]
port 243 nsew signal output
rlabel metal3 s 75170 2688 75570 2744 6 o_ibus_adr[11]
port 244 nsew signal output
rlabel metal3 s 75170 3024 75570 3080 6 o_ibus_adr[12]
port 245 nsew signal output
rlabel metal3 s 75170 3360 75570 3416 6 o_ibus_adr[13]
port 246 nsew signal output
rlabel metal3 s 75170 3696 75570 3752 6 o_ibus_adr[14]
port 247 nsew signal output
rlabel metal3 s 75170 4032 75570 4088 6 o_ibus_adr[15]
port 248 nsew signal output
rlabel metal3 s 75170 4704 75570 4760 6 o_ibus_adr[16]
port 249 nsew signal output
rlabel metal3 s 75170 5376 75570 5432 6 o_ibus_adr[17]
port 250 nsew signal output
rlabel metal3 s 75170 6384 75570 6440 6 o_ibus_adr[18]
port 251 nsew signal output
rlabel metal3 s 75170 7392 75570 7448 6 o_ibus_adr[19]
port 252 nsew signal output
rlabel metal3 s 75170 7728 75570 7784 6 o_ibus_adr[1]
port 253 nsew signal output
rlabel metal3 s 75170 2016 75570 2072 6 o_ibus_adr[20]
port 254 nsew signal output
rlabel metal3 s 75170 7056 75570 7112 6 o_ibus_adr[21]
port 255 nsew signal output
rlabel metal3 s 75170 1680 75570 1736 6 o_ibus_adr[22]
port 256 nsew signal output
rlabel metal3 s 75170 8400 75570 8456 6 o_ibus_adr[23]
port 257 nsew signal output
rlabel metal3 s 75170 9744 75570 9800 6 o_ibus_adr[24]
port 258 nsew signal output
rlabel metal3 s 75170 336 75570 392 6 o_ibus_adr[25]
port 259 nsew signal output
rlabel metal3 s 75170 10752 75570 10808 6 o_ibus_adr[26]
port 260 nsew signal output
rlabel metal3 s 75170 10416 75570 10472 6 o_ibus_adr[27]
port 261 nsew signal output
rlabel metal3 s 75170 10080 75570 10136 6 o_ibus_adr[28]
port 262 nsew signal output
rlabel metal3 s 75170 1008 75570 1064 6 o_ibus_adr[29]
port 263 nsew signal output
rlabel metal3 s 75170 6720 75570 6776 6 o_ibus_adr[2]
port 264 nsew signal output
rlabel metal3 s 75170 9072 75570 9128 6 o_ibus_adr[30]
port 265 nsew signal output
rlabel metal3 s 75170 8736 75570 8792 6 o_ibus_adr[31]
port 266 nsew signal output
rlabel metal3 s 75170 5712 75570 5768 6 o_ibus_adr[3]
port 267 nsew signal output
rlabel metal2 s 64848 0 64904 400 6 o_ibus_adr[4]
port 268 nsew signal output
rlabel metal2 s 65184 0 65240 400 6 o_ibus_adr[5]
port 269 nsew signal output
rlabel metal2 s 65520 0 65576 400 6 o_ibus_adr[6]
port 270 nsew signal output
rlabel metal3 s 75170 4368 75570 4424 6 o_ibus_adr[7]
port 271 nsew signal output
rlabel metal3 s 75170 5040 75570 5096 6 o_ibus_adr[8]
port 272 nsew signal output
rlabel metal3 s 75170 6048 75570 6104 6 o_ibus_adr[9]
port 273 nsew signal output
rlabel metal3 s 75170 11760 75570 11816 6 o_ibus_cyc
port 274 nsew signal output
rlabel metal2 s 57120 76962 57176 77362 6 o_mdu_valid
port 275 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 75570 77362
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15383850
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/serv_rf_top/runs/23_11_05_08_52/results/signoff/serv_rf_top.magic.gds
string GDS_START 468030
<< end >>

