VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_buttons_leds
  CLASS BLOCK ;
  FOREIGN wb_buttons_leds ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 100.000 ;
  PIN buttons[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 12.320 120.000 12.880 ;
    END
  END buttons[0]
  PIN buttons[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 61.600 120.000 62.160 ;
    END
  END buttons[1]
  PIN buttons_enb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 86.240 120.000 86.800 ;
    END
  END buttons_enb[0]
  PIN buttons_enb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 36.960 120.000 37.520 ;
    END
  END buttons_enb[1]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END clk
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END clk2
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 0.000 22.960 4.000 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 4.000 ;
    END
  END i_wb_addr[10]
  PIN i_wb_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END i_wb_addr[11]
  PIN i_wb_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END i_wb_addr[12]
  PIN i_wb_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END i_wb_addr[13]
  PIN i_wb_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END i_wb_addr[14]
  PIN i_wb_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END i_wb_addr[15]
  PIN i_wb_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.280 4.000 ;
    END
  END i_wb_addr[16]
  PIN i_wb_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 4.000 ;
    END
  END i_wb_addr[17]
  PIN i_wb_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END i_wb_addr[18]
  PIN i_wb_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END i_wb_addr[19]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END i_wb_addr[1]
  PIN i_wb_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 4.000 ;
    END
  END i_wb_addr[20]
  PIN i_wb_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END i_wb_addr[21]
  PIN i_wb_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 4.000 ;
    END
  END i_wb_addr[22]
  PIN i_wb_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END i_wb_addr[23]
  PIN i_wb_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END i_wb_addr[24]
  PIN i_wb_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END i_wb_addr[25]
  PIN i_wb_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 4.000 ;
    END
  END i_wb_addr[26]
  PIN i_wb_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END i_wb_addr[27]
  PIN i_wb_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 4.000 ;
    END
  END i_wb_addr[28]
  PIN i_wb_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 4.000 ;
    END
  END i_wb_addr[29]
  PIN i_wb_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 0.000 31.920 4.000 ;
    END
  END i_wb_addr[2]
  PIN i_wb_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END i_wb_addr[30]
  PIN i_wb_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END i_wb_addr[31]
  PIN i_wb_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END i_wb_addr[3]
  PIN i_wb_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 0.000 36.400 4.000 ;
    END
  END i_wb_addr[4]
  PIN i_wb_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END i_wb_addr[5]
  PIN i_wb_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END i_wb_addr[6]
  PIN i_wb_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 0.000 43.120 4.000 ;
    END
  END i_wb_addr[7]
  PIN i_wb_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 0.000 45.360 4.000 ;
    END
  END i_wb_addr[8]
  PIN i_wb_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END i_wb_addr[9]
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 0.000 16.240 4.000 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 0.000 25.200 4.000 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 0.000 29.680 4.000 ;
    END
  END i_wb_data[1]
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 0.000 18.480 4.000 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END i_wb_we
  PIN led_enb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 96.000 66.640 100.000 ;
    END
  END led_enb[0]
  PIN led_enb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 96.000 95.760 100.000 ;
    END
  END led_enb[1]
  PIN leds[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 96.000 81.200 100.000 ;
    END
  END leds[0]
  PIN leds[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 96.000 110.320 100.000 ;
    END
  END leds[1]
  PIN o_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.320 4.000 12.880 ;
    END
  END o_wb_ack
  PIN o_wb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 4.000 17.360 ;
    END
  END o_wb_data[0]
  PIN o_wb_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 4.000 39.760 ;
    END
  END o_wb_data[10]
  PIN o_wb_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 4.000 42.000 ;
    END
  END o_wb_data[11]
  PIN o_wb_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END o_wb_data[12]
  PIN o_wb_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 4.000 46.480 ;
    END
  END o_wb_data[13]
  PIN o_wb_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 4.000 48.720 ;
    END
  END o_wb_data[14]
  PIN o_wb_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 4.000 50.960 ;
    END
  END o_wb_data[15]
  PIN o_wb_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.640 4.000 53.200 ;
    END
  END o_wb_data[16]
  PIN o_wb_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 4.000 55.440 ;
    END
  END o_wb_data[17]
  PIN o_wb_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END o_wb_data[18]
  PIN o_wb_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 4.000 59.920 ;
    END
  END o_wb_data[19]
  PIN o_wb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 4.000 19.600 ;
    END
  END o_wb_data[1]
  PIN o_wb_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 4.000 62.160 ;
    END
  END o_wb_data[20]
  PIN o_wb_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 4.000 64.400 ;
    END
  END o_wb_data[21]
  PIN o_wb_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 4.000 66.640 ;
    END
  END o_wb_data[22]
  PIN o_wb_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 4.000 68.880 ;
    END
  END o_wb_data[23]
  PIN o_wb_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 4.000 71.120 ;
    END
  END o_wb_data[24]
  PIN o_wb_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 4.000 73.360 ;
    END
  END o_wb_data[25]
  PIN o_wb_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.040 4.000 75.600 ;
    END
  END o_wb_data[26]
  PIN o_wb_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END o_wb_data[27]
  PIN o_wb_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.520 4.000 80.080 ;
    END
  END o_wb_data[28]
  PIN o_wb_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.760 4.000 82.320 ;
    END
  END o_wb_data[29]
  PIN o_wb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.280 4.000 21.840 ;
    END
  END o_wb_data[2]
  PIN o_wb_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END o_wb_data[30]
  PIN o_wb_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.240 4.000 86.800 ;
    END
  END o_wb_data[31]
  PIN o_wb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END o_wb_data[3]
  PIN o_wb_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.760 4.000 26.320 ;
    END
  END o_wb_data[4]
  PIN o_wb_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.000 4.000 28.560 ;
    END
  END o_wb_data[5]
  PIN o_wb_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END o_wb_data[6]
  PIN o_wb_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.480 4.000 33.040 ;
    END
  END o_wb_data[7]
  PIN o_wb_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 4.000 35.280 ;
    END
  END o_wb_data[8]
  PIN o_wb_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.960 4.000 37.520 ;
    END
  END o_wb_data[9]
  PIN o_wb_stall
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 14.560 4.000 15.120 ;
    END
  END o_wb_stall
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 0.000 103.600 4.000 ;
    END
  END reset
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.220 15.380 20.820 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 45.820 15.380 47.420 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 72.420 15.380 74.020 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.020 15.380 100.620 82.620 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 32.520 15.380 34.120 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.120 15.380 60.720 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 85.720 15.380 87.320 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.320 15.380 113.920 82.620 ;
    END
  END vss
  PIN xtal_clk[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 96.000 22.960 100.000 ;
    END
  END xtal_clk[0]
  PIN xtal_clk[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 96.000 52.080 100.000 ;
    END
  END xtal_clk[1]
  PIN xtal_clk_enb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 96.000 8.400 100.000 ;
    END
  END xtal_clk_enb[0]
  PIN xtal_clk_enb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 96.000 37.520 100.000 ;
    END
  END xtal_clk_enb[1]
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.150 113.920 82.620 ;
      LAYER Metal2 ;
        RECT 7.420 95.700 7.540 96.000 ;
        RECT 8.700 95.700 22.100 96.000 ;
        RECT 23.260 95.700 36.660 96.000 ;
        RECT 37.820 95.700 51.220 96.000 ;
        RECT 52.380 95.700 65.780 96.000 ;
        RECT 66.940 95.700 80.340 96.000 ;
        RECT 81.500 95.700 94.900 96.000 ;
        RECT 96.060 95.700 109.460 96.000 ;
        RECT 110.620 95.700 113.780 96.000 ;
        RECT 7.420 4.300 113.780 95.700 ;
        RECT 7.420 4.000 15.380 4.300 ;
        RECT 16.540 4.000 17.620 4.300 ;
        RECT 18.780 4.000 19.860 4.300 ;
        RECT 21.020 4.000 22.100 4.300 ;
        RECT 23.260 4.000 24.340 4.300 ;
        RECT 25.500 4.000 26.580 4.300 ;
        RECT 27.740 4.000 28.820 4.300 ;
        RECT 29.980 4.000 31.060 4.300 ;
        RECT 32.220 4.000 33.300 4.300 ;
        RECT 34.460 4.000 35.540 4.300 ;
        RECT 36.700 4.000 37.780 4.300 ;
        RECT 38.940 4.000 40.020 4.300 ;
        RECT 41.180 4.000 42.260 4.300 ;
        RECT 43.420 4.000 44.500 4.300 ;
        RECT 45.660 4.000 46.740 4.300 ;
        RECT 47.900 4.000 48.980 4.300 ;
        RECT 50.140 4.000 51.220 4.300 ;
        RECT 52.380 4.000 53.460 4.300 ;
        RECT 54.620 4.000 55.700 4.300 ;
        RECT 56.860 4.000 57.940 4.300 ;
        RECT 59.100 4.000 60.180 4.300 ;
        RECT 61.340 4.000 62.420 4.300 ;
        RECT 63.580 4.000 64.660 4.300 ;
        RECT 65.820 4.000 66.900 4.300 ;
        RECT 68.060 4.000 69.140 4.300 ;
        RECT 70.300 4.000 71.380 4.300 ;
        RECT 72.540 4.000 73.620 4.300 ;
        RECT 74.780 4.000 75.860 4.300 ;
        RECT 77.020 4.000 78.100 4.300 ;
        RECT 79.260 4.000 80.340 4.300 ;
        RECT 81.500 4.000 82.580 4.300 ;
        RECT 83.740 4.000 84.820 4.300 ;
        RECT 85.980 4.000 87.060 4.300 ;
        RECT 88.220 4.000 89.300 4.300 ;
        RECT 90.460 4.000 91.540 4.300 ;
        RECT 92.700 4.000 93.780 4.300 ;
        RECT 94.940 4.000 96.020 4.300 ;
        RECT 97.180 4.000 98.260 4.300 ;
        RECT 99.420 4.000 100.500 4.300 ;
        RECT 101.660 4.000 102.740 4.300 ;
        RECT 103.900 4.000 113.780 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 85.940 115.700 86.660 ;
        RECT 4.000 84.860 116.000 85.940 ;
        RECT 4.300 83.700 116.000 84.860 ;
        RECT 4.000 82.620 116.000 83.700 ;
        RECT 4.300 81.460 116.000 82.620 ;
        RECT 4.000 80.380 116.000 81.460 ;
        RECT 4.300 79.220 116.000 80.380 ;
        RECT 4.000 78.140 116.000 79.220 ;
        RECT 4.300 76.980 116.000 78.140 ;
        RECT 4.000 75.900 116.000 76.980 ;
        RECT 4.300 74.740 116.000 75.900 ;
        RECT 4.000 73.660 116.000 74.740 ;
        RECT 4.300 72.500 116.000 73.660 ;
        RECT 4.000 71.420 116.000 72.500 ;
        RECT 4.300 70.260 116.000 71.420 ;
        RECT 4.000 69.180 116.000 70.260 ;
        RECT 4.300 68.020 116.000 69.180 ;
        RECT 4.000 66.940 116.000 68.020 ;
        RECT 4.300 65.780 116.000 66.940 ;
        RECT 4.000 64.700 116.000 65.780 ;
        RECT 4.300 63.540 116.000 64.700 ;
        RECT 4.000 62.460 116.000 63.540 ;
        RECT 4.300 61.300 115.700 62.460 ;
        RECT 4.000 60.220 116.000 61.300 ;
        RECT 4.300 59.060 116.000 60.220 ;
        RECT 4.000 57.980 116.000 59.060 ;
        RECT 4.300 56.820 116.000 57.980 ;
        RECT 4.000 55.740 116.000 56.820 ;
        RECT 4.300 54.580 116.000 55.740 ;
        RECT 4.000 53.500 116.000 54.580 ;
        RECT 4.300 52.340 116.000 53.500 ;
        RECT 4.000 51.260 116.000 52.340 ;
        RECT 4.300 50.100 116.000 51.260 ;
        RECT 4.000 49.020 116.000 50.100 ;
        RECT 4.300 47.860 116.000 49.020 ;
        RECT 4.000 46.780 116.000 47.860 ;
        RECT 4.300 45.620 116.000 46.780 ;
        RECT 4.000 44.540 116.000 45.620 ;
        RECT 4.300 43.380 116.000 44.540 ;
        RECT 4.000 42.300 116.000 43.380 ;
        RECT 4.300 41.140 116.000 42.300 ;
        RECT 4.000 40.060 116.000 41.140 ;
        RECT 4.300 38.900 116.000 40.060 ;
        RECT 4.000 37.820 116.000 38.900 ;
        RECT 4.300 36.660 115.700 37.820 ;
        RECT 4.000 35.580 116.000 36.660 ;
        RECT 4.300 34.420 116.000 35.580 ;
        RECT 4.000 33.340 116.000 34.420 ;
        RECT 4.300 32.180 116.000 33.340 ;
        RECT 4.000 31.100 116.000 32.180 ;
        RECT 4.300 29.940 116.000 31.100 ;
        RECT 4.000 28.860 116.000 29.940 ;
        RECT 4.300 27.700 116.000 28.860 ;
        RECT 4.000 26.620 116.000 27.700 ;
        RECT 4.300 25.460 116.000 26.620 ;
        RECT 4.000 24.380 116.000 25.460 ;
        RECT 4.300 23.220 116.000 24.380 ;
        RECT 4.000 22.140 116.000 23.220 ;
        RECT 4.300 20.980 116.000 22.140 ;
        RECT 4.000 19.900 116.000 20.980 ;
        RECT 4.300 18.740 116.000 19.900 ;
        RECT 4.000 17.660 116.000 18.740 ;
        RECT 4.300 16.500 116.000 17.660 ;
        RECT 4.000 15.420 116.000 16.500 ;
        RECT 4.300 14.260 116.000 15.420 ;
        RECT 4.000 13.180 116.000 14.260 ;
        RECT 4.300 12.460 115.700 13.180 ;
      LAYER Metal4 ;
        RECT 9.100 16.330 18.920 60.390 ;
        RECT 21.120 16.330 32.220 60.390 ;
        RECT 34.420 16.330 45.520 60.390 ;
        RECT 47.720 16.330 58.820 60.390 ;
        RECT 61.020 16.330 72.120 60.390 ;
        RECT 74.320 16.330 85.420 60.390 ;
        RECT 87.620 16.330 98.420 60.390 ;
  END
END wb_buttons_leds
END LIBRARY

