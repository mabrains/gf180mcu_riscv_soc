magic
tech gf180mcuD
magscale 1 5
timestamp 1699810877
<< obsm1 >>
rect 672 463 119280 98489
<< metal2 >>
rect 25536 99600 25592 100000
rect 26208 99600 26264 100000
rect 34272 99600 34328 100000
rect 41328 99600 41384 100000
rect 49056 99600 49112 100000
rect 53424 99600 53480 100000
rect 53760 99600 53816 100000
rect 54096 99600 54152 100000
rect 54432 99600 54488 100000
rect 54768 99600 54824 100000
rect 55104 99600 55160 100000
rect 55440 99600 55496 100000
rect 55776 99600 55832 100000
rect 56112 99600 56168 100000
rect 56448 99600 56504 100000
rect 56784 99600 56840 100000
rect 57120 99600 57176 100000
rect 57456 99600 57512 100000
rect 57792 99600 57848 100000
rect 58128 99600 58184 100000
rect 58464 99600 58520 100000
rect 58800 99600 58856 100000
rect 59136 99600 59192 100000
rect 59472 99600 59528 100000
rect 59808 99600 59864 100000
rect 60144 99600 60200 100000
rect 60480 99600 60536 100000
rect 60816 99600 60872 100000
rect 61152 99600 61208 100000
rect 61488 99600 61544 100000
rect 61824 99600 61880 100000
rect 62160 99600 62216 100000
rect 62496 99600 62552 100000
rect 62832 99600 62888 100000
rect 63168 99600 63224 100000
rect 63504 99600 63560 100000
rect 63840 99600 63896 100000
rect 64176 99600 64232 100000
rect 64512 99600 64568 100000
rect 64848 99600 64904 100000
rect 65184 99600 65240 100000
rect 65520 99600 65576 100000
rect 65856 99600 65912 100000
rect 66192 99600 66248 100000
rect 66528 99600 66584 100000
rect 66864 99600 66920 100000
rect 67200 99600 67256 100000
rect 67536 99600 67592 100000
rect 67872 99600 67928 100000
rect 68208 99600 68264 100000
rect 68544 99600 68600 100000
rect 68880 99600 68936 100000
rect 69216 99600 69272 100000
rect 69552 99600 69608 100000
rect 69888 99600 69944 100000
rect 80640 99600 80696 100000
rect 82656 99600 82712 100000
rect 82992 99600 83048 100000
rect 83328 99600 83384 100000
rect 85008 99600 85064 100000
rect 87696 99600 87752 100000
rect 88032 99600 88088 100000
rect 88368 99600 88424 100000
rect 88704 99600 88760 100000
rect 89040 99600 89096 100000
rect 89376 99600 89432 100000
rect 90384 99600 90440 100000
rect 93072 99600 93128 100000
rect 93408 99600 93464 100000
rect 98448 99600 98504 100000
rect 98784 99600 98840 100000
rect 99120 99600 99176 100000
rect 99456 99600 99512 100000
rect 99792 99600 99848 100000
rect 100128 99600 100184 100000
rect 100464 99600 100520 100000
rect 100800 99600 100856 100000
rect 101136 99600 101192 100000
rect 101472 99600 101528 100000
rect 103824 99600 103880 100000
rect 105504 99600 105560 100000
rect 106176 99600 106232 100000
rect 106848 99600 106904 100000
rect 107184 99600 107240 100000
rect 111552 99600 111608 100000
rect 0 0 56 400
rect 336 0 392 400
rect 14448 0 14504 400
rect 14784 0 14840 400
rect 15120 0 15176 400
rect 15456 0 15512 400
rect 15792 0 15848 400
rect 16128 0 16184 400
rect 16464 0 16520 400
rect 16800 0 16856 400
rect 17136 0 17192 400
rect 17472 0 17528 400
rect 17808 0 17864 400
rect 18144 0 18200 400
rect 18480 0 18536 400
rect 18816 0 18872 400
rect 19152 0 19208 400
rect 19488 0 19544 400
rect 19824 0 19880 400
rect 20160 0 20216 400
rect 20496 0 20552 400
rect 20832 0 20888 400
rect 21168 0 21224 400
rect 21504 0 21560 400
rect 21840 0 21896 400
rect 22176 0 22232 400
rect 22512 0 22568 400
rect 22848 0 22904 400
rect 23184 0 23240 400
rect 23520 0 23576 400
rect 23856 0 23912 400
rect 24192 0 24248 400
rect 24528 0 24584 400
rect 24864 0 24920 400
rect 25200 0 25256 400
rect 25536 0 25592 400
rect 25872 0 25928 400
rect 26208 0 26264 400
rect 26544 0 26600 400
rect 26880 0 26936 400
rect 27216 0 27272 400
rect 27552 0 27608 400
rect 27888 0 27944 400
rect 28224 0 28280 400
rect 28560 0 28616 400
rect 28896 0 28952 400
rect 29232 0 29288 400
rect 29568 0 29624 400
rect 29904 0 29960 400
rect 30240 0 30296 400
rect 30576 0 30632 400
rect 30912 0 30968 400
rect 31248 0 31304 400
rect 31584 0 31640 400
rect 31920 0 31976 400
rect 32256 0 32312 400
rect 32592 0 32648 400
rect 32928 0 32984 400
rect 33264 0 33320 400
rect 33600 0 33656 400
rect 33936 0 33992 400
rect 34272 0 34328 400
rect 34608 0 34664 400
rect 34944 0 35000 400
rect 35280 0 35336 400
rect 35616 0 35672 400
rect 35952 0 36008 400
rect 36288 0 36344 400
rect 36624 0 36680 400
rect 36960 0 37016 400
rect 37296 0 37352 400
rect 37632 0 37688 400
rect 37968 0 38024 400
rect 38304 0 38360 400
rect 38640 0 38696 400
rect 38976 0 39032 400
rect 39312 0 39368 400
rect 39648 0 39704 400
rect 39984 0 40040 400
rect 40320 0 40376 400
rect 40656 0 40712 400
rect 40992 0 41048 400
rect 41328 0 41384 400
rect 41664 0 41720 400
rect 42000 0 42056 400
rect 42336 0 42392 400
rect 42672 0 42728 400
rect 43008 0 43064 400
rect 43344 0 43400 400
rect 43680 0 43736 400
rect 44016 0 44072 400
rect 44352 0 44408 400
rect 44688 0 44744 400
rect 45024 0 45080 400
rect 45360 0 45416 400
rect 45696 0 45752 400
rect 46032 0 46088 400
rect 46368 0 46424 400
rect 46704 0 46760 400
rect 47040 0 47096 400
rect 47376 0 47432 400
rect 47712 0 47768 400
rect 48048 0 48104 400
rect 48384 0 48440 400
rect 48720 0 48776 400
rect 49056 0 49112 400
rect 49392 0 49448 400
rect 49728 0 49784 400
rect 50064 0 50120 400
rect 50400 0 50456 400
rect 50736 0 50792 400
rect 51072 0 51128 400
rect 51408 0 51464 400
rect 51744 0 51800 400
rect 52080 0 52136 400
rect 52416 0 52472 400
rect 52752 0 52808 400
rect 53088 0 53144 400
rect 53424 0 53480 400
rect 53760 0 53816 400
rect 54096 0 54152 400
rect 54432 0 54488 400
rect 54768 0 54824 400
rect 55104 0 55160 400
rect 55440 0 55496 400
rect 55776 0 55832 400
rect 56112 0 56168 400
rect 56448 0 56504 400
rect 56784 0 56840 400
rect 57120 0 57176 400
rect 57456 0 57512 400
rect 57792 0 57848 400
rect 58128 0 58184 400
rect 58464 0 58520 400
rect 58800 0 58856 400
rect 59136 0 59192 400
rect 59472 0 59528 400
rect 59808 0 59864 400
rect 60144 0 60200 400
rect 60480 0 60536 400
rect 60816 0 60872 400
rect 61152 0 61208 400
rect 61488 0 61544 400
rect 61824 0 61880 400
rect 62160 0 62216 400
rect 62496 0 62552 400
rect 62832 0 62888 400
rect 63168 0 63224 400
rect 63504 0 63560 400
rect 63840 0 63896 400
rect 64176 0 64232 400
rect 64512 0 64568 400
rect 64848 0 64904 400
rect 65184 0 65240 400
rect 65520 0 65576 400
rect 65856 0 65912 400
rect 66192 0 66248 400
rect 66528 0 66584 400
rect 66864 0 66920 400
rect 67200 0 67256 400
rect 67536 0 67592 400
rect 67872 0 67928 400
rect 68208 0 68264 400
rect 68544 0 68600 400
rect 68880 0 68936 400
rect 69216 0 69272 400
rect 69552 0 69608 400
rect 69888 0 69944 400
rect 70224 0 70280 400
rect 70560 0 70616 400
rect 70896 0 70952 400
rect 71232 0 71288 400
rect 71568 0 71624 400
rect 71904 0 71960 400
rect 72240 0 72296 400
rect 72576 0 72632 400
rect 72912 0 72968 400
rect 73248 0 73304 400
rect 73584 0 73640 400
rect 73920 0 73976 400
rect 74256 0 74312 400
rect 74592 0 74648 400
rect 74928 0 74984 400
rect 75264 0 75320 400
rect 75600 0 75656 400
rect 75936 0 75992 400
rect 76272 0 76328 400
rect 76608 0 76664 400
rect 76944 0 77000 400
rect 77280 0 77336 400
rect 77616 0 77672 400
rect 77952 0 78008 400
rect 78288 0 78344 400
rect 78624 0 78680 400
rect 78960 0 79016 400
rect 79296 0 79352 400
rect 79632 0 79688 400
rect 79968 0 80024 400
rect 80304 0 80360 400
rect 80640 0 80696 400
rect 80976 0 81032 400
rect 81312 0 81368 400
rect 81648 0 81704 400
rect 81984 0 82040 400
rect 82320 0 82376 400
rect 82656 0 82712 400
rect 82992 0 83048 400
rect 83328 0 83384 400
rect 83664 0 83720 400
rect 84000 0 84056 400
rect 84336 0 84392 400
rect 84672 0 84728 400
rect 85008 0 85064 400
rect 85344 0 85400 400
rect 85680 0 85736 400
rect 86016 0 86072 400
rect 86352 0 86408 400
rect 86688 0 86744 400
rect 87024 0 87080 400
rect 87360 0 87416 400
rect 87696 0 87752 400
rect 88032 0 88088 400
rect 90048 0 90104 400
rect 90384 0 90440 400
rect 90720 0 90776 400
rect 95424 0 95480 400
rect 99792 0 99848 400
rect 102144 0 102200 400
rect 102480 0 102536 400
rect 103152 0 103208 400
rect 103824 0 103880 400
rect 104496 0 104552 400
rect 104832 0 104888 400
rect 105504 0 105560 400
rect 110208 0 110264 400
rect 112560 0 112616 400
rect 113904 0 113960 400
<< obsm2 >>
rect 798 99570 25506 99666
rect 25622 99570 26178 99666
rect 26294 99570 34242 99666
rect 34358 99570 41298 99666
rect 41414 99570 49026 99666
rect 49142 99570 53394 99666
rect 53510 99570 53730 99666
rect 53846 99570 54066 99666
rect 54182 99570 54402 99666
rect 54518 99570 54738 99666
rect 54854 99570 55074 99666
rect 55190 99570 55410 99666
rect 55526 99570 55746 99666
rect 55862 99570 56082 99666
rect 56198 99570 56418 99666
rect 56534 99570 56754 99666
rect 56870 99570 57090 99666
rect 57206 99570 57426 99666
rect 57542 99570 57762 99666
rect 57878 99570 58098 99666
rect 58214 99570 58434 99666
rect 58550 99570 58770 99666
rect 58886 99570 59106 99666
rect 59222 99570 59442 99666
rect 59558 99570 59778 99666
rect 59894 99570 60114 99666
rect 60230 99570 60450 99666
rect 60566 99570 60786 99666
rect 60902 99570 61122 99666
rect 61238 99570 61458 99666
rect 61574 99570 61794 99666
rect 61910 99570 62130 99666
rect 62246 99570 62466 99666
rect 62582 99570 62802 99666
rect 62918 99570 63138 99666
rect 63254 99570 63474 99666
rect 63590 99570 63810 99666
rect 63926 99570 64146 99666
rect 64262 99570 64482 99666
rect 64598 99570 64818 99666
rect 64934 99570 65154 99666
rect 65270 99570 65490 99666
rect 65606 99570 65826 99666
rect 65942 99570 66162 99666
rect 66278 99570 66498 99666
rect 66614 99570 66834 99666
rect 66950 99570 67170 99666
rect 67286 99570 67506 99666
rect 67622 99570 67842 99666
rect 67958 99570 68178 99666
rect 68294 99570 68514 99666
rect 68630 99570 68850 99666
rect 68966 99570 69186 99666
rect 69302 99570 69522 99666
rect 69638 99570 69858 99666
rect 69974 99570 80610 99666
rect 80726 99570 82626 99666
rect 82742 99570 82962 99666
rect 83078 99570 83298 99666
rect 83414 99570 84978 99666
rect 85094 99570 87666 99666
rect 87782 99570 88002 99666
rect 88118 99570 88338 99666
rect 88454 99570 88674 99666
rect 88790 99570 89010 99666
rect 89126 99570 89346 99666
rect 89462 99570 90354 99666
rect 90470 99570 93042 99666
rect 93158 99570 93378 99666
rect 93494 99570 98418 99666
rect 98534 99570 98754 99666
rect 98870 99570 99090 99666
rect 99206 99570 99426 99666
rect 99542 99570 99762 99666
rect 99878 99570 100098 99666
rect 100214 99570 100434 99666
rect 100550 99570 100770 99666
rect 100886 99570 101106 99666
rect 101222 99570 101442 99666
rect 101558 99570 103794 99666
rect 103910 99570 105474 99666
rect 105590 99570 106146 99666
rect 106262 99570 106818 99666
rect 106934 99570 107154 99666
rect 107270 99570 111522 99666
rect 111638 99570 119322 99666
rect 798 430 119322 99570
rect 798 350 14418 430
rect 14534 350 14754 430
rect 14870 350 15090 430
rect 15206 350 15426 430
rect 15542 350 15762 430
rect 15878 350 16098 430
rect 16214 350 16434 430
rect 16550 350 16770 430
rect 16886 350 17106 430
rect 17222 350 17442 430
rect 17558 350 17778 430
rect 17894 350 18114 430
rect 18230 350 18450 430
rect 18566 350 18786 430
rect 18902 350 19122 430
rect 19238 350 19458 430
rect 19574 350 19794 430
rect 19910 350 20130 430
rect 20246 350 20466 430
rect 20582 350 20802 430
rect 20918 350 21138 430
rect 21254 350 21474 430
rect 21590 350 21810 430
rect 21926 350 22146 430
rect 22262 350 22482 430
rect 22598 350 22818 430
rect 22934 350 23154 430
rect 23270 350 23490 430
rect 23606 350 23826 430
rect 23942 350 24162 430
rect 24278 350 24498 430
rect 24614 350 24834 430
rect 24950 350 25170 430
rect 25286 350 25506 430
rect 25622 350 25842 430
rect 25958 350 26178 430
rect 26294 350 26514 430
rect 26630 350 26850 430
rect 26966 350 27186 430
rect 27302 350 27522 430
rect 27638 350 27858 430
rect 27974 350 28194 430
rect 28310 350 28530 430
rect 28646 350 28866 430
rect 28982 350 29202 430
rect 29318 350 29538 430
rect 29654 350 29874 430
rect 29990 350 30210 430
rect 30326 350 30546 430
rect 30662 350 30882 430
rect 30998 350 31218 430
rect 31334 350 31554 430
rect 31670 350 31890 430
rect 32006 350 32226 430
rect 32342 350 32562 430
rect 32678 350 32898 430
rect 33014 350 33234 430
rect 33350 350 33570 430
rect 33686 350 33906 430
rect 34022 350 34242 430
rect 34358 350 34578 430
rect 34694 350 34914 430
rect 35030 350 35250 430
rect 35366 350 35586 430
rect 35702 350 35922 430
rect 36038 350 36258 430
rect 36374 350 36594 430
rect 36710 350 36930 430
rect 37046 350 37266 430
rect 37382 350 37602 430
rect 37718 350 37938 430
rect 38054 350 38274 430
rect 38390 350 38610 430
rect 38726 350 38946 430
rect 39062 350 39282 430
rect 39398 350 39618 430
rect 39734 350 39954 430
rect 40070 350 40290 430
rect 40406 350 40626 430
rect 40742 350 40962 430
rect 41078 350 41298 430
rect 41414 350 41634 430
rect 41750 350 41970 430
rect 42086 350 42306 430
rect 42422 350 42642 430
rect 42758 350 42978 430
rect 43094 350 43314 430
rect 43430 350 43650 430
rect 43766 350 43986 430
rect 44102 350 44322 430
rect 44438 350 44658 430
rect 44774 350 44994 430
rect 45110 350 45330 430
rect 45446 350 45666 430
rect 45782 350 46002 430
rect 46118 350 46338 430
rect 46454 350 46674 430
rect 46790 350 47010 430
rect 47126 350 47346 430
rect 47462 350 47682 430
rect 47798 350 48018 430
rect 48134 350 48354 430
rect 48470 350 48690 430
rect 48806 350 49026 430
rect 49142 350 49362 430
rect 49478 350 49698 430
rect 49814 350 50034 430
rect 50150 350 50370 430
rect 50486 350 50706 430
rect 50822 350 51042 430
rect 51158 350 51378 430
rect 51494 350 51714 430
rect 51830 350 52050 430
rect 52166 350 52386 430
rect 52502 350 52722 430
rect 52838 350 53058 430
rect 53174 350 53394 430
rect 53510 350 53730 430
rect 53846 350 54066 430
rect 54182 350 54402 430
rect 54518 350 54738 430
rect 54854 350 55074 430
rect 55190 350 55410 430
rect 55526 350 55746 430
rect 55862 350 56082 430
rect 56198 350 56418 430
rect 56534 350 56754 430
rect 56870 350 57090 430
rect 57206 350 57426 430
rect 57542 350 57762 430
rect 57878 350 58098 430
rect 58214 350 58434 430
rect 58550 350 58770 430
rect 58886 350 59106 430
rect 59222 350 59442 430
rect 59558 350 59778 430
rect 59894 350 60114 430
rect 60230 350 60450 430
rect 60566 350 60786 430
rect 60902 350 61122 430
rect 61238 350 61458 430
rect 61574 350 61794 430
rect 61910 350 62130 430
rect 62246 350 62466 430
rect 62582 350 62802 430
rect 62918 350 63138 430
rect 63254 350 63474 430
rect 63590 350 63810 430
rect 63926 350 64146 430
rect 64262 350 64482 430
rect 64598 350 64818 430
rect 64934 350 65154 430
rect 65270 350 65490 430
rect 65606 350 65826 430
rect 65942 350 66162 430
rect 66278 350 66498 430
rect 66614 350 66834 430
rect 66950 350 67170 430
rect 67286 350 67506 430
rect 67622 350 67842 430
rect 67958 350 68178 430
rect 68294 350 68514 430
rect 68630 350 68850 430
rect 68966 350 69186 430
rect 69302 350 69522 430
rect 69638 350 69858 430
rect 69974 350 70194 430
rect 70310 350 70530 430
rect 70646 350 70866 430
rect 70982 350 71202 430
rect 71318 350 71538 430
rect 71654 350 71874 430
rect 71990 350 72210 430
rect 72326 350 72546 430
rect 72662 350 72882 430
rect 72998 350 73218 430
rect 73334 350 73554 430
rect 73670 350 73890 430
rect 74006 350 74226 430
rect 74342 350 74562 430
rect 74678 350 74898 430
rect 75014 350 75234 430
rect 75350 350 75570 430
rect 75686 350 75906 430
rect 76022 350 76242 430
rect 76358 350 76578 430
rect 76694 350 76914 430
rect 77030 350 77250 430
rect 77366 350 77586 430
rect 77702 350 77922 430
rect 78038 350 78258 430
rect 78374 350 78594 430
rect 78710 350 78930 430
rect 79046 350 79266 430
rect 79382 350 79602 430
rect 79718 350 79938 430
rect 80054 350 80274 430
rect 80390 350 80610 430
rect 80726 350 80946 430
rect 81062 350 81282 430
rect 81398 350 81618 430
rect 81734 350 81954 430
rect 82070 350 82290 430
rect 82406 350 82626 430
rect 82742 350 82962 430
rect 83078 350 83298 430
rect 83414 350 83634 430
rect 83750 350 83970 430
rect 84086 350 84306 430
rect 84422 350 84642 430
rect 84758 350 84978 430
rect 85094 350 85314 430
rect 85430 350 85650 430
rect 85766 350 85986 430
rect 86102 350 86322 430
rect 86438 350 86658 430
rect 86774 350 86994 430
rect 87110 350 87330 430
rect 87446 350 87666 430
rect 87782 350 88002 430
rect 88118 350 90018 430
rect 90134 350 90354 430
rect 90470 350 90690 430
rect 90806 350 95394 430
rect 95510 350 99762 430
rect 99878 350 102114 430
rect 102230 350 102450 430
rect 102566 350 103122 430
rect 103238 350 103794 430
rect 103910 350 104466 430
rect 104582 350 104802 430
rect 104918 350 105474 430
rect 105590 350 110178 430
rect 110294 350 112530 430
rect 112646 350 113874 430
rect 113990 350 119322 430
<< metal3 >>
rect 119600 98112 120000 98168
rect 0 97776 400 97832
rect 119600 97776 120000 97832
rect 119600 97440 120000 97496
rect 119600 95760 120000 95816
rect 119600 95424 120000 95480
rect 119600 95088 120000 95144
rect 119600 94752 120000 94808
rect 119600 93408 120000 93464
rect 119600 93072 120000 93128
rect 119600 90048 120000 90104
rect 119600 89712 120000 89768
rect 119600 89376 120000 89432
rect 119600 87696 120000 87752
rect 0 87360 400 87416
rect 0 86352 400 86408
rect 0 84336 400 84392
rect 119600 83328 120000 83384
rect 119600 82992 120000 83048
rect 0 82656 400 82712
rect 0 82320 400 82376
rect 0 81984 400 82040
rect 0 81648 400 81704
rect 119600 81648 120000 81704
rect 0 81312 400 81368
rect 119600 81312 120000 81368
rect 0 80976 400 81032
rect 0 80640 400 80696
rect 0 80304 400 80360
rect 0 79968 400 80024
rect 0 79632 400 79688
rect 0 79296 400 79352
rect 0 78960 400 79016
rect 0 78624 400 78680
rect 0 78288 400 78344
rect 0 77952 400 78008
rect 0 77616 400 77672
rect 0 77280 400 77336
rect 0 76944 400 77000
rect 0 76608 400 76664
rect 0 76272 400 76328
rect 0 75936 400 75992
rect 0 75600 400 75656
rect 0 75264 400 75320
rect 0 74928 400 74984
rect 0 74592 400 74648
rect 0 74256 400 74312
rect 0 73920 400 73976
rect 0 73584 400 73640
rect 0 73248 400 73304
rect 0 72912 400 72968
rect 0 72576 400 72632
rect 0 72240 400 72296
rect 0 71904 400 71960
rect 0 71568 400 71624
rect 0 71232 400 71288
rect 0 70896 400 70952
rect 0 70560 400 70616
rect 0 70224 400 70280
rect 0 69888 400 69944
rect 0 69552 400 69608
rect 0 69216 400 69272
rect 0 68880 400 68936
rect 0 68544 400 68600
rect 0 68208 400 68264
rect 0 67872 400 67928
rect 0 67536 400 67592
rect 0 67200 400 67256
rect 0 66864 400 66920
rect 0 66528 400 66584
rect 0 66192 400 66248
rect 0 65856 400 65912
rect 0 65520 400 65576
rect 0 65184 400 65240
rect 0 64848 400 64904
rect 0 64512 400 64568
rect 0 64176 400 64232
rect 0 63840 400 63896
rect 0 63504 400 63560
rect 0 63168 400 63224
rect 0 62832 400 62888
rect 0 62496 400 62552
rect 0 62160 400 62216
rect 0 61824 400 61880
rect 0 61488 400 61544
rect 0 61152 400 61208
rect 0 60816 400 60872
rect 0 60480 400 60536
rect 0 60144 400 60200
rect 0 59808 400 59864
rect 0 59472 400 59528
rect 0 59136 400 59192
rect 0 58800 400 58856
rect 0 58464 400 58520
rect 0 58128 400 58184
rect 0 57792 400 57848
rect 0 57456 400 57512
rect 0 57120 400 57176
rect 0 56784 400 56840
rect 0 56448 400 56504
rect 0 56112 400 56168
rect 0 55776 400 55832
rect 0 55440 400 55496
rect 0 55104 400 55160
rect 0 54768 400 54824
rect 0 54432 400 54488
rect 0 54096 400 54152
rect 0 53760 400 53816
rect 0 53424 400 53480
rect 0 53088 400 53144
rect 0 52752 400 52808
rect 0 52416 400 52472
rect 0 52080 400 52136
rect 0 51744 400 51800
rect 0 51408 400 51464
rect 0 51072 400 51128
rect 0 50736 400 50792
rect 0 50400 400 50456
rect 0 50064 400 50120
rect 0 49728 400 49784
rect 0 49392 400 49448
rect 0 49056 400 49112
rect 0 48720 400 48776
rect 0 48384 400 48440
rect 0 48048 400 48104
rect 0 47712 400 47768
rect 0 47376 400 47432
rect 0 47040 400 47096
rect 0 46704 400 46760
rect 0 46368 400 46424
rect 0 46032 400 46088
rect 0 45696 400 45752
rect 119600 45696 120000 45752
rect 0 45360 400 45416
rect 0 45024 400 45080
rect 0 44688 400 44744
rect 0 44352 400 44408
rect 0 44016 400 44072
rect 0 43680 400 43736
rect 0 43344 400 43400
rect 0 43008 400 43064
rect 0 42672 400 42728
rect 0 42336 400 42392
rect 0 42000 400 42056
rect 0 41664 400 41720
rect 0 41328 400 41384
rect 0 40992 400 41048
rect 0 40656 400 40712
rect 0 40320 400 40376
rect 0 39984 400 40040
rect 0 39648 400 39704
rect 0 39312 400 39368
rect 119600 39312 120000 39368
rect 0 38976 400 39032
rect 0 38640 400 38696
rect 0 38304 400 38360
rect 119600 38304 120000 38360
rect 0 37968 400 38024
rect 119600 37968 120000 38024
rect 0 37632 400 37688
rect 119600 37632 120000 37688
rect 0 37296 400 37352
rect 119600 37296 120000 37352
rect 0 36960 400 37016
rect 0 36624 400 36680
rect 119600 36624 120000 36680
rect 0 36288 400 36344
rect 119600 36288 120000 36344
rect 0 35952 400 36008
rect 0 35616 400 35672
rect 0 35280 400 35336
rect 0 34944 400 35000
rect 0 34608 400 34664
rect 0 34272 400 34328
rect 119600 34272 120000 34328
rect 119600 33936 120000 33992
rect 119600 33264 120000 33320
rect 119600 32928 120000 32984
rect 0 32592 400 32648
rect 0 32256 400 32312
rect 119600 32256 120000 32312
rect 0 31920 400 31976
rect 0 31584 400 31640
rect 0 31248 400 31304
rect 119600 31248 120000 31304
rect 0 30912 400 30968
rect 119600 30912 120000 30968
rect 0 30576 400 30632
rect 119600 30576 120000 30632
rect 0 30240 400 30296
rect 0 29904 400 29960
rect 119600 29904 120000 29960
rect 0 29568 400 29624
rect 0 29232 400 29288
rect 0 28896 400 28952
rect 0 28560 400 28616
rect 119600 28560 120000 28616
rect 0 28224 400 28280
rect 0 27888 400 27944
rect 0 27552 400 27608
rect 0 27216 400 27272
rect 119600 27216 120000 27272
rect 0 26880 400 26936
rect 0 26544 400 26600
rect 0 26208 400 26264
rect 119600 26208 120000 26264
rect 0 25872 400 25928
rect 119600 25872 120000 25928
rect 0 25536 400 25592
rect 119600 25536 120000 25592
rect 0 25200 400 25256
rect 0 24864 400 24920
rect 0 24528 400 24584
rect 119600 24528 120000 24584
rect 0 24192 400 24248
rect 119600 24192 120000 24248
rect 0 23856 400 23912
rect 0 23520 400 23576
rect 0 23184 400 23240
rect 0 22848 400 22904
rect 0 22512 400 22568
rect 0 22176 400 22232
rect 0 21840 400 21896
rect 0 21504 400 21560
rect 0 21168 400 21224
rect 0 20832 400 20888
rect 0 20496 400 20552
rect 0 20160 400 20216
rect 0 19824 400 19880
rect 0 19488 400 19544
rect 0 19152 400 19208
<< obsm3 >>
rect 400 98198 119658 98406
rect 400 98082 119570 98198
rect 400 97862 119658 98082
rect 430 97746 119570 97862
rect 400 97526 119658 97746
rect 400 97410 119570 97526
rect 400 95846 119658 97410
rect 400 95730 119570 95846
rect 400 95510 119658 95730
rect 400 95394 119570 95510
rect 400 95174 119658 95394
rect 400 95058 119570 95174
rect 400 94838 119658 95058
rect 400 94722 119570 94838
rect 400 93494 119658 94722
rect 400 93378 119570 93494
rect 400 93158 119658 93378
rect 400 93042 119570 93158
rect 400 90134 119658 93042
rect 400 90018 119570 90134
rect 400 89798 119658 90018
rect 400 89682 119570 89798
rect 400 89462 119658 89682
rect 400 89346 119570 89462
rect 400 87782 119658 89346
rect 400 87666 119570 87782
rect 400 87446 119658 87666
rect 430 87330 119658 87446
rect 400 86438 119658 87330
rect 430 86322 119658 86438
rect 400 84422 119658 86322
rect 430 84306 119658 84422
rect 400 83414 119658 84306
rect 400 83298 119570 83414
rect 400 83078 119658 83298
rect 400 82962 119570 83078
rect 400 82742 119658 82962
rect 430 82626 119658 82742
rect 400 82406 119658 82626
rect 430 82290 119658 82406
rect 400 82070 119658 82290
rect 430 81954 119658 82070
rect 400 81734 119658 81954
rect 430 81618 119570 81734
rect 400 81398 119658 81618
rect 430 81282 119570 81398
rect 400 81062 119658 81282
rect 430 80946 119658 81062
rect 400 80726 119658 80946
rect 430 80610 119658 80726
rect 400 80390 119658 80610
rect 430 80274 119658 80390
rect 400 80054 119658 80274
rect 430 79938 119658 80054
rect 400 79718 119658 79938
rect 430 79602 119658 79718
rect 400 79382 119658 79602
rect 430 79266 119658 79382
rect 400 79046 119658 79266
rect 430 78930 119658 79046
rect 400 78710 119658 78930
rect 430 78594 119658 78710
rect 400 78374 119658 78594
rect 430 78258 119658 78374
rect 400 78038 119658 78258
rect 430 77922 119658 78038
rect 400 77702 119658 77922
rect 430 77586 119658 77702
rect 400 77366 119658 77586
rect 430 77250 119658 77366
rect 400 77030 119658 77250
rect 430 76914 119658 77030
rect 400 76694 119658 76914
rect 430 76578 119658 76694
rect 400 76358 119658 76578
rect 430 76242 119658 76358
rect 400 76022 119658 76242
rect 430 75906 119658 76022
rect 400 75686 119658 75906
rect 430 75570 119658 75686
rect 400 75350 119658 75570
rect 430 75234 119658 75350
rect 400 75014 119658 75234
rect 430 74898 119658 75014
rect 400 74678 119658 74898
rect 430 74562 119658 74678
rect 400 74342 119658 74562
rect 430 74226 119658 74342
rect 400 74006 119658 74226
rect 430 73890 119658 74006
rect 400 73670 119658 73890
rect 430 73554 119658 73670
rect 400 73334 119658 73554
rect 430 73218 119658 73334
rect 400 72998 119658 73218
rect 430 72882 119658 72998
rect 400 72662 119658 72882
rect 430 72546 119658 72662
rect 400 72326 119658 72546
rect 430 72210 119658 72326
rect 400 71990 119658 72210
rect 430 71874 119658 71990
rect 400 71654 119658 71874
rect 430 71538 119658 71654
rect 400 71318 119658 71538
rect 430 71202 119658 71318
rect 400 70982 119658 71202
rect 430 70866 119658 70982
rect 400 70646 119658 70866
rect 430 70530 119658 70646
rect 400 70310 119658 70530
rect 430 70194 119658 70310
rect 400 69974 119658 70194
rect 430 69858 119658 69974
rect 400 69638 119658 69858
rect 430 69522 119658 69638
rect 400 69302 119658 69522
rect 430 69186 119658 69302
rect 400 68966 119658 69186
rect 430 68850 119658 68966
rect 400 68630 119658 68850
rect 430 68514 119658 68630
rect 400 68294 119658 68514
rect 430 68178 119658 68294
rect 400 67958 119658 68178
rect 430 67842 119658 67958
rect 400 67622 119658 67842
rect 430 67506 119658 67622
rect 400 67286 119658 67506
rect 430 67170 119658 67286
rect 400 66950 119658 67170
rect 430 66834 119658 66950
rect 400 66614 119658 66834
rect 430 66498 119658 66614
rect 400 66278 119658 66498
rect 430 66162 119658 66278
rect 400 65942 119658 66162
rect 430 65826 119658 65942
rect 400 65606 119658 65826
rect 430 65490 119658 65606
rect 400 65270 119658 65490
rect 430 65154 119658 65270
rect 400 64934 119658 65154
rect 430 64818 119658 64934
rect 400 64598 119658 64818
rect 430 64482 119658 64598
rect 400 64262 119658 64482
rect 430 64146 119658 64262
rect 400 63926 119658 64146
rect 430 63810 119658 63926
rect 400 63590 119658 63810
rect 430 63474 119658 63590
rect 400 63254 119658 63474
rect 430 63138 119658 63254
rect 400 62918 119658 63138
rect 430 62802 119658 62918
rect 400 62582 119658 62802
rect 430 62466 119658 62582
rect 400 62246 119658 62466
rect 430 62130 119658 62246
rect 400 61910 119658 62130
rect 430 61794 119658 61910
rect 400 61574 119658 61794
rect 430 61458 119658 61574
rect 400 61238 119658 61458
rect 430 61122 119658 61238
rect 400 60902 119658 61122
rect 430 60786 119658 60902
rect 400 60566 119658 60786
rect 430 60450 119658 60566
rect 400 60230 119658 60450
rect 430 60114 119658 60230
rect 400 59894 119658 60114
rect 430 59778 119658 59894
rect 400 59558 119658 59778
rect 430 59442 119658 59558
rect 400 59222 119658 59442
rect 430 59106 119658 59222
rect 400 58886 119658 59106
rect 430 58770 119658 58886
rect 400 58550 119658 58770
rect 430 58434 119658 58550
rect 400 58214 119658 58434
rect 430 58098 119658 58214
rect 400 57878 119658 58098
rect 430 57762 119658 57878
rect 400 57542 119658 57762
rect 430 57426 119658 57542
rect 400 57206 119658 57426
rect 430 57090 119658 57206
rect 400 56870 119658 57090
rect 430 56754 119658 56870
rect 400 56534 119658 56754
rect 430 56418 119658 56534
rect 400 56198 119658 56418
rect 430 56082 119658 56198
rect 400 55862 119658 56082
rect 430 55746 119658 55862
rect 400 55526 119658 55746
rect 430 55410 119658 55526
rect 400 55190 119658 55410
rect 430 55074 119658 55190
rect 400 54854 119658 55074
rect 430 54738 119658 54854
rect 400 54518 119658 54738
rect 430 54402 119658 54518
rect 400 54182 119658 54402
rect 430 54066 119658 54182
rect 400 53846 119658 54066
rect 430 53730 119658 53846
rect 400 53510 119658 53730
rect 430 53394 119658 53510
rect 400 53174 119658 53394
rect 430 53058 119658 53174
rect 400 52838 119658 53058
rect 430 52722 119658 52838
rect 400 52502 119658 52722
rect 430 52386 119658 52502
rect 400 52166 119658 52386
rect 430 52050 119658 52166
rect 400 51830 119658 52050
rect 430 51714 119658 51830
rect 400 51494 119658 51714
rect 430 51378 119658 51494
rect 400 51158 119658 51378
rect 430 51042 119658 51158
rect 400 50822 119658 51042
rect 430 50706 119658 50822
rect 400 50486 119658 50706
rect 430 50370 119658 50486
rect 400 50150 119658 50370
rect 430 50034 119658 50150
rect 400 49814 119658 50034
rect 430 49698 119658 49814
rect 400 49478 119658 49698
rect 430 49362 119658 49478
rect 400 49142 119658 49362
rect 430 49026 119658 49142
rect 400 48806 119658 49026
rect 430 48690 119658 48806
rect 400 48470 119658 48690
rect 430 48354 119658 48470
rect 400 48134 119658 48354
rect 430 48018 119658 48134
rect 400 47798 119658 48018
rect 430 47682 119658 47798
rect 400 47462 119658 47682
rect 430 47346 119658 47462
rect 400 47126 119658 47346
rect 430 47010 119658 47126
rect 400 46790 119658 47010
rect 430 46674 119658 46790
rect 400 46454 119658 46674
rect 430 46338 119658 46454
rect 400 46118 119658 46338
rect 430 46002 119658 46118
rect 400 45782 119658 46002
rect 430 45666 119570 45782
rect 400 45446 119658 45666
rect 430 45330 119658 45446
rect 400 45110 119658 45330
rect 430 44994 119658 45110
rect 400 44774 119658 44994
rect 430 44658 119658 44774
rect 400 44438 119658 44658
rect 430 44322 119658 44438
rect 400 44102 119658 44322
rect 430 43986 119658 44102
rect 400 43766 119658 43986
rect 430 43650 119658 43766
rect 400 43430 119658 43650
rect 430 43314 119658 43430
rect 400 43094 119658 43314
rect 430 42978 119658 43094
rect 400 42758 119658 42978
rect 430 42642 119658 42758
rect 400 42422 119658 42642
rect 430 42306 119658 42422
rect 400 42086 119658 42306
rect 430 41970 119658 42086
rect 400 41750 119658 41970
rect 430 41634 119658 41750
rect 400 41414 119658 41634
rect 430 41298 119658 41414
rect 400 41078 119658 41298
rect 430 40962 119658 41078
rect 400 40742 119658 40962
rect 430 40626 119658 40742
rect 400 40406 119658 40626
rect 430 40290 119658 40406
rect 400 40070 119658 40290
rect 430 39954 119658 40070
rect 400 39734 119658 39954
rect 430 39618 119658 39734
rect 400 39398 119658 39618
rect 430 39282 119570 39398
rect 400 39062 119658 39282
rect 430 38946 119658 39062
rect 400 38726 119658 38946
rect 430 38610 119658 38726
rect 400 38390 119658 38610
rect 430 38274 119570 38390
rect 400 38054 119658 38274
rect 430 37938 119570 38054
rect 400 37718 119658 37938
rect 430 37602 119570 37718
rect 400 37382 119658 37602
rect 430 37266 119570 37382
rect 400 37046 119658 37266
rect 430 36930 119658 37046
rect 400 36710 119658 36930
rect 430 36594 119570 36710
rect 400 36374 119658 36594
rect 430 36258 119570 36374
rect 400 36038 119658 36258
rect 430 35922 119658 36038
rect 400 35702 119658 35922
rect 430 35586 119658 35702
rect 400 35366 119658 35586
rect 430 35250 119658 35366
rect 400 35030 119658 35250
rect 430 34914 119658 35030
rect 400 34694 119658 34914
rect 430 34578 119658 34694
rect 400 34358 119658 34578
rect 430 34242 119570 34358
rect 400 34022 119658 34242
rect 400 33906 119570 34022
rect 400 33350 119658 33906
rect 400 33234 119570 33350
rect 400 33014 119658 33234
rect 400 32898 119570 33014
rect 400 32678 119658 32898
rect 430 32562 119658 32678
rect 400 32342 119658 32562
rect 430 32226 119570 32342
rect 400 32006 119658 32226
rect 430 31890 119658 32006
rect 400 31670 119658 31890
rect 430 31554 119658 31670
rect 400 31334 119658 31554
rect 430 31218 119570 31334
rect 400 30998 119658 31218
rect 430 30882 119570 30998
rect 400 30662 119658 30882
rect 430 30546 119570 30662
rect 400 30326 119658 30546
rect 430 30210 119658 30326
rect 400 29990 119658 30210
rect 430 29874 119570 29990
rect 400 29654 119658 29874
rect 430 29538 119658 29654
rect 400 29318 119658 29538
rect 430 29202 119658 29318
rect 400 28982 119658 29202
rect 430 28866 119658 28982
rect 400 28646 119658 28866
rect 430 28530 119570 28646
rect 400 28310 119658 28530
rect 430 28194 119658 28310
rect 400 27974 119658 28194
rect 430 27858 119658 27974
rect 400 27638 119658 27858
rect 430 27522 119658 27638
rect 400 27302 119658 27522
rect 430 27186 119570 27302
rect 400 26966 119658 27186
rect 430 26850 119658 26966
rect 400 26630 119658 26850
rect 430 26514 119658 26630
rect 400 26294 119658 26514
rect 430 26178 119570 26294
rect 400 25958 119658 26178
rect 430 25842 119570 25958
rect 400 25622 119658 25842
rect 430 25506 119570 25622
rect 400 25286 119658 25506
rect 430 25170 119658 25286
rect 400 24950 119658 25170
rect 430 24834 119658 24950
rect 400 24614 119658 24834
rect 430 24498 119570 24614
rect 400 24278 119658 24498
rect 430 24162 119570 24278
rect 400 23942 119658 24162
rect 430 23826 119658 23942
rect 400 23606 119658 23826
rect 430 23490 119658 23606
rect 400 23270 119658 23490
rect 430 23154 119658 23270
rect 400 22934 119658 23154
rect 430 22818 119658 22934
rect 400 22598 119658 22818
rect 430 22482 119658 22598
rect 400 22262 119658 22482
rect 430 22146 119658 22262
rect 400 21926 119658 22146
rect 430 21810 119658 21926
rect 400 21590 119658 21810
rect 430 21474 119658 21590
rect 400 21254 119658 21474
rect 430 21138 119658 21254
rect 400 20918 119658 21138
rect 430 20802 119658 20918
rect 400 20582 119658 20802
rect 430 20466 119658 20582
rect 400 20246 119658 20466
rect 430 20130 119658 20246
rect 400 19910 119658 20130
rect 430 19794 119658 19910
rect 400 19574 119658 19794
rect 430 19458 119658 19574
rect 400 19238 119658 19458
rect 430 19122 119658 19238
rect 400 462 119658 19122
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
rect 94384 1538 94544 98422
rect 102064 1538 102224 98422
rect 109744 1538 109904 98422
rect 117424 1538 117584 98422
<< obsm4 >>
rect 1470 1508 2194 98215
rect 2414 1508 9874 98215
rect 10094 1508 17554 98215
rect 17774 1508 25234 98215
rect 25454 1508 32914 98215
rect 33134 1508 40594 98215
rect 40814 1508 48274 98215
rect 48494 1508 55954 98215
rect 56174 1508 63634 98215
rect 63854 1508 71314 98215
rect 71534 1508 78994 98215
rect 79214 1508 86674 98215
rect 86894 1508 94354 98215
rect 94574 1508 102034 98215
rect 102254 1508 109714 98215
rect 109934 1508 117394 98215
rect 117614 1508 118762 98215
rect 1470 457 118762 1508
<< obsm5 >>
rect 1462 2093 118770 87997
<< labels >>
rlabel metal4 s 2224 1538 2384 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 103152 0 103208 400 6 cfg_cska_pinmux[0]
port 3 nsew signal input
rlabel metal2 s 103824 0 103880 400 6 cfg_cska_pinmux[1]
port 4 nsew signal input
rlabel metal2 s 104832 0 104888 400 6 cfg_cska_pinmux[2]
port 5 nsew signal input
rlabel metal2 s 104496 0 104552 400 6 cfg_cska_pinmux[3]
port 6 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 cfg_dc_trim[0]
port 7 nsew signal output
rlabel metal3 s 0 19152 400 19208 6 cfg_dc_trim[10]
port 8 nsew signal output
rlabel metal3 s 0 22512 400 22568 6 cfg_dc_trim[11]
port 9 nsew signal output
rlabel metal3 s 0 24528 400 24584 6 cfg_dc_trim[12]
port 10 nsew signal output
rlabel metal3 s 0 32256 400 32312 6 cfg_dc_trim[13]
port 11 nsew signal output
rlabel metal3 s 0 31584 400 31640 6 cfg_dc_trim[14]
port 12 nsew signal output
rlabel metal3 s 0 30240 400 30296 6 cfg_dc_trim[15]
port 13 nsew signal output
rlabel metal2 s 87696 0 87752 400 6 cfg_dc_trim[16]
port 14 nsew signal output
rlabel metal2 s 87360 0 87416 400 6 cfg_dc_trim[17]
port 15 nsew signal output
rlabel metal2 s 86352 0 86408 400 6 cfg_dc_trim[18]
port 16 nsew signal output
rlabel metal2 s 72240 0 72296 400 6 cfg_dc_trim[19]
port 17 nsew signal output
rlabel metal2 s 51408 0 51464 400 6 cfg_dc_trim[1]
port 18 nsew signal output
rlabel metal2 s 75600 0 75656 400 6 cfg_dc_trim[20]
port 19 nsew signal output
rlabel metal2 s 72576 0 72632 400 6 cfg_dc_trim[21]
port 20 nsew signal output
rlabel metal2 s 82320 0 82376 400 6 cfg_dc_trim[22]
port 21 nsew signal output
rlabel metal2 s 76608 0 76664 400 6 cfg_dc_trim[23]
port 22 nsew signal output
rlabel metal2 s 76272 0 76328 400 6 cfg_dc_trim[24]
port 23 nsew signal output
rlabel metal2 s 78624 0 78680 400 6 cfg_dc_trim[25]
port 24 nsew signal output
rlabel metal2 s 17808 0 17864 400 6 cfg_dc_trim[2]
port 25 nsew signal output
rlabel metal2 s 49392 0 49448 400 6 cfg_dc_trim[3]
port 26 nsew signal output
rlabel metal2 s 51744 0 51800 400 6 cfg_dc_trim[4]
port 27 nsew signal output
rlabel metal2 s 19152 0 19208 400 6 cfg_dc_trim[5]
port 28 nsew signal output
rlabel metal2 s 18816 0 18872 400 6 cfg_dc_trim[6]
port 29 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 cfg_dc_trim[7]
port 30 nsew signal output
rlabel metal3 s 0 24192 400 24248 6 cfg_dc_trim[8]
port 31 nsew signal output
rlabel metal3 s 0 28224 400 28280 6 cfg_dc_trim[9]
port 32 nsew signal output
rlabel metal2 s 73248 0 73304 400 6 cfg_dco_mode
port 33 nsew signal output
rlabel metal3 s 119600 37632 120000 37688 6 cfg_pll_enb
port 34 nsew signal output
rlabel metal2 s 70896 0 70952 400 6 cfg_pll_fed_div[0]
port 35 nsew signal output
rlabel metal2 s 68544 0 68600 400 6 cfg_pll_fed_div[1]
port 36 nsew signal output
rlabel metal2 s 71232 0 71288 400 6 cfg_pll_fed_div[2]
port 37 nsew signal output
rlabel metal2 s 69552 0 69608 400 6 cfg_pll_fed_div[3]
port 38 nsew signal output
rlabel metal2 s 74256 0 74312 400 6 cfg_pll_fed_div[4]
port 39 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 cfg_riscv_ctrl[0]
port 40 nsew signal output
rlabel metal2 s 22176 0 22232 400 6 cfg_riscv_ctrl[10]
port 41 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 cfg_riscv_ctrl[11]
port 42 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 cfg_riscv_ctrl[12]
port 43 nsew signal output
rlabel metal2 s 45360 0 45416 400 6 cfg_riscv_ctrl[13]
port 44 nsew signal output
rlabel metal2 s 38976 0 39032 400 6 cfg_riscv_ctrl[14]
port 45 nsew signal output
rlabel metal2 s 55104 0 55160 400 6 cfg_riscv_ctrl[15]
port 46 nsew signal output
rlabel metal2 s 22848 0 22904 400 6 cfg_riscv_ctrl[1]
port 47 nsew signal output
rlabel metal2 s 20160 0 20216 400 6 cfg_riscv_ctrl[2]
port 48 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 cfg_riscv_ctrl[3]
port 49 nsew signal output
rlabel metal2 s 20496 0 20552 400 6 cfg_riscv_ctrl[4]
port 50 nsew signal output
rlabel metal2 s 54432 0 54488 400 6 cfg_riscv_ctrl[5]
port 51 nsew signal output
rlabel metal2 s 66192 0 66248 400 6 cfg_riscv_ctrl[6]
port 52 nsew signal output
rlabel metal2 s 44016 0 44072 400 6 cfg_riscv_ctrl[7]
port 53 nsew signal output
rlabel metal2 s 43008 0 43064 400 6 cfg_riscv_ctrl[8]
port 54 nsew signal output
rlabel metal2 s 53088 0 53144 400 6 cfg_riscv_ctrl[9]
port 55 nsew signal output
rlabel metal3 s 0 34608 400 34664 6 cfg_strap_pad_ctrl
port 56 nsew signal input
rlabel metal2 s 52416 0 52472 400 6 cpu_clk
port 57 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 cpu_core_rst_n[0]
port 58 nsew signal output
rlabel metal2 s 24528 0 24584 400 6 cpu_core_rst_n[1]
port 59 nsew signal output
rlabel metal3 s 0 19488 400 19544 6 cpu_core_rst_n[2]
port 60 nsew signal output
rlabel metal3 s 0 30912 400 30968 6 cpu_core_rst_n[3]
port 61 nsew signal output
rlabel metal2 s 43344 0 43400 400 6 cpu_intf_rst_n
port 62 nsew signal output
rlabel metal2 s 25536 99600 25592 100000 6 digital_io_in[0]
port 63 nsew signal input
rlabel metal3 s 0 82656 400 82712 6 digital_io_in[10]
port 64 nsew signal input
rlabel metal3 s 0 27216 400 27272 6 digital_io_in[11]
port 65 nsew signal input
rlabel metal3 s 0 73584 400 73640 6 digital_io_in[12]
port 66 nsew signal input
rlabel metal3 s 0 45024 400 45080 6 digital_io_in[13]
port 67 nsew signal input
rlabel metal3 s 0 29568 400 29624 6 digital_io_in[14]
port 68 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 digital_io_in[15]
port 69 nsew signal input
rlabel metal3 s 0 26880 400 26936 6 digital_io_in[16]
port 70 nsew signal input
rlabel metal3 s 0 29904 400 29960 6 digital_io_in[17]
port 71 nsew signal input
rlabel metal3 s 0 41328 400 41384 6 digital_io_in[18]
port 72 nsew signal input
rlabel metal3 s 0 37968 400 38024 6 digital_io_in[19]
port 73 nsew signal input
rlabel metal3 s 0 71568 400 71624 6 digital_io_in[1]
port 74 nsew signal input
rlabel metal3 s 0 36288 400 36344 6 digital_io_in[20]
port 75 nsew signal input
rlabel metal3 s 0 56784 400 56840 6 digital_io_in[21]
port 76 nsew signal input
rlabel metal2 s 41328 99600 41384 100000 6 digital_io_in[22]
port 77 nsew signal input
rlabel metal2 s 34272 99600 34328 100000 6 digital_io_in[23]
port 78 nsew signal input
rlabel metal3 s 0 71232 400 71288 6 digital_io_in[24]
port 79 nsew signal input
rlabel metal3 s 0 70560 400 70616 6 digital_io_in[25]
port 80 nsew signal input
rlabel metal3 s 0 51072 400 51128 6 digital_io_in[26]
port 81 nsew signal input
rlabel metal3 s 0 42336 400 42392 6 digital_io_in[27]
port 82 nsew signal input
rlabel metal2 s 0 0 56 400 6 digital_io_in[28]
port 83 nsew signal input
rlabel metal3 s 0 25200 400 25256 6 digital_io_in[29]
port 84 nsew signal input
rlabel metal3 s 0 71904 400 71960 6 digital_io_in[2]
port 85 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 digital_io_in[30]
port 86 nsew signal input
rlabel metal2 s 25536 0 25592 400 6 digital_io_in[31]
port 87 nsew signal input
rlabel metal2 s 29904 0 29960 400 6 digital_io_in[32]
port 88 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 digital_io_in[33]
port 89 nsew signal input
rlabel metal3 s 0 20832 400 20888 6 digital_io_in[34]
port 90 nsew signal input
rlabel metal3 s 0 21504 400 21560 6 digital_io_in[35]
port 91 nsew signal input
rlabel metal3 s 0 20160 400 20216 6 digital_io_in[36]
port 92 nsew signal input
rlabel metal2 s 336 0 392 400 6 digital_io_in[37]
port 93 nsew signal input
rlabel metal3 s 0 72576 400 72632 6 digital_io_in[3]
port 94 nsew signal input
rlabel metal3 s 0 76944 400 77000 6 digital_io_in[4]
port 95 nsew signal input
rlabel metal3 s 0 46704 400 46760 6 digital_io_in[5]
port 96 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 digital_io_in[6]
port 97 nsew signal input
rlabel metal3 s 0 60816 400 60872 6 digital_io_in[7]
port 98 nsew signal input
rlabel metal3 s 0 47040 400 47096 6 digital_io_in[8]
port 99 nsew signal input
rlabel metal3 s 0 63504 400 63560 6 digital_io_in[9]
port 100 nsew signal input
rlabel metal3 s 0 77280 400 77336 6 digital_io_oen[0]
port 101 nsew signal output
rlabel metal3 s 0 54768 400 54824 6 digital_io_oen[10]
port 102 nsew signal output
rlabel metal3 s 0 61152 400 61208 6 digital_io_oen[11]
port 103 nsew signal output
rlabel metal3 s 0 60480 400 60536 6 digital_io_oen[12]
port 104 nsew signal output
rlabel metal2 s 23856 0 23912 400 6 digital_io_oen[13]
port 105 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 digital_io_oen[14]
port 106 nsew signal output
rlabel metal2 s 40656 0 40712 400 6 digital_io_oen[15]
port 107 nsew signal output
rlabel metal3 s 0 55104 400 55160 6 digital_io_oen[16]
port 108 nsew signal output
rlabel metal3 s 0 34944 400 35000 6 digital_io_oen[17]
port 109 nsew signal output
rlabel metal3 s 0 35952 400 36008 6 digital_io_oen[18]
port 110 nsew signal output
rlabel metal3 s 0 39312 400 39368 6 digital_io_oen[19]
port 111 nsew signal output
rlabel metal3 s 0 74592 400 74648 6 digital_io_oen[1]
port 112 nsew signal output
rlabel metal3 s 0 56112 400 56168 6 digital_io_oen[20]
port 113 nsew signal output
rlabel metal3 s 0 81312 400 81368 6 digital_io_oen[21]
port 114 nsew signal output
rlabel metal3 s 0 68880 400 68936 6 digital_io_oen[22]
port 115 nsew signal output
rlabel metal3 s 0 69216 400 69272 6 digital_io_oen[23]
port 116 nsew signal output
rlabel metal3 s 0 75936 400 75992 6 digital_io_oen[24]
port 117 nsew signal output
rlabel metal3 s 0 78960 400 79016 6 digital_io_oen[25]
port 118 nsew signal output
rlabel metal3 s 0 59472 400 59528 6 digital_io_oen[26]
port 119 nsew signal output
rlabel metal3 s 0 48720 400 48776 6 digital_io_oen[27]
port 120 nsew signal output
rlabel metal3 s 0 40656 400 40712 6 digital_io_oen[28]
port 121 nsew signal output
rlabel metal3 s 0 40992 400 41048 6 digital_io_oen[29]
port 122 nsew signal output
rlabel metal3 s 0 64848 400 64904 6 digital_io_oen[2]
port 123 nsew signal output
rlabel metal3 s 0 48384 400 48440 6 digital_io_oen[30]
port 124 nsew signal output
rlabel metal3 s 0 45696 400 45752 6 digital_io_oen[31]
port 125 nsew signal output
rlabel metal3 s 0 43680 400 43736 6 digital_io_oen[32]
port 126 nsew signal output
rlabel metal3 s 0 44352 400 44408 6 digital_io_oen[33]
port 127 nsew signal output
rlabel metal3 s 0 38640 400 38696 6 digital_io_oen[34]
port 128 nsew signal output
rlabel metal3 s 0 38304 400 38360 6 digital_io_oen[35]
port 129 nsew signal output
rlabel metal3 s 0 44688 400 44744 6 digital_io_oen[36]
port 130 nsew signal output
rlabel metal3 s 0 47712 400 47768 6 digital_io_oen[37]
port 131 nsew signal output
rlabel metal3 s 0 77616 400 77672 6 digital_io_oen[3]
port 132 nsew signal output
rlabel metal3 s 0 72912 400 72968 6 digital_io_oen[4]
port 133 nsew signal output
rlabel metal3 s 0 58128 400 58184 6 digital_io_oen[5]
port 134 nsew signal output
rlabel metal3 s 0 50736 400 50792 6 digital_io_oen[6]
port 135 nsew signal output
rlabel metal2 s 46704 0 46760 400 6 digital_io_oen[7]
port 136 nsew signal output
rlabel metal2 s 48384 0 48440 400 6 digital_io_oen[8]
port 137 nsew signal output
rlabel metal2 s 20832 0 20888 400 6 digital_io_oen[9]
port 138 nsew signal output
rlabel metal3 s 0 79968 400 80024 6 digital_io_out[0]
port 139 nsew signal output
rlabel metal3 s 0 45360 400 45416 6 digital_io_out[10]
port 140 nsew signal output
rlabel metal3 s 0 58800 400 58856 6 digital_io_out[11]
port 141 nsew signal output
rlabel metal3 s 0 59808 400 59864 6 digital_io_out[12]
port 142 nsew signal output
rlabel metal2 s 32592 0 32648 400 6 digital_io_out[13]
port 143 nsew signal output
rlabel metal2 s 37296 0 37352 400 6 digital_io_out[14]
port 144 nsew signal output
rlabel metal2 s 21840 0 21896 400 6 digital_io_out[15]
port 145 nsew signal output
rlabel metal3 s 0 53424 400 53480 6 digital_io_out[16]
port 146 nsew signal output
rlabel metal3 s 0 50400 400 50456 6 digital_io_out[17]
port 147 nsew signal output
rlabel metal3 s 0 42000 400 42056 6 digital_io_out[18]
port 148 nsew signal output
rlabel metal3 s 0 43008 400 43064 6 digital_io_out[19]
port 149 nsew signal output
rlabel metal3 s 0 76272 400 76328 6 digital_io_out[1]
port 150 nsew signal output
rlabel metal3 s 0 53088 400 53144 6 digital_io_out[20]
port 151 nsew signal output
rlabel metal3 s 0 59136 400 59192 6 digital_io_out[21]
port 152 nsew signal output
rlabel metal3 s 0 68544 400 68600 6 digital_io_out[22]
port 153 nsew signal output
rlabel metal3 s 0 67536 400 67592 6 digital_io_out[23]
port 154 nsew signal output
rlabel metal3 s 0 75264 400 75320 6 digital_io_out[24]
port 155 nsew signal output
rlabel metal3 s 0 79296 400 79352 6 digital_io_out[25]
port 156 nsew signal output
rlabel metal3 s 0 80640 400 80696 6 digital_io_out[26]
port 157 nsew signal output
rlabel metal3 s 0 57792 400 57848 6 digital_io_out[27]
port 158 nsew signal output
rlabel metal2 s 89376 99600 89432 100000 6 digital_io_out[28]
port 159 nsew signal output
rlabel metal2 s 64848 0 64904 400 6 digital_io_out[29]
port 160 nsew signal output
rlabel metal3 s 0 66192 400 66248 6 digital_io_out[2]
port 161 nsew signal output
rlabel metal3 s 119600 93408 120000 93464 6 digital_io_out[30]
port 162 nsew signal output
rlabel metal2 s 99120 99600 99176 100000 6 digital_io_out[31]
port 163 nsew signal output
rlabel metal2 s 102480 0 102536 400 6 digital_io_out[32]
port 164 nsew signal output
rlabel metal3 s 119600 95424 120000 95480 6 digital_io_out[33]
port 165 nsew signal output
rlabel metal2 s 100464 99600 100520 100000 6 digital_io_out[34]
port 166 nsew signal output
rlabel metal3 s 119600 90048 120000 90104 6 digital_io_out[35]
port 167 nsew signal output
rlabel metal2 s 87024 0 87080 400 6 digital_io_out[36]
port 168 nsew signal output
rlabel metal2 s 75936 0 75992 400 6 digital_io_out[37]
port 169 nsew signal output
rlabel metal3 s 0 78624 400 78680 6 digital_io_out[3]
port 170 nsew signal output
rlabel metal3 s 0 67872 400 67928 6 digital_io_out[4]
port 171 nsew signal output
rlabel metal3 s 0 38976 400 39032 6 digital_io_out[5]
port 172 nsew signal output
rlabel metal3 s 0 49392 400 49448 6 digital_io_out[6]
port 173 nsew signal output
rlabel metal2 s 16800 0 16856 400 6 digital_io_out[7]
port 174 nsew signal output
rlabel metal3 s 0 39648 400 39704 6 digital_io_out[8]
port 175 nsew signal output
rlabel metal3 s 0 46368 400 46424 6 digital_io_out[9]
port 176 nsew signal output
rlabel metal2 s 17136 0 17192 400 6 e_reset_n
port 177 nsew signal input
rlabel metal3 s 0 47376 400 47432 6 i2cm_clk_i
port 178 nsew signal output
rlabel metal3 s 0 56448 400 56504 6 i2cm_clk_o
port 179 nsew signal input
rlabel metal3 s 0 46032 400 46088 6 i2cm_clk_oen
port 180 nsew signal input
rlabel metal3 s 0 40320 400 40376 6 i2cm_data_i
port 181 nsew signal output
rlabel metal3 s 0 80304 400 80360 6 i2cm_data_o
port 182 nsew signal input
rlabel metal3 s 0 80976 400 81032 6 i2cm_data_oen
port 183 nsew signal input
rlabel metal2 s 50064 0 50120 400 6 i2cm_intr
port 184 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 i2cm_rst_n
port 185 nsew signal output
rlabel metal2 s 49056 0 49112 400 6 int_pll_clock
port 186 nsew signal input
rlabel metal2 s 45024 0 45080 400 6 ir_intr
port 187 nsew signal input
rlabel metal3 s 0 69888 400 69944 6 ir_rx
port 188 nsew signal output
rlabel metal2 s 21504 0 21560 400 6 ir_tx
port 189 nsew signal input
rlabel metal2 s 48048 0 48104 400 6 irq_lines[0]
port 190 nsew signal output
rlabel metal3 s 0 41664 400 41720 6 irq_lines[10]
port 191 nsew signal output
rlabel metal3 s 0 23520 400 23576 6 irq_lines[11]
port 192 nsew signal output
rlabel metal3 s 0 30576 400 30632 6 irq_lines[12]
port 193 nsew signal output
rlabel metal3 s 0 26208 400 26264 6 irq_lines[13]
port 194 nsew signal output
rlabel metal3 s 0 31248 400 31304 6 irq_lines[14]
port 195 nsew signal output
rlabel metal3 s 0 39984 400 40040 6 irq_lines[15]
port 196 nsew signal output
rlabel metal3 s 119600 29904 120000 29960 6 irq_lines[16]
port 197 nsew signal output
rlabel metal3 s 119600 30576 120000 30632 6 irq_lines[17]
port 198 nsew signal output
rlabel metal3 s 119600 34272 120000 34328 6 irq_lines[18]
port 199 nsew signal output
rlabel metal2 s 68208 0 68264 400 6 irq_lines[19]
port 200 nsew signal output
rlabel metal2 s 59136 0 59192 400 6 irq_lines[1]
port 201 nsew signal output
rlabel metal3 s 119600 33264 120000 33320 6 irq_lines[20]
port 202 nsew signal output
rlabel metal2 s 70224 0 70280 400 6 irq_lines[21]
port 203 nsew signal output
rlabel metal2 s 71568 0 71624 400 6 irq_lines[22]
port 204 nsew signal output
rlabel metal3 s 119600 33936 120000 33992 6 irq_lines[23]
port 205 nsew signal output
rlabel metal2 s 71904 0 71960 400 6 irq_lines[24]
port 206 nsew signal output
rlabel metal2 s 57120 0 57176 400 6 irq_lines[25]
port 207 nsew signal output
rlabel metal2 s 67536 0 67592 400 6 irq_lines[26]
port 208 nsew signal output
rlabel metal2 s 58464 0 58520 400 6 irq_lines[27]
port 209 nsew signal output
rlabel metal2 s 63168 0 63224 400 6 irq_lines[28]
port 210 nsew signal output
rlabel metal2 s 61488 0 61544 400 6 irq_lines[29]
port 211 nsew signal output
rlabel metal2 s 60144 0 60200 400 6 irq_lines[2]
port 212 nsew signal output
rlabel metal2 s 63840 0 63896 400 6 irq_lines[30]
port 213 nsew signal output
rlabel metal2 s 56784 0 56840 400 6 irq_lines[31]
port 214 nsew signal output
rlabel metal2 s 55440 0 55496 400 6 irq_lines[3]
port 215 nsew signal output
rlabel metal2 s 52752 0 52808 400 6 irq_lines[4]
port 216 nsew signal output
rlabel metal2 s 55776 0 55832 400 6 irq_lines[5]
port 217 nsew signal output
rlabel metal2 s 47376 0 47432 400 6 irq_lines[6]
port 218 nsew signal output
rlabel metal2 s 47040 0 47096 400 6 irq_lines[7]
port 219 nsew signal output
rlabel metal3 s 0 27888 400 27944 6 irq_lines[8]
port 220 nsew signal output
rlabel metal3 s 0 25872 400 25928 6 irq_lines[9]
port 221 nsew signal output
rlabel metal3 s 0 97776 400 97832 6 mclk
port 222 nsew signal input
rlabel metal2 s 75264 0 75320 400 6 p_reset_n
port 223 nsew signal input
rlabel metal2 s 100800 99600 100856 100000 6 pinmux_debug[0]
port 224 nsew signal output
rlabel metal3 s 119600 95760 120000 95816 6 pinmux_debug[10]
port 225 nsew signal output
rlabel metal2 s 88032 99600 88088 100000 6 pinmux_debug[11]
port 226 nsew signal output
rlabel metal2 s 93072 99600 93128 100000 6 pinmux_debug[12]
port 227 nsew signal output
rlabel metal2 s 88368 99600 88424 100000 6 pinmux_debug[13]
port 228 nsew signal output
rlabel metal2 s 90720 0 90776 400 6 pinmux_debug[14]
port 229 nsew signal output
rlabel metal3 s 119600 97776 120000 97832 6 pinmux_debug[15]
port 230 nsew signal output
rlabel metal2 s 61152 0 61208 400 6 pinmux_debug[16]
port 231 nsew signal output
rlabel metal2 s 85008 99600 85064 100000 6 pinmux_debug[17]
port 232 nsew signal output
rlabel metal2 s 49056 99600 49112 100000 6 pinmux_debug[18]
port 233 nsew signal output
rlabel metal2 s 105504 99600 105560 100000 6 pinmux_debug[19]
port 234 nsew signal output
rlabel metal2 s 101136 99600 101192 100000 6 pinmux_debug[1]
port 235 nsew signal output
rlabel metal2 s 85008 0 85064 400 6 pinmux_debug[20]
port 236 nsew signal output
rlabel metal2 s 72912 0 72968 400 6 pinmux_debug[21]
port 237 nsew signal output
rlabel metal3 s 119600 94752 120000 94808 6 pinmux_debug[22]
port 238 nsew signal output
rlabel metal2 s 62496 0 62552 400 6 pinmux_debug[23]
port 239 nsew signal output
rlabel metal3 s 119600 98112 120000 98168 6 pinmux_debug[24]
port 240 nsew signal output
rlabel metal2 s 62160 0 62216 400 6 pinmux_debug[25]
port 241 nsew signal output
rlabel metal2 s 99792 99600 99848 100000 6 pinmux_debug[26]
port 242 nsew signal output
rlabel metal2 s 53424 0 53480 400 6 pinmux_debug[27]
port 243 nsew signal output
rlabel metal2 s 83328 99600 83384 100000 6 pinmux_debug[28]
port 244 nsew signal output
rlabel metal2 s 95424 0 95480 400 6 pinmux_debug[29]
port 245 nsew signal output
rlabel metal2 s 113904 0 113960 400 6 pinmux_debug[2]
port 246 nsew signal output
rlabel metal2 s 110208 0 110264 400 6 pinmux_debug[30]
port 247 nsew signal output
rlabel metal3 s 119600 82992 120000 83048 6 pinmux_debug[31]
port 248 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 pinmux_debug[3]
port 249 nsew signal output
rlabel metal3 s 119600 83328 120000 83384 6 pinmux_debug[4]
port 250 nsew signal output
rlabel metal2 s 103824 99600 103880 100000 6 pinmux_debug[5]
port 251 nsew signal output
rlabel metal3 s 119600 97440 120000 97496 6 pinmux_debug[6]
port 252 nsew signal output
rlabel metal2 s 51072 0 51128 400 6 pinmux_debug[7]
port 253 nsew signal output
rlabel metal2 s 89040 99600 89096 100000 6 pinmux_debug[8]
port 254 nsew signal output
rlabel metal2 s 112560 0 112616 400 6 pinmux_debug[9]
port 255 nsew signal output
rlabel metal3 s 119600 38304 120000 38360 6 pll_ref_clk
port 256 nsew signal output
rlabel metal2 s 53424 99600 53480 100000 6 pulse1m_mclk
port 257 nsew signal output
rlabel metal2 s 35616 0 35672 400 6 qspim_rst_n
port 258 nsew signal output
rlabel metal3 s 0 61488 400 61544 6 reg_ack
port 259 nsew signal output
rlabel metal2 s 90048 0 90104 400 6 reg_addr[0]
port 260 nsew signal input
rlabel metal2 s 69888 99600 69944 100000 6 reg_addr[10]
port 261 nsew signal input
rlabel metal2 s 84672 0 84728 400 6 reg_addr[1]
port 262 nsew signal input
rlabel metal2 s 90384 99600 90440 100000 6 reg_addr[2]
port 263 nsew signal input
rlabel metal2 s 93408 99600 93464 100000 6 reg_addr[3]
port 264 nsew signal input
rlabel metal2 s 82992 99600 83048 100000 6 reg_addr[4]
port 265 nsew signal input
rlabel metal2 s 82656 99600 82712 100000 6 reg_addr[5]
port 266 nsew signal input
rlabel metal3 s 119600 31248 120000 31304 6 reg_addr[6]
port 267 nsew signal input
rlabel metal2 s 67200 99600 67256 100000 6 reg_addr[7]
port 268 nsew signal input
rlabel metal2 s 67872 99600 67928 100000 6 reg_addr[8]
port 269 nsew signal input
rlabel metal2 s 67536 99600 67592 100000 6 reg_addr[9]
port 270 nsew signal input
rlabel metal3 s 119600 25872 120000 25928 6 reg_be[0]
port 271 nsew signal input
rlabel metal2 s 98784 99600 98840 100000 6 reg_be[1]
port 272 nsew signal input
rlabel metal2 s 88032 0 88088 400 6 reg_be[2]
port 273 nsew signal input
rlabel metal2 s 33600 0 33656 400 6 reg_be[3]
port 274 nsew signal input
rlabel metal2 s 68208 99600 68264 100000 6 reg_cs
port 275 nsew signal input
rlabel metal2 s 68880 99600 68936 100000 6 reg_peri_ack
port 276 nsew signal input
rlabel metal2 s 90384 0 90440 400 6 reg_peri_addr[0]
port 277 nsew signal output
rlabel metal2 s 65520 99600 65576 100000 6 reg_peri_addr[10]
port 278 nsew signal output
rlabel metal2 s 82656 0 82712 400 6 reg_peri_addr[1]
port 279 nsew signal output
rlabel metal3 s 119600 32928 120000 32984 6 reg_peri_addr[2]
port 280 nsew signal output
rlabel metal2 s 79968 0 80024 400 6 reg_peri_addr[3]
port 281 nsew signal output
rlabel metal3 s 119600 32256 120000 32312 6 reg_peri_addr[4]
port 282 nsew signal output
rlabel metal2 s 83328 0 83384 400 6 reg_peri_addr[5]
port 283 nsew signal output
rlabel metal2 s 66864 99600 66920 100000 6 reg_peri_addr[6]
port 284 nsew signal output
rlabel metal2 s 65184 99600 65240 100000 6 reg_peri_addr[7]
port 285 nsew signal output
rlabel metal2 s 64512 99600 64568 100000 6 reg_peri_addr[8]
port 286 nsew signal output
rlabel metal2 s 65856 99600 65912 100000 6 reg_peri_addr[9]
port 287 nsew signal output
rlabel metal2 s 81984 0 82040 400 6 reg_peri_be[0]
port 288 nsew signal output
rlabel metal2 s 80304 0 80360 400 6 reg_peri_be[1]
port 289 nsew signal output
rlabel metal2 s 85344 0 85400 400 6 reg_peri_be[2]
port 290 nsew signal output
rlabel metal3 s 119600 45696 120000 45752 6 reg_peri_be[3]
port 291 nsew signal output
rlabel metal2 s 66528 99600 66584 100000 6 reg_peri_cs
port 292 nsew signal output
rlabel metal2 s 53760 99600 53816 100000 6 reg_peri_rdata[0]
port 293 nsew signal input
rlabel metal2 s 55440 99600 55496 100000 6 reg_peri_rdata[10]
port 294 nsew signal input
rlabel metal2 s 59808 99600 59864 100000 6 reg_peri_rdata[11]
port 295 nsew signal input
rlabel metal2 s 60816 99600 60872 100000 6 reg_peri_rdata[12]
port 296 nsew signal input
rlabel metal2 s 58128 99600 58184 100000 6 reg_peri_rdata[13]
port 297 nsew signal input
rlabel metal2 s 63168 99600 63224 100000 6 reg_peri_rdata[14]
port 298 nsew signal input
rlabel metal2 s 60144 99600 60200 100000 6 reg_peri_rdata[15]
port 299 nsew signal input
rlabel metal2 s 64848 99600 64904 100000 6 reg_peri_rdata[16]
port 300 nsew signal input
rlabel metal2 s 64176 99600 64232 100000 6 reg_peri_rdata[17]
port 301 nsew signal input
rlabel metal2 s 62160 99600 62216 100000 6 reg_peri_rdata[18]
port 302 nsew signal input
rlabel metal2 s 58464 99600 58520 100000 6 reg_peri_rdata[19]
port 303 nsew signal input
rlabel metal2 s 55776 99600 55832 100000 6 reg_peri_rdata[1]
port 304 nsew signal input
rlabel metal3 s 0 72240 400 72296 6 reg_peri_rdata[20]
port 305 nsew signal input
rlabel metal2 s 60480 99600 60536 100000 6 reg_peri_rdata[21]
port 306 nsew signal input
rlabel metal3 s 0 73248 400 73304 6 reg_peri_rdata[22]
port 307 nsew signal input
rlabel metal3 s 0 75600 400 75656 6 reg_peri_rdata[23]
port 308 nsew signal input
rlabel metal2 s 54768 99600 54824 100000 6 reg_peri_rdata[24]
port 309 nsew signal input
rlabel metal3 s 0 35616 400 35672 6 reg_peri_rdata[25]
port 310 nsew signal input
rlabel metal2 s 63840 99600 63896 100000 6 reg_peri_rdata[26]
port 311 nsew signal input
rlabel metal3 s 0 36624 400 36680 6 reg_peri_rdata[27]
port 312 nsew signal input
rlabel metal3 s 0 60144 400 60200 6 reg_peri_rdata[28]
port 313 nsew signal input
rlabel metal2 s 69216 99600 69272 100000 6 reg_peri_rdata[29]
port 314 nsew signal input
rlabel metal2 s 57792 99600 57848 100000 6 reg_peri_rdata[2]
port 315 nsew signal input
rlabel metal2 s 54432 99600 54488 100000 6 reg_peri_rdata[30]
port 316 nsew signal input
rlabel metal3 s 0 35280 400 35336 6 reg_peri_rdata[31]
port 317 nsew signal input
rlabel metal2 s 55104 99600 55160 100000 6 reg_peri_rdata[3]
port 318 nsew signal input
rlabel metal2 s 57120 99600 57176 100000 6 reg_peri_rdata[4]
port 319 nsew signal input
rlabel metal2 s 57456 99600 57512 100000 6 reg_peri_rdata[5]
port 320 nsew signal input
rlabel metal2 s 56784 99600 56840 100000 6 reg_peri_rdata[6]
port 321 nsew signal input
rlabel metal2 s 54096 99600 54152 100000 6 reg_peri_rdata[7]
port 322 nsew signal input
rlabel metal2 s 58800 99600 58856 100000 6 reg_peri_rdata[8]
port 323 nsew signal input
rlabel metal2 s 56112 99600 56168 100000 6 reg_peri_rdata[9]
port 324 nsew signal input
rlabel metal2 s 66192 99600 66248 100000 6 reg_peri_wdata[0]
port 325 nsew signal output
rlabel metal2 s 81312 0 81368 400 6 reg_peri_wdata[10]
port 326 nsew signal output
rlabel metal2 s 80976 0 81032 400 6 reg_peri_wdata[11]
port 327 nsew signal output
rlabel metal2 s 79632 0 79688 400 6 reg_peri_wdata[12]
port 328 nsew signal output
rlabel metal2 s 81648 0 81704 400 6 reg_peri_wdata[13]
port 329 nsew signal output
rlabel metal2 s 86016 0 86072 400 6 reg_peri_wdata[14]
port 330 nsew signal output
rlabel metal2 s 84000 0 84056 400 6 reg_peri_wdata[15]
port 331 nsew signal output
rlabel metal2 s 80640 0 80696 400 6 reg_peri_wdata[16]
port 332 nsew signal output
rlabel metal2 s 83664 0 83720 400 6 reg_peri_wdata[17]
port 333 nsew signal output
rlabel metal2 s 82992 0 83048 400 6 reg_peri_wdata[18]
port 334 nsew signal output
rlabel metal2 s 78288 0 78344 400 6 reg_peri_wdata[19]
port 335 nsew signal output
rlabel metal3 s 119600 81312 120000 81368 6 reg_peri_wdata[1]
port 336 nsew signal output
rlabel metal2 s 73920 0 73976 400 6 reg_peri_wdata[20]
port 337 nsew signal output
rlabel metal2 s 77952 0 78008 400 6 reg_peri_wdata[21]
port 338 nsew signal output
rlabel metal2 s 77280 0 77336 400 6 reg_peri_wdata[22]
port 339 nsew signal output
rlabel metal2 s 74592 0 74648 400 6 reg_peri_wdata[23]
port 340 nsew signal output
rlabel metal2 s 74928 0 74984 400 6 reg_peri_wdata[24]
port 341 nsew signal output
rlabel metal2 s 73584 0 73640 400 6 reg_peri_wdata[25]
port 342 nsew signal output
rlabel metal2 s 65856 0 65912 400 6 reg_peri_wdata[26]
port 343 nsew signal output
rlabel metal2 s 76944 0 77000 400 6 reg_peri_wdata[27]
port 344 nsew signal output
rlabel metal2 s 67872 0 67928 400 6 reg_peri_wdata[28]
port 345 nsew signal output
rlabel metal2 s 85680 0 85736 400 6 reg_peri_wdata[29]
port 346 nsew signal output
rlabel metal3 s 119600 81648 120000 81704 6 reg_peri_wdata[2]
port 347 nsew signal output
rlabel metal2 s 78960 0 79016 400 6 reg_peri_wdata[30]
port 348 nsew signal output
rlabel metal2 s 77616 0 77672 400 6 reg_peri_wdata[31]
port 349 nsew signal output
rlabel metal3 s 119600 87696 120000 87752 6 reg_peri_wdata[3]
port 350 nsew signal output
rlabel metal2 s 61488 99600 61544 100000 6 reg_peri_wdata[4]
port 351 nsew signal output
rlabel metal3 s 119600 89376 120000 89432 6 reg_peri_wdata[5]
port 352 nsew signal output
rlabel metal3 s 119600 30912 120000 30968 6 reg_peri_wdata[6]
port 353 nsew signal output
rlabel metal3 s 119600 39312 120000 39368 6 reg_peri_wdata[7]
port 354 nsew signal output
rlabel metal2 s 80640 99600 80696 100000 6 reg_peri_wdata[8]
port 355 nsew signal output
rlabel metal2 s 79296 0 79352 400 6 reg_peri_wdata[9]
port 356 nsew signal output
rlabel metal2 s 84336 0 84392 400 6 reg_peri_wr
port 357 nsew signal output
rlabel metal3 s 0 64512 400 64568 6 reg_rdata[0]
port 358 nsew signal output
rlabel metal3 s 0 54096 400 54152 6 reg_rdata[10]
port 359 nsew signal output
rlabel metal3 s 0 55440 400 55496 6 reg_rdata[11]
port 360 nsew signal output
rlabel metal3 s 0 57456 400 57512 6 reg_rdata[12]
port 361 nsew signal output
rlabel metal3 s 0 62832 400 62888 6 reg_rdata[13]
port 362 nsew signal output
rlabel metal3 s 0 58464 400 58520 6 reg_rdata[14]
port 363 nsew signal output
rlabel metal3 s 0 62160 400 62216 6 reg_rdata[15]
port 364 nsew signal output
rlabel metal2 s 63504 99600 63560 100000 6 reg_rdata[16]
port 365 nsew signal output
rlabel metal2 s 68544 99600 68600 100000 6 reg_rdata[17]
port 366 nsew signal output
rlabel metal2 s 61824 99600 61880 100000 6 reg_rdata[18]
port 367 nsew signal output
rlabel metal3 s 0 74928 400 74984 6 reg_rdata[19]
port 368 nsew signal output
rlabel metal2 s 69552 99600 69608 100000 6 reg_rdata[1]
port 369 nsew signal output
rlabel metal3 s 0 61824 400 61880 6 reg_rdata[20]
port 370 nsew signal output
rlabel metal2 s 59472 99600 59528 100000 6 reg_rdata[21]
port 371 nsew signal output
rlabel metal3 s 0 81984 400 82040 6 reg_rdata[22]
port 372 nsew signal output
rlabel metal3 s 0 62496 400 62552 6 reg_rdata[23]
port 373 nsew signal output
rlabel metal2 s 61152 99600 61208 100000 6 reg_rdata[24]
port 374 nsew signal output
rlabel metal3 s 0 49728 400 49784 6 reg_rdata[25]
port 375 nsew signal output
rlabel metal2 s 62832 99600 62888 100000 6 reg_rdata[26]
port 376 nsew signal output
rlabel metal3 s 0 54432 400 54488 6 reg_rdata[27]
port 377 nsew signal output
rlabel metal3 s 0 81648 400 81704 6 reg_rdata[28]
port 378 nsew signal output
rlabel metal2 s 59136 99600 59192 100000 6 reg_rdata[29]
port 379 nsew signal output
rlabel metal2 s 62496 99600 62552 100000 6 reg_rdata[2]
port 380 nsew signal output
rlabel metal2 s 56448 99600 56504 100000 6 reg_rdata[30]
port 381 nsew signal output
rlabel metal3 s 0 52080 400 52136 6 reg_rdata[31]
port 382 nsew signal output
rlabel metal3 s 0 77952 400 78008 6 reg_rdata[3]
port 383 nsew signal output
rlabel metal3 s 0 74256 400 74312 6 reg_rdata[4]
port 384 nsew signal output
rlabel metal3 s 0 65520 400 65576 6 reg_rdata[5]
port 385 nsew signal output
rlabel metal3 s 0 65856 400 65912 6 reg_rdata[6]
port 386 nsew signal output
rlabel metal3 s 0 65184 400 65240 6 reg_rdata[7]
port 387 nsew signal output
rlabel metal3 s 0 51408 400 51464 6 reg_rdata[8]
port 388 nsew signal output
rlabel metal3 s 0 37632 400 37688 6 reg_rdata[9]
port 389 nsew signal output
rlabel metal3 s 119600 26208 120000 26264 6 reg_wdata[0]
port 390 nsew signal input
rlabel metal2 s 106176 99600 106232 100000 6 reg_wdata[10]
port 391 nsew signal input
rlabel metal2 s 98448 99600 98504 100000 6 reg_wdata[11]
port 392 nsew signal input
rlabel metal3 s 0 87360 400 87416 6 reg_wdata[12]
port 393 nsew signal input
rlabel metal3 s 0 86352 400 86408 6 reg_wdata[13]
port 394 nsew signal input
rlabel metal3 s 0 34272 400 34328 6 reg_wdata[14]
port 395 nsew signal input
rlabel metal3 s 0 84336 400 84392 6 reg_wdata[15]
port 396 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 reg_wdata[16]
port 397 nsew signal input
rlabel metal2 s 24192 0 24248 400 6 reg_wdata[17]
port 398 nsew signal input
rlabel metal2 s 25872 0 25928 400 6 reg_wdata[18]
port 399 nsew signal input
rlabel metal2 s 28224 0 28280 400 6 reg_wdata[19]
port 400 nsew signal input
rlabel metal3 s 119600 24528 120000 24584 6 reg_wdata[1]
port 401 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 reg_wdata[20]
port 402 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 reg_wdata[21]
port 403 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 reg_wdata[22]
port 404 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 reg_wdata[23]
port 405 nsew signal input
rlabel metal2 s 66864 0 66920 400 6 reg_wdata[24]
port 406 nsew signal input
rlabel metal2 s 66528 0 66584 400 6 reg_wdata[25]
port 407 nsew signal input
rlabel metal2 s 14784 0 14840 400 6 reg_wdata[26]
port 408 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 reg_wdata[27]
port 409 nsew signal input
rlabel metal2 s 34944 0 35000 400 6 reg_wdata[28]
port 410 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 reg_wdata[29]
port 411 nsew signal input
rlabel metal3 s 119600 28560 120000 28616 6 reg_wdata[2]
port 412 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 reg_wdata[30]
port 413 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 reg_wdata[31]
port 414 nsew signal input
rlabel metal3 s 119600 24192 120000 24248 6 reg_wdata[3]
port 415 nsew signal input
rlabel metal3 s 119600 27216 120000 27272 6 reg_wdata[4]
port 416 nsew signal input
rlabel metal3 s 119600 25536 120000 25592 6 reg_wdata[5]
port 417 nsew signal input
rlabel metal2 s 111552 99600 111608 100000 6 reg_wdata[6]
port 418 nsew signal input
rlabel metal2 s 107184 99600 107240 100000 6 reg_wdata[7]
port 419 nsew signal input
rlabel metal2 s 106848 99600 106904 100000 6 reg_wdata[8]
port 420 nsew signal input
rlabel metal2 s 101472 99600 101528 100000 6 reg_wdata[9]
port 421 nsew signal input
rlabel metal2 s 87696 99600 87752 100000 6 reg_wr
port 422 nsew signal input
rlabel metal3 s 0 70896 400 70952 6 riscv_tck
port 423 nsew signal output
rlabel metal3 s 0 66864 400 66920 6 riscv_tdi
port 424 nsew signal output
rlabel metal3 s 0 67200 400 67256 6 riscv_tdo
port 425 nsew signal input
rlabel metal3 s 0 66528 400 66584 6 riscv_tdo_en
port 426 nsew signal input
rlabel metal3 s 0 68208 400 68264 6 riscv_tms
port 427 nsew signal output
rlabel metal2 s 26208 99600 26264 100000 6 riscv_trst_n
port 428 nsew signal output
rlabel metal2 s 64512 0 64568 400 6 rtc_clk
port 429 nsew signal output
rlabel metal2 s 18144 0 18200 400 6 rtc_intr
port 430 nsew signal input
rlabel metal2 s 69216 0 69272 400 6 s_reset_n
port 431 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 sflash_di[0]
port 432 nsew signal output
rlabel metal3 s 0 21168 400 21224 6 sflash_di[1]
port 433 nsew signal output
rlabel metal3 s 0 21840 400 21896 6 sflash_di[2]
port 434 nsew signal output
rlabel metal3 s 0 20496 400 20552 6 sflash_di[3]
port 435 nsew signal output
rlabel metal3 s 119600 95088 120000 95144 6 sflash_do[0]
port 436 nsew signal input
rlabel metal2 s 100128 99600 100184 100000 6 sflash_do[1]
port 437 nsew signal input
rlabel metal3 s 119600 89712 120000 89768 6 sflash_do[2]
port 438 nsew signal input
rlabel metal2 s 86688 0 86744 400 6 sflash_do[3]
port 439 nsew signal input
rlabel metal3 s 0 43344 400 43400 6 sflash_oen[0]
port 440 nsew signal input
rlabel metal3 s 0 37296 400 37352 6 sflash_oen[1]
port 441 nsew signal input
rlabel metal3 s 0 48048 400 48104 6 sflash_oen[2]
port 442 nsew signal input
rlabel metal3 s 0 42672 400 42728 6 sflash_oen[3]
port 443 nsew signal input
rlabel metal2 s 88704 99600 88760 100000 6 sflash_sck
port 444 nsew signal input
rlabel metal2 s 65184 0 65240 400 6 sflash_ss[0]
port 445 nsew signal input
rlabel metal3 s 119600 93072 120000 93128 6 sflash_ss[1]
port 446 nsew signal input
rlabel metal2 s 99456 99600 99512 100000 6 sflash_ss[2]
port 447 nsew signal input
rlabel metal2 s 102144 0 102200 400 6 sflash_ss[3]
port 448 nsew signal input
rlabel metal3 s 0 79632 400 79688 6 sm_a1
port 449 nsew signal input
rlabel metal3 s 0 76608 400 76664 6 sm_a2
port 450 nsew signal input
rlabel metal3 s 0 73920 400 73976 6 sm_b1
port 451 nsew signal input
rlabel metal3 s 0 78288 400 78344 6 sm_b2
port 452 nsew signal input
rlabel metal2 s 57792 0 57848 400 6 soft_irq
port 453 nsew signal output
rlabel metal3 s 0 53760 400 53816 6 spim_miso
port 454 nsew signal input
rlabel metal3 s 0 44016 400 44072 6 spim_mosi
port 455 nsew signal output
rlabel metal3 s 0 82320 400 82376 6 spim_sck
port 456 nsew signal input
rlabel metal3 s 0 50064 400 50120 6 spim_ssn[0]
port 457 nsew signal input
rlabel metal3 s 0 49056 400 49112 6 spim_ssn[1]
port 458 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 spim_ssn[2]
port 459 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 spim_ssn[3]
port 460 nsew signal input
rlabel metal3 s 0 52752 400 52808 6 spis_miso
port 461 nsew signal input
rlabel metal3 s 0 52416 400 52472 6 spis_mosi
port 462 nsew signal output
rlabel metal3 s 0 57120 400 57176 6 spis_sck
port 463 nsew signal output
rlabel metal3 s 0 51744 400 51800 6 spis_ssn
port 464 nsew signal output
rlabel metal2 s 41328 0 41384 400 6 sspim_rst_n
port 465 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 strap_sticky[0]
port 466 nsew signal output
rlabel metal2 s 26208 0 26264 400 6 strap_sticky[10]
port 467 nsew signal output
rlabel metal3 s 0 26544 400 26600 6 strap_sticky[11]
port 468 nsew signal output
rlabel metal2 s 26544 0 26600 400 6 strap_sticky[12]
port 469 nsew signal output
rlabel metal3 s 0 24864 400 24920 6 strap_sticky[13]
port 470 nsew signal output
rlabel metal3 s 0 23856 400 23912 6 strap_sticky[14]
port 471 nsew signal output
rlabel metal3 s 0 22848 400 22904 6 strap_sticky[15]
port 472 nsew signal output
rlabel metal2 s 36960 0 37016 400 6 strap_sticky[16]
port 473 nsew signal output
rlabel metal2 s 40320 0 40376 400 6 strap_sticky[17]
port 474 nsew signal output
rlabel metal2 s 36288 0 36344 400 6 strap_sticky[18]
port 475 nsew signal output
rlabel metal2 s 16464 0 16520 400 6 strap_sticky[19]
port 476 nsew signal output
rlabel metal2 s 27552 0 27608 400 6 strap_sticky[1]
port 477 nsew signal output
rlabel metal2 s 39648 0 39704 400 6 strap_sticky[20]
port 478 nsew signal output
rlabel metal2 s 45696 0 45752 400 6 strap_sticky[21]
port 479 nsew signal output
rlabel metal2 s 46368 0 46424 400 6 strap_sticky[22]
port 480 nsew signal output
rlabel metal2 s 41664 0 41720 400 6 strap_sticky[23]
port 481 nsew signal output
rlabel metal2 s 42000 0 42056 400 6 strap_sticky[24]
port 482 nsew signal output
rlabel metal2 s 46032 0 46088 400 6 strap_sticky[25]
port 483 nsew signal output
rlabel metal2 s 22512 0 22568 400 6 strap_sticky[26]
port 484 nsew signal output
rlabel metal2 s 37968 0 38024 400 6 strap_sticky[27]
port 485 nsew signal output
rlabel metal2 s 40992 0 41048 400 6 strap_sticky[28]
port 486 nsew signal output
rlabel metal2 s 42336 0 42392 400 6 strap_sticky[29]
port 487 nsew signal output
rlabel metal2 s 31248 0 31304 400 6 strap_sticky[2]
port 488 nsew signal output
rlabel metal2 s 38304 0 38360 400 6 strap_sticky[30]
port 489 nsew signal output
rlabel metal2 s 37632 0 37688 400 6 strap_sticky[31]
port 490 nsew signal output
rlabel metal2 s 35280 0 35336 400 6 strap_sticky[3]
port 491 nsew signal output
rlabel metal2 s 33936 0 33992 400 6 strap_sticky[4]
port 492 nsew signal output
rlabel metal2 s 28896 0 28952 400 6 strap_sticky[5]
port 493 nsew signal output
rlabel metal2 s 29232 0 29288 400 6 strap_sticky[6]
port 494 nsew signal output
rlabel metal2 s 35952 0 36008 400 6 strap_sticky[7]
port 495 nsew signal output
rlabel metal3 s 0 27552 400 27608 6 strap_sticky[8]
port 496 nsew signal output
rlabel metal2 s 26880 0 26936 400 6 strap_sticky[9]
port 497 nsew signal output
rlabel metal3 s 0 19824 400 19880 6 strap_uartm[0]
port 498 nsew signal output
rlabel metal3 s 0 22176 400 22232 6 strap_uartm[1]
port 499 nsew signal output
rlabel metal2 s 50736 0 50792 400 6 system_strap[0]
port 500 nsew signal input
rlabel metal3 s 0 25536 400 25592 6 system_strap[10]
port 501 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 system_strap[11]
port 502 nsew signal input
rlabel metal3 s 0 29232 400 29288 6 system_strap[12]
port 503 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 system_strap[13]
port 504 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 system_strap[14]
port 505 nsew signal input
rlabel metal3 s 0 28896 400 28952 6 system_strap[15]
port 506 nsew signal input
rlabel metal2 s 70560 0 70616 400 6 system_strap[16]
port 507 nsew signal input
rlabel metal2 s 69888 0 69944 400 6 system_strap[17]
port 508 nsew signal input
rlabel metal2 s 68880 0 68936 400 6 system_strap[18]
port 509 nsew signal input
rlabel metal2 s 60816 0 60872 400 6 system_strap[19]
port 510 nsew signal input
rlabel metal3 s 119600 36288 120000 36344 6 system_strap[1]
port 511 nsew signal input
rlabel metal2 s 67200 0 67256 400 6 system_strap[20]
port 512 nsew signal input
rlabel metal2 s 59472 0 59528 400 6 system_strap[21]
port 513 nsew signal input
rlabel metal2 s 59808 0 59864 400 6 system_strap[22]
port 514 nsew signal input
rlabel metal2 s 62832 0 62888 400 6 system_strap[23]
port 515 nsew signal input
rlabel metal2 s 64176 0 64232 400 6 system_strap[24]
port 516 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 system_strap[25]
port 517 nsew signal input
rlabel metal2 s 63504 0 63560 400 6 system_strap[26]
port 518 nsew signal input
rlabel metal2 s 56112 0 56168 400 6 system_strap[27]
port 519 nsew signal input
rlabel metal2 s 60480 0 60536 400 6 system_strap[28]
port 520 nsew signal input
rlabel metal2 s 58800 0 58856 400 6 system_strap[29]
port 521 nsew signal input
rlabel metal3 s 119600 37296 120000 37352 6 system_strap[2]
port 522 nsew signal input
rlabel metal2 s 65520 0 65576 400 6 system_strap[30]
port 523 nsew signal input
rlabel metal2 s 56448 0 56504 400 6 system_strap[31]
port 524 nsew signal input
rlabel metal3 s 119600 37968 120000 38024 6 system_strap[3]
port 525 nsew signal input
rlabel metal2 s 53760 0 53816 400 6 system_strap[4]
port 526 nsew signal input
rlabel metal2 s 58128 0 58184 400 6 system_strap[5]
port 527 nsew signal input
rlabel metal2 s 47712 0 47768 400 6 system_strap[6]
port 528 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 system_strap[7]
port 529 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 system_strap[8]
port 530 nsew signal input
rlabel metal3 s 0 31920 400 31976 6 system_strap[9]
port 531 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 uart_rst_n[0]
port 532 nsew signal output
rlabel metal2 s 42672 0 42728 400 6 uart_rst_n[1]
port 533 nsew signal output
rlabel metal2 s 43680 0 43736 400 6 uart_rxd[0]
port 534 nsew signal output
rlabel metal3 s 0 36960 400 37016 6 uart_rxd[1]
port 535 nsew signal output
rlabel metal2 s 44688 0 44744 400 6 uart_txd[0]
port 536 nsew signal input
rlabel metal3 s 0 55776 400 55832 6 uart_txd[1]
port 537 nsew signal input
rlabel metal2 s 44352 0 44408 400 6 uartm_rxd
port 538 nsew signal output
rlabel metal2 s 17472 0 17528 400 6 uartm_txd
port 539 nsew signal input
rlabel metal3 s 0 23184 400 23240 6 usb_clk
port 540 nsew signal output
rlabel metal3 s 0 70224 400 70280 6 usb_dn_i
port 541 nsew signal output
rlabel metal3 s 0 63168 400 63224 6 usb_dn_o
port 542 nsew signal input
rlabel metal3 s 0 69552 400 69608 6 usb_dp_i
port 543 nsew signal output
rlabel metal3 s 0 64176 400 64232 6 usb_dp_o
port 544 nsew signal input
rlabel metal2 s 48720 0 48776 400 6 usb_intr
port 545 nsew signal input
rlabel metal3 s 0 63840 400 63896 6 usb_oen
port 546 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 usb_rst_n
port 547 nsew signal output
rlabel metal3 s 119600 36624 120000 36680 6 user_clock1
port 548 nsew signal input
rlabel metal2 s 50400 0 50456 400 6 user_clock2
port 549 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 user_irq[0]
port 550 nsew signal output
rlabel metal2 s 54096 0 54152 400 6 user_irq[1]
port 551 nsew signal output
rlabel metal2 s 61824 0 61880 400 6 user_irq[2]
port 552 nsew signal output
rlabel metal2 s 99792 0 99848 400 6 wbd_clk_int
port 553 nsew signal input
rlabel metal2 s 105504 0 105560 400 6 wbd_clk_pinmux
port 554 nsew signal output
rlabel metal3 s 0 32592 400 32648 6 xtal_clk
port 555 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 36320770
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/pinmux_top/runs/23_11_12_19_15/results/signoff/pinmux_top.magic.gds
string GDS_START 649652
<< end >>

