VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO peri_top
  CLASS BLOCK ;
  FOREIGN peri_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 500.000 ;
  PIN mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END mclk
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.000 4.000 476.560 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 89.600 4.000 90.160 ;
    END
  END reg_addr[0]
  PIN reg_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END reg_addr[10]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 4.000 73.360 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 4.000 67.760 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 4.000 62.160 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 4.000 56.560 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 4.000 50.960 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.800 4.000 45.360 ;
    END
  END reg_addr[8]
  PIN reg_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 4.000 39.760 ;
    END
  END reg_addr[9]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.000 4.000 112.560 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 4.000 106.960 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.200 4.000 95.760 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.400 4.000 22.960 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.400 4.000 470.960 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 414.400 4.000 414.960 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 403.200 4.000 403.760 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 397.600 4.000 398.160 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.000 4.000 392.560 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.200 4.000 375.760 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.600 4.000 370.160 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.000 4.000 364.560 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 464.800 4.000 465.360 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.400 4.000 358.960 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.800 4.000 353.360 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.200 4.000 347.760 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 341.600 4.000 342.160 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.000 4.000 336.560 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.400 4.000 330.960 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.200 4.000 319.760 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.600 4.000 314.160 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.000 4.000 308.560 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 459.200 4.000 459.760 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 296.800 4.000 297.360 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.400 4.000 442.960 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 436.800 4.000 437.360 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 431.200 4.000 431.760 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.600 4.000 426.160 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.000 4.000 420.560 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.200 4.000 291.760 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.200 4.000 235.760 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 4.000 230.160 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.000 4.000 224.560 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 4.000 196.560 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.400 4.000 190.960 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 4.000 286.160 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.200 4.000 179.760 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 4.000 174.160 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 4.000 162.960 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 156.800 4.000 157.360 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.600 4.000 146.160 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 4.000 129.360 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.000 4.000 280.560 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 4.000 274.960 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.800 4.000 269.360 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.400 4.000 246.960 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 4.000 241.360 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.000 4.000 28.560 ;
    END
  END reg_wr
  PIN rtc_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 496.000 49.840 500.000 ;
    END
  END rtc_clk
  PIN rtc_intr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 496.000 149.520 500.000 ;
    END
  END rtc_intr
  PIN s_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.498000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 4.000 ;
    END
  END s_reset_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.940 15.380 26.140 482.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.940 15.380 126.140 482.460 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 69.940 15.380 76.140 482.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.940 15.380 176.140 482.460 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 193.200 482.460 ;
      LAYER Metal2 ;
        RECT 7.980 495.700 48.980 496.000 ;
        RECT 50.140 495.700 148.660 496.000 ;
        RECT 149.820 495.700 191.940 496.000 ;
        RECT 7.980 4.300 191.940 495.700 ;
        RECT 7.980 4.000 48.980 4.300 ;
        RECT 50.140 4.000 148.660 4.300 ;
        RECT 149.820 4.000 191.940 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 476.860 191.990 482.300 ;
        RECT 4.300 475.700 191.990 476.860 ;
        RECT 4.000 471.260 191.990 475.700 ;
        RECT 4.300 470.100 191.990 471.260 ;
        RECT 4.000 465.660 191.990 470.100 ;
        RECT 4.300 464.500 191.990 465.660 ;
        RECT 4.000 460.060 191.990 464.500 ;
        RECT 4.300 458.900 191.990 460.060 ;
        RECT 4.000 454.460 191.990 458.900 ;
        RECT 4.300 453.300 191.990 454.460 ;
        RECT 4.000 448.860 191.990 453.300 ;
        RECT 4.300 447.700 191.990 448.860 ;
        RECT 4.000 443.260 191.990 447.700 ;
        RECT 4.300 442.100 191.990 443.260 ;
        RECT 4.000 437.660 191.990 442.100 ;
        RECT 4.300 436.500 191.990 437.660 ;
        RECT 4.000 432.060 191.990 436.500 ;
        RECT 4.300 430.900 191.990 432.060 ;
        RECT 4.000 426.460 191.990 430.900 ;
        RECT 4.300 425.300 191.990 426.460 ;
        RECT 4.000 420.860 191.990 425.300 ;
        RECT 4.300 419.700 191.990 420.860 ;
        RECT 4.000 415.260 191.990 419.700 ;
        RECT 4.300 414.100 191.990 415.260 ;
        RECT 4.000 409.660 191.990 414.100 ;
        RECT 4.300 408.500 191.990 409.660 ;
        RECT 4.000 404.060 191.990 408.500 ;
        RECT 4.300 402.900 191.990 404.060 ;
        RECT 4.000 398.460 191.990 402.900 ;
        RECT 4.300 397.300 191.990 398.460 ;
        RECT 4.000 392.860 191.990 397.300 ;
        RECT 4.300 391.700 191.990 392.860 ;
        RECT 4.000 387.260 191.990 391.700 ;
        RECT 4.300 386.100 191.990 387.260 ;
        RECT 4.000 381.660 191.990 386.100 ;
        RECT 4.300 380.500 191.990 381.660 ;
        RECT 4.000 376.060 191.990 380.500 ;
        RECT 4.300 374.900 191.990 376.060 ;
        RECT 4.000 370.460 191.990 374.900 ;
        RECT 4.300 369.300 191.990 370.460 ;
        RECT 4.000 364.860 191.990 369.300 ;
        RECT 4.300 363.700 191.990 364.860 ;
        RECT 4.000 359.260 191.990 363.700 ;
        RECT 4.300 358.100 191.990 359.260 ;
        RECT 4.000 353.660 191.990 358.100 ;
        RECT 4.300 352.500 191.990 353.660 ;
        RECT 4.000 348.060 191.990 352.500 ;
        RECT 4.300 346.900 191.990 348.060 ;
        RECT 4.000 342.460 191.990 346.900 ;
        RECT 4.300 341.300 191.990 342.460 ;
        RECT 4.000 336.860 191.990 341.300 ;
        RECT 4.300 335.700 191.990 336.860 ;
        RECT 4.000 331.260 191.990 335.700 ;
        RECT 4.300 330.100 191.990 331.260 ;
        RECT 4.000 325.660 191.990 330.100 ;
        RECT 4.300 324.500 191.990 325.660 ;
        RECT 4.000 320.060 191.990 324.500 ;
        RECT 4.300 318.900 191.990 320.060 ;
        RECT 4.000 314.460 191.990 318.900 ;
        RECT 4.300 313.300 191.990 314.460 ;
        RECT 4.000 308.860 191.990 313.300 ;
        RECT 4.300 307.700 191.990 308.860 ;
        RECT 4.000 303.260 191.990 307.700 ;
        RECT 4.300 302.100 191.990 303.260 ;
        RECT 4.000 297.660 191.990 302.100 ;
        RECT 4.300 296.500 191.990 297.660 ;
        RECT 4.000 292.060 191.990 296.500 ;
        RECT 4.300 290.900 191.990 292.060 ;
        RECT 4.000 286.460 191.990 290.900 ;
        RECT 4.300 285.300 191.990 286.460 ;
        RECT 4.000 280.860 191.990 285.300 ;
        RECT 4.300 279.700 191.990 280.860 ;
        RECT 4.000 275.260 191.990 279.700 ;
        RECT 4.300 274.100 191.990 275.260 ;
        RECT 4.000 269.660 191.990 274.100 ;
        RECT 4.300 268.500 191.990 269.660 ;
        RECT 4.000 264.060 191.990 268.500 ;
        RECT 4.300 262.900 191.990 264.060 ;
        RECT 4.000 258.460 191.990 262.900 ;
        RECT 4.300 257.300 191.990 258.460 ;
        RECT 4.000 252.860 191.990 257.300 ;
        RECT 4.300 251.700 191.990 252.860 ;
        RECT 4.000 247.260 191.990 251.700 ;
        RECT 4.300 246.100 191.990 247.260 ;
        RECT 4.000 241.660 191.990 246.100 ;
        RECT 4.300 240.500 191.990 241.660 ;
        RECT 4.000 236.060 191.990 240.500 ;
        RECT 4.300 234.900 191.990 236.060 ;
        RECT 4.000 230.460 191.990 234.900 ;
        RECT 4.300 229.300 191.990 230.460 ;
        RECT 4.000 224.860 191.990 229.300 ;
        RECT 4.300 223.700 191.990 224.860 ;
        RECT 4.000 219.260 191.990 223.700 ;
        RECT 4.300 218.100 191.990 219.260 ;
        RECT 4.000 213.660 191.990 218.100 ;
        RECT 4.300 212.500 191.990 213.660 ;
        RECT 4.000 208.060 191.990 212.500 ;
        RECT 4.300 206.900 191.990 208.060 ;
        RECT 4.000 202.460 191.990 206.900 ;
        RECT 4.300 201.300 191.990 202.460 ;
        RECT 4.000 196.860 191.990 201.300 ;
        RECT 4.300 195.700 191.990 196.860 ;
        RECT 4.000 191.260 191.990 195.700 ;
        RECT 4.300 190.100 191.990 191.260 ;
        RECT 4.000 185.660 191.990 190.100 ;
        RECT 4.300 184.500 191.990 185.660 ;
        RECT 4.000 180.060 191.990 184.500 ;
        RECT 4.300 178.900 191.990 180.060 ;
        RECT 4.000 174.460 191.990 178.900 ;
        RECT 4.300 173.300 191.990 174.460 ;
        RECT 4.000 168.860 191.990 173.300 ;
        RECT 4.300 167.700 191.990 168.860 ;
        RECT 4.000 163.260 191.990 167.700 ;
        RECT 4.300 162.100 191.990 163.260 ;
        RECT 4.000 157.660 191.990 162.100 ;
        RECT 4.300 156.500 191.990 157.660 ;
        RECT 4.000 152.060 191.990 156.500 ;
        RECT 4.300 150.900 191.990 152.060 ;
        RECT 4.000 146.460 191.990 150.900 ;
        RECT 4.300 145.300 191.990 146.460 ;
        RECT 4.000 140.860 191.990 145.300 ;
        RECT 4.300 139.700 191.990 140.860 ;
        RECT 4.000 135.260 191.990 139.700 ;
        RECT 4.300 134.100 191.990 135.260 ;
        RECT 4.000 129.660 191.990 134.100 ;
        RECT 4.300 128.500 191.990 129.660 ;
        RECT 4.000 124.060 191.990 128.500 ;
        RECT 4.300 122.900 191.990 124.060 ;
        RECT 4.000 118.460 191.990 122.900 ;
        RECT 4.300 117.300 191.990 118.460 ;
        RECT 4.000 112.860 191.990 117.300 ;
        RECT 4.300 111.700 191.990 112.860 ;
        RECT 4.000 107.260 191.990 111.700 ;
        RECT 4.300 106.100 191.990 107.260 ;
        RECT 4.000 101.660 191.990 106.100 ;
        RECT 4.300 100.500 191.990 101.660 ;
        RECT 4.000 96.060 191.990 100.500 ;
        RECT 4.300 94.900 191.990 96.060 ;
        RECT 4.000 90.460 191.990 94.900 ;
        RECT 4.300 89.300 191.990 90.460 ;
        RECT 4.000 84.860 191.990 89.300 ;
        RECT 4.300 83.700 191.990 84.860 ;
        RECT 4.000 79.260 191.990 83.700 ;
        RECT 4.300 78.100 191.990 79.260 ;
        RECT 4.000 73.660 191.990 78.100 ;
        RECT 4.300 72.500 191.990 73.660 ;
        RECT 4.000 68.060 191.990 72.500 ;
        RECT 4.300 66.900 191.990 68.060 ;
        RECT 4.000 62.460 191.990 66.900 ;
        RECT 4.300 61.300 191.990 62.460 ;
        RECT 4.000 56.860 191.990 61.300 ;
        RECT 4.300 55.700 191.990 56.860 ;
        RECT 4.000 51.260 191.990 55.700 ;
        RECT 4.300 50.100 191.990 51.260 ;
        RECT 4.000 45.660 191.990 50.100 ;
        RECT 4.300 44.500 191.990 45.660 ;
        RECT 4.000 40.060 191.990 44.500 ;
        RECT 4.300 38.900 191.990 40.060 ;
        RECT 4.000 34.460 191.990 38.900 ;
        RECT 4.300 33.300 191.990 34.460 ;
        RECT 4.000 28.860 191.990 33.300 ;
        RECT 4.300 27.700 191.990 28.860 ;
        RECT 4.000 23.260 191.990 27.700 ;
        RECT 4.300 22.100 191.990 23.260 ;
        RECT 4.000 15.540 191.990 22.100 ;
      LAYER Metal4 ;
        RECT 9.100 57.210 19.640 433.350 ;
        RECT 26.440 57.210 69.640 433.350 ;
        RECT 76.440 57.210 119.640 433.350 ;
        RECT 126.440 57.210 169.640 433.350 ;
        RECT 176.440 57.210 176.820 433.350 ;
  END
END peri_top
END LIBRARY

