* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuD

* Black-box entry subcircuit for serv_rf_top abstract view
.subckt serv_rf_top clk i_dbus_ack i_dbus_rdt[0] i_dbus_rdt[10] i_dbus_rdt[11] i_dbus_rdt[12]
+ i_dbus_rdt[13] i_dbus_rdt[14] i_dbus_rdt[15] i_dbus_rdt[16] i_dbus_rdt[17] i_dbus_rdt[18]
+ i_dbus_rdt[19] i_dbus_rdt[1] i_dbus_rdt[20] i_dbus_rdt[21] i_dbus_rdt[22] i_dbus_rdt[23]
+ i_dbus_rdt[24] i_dbus_rdt[25] i_dbus_rdt[26] i_dbus_rdt[27] i_dbus_rdt[28] i_dbus_rdt[29]
+ i_dbus_rdt[2] i_dbus_rdt[30] i_dbus_rdt[31] i_dbus_rdt[3] i_dbus_rdt[4] i_dbus_rdt[5]
+ i_dbus_rdt[6] i_dbus_rdt[7] i_dbus_rdt[8] i_dbus_rdt[9] i_ext_rd[0] i_ext_rd[10]
+ i_ext_rd[11] i_ext_rd[12] i_ext_rd[13] i_ext_rd[14] i_ext_rd[15] i_ext_rd[16] i_ext_rd[17]
+ i_ext_rd[18] i_ext_rd[19] i_ext_rd[1] i_ext_rd[20] i_ext_rd[21] i_ext_rd[22] i_ext_rd[23]
+ i_ext_rd[24] i_ext_rd[25] i_ext_rd[26] i_ext_rd[27] i_ext_rd[28] i_ext_rd[29] i_ext_rd[2]
+ i_ext_rd[30] i_ext_rd[31] i_ext_rd[3] i_ext_rd[4] i_ext_rd[5] i_ext_rd[6] i_ext_rd[7]
+ i_ext_rd[8] i_ext_rd[9] i_ext_ready i_ibus_ack i_ibus_rdt[0] i_ibus_rdt[10] i_ibus_rdt[11]
+ i_ibus_rdt[12] i_ibus_rdt[13] i_ibus_rdt[14] i_ibus_rdt[15] i_ibus_rdt[16] i_ibus_rdt[17]
+ i_ibus_rdt[18] i_ibus_rdt[19] i_ibus_rdt[1] i_ibus_rdt[20] i_ibus_rdt[21] i_ibus_rdt[22]
+ i_ibus_rdt[23] i_ibus_rdt[24] i_ibus_rdt[25] i_ibus_rdt[26] i_ibus_rdt[27] i_ibus_rdt[28]
+ i_ibus_rdt[29] i_ibus_rdt[2] i_ibus_rdt[30] i_ibus_rdt[31] i_ibus_rdt[3] i_ibus_rdt[4]
+ i_ibus_rdt[5] i_ibus_rdt[6] i_ibus_rdt[7] i_ibus_rdt[8] i_ibus_rdt[9] i_rst i_timer_irq
+ o_dbus_adr[0] o_dbus_adr[10] o_dbus_adr[11] o_dbus_adr[12] o_dbus_adr[13] o_dbus_adr[14]
+ o_dbus_adr[15] o_dbus_adr[16] o_dbus_adr[17] o_dbus_adr[18] o_dbus_adr[19] o_dbus_adr[1]
+ o_dbus_adr[20] o_dbus_adr[21] o_dbus_adr[22] o_dbus_adr[23] o_dbus_adr[24] o_dbus_adr[25]
+ o_dbus_adr[26] o_dbus_adr[27] o_dbus_adr[28] o_dbus_adr[29] o_dbus_adr[2] o_dbus_adr[30]
+ o_dbus_adr[31] o_dbus_adr[3] o_dbus_adr[4] o_dbus_adr[5] o_dbus_adr[6] o_dbus_adr[7]
+ o_dbus_adr[8] o_dbus_adr[9] o_dbus_cyc o_dbus_dat[0] o_dbus_dat[10] o_dbus_dat[11]
+ o_dbus_dat[12] o_dbus_dat[13] o_dbus_dat[14] o_dbus_dat[15] o_dbus_dat[16] o_dbus_dat[17]
+ o_dbus_dat[18] o_dbus_dat[19] o_dbus_dat[1] o_dbus_dat[20] o_dbus_dat[21] o_dbus_dat[22]
+ o_dbus_dat[23] o_dbus_dat[24] o_dbus_dat[25] o_dbus_dat[26] o_dbus_dat[27] o_dbus_dat[28]
+ o_dbus_dat[29] o_dbus_dat[2] o_dbus_dat[30] o_dbus_dat[31] o_dbus_dat[3] o_dbus_dat[4]
+ o_dbus_dat[5] o_dbus_dat[6] o_dbus_dat[7] o_dbus_dat[8] o_dbus_dat[9] o_dbus_sel[0]
+ o_dbus_sel[1] o_dbus_sel[2] o_dbus_sel[3] o_dbus_we o_ext_funct3[0] o_ext_funct3[1]
+ o_ext_funct3[2] o_ext_rs1[0] o_ext_rs1[10] o_ext_rs1[11] o_ext_rs1[12] o_ext_rs1[13]
+ o_ext_rs1[14] o_ext_rs1[15] o_ext_rs1[16] o_ext_rs1[17] o_ext_rs1[18] o_ext_rs1[19]
+ o_ext_rs1[1] o_ext_rs1[20] o_ext_rs1[21] o_ext_rs1[22] o_ext_rs1[23] o_ext_rs1[24]
+ o_ext_rs1[25] o_ext_rs1[26] o_ext_rs1[27] o_ext_rs1[28] o_ext_rs1[29] o_ext_rs1[2]
+ o_ext_rs1[30] o_ext_rs1[31] o_ext_rs1[3] o_ext_rs1[4] o_ext_rs1[5] o_ext_rs1[6]
+ o_ext_rs1[7] o_ext_rs1[8] o_ext_rs1[9] o_ext_rs2[0] o_ext_rs2[10] o_ext_rs2[11]
+ o_ext_rs2[12] o_ext_rs2[13] o_ext_rs2[14] o_ext_rs2[15] o_ext_rs2[16] o_ext_rs2[17]
+ o_ext_rs2[18] o_ext_rs2[19] o_ext_rs2[1] o_ext_rs2[20] o_ext_rs2[21] o_ext_rs2[22]
+ o_ext_rs2[23] o_ext_rs2[24] o_ext_rs2[25] o_ext_rs2[26] o_ext_rs2[27] o_ext_rs2[28]
+ o_ext_rs2[29] o_ext_rs2[2] o_ext_rs2[30] o_ext_rs2[31] o_ext_rs2[3] o_ext_rs2[4]
+ o_ext_rs2[5] o_ext_rs2[6] o_ext_rs2[7] o_ext_rs2[8] o_ext_rs2[9] o_ibus_adr[0] o_ibus_adr[10]
+ o_ibus_adr[11] o_ibus_adr[12] o_ibus_adr[13] o_ibus_adr[14] o_ibus_adr[15] o_ibus_adr[16]
+ o_ibus_adr[17] o_ibus_adr[18] o_ibus_adr[19] o_ibus_adr[1] o_ibus_adr[20] o_ibus_adr[21]
+ o_ibus_adr[22] o_ibus_adr[23] o_ibus_adr[24] o_ibus_adr[25] o_ibus_adr[26] o_ibus_adr[27]
+ o_ibus_adr[28] o_ibus_adr[29] o_ibus_adr[2] o_ibus_adr[30] o_ibus_adr[31] o_ibus_adr[3]
+ o_ibus_adr[4] o_ibus_adr[5] o_ibus_adr[6] o_ibus_adr[7] o_ibus_adr[8] o_ibus_adr[9]
+ o_ibus_cyc o_mdu_valid vdd vss
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xserv_rf_top wb_clk_i serv_rf_top/i_dbus_ack serv_rf_top/i_dbus_rdt[0] serv_rf_top/i_dbus_rdt[10]
+ serv_rf_top/i_dbus_rdt[11] serv_rf_top/i_dbus_rdt[12] serv_rf_top/i_dbus_rdt[13]
+ serv_rf_top/i_dbus_rdt[14] serv_rf_top/i_dbus_rdt[15] serv_rf_top/i_dbus_rdt[16]
+ serv_rf_top/i_dbus_rdt[17] serv_rf_top/i_dbus_rdt[18] serv_rf_top/i_dbus_rdt[19]
+ serv_rf_top/i_dbus_rdt[1] serv_rf_top/i_dbus_rdt[20] serv_rf_top/i_dbus_rdt[21]
+ serv_rf_top/i_dbus_rdt[22] serv_rf_top/i_dbus_rdt[23] serv_rf_top/i_dbus_rdt[24]
+ serv_rf_top/i_dbus_rdt[25] serv_rf_top/i_dbus_rdt[26] serv_rf_top/i_dbus_rdt[27]
+ serv_rf_top/i_dbus_rdt[28] serv_rf_top/i_dbus_rdt[29] serv_rf_top/i_dbus_rdt[2]
+ serv_rf_top/i_dbus_rdt[30] serv_rf_top/i_dbus_rdt[31] serv_rf_top/i_dbus_rdt[3]
+ serv_rf_top/i_dbus_rdt[4] serv_rf_top/i_dbus_rdt[5] serv_rf_top/i_dbus_rdt[6] serv_rf_top/i_dbus_rdt[7]
+ serv_rf_top/i_dbus_rdt[8] serv_rf_top/i_dbus_rdt[9] serv_rf_top/i_ext_rd[0] serv_rf_top/i_ext_rd[10]
+ serv_rf_top/i_ext_rd[11] serv_rf_top/i_ext_rd[12] serv_rf_top/i_ext_rd[13] serv_rf_top/i_ext_rd[14]
+ serv_rf_top/i_ext_rd[15] serv_rf_top/i_ext_rd[16] serv_rf_top/i_ext_rd[17] serv_rf_top/i_ext_rd[18]
+ serv_rf_top/i_ext_rd[19] serv_rf_top/i_ext_rd[1] serv_rf_top/i_ext_rd[20] serv_rf_top/i_ext_rd[21]
+ serv_rf_top/i_ext_rd[22] serv_rf_top/i_ext_rd[23] serv_rf_top/i_ext_rd[24] serv_rf_top/i_ext_rd[25]
+ serv_rf_top/i_ext_rd[26] serv_rf_top/i_ext_rd[27] serv_rf_top/i_ext_rd[28] serv_rf_top/i_ext_rd[29]
+ serv_rf_top/i_ext_rd[2] serv_rf_top/i_ext_rd[30] serv_rf_top/i_ext_rd[31] serv_rf_top/i_ext_rd[3]
+ serv_rf_top/i_ext_rd[4] serv_rf_top/i_ext_rd[5] serv_rf_top/i_ext_rd[6] serv_rf_top/i_ext_rd[7]
+ serv_rf_top/i_ext_rd[8] serv_rf_top/i_ext_rd[9] serv_rf_top/i_ext_ready serv_rf_top/i_ibus_ack
+ serv_rf_top/i_ibus_rdt[0] serv_rf_top/i_ibus_rdt[10] serv_rf_top/i_ibus_rdt[11]
+ serv_rf_top/i_ibus_rdt[12] serv_rf_top/i_ibus_rdt[13] serv_rf_top/i_ibus_rdt[14]
+ serv_rf_top/i_ibus_rdt[15] serv_rf_top/i_ibus_rdt[16] serv_rf_top/i_ibus_rdt[17]
+ serv_rf_top/i_ibus_rdt[18] serv_rf_top/i_ibus_rdt[19] serv_rf_top/i_ibus_rdt[1]
+ serv_rf_top/i_ibus_rdt[20] serv_rf_top/i_ibus_rdt[21] serv_rf_top/i_ibus_rdt[22]
+ serv_rf_top/i_ibus_rdt[23] serv_rf_top/i_ibus_rdt[24] serv_rf_top/i_ibus_rdt[25]
+ serv_rf_top/i_ibus_rdt[26] serv_rf_top/i_ibus_rdt[27] serv_rf_top/i_ibus_rdt[28]
+ serv_rf_top/i_ibus_rdt[29] serv_rf_top/i_ibus_rdt[2] serv_rf_top/i_ibus_rdt[30]
+ serv_rf_top/i_ibus_rdt[31] serv_rf_top/i_ibus_rdt[3] serv_rf_top/i_ibus_rdt[4] serv_rf_top/i_ibus_rdt[5]
+ serv_rf_top/i_ibus_rdt[6] serv_rf_top/i_ibus_rdt[7] serv_rf_top/i_ibus_rdt[8] serv_rf_top/i_ibus_rdt[9]
+ wb_rst_i user_irq[0] serv_rf_top/o_dbus_adr[0] serv_rf_top/o_dbus_adr[10] serv_rf_top/o_dbus_adr[11]
+ serv_rf_top/o_dbus_adr[12] serv_rf_top/o_dbus_adr[13] serv_rf_top/o_dbus_adr[14]
+ serv_rf_top/o_dbus_adr[15] serv_rf_top/o_dbus_adr[16] serv_rf_top/o_dbus_adr[17]
+ serv_rf_top/o_dbus_adr[18] serv_rf_top/o_dbus_adr[19] serv_rf_top/o_dbus_adr[1]
+ serv_rf_top/o_dbus_adr[20] serv_rf_top/o_dbus_adr[21] serv_rf_top/o_dbus_adr[22]
+ serv_rf_top/o_dbus_adr[23] serv_rf_top/o_dbus_adr[24] serv_rf_top/o_dbus_adr[25]
+ serv_rf_top/o_dbus_adr[26] serv_rf_top/o_dbus_adr[27] serv_rf_top/o_dbus_adr[28]
+ serv_rf_top/o_dbus_adr[29] serv_rf_top/o_dbus_adr[2] serv_rf_top/o_dbus_adr[30]
+ serv_rf_top/o_dbus_adr[31] serv_rf_top/o_dbus_adr[3] serv_rf_top/o_dbus_adr[4] serv_rf_top/o_dbus_adr[5]
+ serv_rf_top/o_dbus_adr[6] serv_rf_top/o_dbus_adr[7] serv_rf_top/o_dbus_adr[8] serv_rf_top/o_dbus_adr[9]
+ serv_rf_top/o_dbus_cyc serv_rf_top/o_dbus_dat[0] serv_rf_top/o_dbus_dat[10] serv_rf_top/o_dbus_dat[11]
+ serv_rf_top/o_dbus_dat[12] serv_rf_top/o_dbus_dat[13] serv_rf_top/o_dbus_dat[14]
+ serv_rf_top/o_dbus_dat[15] serv_rf_top/o_dbus_dat[16] serv_rf_top/o_dbus_dat[17]
+ serv_rf_top/o_dbus_dat[18] serv_rf_top/o_dbus_dat[19] serv_rf_top/o_dbus_dat[1]
+ serv_rf_top/o_dbus_dat[20] serv_rf_top/o_dbus_dat[21] serv_rf_top/o_dbus_dat[22]
+ serv_rf_top/o_dbus_dat[23] serv_rf_top/o_dbus_dat[24] serv_rf_top/o_dbus_dat[25]
+ serv_rf_top/o_dbus_dat[26] serv_rf_top/o_dbus_dat[27] serv_rf_top/o_dbus_dat[28]
+ serv_rf_top/o_dbus_dat[29] serv_rf_top/o_dbus_dat[2] serv_rf_top/o_dbus_dat[30]
+ serv_rf_top/o_dbus_dat[31] serv_rf_top/o_dbus_dat[3] serv_rf_top/o_dbus_dat[4] serv_rf_top/o_dbus_dat[5]
+ serv_rf_top/o_dbus_dat[6] serv_rf_top/o_dbus_dat[7] serv_rf_top/o_dbus_dat[8] serv_rf_top/o_dbus_dat[9]
+ serv_rf_top/o_dbus_sel[0] serv_rf_top/o_dbus_sel[1] serv_rf_top/o_dbus_sel[2] serv_rf_top/o_dbus_sel[3]
+ serv_rf_top/o_dbus_we serv_rf_top/o_ext_funct3[0] serv_rf_top/o_ext_funct3[1] serv_rf_top/o_ext_funct3[2]
+ serv_rf_top/o_ext_rs1[0] serv_rf_top/o_ext_rs1[10] serv_rf_top/o_ext_rs1[11] serv_rf_top/o_ext_rs1[12]
+ serv_rf_top/o_ext_rs1[13] serv_rf_top/o_ext_rs1[14] serv_rf_top/o_ext_rs1[15] serv_rf_top/o_ext_rs1[16]
+ serv_rf_top/o_ext_rs1[17] serv_rf_top/o_ext_rs1[18] serv_rf_top/o_ext_rs1[19] serv_rf_top/o_ext_rs1[1]
+ serv_rf_top/o_ext_rs1[20] serv_rf_top/o_ext_rs1[21] serv_rf_top/o_ext_rs1[22] serv_rf_top/o_ext_rs1[23]
+ serv_rf_top/o_ext_rs1[24] serv_rf_top/o_ext_rs1[25] serv_rf_top/o_ext_rs1[26] serv_rf_top/o_ext_rs1[27]
+ serv_rf_top/o_ext_rs1[28] serv_rf_top/o_ext_rs1[29] serv_rf_top/o_ext_rs1[2] serv_rf_top/o_ext_rs1[30]
+ serv_rf_top/o_ext_rs1[31] serv_rf_top/o_ext_rs1[3] serv_rf_top/o_ext_rs1[4] serv_rf_top/o_ext_rs1[5]
+ serv_rf_top/o_ext_rs1[6] serv_rf_top/o_ext_rs1[7] serv_rf_top/o_ext_rs1[8] serv_rf_top/o_ext_rs1[9]
+ serv_rf_top/o_ext_rs2[0] serv_rf_top/o_ext_rs2[10] serv_rf_top/o_ext_rs2[11] serv_rf_top/o_ext_rs2[12]
+ serv_rf_top/o_ext_rs2[13] serv_rf_top/o_ext_rs2[14] serv_rf_top/o_ext_rs2[15] serv_rf_top/o_ext_rs2[16]
+ serv_rf_top/o_ext_rs2[17] serv_rf_top/o_ext_rs2[18] serv_rf_top/o_ext_rs2[19] serv_rf_top/o_ext_rs2[1]
+ serv_rf_top/o_ext_rs2[20] serv_rf_top/o_ext_rs2[21] serv_rf_top/o_ext_rs2[22] serv_rf_top/o_ext_rs2[23]
+ serv_rf_top/o_ext_rs2[24] serv_rf_top/o_ext_rs2[25] serv_rf_top/o_ext_rs2[26] serv_rf_top/o_ext_rs2[27]
+ serv_rf_top/o_ext_rs2[28] serv_rf_top/o_ext_rs2[29] serv_rf_top/o_ext_rs2[2] serv_rf_top/o_ext_rs2[30]
+ serv_rf_top/o_ext_rs2[31] serv_rf_top/o_ext_rs2[3] serv_rf_top/o_ext_rs2[4] serv_rf_top/o_ext_rs2[5]
+ serv_rf_top/o_ext_rs2[6] serv_rf_top/o_ext_rs2[7] serv_rf_top/o_ext_rs2[8] serv_rf_top/o_ext_rs2[9]
+ serv_rf_top/o_ibus_adr[0] serv_rf_top/o_ibus_adr[10] serv_rf_top/o_ibus_adr[11]
+ serv_rf_top/o_ibus_adr[12] serv_rf_top/o_ibus_adr[13] serv_rf_top/o_ibus_adr[14]
+ serv_rf_top/o_ibus_adr[15] serv_rf_top/o_ibus_adr[16] serv_rf_top/o_ibus_adr[17]
+ serv_rf_top/o_ibus_adr[18] serv_rf_top/o_ibus_adr[19] serv_rf_top/o_ibus_adr[1]
+ serv_rf_top/o_ibus_adr[20] serv_rf_top/o_ibus_adr[21] serv_rf_top/o_ibus_adr[22]
+ serv_rf_top/o_ibus_adr[23] serv_rf_top/o_ibus_adr[24] serv_rf_top/o_ibus_adr[25]
+ serv_rf_top/o_ibus_adr[26] serv_rf_top/o_ibus_adr[27] serv_rf_top/o_ibus_adr[28]
+ serv_rf_top/o_ibus_adr[29] serv_rf_top/o_ibus_adr[2] serv_rf_top/o_ibus_adr[30]
+ serv_rf_top/o_ibus_adr[31] serv_rf_top/o_ibus_adr[3] serv_rf_top/o_ibus_adr[4] serv_rf_top/o_ibus_adr[5]
+ serv_rf_top/o_ibus_adr[6] serv_rf_top/o_ibus_adr[7] serv_rf_top/o_ibus_adr[8] serv_rf_top/o_ibus_adr[9]
+ serv_rf_top/o_ibus_cyc serv_rf_top/o_mdu_valid vdd vss serv_rf_top
.ends

