magic
tech gf180mcuD
magscale 1 5
timestamp 1700578260
<< obsm1 >>
rect 672 1538 19320 48246
<< metal2 >>
rect 4928 49600 4984 50000
rect 14896 49600 14952 50000
rect 4928 0 4984 400
rect 14896 0 14952 400
<< obsm2 >>
rect 798 49570 4898 49600
rect 5014 49570 14866 49600
rect 14982 49570 19194 49600
rect 798 430 19194 49570
rect 798 400 4898 430
rect 5014 400 14866 430
rect 14982 400 19194 430
<< metal3 >>
rect 0 47600 400 47656
rect 0 47040 400 47096
rect 0 46480 400 46536
rect 0 45920 400 45976
rect 0 45360 400 45416
rect 0 44800 400 44856
rect 0 44240 400 44296
rect 0 43680 400 43736
rect 0 43120 400 43176
rect 0 42560 400 42616
rect 0 42000 400 42056
rect 0 41440 400 41496
rect 0 40880 400 40936
rect 0 40320 400 40376
rect 0 39760 400 39816
rect 0 39200 400 39256
rect 0 38640 400 38696
rect 0 38080 400 38136
rect 0 37520 400 37576
rect 0 36960 400 37016
rect 0 36400 400 36456
rect 0 35840 400 35896
rect 0 35280 400 35336
rect 0 34720 400 34776
rect 0 34160 400 34216
rect 0 33600 400 33656
rect 0 33040 400 33096
rect 0 32480 400 32536
rect 0 31920 400 31976
rect 0 31360 400 31416
rect 0 30800 400 30856
rect 0 30240 400 30296
rect 0 29680 400 29736
rect 0 29120 400 29176
rect 0 28560 400 28616
rect 0 28000 400 28056
rect 0 27440 400 27496
rect 0 26880 400 26936
rect 0 26320 400 26376
rect 0 25760 400 25816
rect 0 25200 400 25256
rect 0 24640 400 24696
rect 0 24080 400 24136
rect 0 23520 400 23576
rect 0 22960 400 23016
rect 0 22400 400 22456
rect 0 21840 400 21896
rect 0 21280 400 21336
rect 0 20720 400 20776
rect 0 20160 400 20216
rect 0 19600 400 19656
rect 0 19040 400 19096
rect 0 18480 400 18536
rect 0 17920 400 17976
rect 0 17360 400 17416
rect 0 16800 400 16856
rect 0 16240 400 16296
rect 0 15680 400 15736
rect 0 15120 400 15176
rect 0 14560 400 14616
rect 0 14000 400 14056
rect 0 13440 400 13496
rect 0 12880 400 12936
rect 0 12320 400 12376
rect 0 11760 400 11816
rect 0 11200 400 11256
rect 0 10640 400 10696
rect 0 10080 400 10136
rect 0 9520 400 9576
rect 0 8960 400 9016
rect 0 8400 400 8456
rect 0 7840 400 7896
rect 0 7280 400 7336
rect 0 6720 400 6776
rect 0 6160 400 6216
rect 0 5600 400 5656
rect 0 5040 400 5096
rect 0 4480 400 4536
rect 0 3920 400 3976
rect 0 3360 400 3416
rect 0 2800 400 2856
rect 0 2240 400 2296
<< obsm3 >>
rect 400 47686 19199 48230
rect 430 47570 19199 47686
rect 400 47126 19199 47570
rect 430 47010 19199 47126
rect 400 46566 19199 47010
rect 430 46450 19199 46566
rect 400 46006 19199 46450
rect 430 45890 19199 46006
rect 400 45446 19199 45890
rect 430 45330 19199 45446
rect 400 44886 19199 45330
rect 430 44770 19199 44886
rect 400 44326 19199 44770
rect 430 44210 19199 44326
rect 400 43766 19199 44210
rect 430 43650 19199 43766
rect 400 43206 19199 43650
rect 430 43090 19199 43206
rect 400 42646 19199 43090
rect 430 42530 19199 42646
rect 400 42086 19199 42530
rect 430 41970 19199 42086
rect 400 41526 19199 41970
rect 430 41410 19199 41526
rect 400 40966 19199 41410
rect 430 40850 19199 40966
rect 400 40406 19199 40850
rect 430 40290 19199 40406
rect 400 39846 19199 40290
rect 430 39730 19199 39846
rect 400 39286 19199 39730
rect 430 39170 19199 39286
rect 400 38726 19199 39170
rect 430 38610 19199 38726
rect 400 38166 19199 38610
rect 430 38050 19199 38166
rect 400 37606 19199 38050
rect 430 37490 19199 37606
rect 400 37046 19199 37490
rect 430 36930 19199 37046
rect 400 36486 19199 36930
rect 430 36370 19199 36486
rect 400 35926 19199 36370
rect 430 35810 19199 35926
rect 400 35366 19199 35810
rect 430 35250 19199 35366
rect 400 34806 19199 35250
rect 430 34690 19199 34806
rect 400 34246 19199 34690
rect 430 34130 19199 34246
rect 400 33686 19199 34130
rect 430 33570 19199 33686
rect 400 33126 19199 33570
rect 430 33010 19199 33126
rect 400 32566 19199 33010
rect 430 32450 19199 32566
rect 400 32006 19199 32450
rect 430 31890 19199 32006
rect 400 31446 19199 31890
rect 430 31330 19199 31446
rect 400 30886 19199 31330
rect 430 30770 19199 30886
rect 400 30326 19199 30770
rect 430 30210 19199 30326
rect 400 29766 19199 30210
rect 430 29650 19199 29766
rect 400 29206 19199 29650
rect 430 29090 19199 29206
rect 400 28646 19199 29090
rect 430 28530 19199 28646
rect 400 28086 19199 28530
rect 430 27970 19199 28086
rect 400 27526 19199 27970
rect 430 27410 19199 27526
rect 400 26966 19199 27410
rect 430 26850 19199 26966
rect 400 26406 19199 26850
rect 430 26290 19199 26406
rect 400 25846 19199 26290
rect 430 25730 19199 25846
rect 400 25286 19199 25730
rect 430 25170 19199 25286
rect 400 24726 19199 25170
rect 430 24610 19199 24726
rect 400 24166 19199 24610
rect 430 24050 19199 24166
rect 400 23606 19199 24050
rect 430 23490 19199 23606
rect 400 23046 19199 23490
rect 430 22930 19199 23046
rect 400 22486 19199 22930
rect 430 22370 19199 22486
rect 400 21926 19199 22370
rect 430 21810 19199 21926
rect 400 21366 19199 21810
rect 430 21250 19199 21366
rect 400 20806 19199 21250
rect 430 20690 19199 20806
rect 400 20246 19199 20690
rect 430 20130 19199 20246
rect 400 19686 19199 20130
rect 430 19570 19199 19686
rect 400 19126 19199 19570
rect 430 19010 19199 19126
rect 400 18566 19199 19010
rect 430 18450 19199 18566
rect 400 18006 19199 18450
rect 430 17890 19199 18006
rect 400 17446 19199 17890
rect 430 17330 19199 17446
rect 400 16886 19199 17330
rect 430 16770 19199 16886
rect 400 16326 19199 16770
rect 430 16210 19199 16326
rect 400 15766 19199 16210
rect 430 15650 19199 15766
rect 400 15206 19199 15650
rect 430 15090 19199 15206
rect 400 14646 19199 15090
rect 430 14530 19199 14646
rect 400 14086 19199 14530
rect 430 13970 19199 14086
rect 400 13526 19199 13970
rect 430 13410 19199 13526
rect 400 12966 19199 13410
rect 430 12850 19199 12966
rect 400 12406 19199 12850
rect 430 12290 19199 12406
rect 400 11846 19199 12290
rect 430 11730 19199 11846
rect 400 11286 19199 11730
rect 430 11170 19199 11286
rect 400 10726 19199 11170
rect 430 10610 19199 10726
rect 400 10166 19199 10610
rect 430 10050 19199 10166
rect 400 9606 19199 10050
rect 430 9490 19199 9606
rect 400 9046 19199 9490
rect 430 8930 19199 9046
rect 400 8486 19199 8930
rect 430 8370 19199 8486
rect 400 7926 19199 8370
rect 430 7810 19199 7926
rect 400 7366 19199 7810
rect 430 7250 19199 7366
rect 400 6806 19199 7250
rect 430 6690 19199 6806
rect 400 6246 19199 6690
rect 430 6130 19199 6246
rect 400 5686 19199 6130
rect 430 5570 19199 5686
rect 400 5126 19199 5570
rect 430 5010 19199 5126
rect 400 4566 19199 5010
rect 430 4450 19199 4566
rect 400 4006 19199 4450
rect 430 3890 19199 4006
rect 400 3446 19199 3890
rect 430 3330 19199 3446
rect 400 2886 19199 3330
rect 430 2770 19199 2886
rect 400 2326 19199 2770
rect 430 2210 19199 2326
rect 400 1554 19199 2210
<< metal4 >>
rect 1994 1538 2614 48246
rect 6994 1538 7614 48246
rect 11994 1538 12614 48246
rect 16994 1538 17614 48246
<< obsm4 >>
rect 910 5721 1964 43335
rect 2644 5721 6964 43335
rect 7644 5721 11964 43335
rect 12644 5721 16964 43335
rect 17644 5721 17682 43335
<< labels >>
rlabel metal4 s 1994 1538 2614 48246 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 11994 1538 12614 48246 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 6994 1538 7614 48246 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 16994 1538 17614 48246 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 14896 0 14952 400 6 mclk
port 3 nsew signal input
rlabel metal3 s 0 47600 400 47656 6 reg_ack
port 4 nsew signal output
rlabel metal3 s 0 8960 400 9016 6 reg_addr[0]
port 5 nsew signal input
rlabel metal3 s 0 3360 400 3416 6 reg_addr[10]
port 6 nsew signal input
rlabel metal3 s 0 8400 400 8456 6 reg_addr[1]
port 7 nsew signal input
rlabel metal3 s 0 7840 400 7896 6 reg_addr[2]
port 8 nsew signal input
rlabel metal3 s 0 7280 400 7336 6 reg_addr[3]
port 9 nsew signal input
rlabel metal3 s 0 6720 400 6776 6 reg_addr[4]
port 10 nsew signal input
rlabel metal3 s 0 6160 400 6216 6 reg_addr[5]
port 11 nsew signal input
rlabel metal3 s 0 5600 400 5656 6 reg_addr[6]
port 12 nsew signal input
rlabel metal3 s 0 5040 400 5096 6 reg_addr[7]
port 13 nsew signal input
rlabel metal3 s 0 4480 400 4536 6 reg_addr[8]
port 14 nsew signal input
rlabel metal3 s 0 3920 400 3976 6 reg_addr[9]
port 15 nsew signal input
rlabel metal3 s 0 11200 400 11256 6 reg_be[0]
port 16 nsew signal input
rlabel metal3 s 0 10640 400 10696 6 reg_be[1]
port 17 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 reg_be[2]
port 18 nsew signal input
rlabel metal3 s 0 9520 400 9576 6 reg_be[3]
port 19 nsew signal input
rlabel metal3 s 0 2240 400 2296 6 reg_cs
port 20 nsew signal input
rlabel metal3 s 0 47040 400 47096 6 reg_rdata[0]
port 21 nsew signal output
rlabel metal3 s 0 41440 400 41496 6 reg_rdata[10]
port 22 nsew signal output
rlabel metal3 s 0 40880 400 40936 6 reg_rdata[11]
port 23 nsew signal output
rlabel metal3 s 0 40320 400 40376 6 reg_rdata[12]
port 24 nsew signal output
rlabel metal3 s 0 39760 400 39816 6 reg_rdata[13]
port 25 nsew signal output
rlabel metal3 s 0 39200 400 39256 6 reg_rdata[14]
port 26 nsew signal output
rlabel metal3 s 0 38640 400 38696 6 reg_rdata[15]
port 27 nsew signal output
rlabel metal3 s 0 38080 400 38136 6 reg_rdata[16]
port 28 nsew signal output
rlabel metal3 s 0 37520 400 37576 6 reg_rdata[17]
port 29 nsew signal output
rlabel metal3 s 0 36960 400 37016 6 reg_rdata[18]
port 30 nsew signal output
rlabel metal3 s 0 36400 400 36456 6 reg_rdata[19]
port 31 nsew signal output
rlabel metal3 s 0 46480 400 46536 6 reg_rdata[1]
port 32 nsew signal output
rlabel metal3 s 0 35840 400 35896 6 reg_rdata[20]
port 33 nsew signal output
rlabel metal3 s 0 35280 400 35336 6 reg_rdata[21]
port 34 nsew signal output
rlabel metal3 s 0 34720 400 34776 6 reg_rdata[22]
port 35 nsew signal output
rlabel metal3 s 0 34160 400 34216 6 reg_rdata[23]
port 36 nsew signal output
rlabel metal3 s 0 33600 400 33656 6 reg_rdata[24]
port 37 nsew signal output
rlabel metal3 s 0 33040 400 33096 6 reg_rdata[25]
port 38 nsew signal output
rlabel metal3 s 0 32480 400 32536 6 reg_rdata[26]
port 39 nsew signal output
rlabel metal3 s 0 31920 400 31976 6 reg_rdata[27]
port 40 nsew signal output
rlabel metal3 s 0 31360 400 31416 6 reg_rdata[28]
port 41 nsew signal output
rlabel metal3 s 0 30800 400 30856 6 reg_rdata[29]
port 42 nsew signal output
rlabel metal3 s 0 45920 400 45976 6 reg_rdata[2]
port 43 nsew signal output
rlabel metal3 s 0 30240 400 30296 6 reg_rdata[30]
port 44 nsew signal output
rlabel metal3 s 0 29680 400 29736 6 reg_rdata[31]
port 45 nsew signal output
rlabel metal3 s 0 45360 400 45416 6 reg_rdata[3]
port 46 nsew signal output
rlabel metal3 s 0 44800 400 44856 6 reg_rdata[4]
port 47 nsew signal output
rlabel metal3 s 0 44240 400 44296 6 reg_rdata[5]
port 48 nsew signal output
rlabel metal3 s 0 43680 400 43736 6 reg_rdata[6]
port 49 nsew signal output
rlabel metal3 s 0 43120 400 43176 6 reg_rdata[7]
port 50 nsew signal output
rlabel metal3 s 0 42560 400 42616 6 reg_rdata[8]
port 51 nsew signal output
rlabel metal3 s 0 42000 400 42056 6 reg_rdata[9]
port 52 nsew signal output
rlabel metal3 s 0 29120 400 29176 6 reg_wdata[0]
port 53 nsew signal input
rlabel metal3 s 0 23520 400 23576 6 reg_wdata[10]
port 54 nsew signal input
rlabel metal3 s 0 22960 400 23016 6 reg_wdata[11]
port 55 nsew signal input
rlabel metal3 s 0 22400 400 22456 6 reg_wdata[12]
port 56 nsew signal input
rlabel metal3 s 0 21840 400 21896 6 reg_wdata[13]
port 57 nsew signal input
rlabel metal3 s 0 21280 400 21336 6 reg_wdata[14]
port 58 nsew signal input
rlabel metal3 s 0 20720 400 20776 6 reg_wdata[15]
port 59 nsew signal input
rlabel metal3 s 0 20160 400 20216 6 reg_wdata[16]
port 60 nsew signal input
rlabel metal3 s 0 19600 400 19656 6 reg_wdata[17]
port 61 nsew signal input
rlabel metal3 s 0 19040 400 19096 6 reg_wdata[18]
port 62 nsew signal input
rlabel metal3 s 0 18480 400 18536 6 reg_wdata[19]
port 63 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 reg_wdata[1]
port 64 nsew signal input
rlabel metal3 s 0 17920 400 17976 6 reg_wdata[20]
port 65 nsew signal input
rlabel metal3 s 0 17360 400 17416 6 reg_wdata[21]
port 66 nsew signal input
rlabel metal3 s 0 16800 400 16856 6 reg_wdata[22]
port 67 nsew signal input
rlabel metal3 s 0 16240 400 16296 6 reg_wdata[23]
port 68 nsew signal input
rlabel metal3 s 0 15680 400 15736 6 reg_wdata[24]
port 69 nsew signal input
rlabel metal3 s 0 15120 400 15176 6 reg_wdata[25]
port 70 nsew signal input
rlabel metal3 s 0 14560 400 14616 6 reg_wdata[26]
port 71 nsew signal input
rlabel metal3 s 0 14000 400 14056 6 reg_wdata[27]
port 72 nsew signal input
rlabel metal3 s 0 13440 400 13496 6 reg_wdata[28]
port 73 nsew signal input
rlabel metal3 s 0 12880 400 12936 6 reg_wdata[29]
port 74 nsew signal input
rlabel metal3 s 0 28000 400 28056 6 reg_wdata[2]
port 75 nsew signal input
rlabel metal3 s 0 12320 400 12376 6 reg_wdata[30]
port 76 nsew signal input
rlabel metal3 s 0 11760 400 11816 6 reg_wdata[31]
port 77 nsew signal input
rlabel metal3 s 0 27440 400 27496 6 reg_wdata[3]
port 78 nsew signal input
rlabel metal3 s 0 26880 400 26936 6 reg_wdata[4]
port 79 nsew signal input
rlabel metal3 s 0 26320 400 26376 6 reg_wdata[5]
port 80 nsew signal input
rlabel metal3 s 0 25760 400 25816 6 reg_wdata[6]
port 81 nsew signal input
rlabel metal3 s 0 25200 400 25256 6 reg_wdata[7]
port 82 nsew signal input
rlabel metal3 s 0 24640 400 24696 6 reg_wdata[8]
port 83 nsew signal input
rlabel metal3 s 0 24080 400 24136 6 reg_wdata[9]
port 84 nsew signal input
rlabel metal3 s 0 2800 400 2856 6 reg_wr
port 85 nsew signal input
rlabel metal2 s 4928 49600 4984 50000 6 rtc_clk
port 86 nsew signal input
rlabel metal2 s 14896 49600 14952 50000 6 rtc_intr
port 87 nsew signal output
rlabel metal2 s 4928 0 4984 400 6 s_reset_n
port 88 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3338868
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/peri_top/runs/23_11_21_16_46/results/signoff/peri_top.magic.gds
string GDS_START 424868
<< end >>

