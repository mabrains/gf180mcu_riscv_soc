magic
tech gf180mcuD
magscale 1 10
timestamp 1700584328
<< metal1 >>
rect 2482 12686 2494 12738
rect 2546 12735 2558 12738
rect 3042 12735 3054 12738
rect 2546 12689 3054 12735
rect 2546 12686 2558 12689
rect 3042 12686 3054 12689
rect 3106 12686 3118 12738
rect 17154 12686 17166 12738
rect 17218 12735 17230 12738
rect 19170 12735 19182 12738
rect 17218 12689 19182 12735
rect 17218 12686 17230 12689
rect 19170 12686 19182 12689
rect 19234 12686 19246 12738
rect 1344 12570 18752 12604
rect 1344 12518 5526 12570
rect 5578 12518 5630 12570
rect 5682 12518 5734 12570
rect 5786 12518 9838 12570
rect 9890 12518 9942 12570
rect 9994 12518 10046 12570
rect 10098 12518 14150 12570
rect 14202 12518 14254 12570
rect 14306 12518 14358 12570
rect 14410 12518 18462 12570
rect 18514 12518 18566 12570
rect 18618 12518 18670 12570
rect 18722 12518 18752 12570
rect 1344 12484 18752 12518
rect 4286 12402 4338 12414
rect 4286 12338 4338 12350
rect 4734 12402 4786 12414
rect 4734 12338 4786 12350
rect 7646 12402 7698 12414
rect 7646 12338 7698 12350
rect 16382 12402 16434 12414
rect 16382 12338 16434 12350
rect 1710 12290 1762 12302
rect 1710 12226 1762 12238
rect 2158 12290 2210 12302
rect 15822 12290 15874 12302
rect 17838 12290 17890 12302
rect 3042 12238 3054 12290
rect 3106 12238 3118 12290
rect 17154 12238 17166 12290
rect 17218 12238 17230 12290
rect 2158 12226 2210 12238
rect 15822 12226 15874 12238
rect 17838 12226 17890 12238
rect 14926 12178 14978 12190
rect 3938 12126 3950 12178
rect 4002 12126 4014 12178
rect 13234 12126 13246 12178
rect 13298 12126 13310 12178
rect 14926 12114 14978 12126
rect 17502 12178 17554 12190
rect 18050 12126 18062 12178
rect 18114 12126 18126 12178
rect 17502 12114 17554 12126
rect 5630 12066 5682 12078
rect 5630 12002 5682 12014
rect 6078 12066 6130 12078
rect 6078 12002 6130 12014
rect 6638 12066 6690 12078
rect 6638 12002 6690 12014
rect 12238 12066 12290 12078
rect 12238 12002 12290 12014
rect 12686 12066 12738 12078
rect 14478 12066 14530 12078
rect 13570 12014 13582 12066
rect 13634 12014 13646 12066
rect 12686 12002 12738 12014
rect 14478 12002 14530 12014
rect 15374 12066 15426 12078
rect 15374 12002 15426 12014
rect 1344 11786 18592 11820
rect 1344 11734 3370 11786
rect 3422 11734 3474 11786
rect 3526 11734 3578 11786
rect 3630 11734 7682 11786
rect 7734 11734 7786 11786
rect 7838 11734 7890 11786
rect 7942 11734 11994 11786
rect 12046 11734 12098 11786
rect 12150 11734 12202 11786
rect 12254 11734 16306 11786
rect 16358 11734 16410 11786
rect 16462 11734 16514 11786
rect 16566 11734 18592 11786
rect 1344 11700 18592 11734
rect 16818 11454 16830 11506
rect 16882 11454 16894 11506
rect 14814 11394 14866 11406
rect 16930 11342 16942 11394
rect 16994 11342 17006 11394
rect 14814 11330 14866 11342
rect 2158 11282 2210 11294
rect 2158 11218 2210 11230
rect 2606 11282 2658 11294
rect 2606 11218 2658 11230
rect 3054 11282 3106 11294
rect 3054 11218 3106 11230
rect 3502 11282 3554 11294
rect 3502 11218 3554 11230
rect 13694 11282 13746 11294
rect 13694 11218 13746 11230
rect 16046 11282 16098 11294
rect 16046 11218 16098 11230
rect 16382 11282 16434 11294
rect 16382 11218 16434 11230
rect 17726 11282 17778 11294
rect 17726 11218 17778 11230
rect 18062 11282 18114 11294
rect 18062 11218 18114 11230
rect 1710 11170 1762 11182
rect 1710 11106 1762 11118
rect 4510 11170 4562 11182
rect 4510 11106 4562 11118
rect 4958 11170 5010 11182
rect 4958 11106 5010 11118
rect 5854 11170 5906 11182
rect 5854 11106 5906 11118
rect 6302 11170 6354 11182
rect 6302 11106 6354 11118
rect 6638 11170 6690 11182
rect 6638 11106 6690 11118
rect 7086 11170 7138 11182
rect 7086 11106 7138 11118
rect 7534 11170 7586 11182
rect 7534 11106 7586 11118
rect 11678 11170 11730 11182
rect 11678 11106 11730 11118
rect 12126 11170 12178 11182
rect 12126 11106 12178 11118
rect 12574 11170 12626 11182
rect 12574 11106 12626 11118
rect 13022 11170 13074 11182
rect 13022 11106 13074 11118
rect 14142 11170 14194 11182
rect 14142 11106 14194 11118
rect 15150 11170 15202 11182
rect 15698 11118 15710 11170
rect 15762 11118 15774 11170
rect 15150 11106 15202 11118
rect 1344 11002 18752 11036
rect 1344 10950 5526 11002
rect 5578 10950 5630 11002
rect 5682 10950 5734 11002
rect 5786 10950 9838 11002
rect 9890 10950 9942 11002
rect 9994 10950 10046 11002
rect 10098 10950 14150 11002
rect 14202 10950 14254 11002
rect 14306 10950 14358 11002
rect 14410 10950 18462 11002
rect 18514 10950 18566 11002
rect 18618 10950 18670 11002
rect 18722 10950 18752 11002
rect 1344 10916 18752 10950
rect 2158 10834 2210 10846
rect 2158 10770 2210 10782
rect 13694 10834 13746 10846
rect 13694 10770 13746 10782
rect 17390 10834 17442 10846
rect 17390 10770 17442 10782
rect 1710 10722 1762 10734
rect 1710 10658 1762 10670
rect 2606 10722 2658 10734
rect 2606 10658 2658 10670
rect 3054 10722 3106 10734
rect 3054 10658 3106 10670
rect 3502 10722 3554 10734
rect 3502 10658 3554 10670
rect 8990 10722 9042 10734
rect 8990 10658 9042 10670
rect 10670 10722 10722 10734
rect 10670 10658 10722 10670
rect 14702 10722 14754 10734
rect 14702 10658 14754 10670
rect 15374 10722 15426 10734
rect 15374 10658 15426 10670
rect 16158 10722 16210 10734
rect 16158 10658 16210 10670
rect 16830 10722 16882 10734
rect 16830 10658 16882 10670
rect 8206 10610 8258 10622
rect 6850 10558 6862 10610
rect 6914 10558 6926 10610
rect 8206 10546 8258 10558
rect 11678 10610 11730 10622
rect 11678 10546 11730 10558
rect 13134 10610 13186 10622
rect 13134 10546 13186 10558
rect 13582 10610 13634 10622
rect 13582 10546 13634 10558
rect 13806 10610 13858 10622
rect 13806 10546 13858 10558
rect 14366 10610 14418 10622
rect 14366 10546 14418 10558
rect 15038 10610 15090 10622
rect 15038 10546 15090 10558
rect 15822 10610 15874 10622
rect 17726 10610 17778 10622
rect 16594 10558 16606 10610
rect 16658 10558 16670 10610
rect 15822 10546 15874 10558
rect 17726 10546 17778 10558
rect 7310 10498 7362 10510
rect 3938 10446 3950 10498
rect 4002 10446 4014 10498
rect 6066 10446 6078 10498
rect 6130 10446 6142 10498
rect 7310 10434 7362 10446
rect 7758 10498 7810 10510
rect 7758 10434 7810 10446
rect 11230 10498 11282 10510
rect 11230 10434 11282 10446
rect 12126 10498 12178 10510
rect 12126 10434 12178 10446
rect 12574 10498 12626 10510
rect 12574 10434 12626 10446
rect 13022 10498 13074 10510
rect 13022 10434 13074 10446
rect 18174 10498 18226 10510
rect 18174 10434 18226 10446
rect 1344 10218 18592 10252
rect 1344 10166 3370 10218
rect 3422 10166 3474 10218
rect 3526 10166 3578 10218
rect 3630 10166 7682 10218
rect 7734 10166 7786 10218
rect 7838 10166 7890 10218
rect 7942 10166 11994 10218
rect 12046 10166 12098 10218
rect 12150 10166 12202 10218
rect 12254 10166 16306 10218
rect 16358 10166 16410 10218
rect 16462 10166 16514 10218
rect 16566 10166 18592 10218
rect 1344 10132 18592 10166
rect 11454 10050 11506 10062
rect 11454 9986 11506 9998
rect 10222 9938 10274 9950
rect 18162 9886 18174 9938
rect 18226 9886 18238 9938
rect 10222 9874 10274 9886
rect 9886 9826 9938 9838
rect 9886 9762 9938 9774
rect 12126 9826 12178 9838
rect 13806 9826 13858 9838
rect 13682 9774 13694 9826
rect 13746 9774 13758 9826
rect 14018 9774 14030 9826
rect 14082 9774 14094 9826
rect 14690 9774 14702 9826
rect 14754 9774 14766 9826
rect 15362 9774 15374 9826
rect 15426 9774 15438 9826
rect 12126 9762 12178 9774
rect 13806 9762 13858 9774
rect 1710 9714 1762 9726
rect 1710 9650 1762 9662
rect 10558 9714 10610 9726
rect 10558 9650 10610 9662
rect 10670 9714 10722 9726
rect 10670 9650 10722 9662
rect 11342 9714 11394 9726
rect 11342 9650 11394 9662
rect 12462 9714 12514 9726
rect 12462 9650 12514 9662
rect 14254 9714 14306 9726
rect 16034 9662 16046 9714
rect 16098 9662 16110 9714
rect 14254 9650 14306 9662
rect 2158 9602 2210 9614
rect 2158 9538 2210 9550
rect 2606 9602 2658 9614
rect 2606 9538 2658 9550
rect 3054 9602 3106 9614
rect 3054 9538 3106 9550
rect 3502 9602 3554 9614
rect 3502 9538 3554 9550
rect 3950 9602 4002 9614
rect 3950 9538 4002 9550
rect 4398 9602 4450 9614
rect 4398 9538 4450 9550
rect 5070 9602 5122 9614
rect 5070 9538 5122 9550
rect 5742 9602 5794 9614
rect 5742 9538 5794 9550
rect 6302 9602 6354 9614
rect 6302 9538 6354 9550
rect 6750 9602 6802 9614
rect 6750 9538 6802 9550
rect 7198 9602 7250 9614
rect 7198 9538 7250 9550
rect 7534 9602 7586 9614
rect 7534 9538 7586 9550
rect 7982 9602 8034 9614
rect 7982 9538 8034 9550
rect 8430 9602 8482 9614
rect 8430 9538 8482 9550
rect 8878 9602 8930 9614
rect 8878 9538 8930 9550
rect 9438 9602 9490 9614
rect 9438 9538 9490 9550
rect 10894 9602 10946 9614
rect 10894 9538 10946 9550
rect 11454 9602 11506 9614
rect 11454 9538 11506 9550
rect 11790 9602 11842 9614
rect 11790 9538 11842 9550
rect 12014 9602 12066 9614
rect 12014 9538 12066 9550
rect 12574 9602 12626 9614
rect 12574 9538 12626 9550
rect 12798 9602 12850 9614
rect 14926 9602 14978 9614
rect 13794 9550 13806 9602
rect 13858 9550 13870 9602
rect 12798 9538 12850 9550
rect 14926 9538 14978 9550
rect 1344 9434 18752 9468
rect 1344 9382 5526 9434
rect 5578 9382 5630 9434
rect 5682 9382 5734 9434
rect 5786 9382 9838 9434
rect 9890 9382 9942 9434
rect 9994 9382 10046 9434
rect 10098 9382 14150 9434
rect 14202 9382 14254 9434
rect 14306 9382 14358 9434
rect 14410 9382 18462 9434
rect 18514 9382 18566 9434
rect 18618 9382 18670 9434
rect 18722 9382 18752 9434
rect 1344 9348 18752 9382
rect 1710 9154 1762 9166
rect 1710 9090 1762 9102
rect 2158 9154 2210 9166
rect 2158 9090 2210 9102
rect 2606 9154 2658 9166
rect 2606 9090 2658 9102
rect 3054 9154 3106 9166
rect 3054 9090 3106 9102
rect 3502 9154 3554 9166
rect 3502 9090 3554 9102
rect 3950 9154 4002 9166
rect 3950 9090 4002 9102
rect 4398 9154 4450 9166
rect 8318 9154 8370 9166
rect 5282 9102 5294 9154
rect 5346 9102 5358 9154
rect 4398 9090 4450 9102
rect 8318 9090 8370 9102
rect 10110 9154 10162 9166
rect 17390 9154 17442 9166
rect 13234 9102 13246 9154
rect 13298 9102 13310 9154
rect 10110 9090 10162 9102
rect 17390 9090 17442 9102
rect 5170 8990 5182 9042
rect 5234 8990 5246 9042
rect 7186 8990 7198 9042
rect 7250 8990 7262 9042
rect 9538 8990 9550 9042
rect 9602 8990 9614 9042
rect 11554 8990 11566 9042
rect 11618 8990 11630 9042
rect 16706 8990 16718 9042
rect 16770 8990 16782 9042
rect 17602 8990 17614 9042
rect 17666 8990 17678 9042
rect 18174 8930 18226 8942
rect 8194 8878 8206 8930
rect 8258 8878 8270 8930
rect 12898 8878 12910 8930
rect 12962 8878 12974 8930
rect 13906 8878 13918 8930
rect 13970 8878 13982 8930
rect 16034 8878 16046 8930
rect 16098 8878 16110 8930
rect 18174 8866 18226 8878
rect 17938 8766 17950 8818
rect 18002 8815 18014 8818
rect 18274 8815 18286 8818
rect 18002 8769 18286 8815
rect 18002 8766 18014 8769
rect 18274 8766 18286 8769
rect 18338 8766 18350 8818
rect 1344 8650 18592 8684
rect 1344 8598 3370 8650
rect 3422 8598 3474 8650
rect 3526 8598 3578 8650
rect 3630 8598 7682 8650
rect 7734 8598 7786 8650
rect 7838 8598 7890 8650
rect 7942 8598 11994 8650
rect 12046 8598 12098 8650
rect 12150 8598 12202 8650
rect 12254 8598 16306 8650
rect 16358 8598 16410 8650
rect 16462 8598 16514 8650
rect 16566 8598 18592 8650
rect 1344 8564 18592 8598
rect 16830 8370 16882 8382
rect 13458 8318 13470 8370
rect 13522 8318 13534 8370
rect 16830 8306 16882 8318
rect 2146 8206 2158 8258
rect 2210 8206 2222 8258
rect 7186 8206 7198 8258
rect 7250 8206 7262 8258
rect 12114 8206 12126 8258
rect 12178 8206 12190 8258
rect 16258 8206 16270 8258
rect 16322 8206 16334 8258
rect 2382 8146 2434 8158
rect 2382 8082 2434 8094
rect 4174 8146 4226 8158
rect 4174 8082 4226 8094
rect 4622 8146 4674 8158
rect 4622 8082 4674 8094
rect 5630 8146 5682 8158
rect 16718 8146 16770 8158
rect 7858 8094 7870 8146
rect 7922 8094 7934 8146
rect 15586 8094 15598 8146
rect 15650 8094 15662 8146
rect 5630 8082 5682 8094
rect 16718 8082 16770 8094
rect 17054 8146 17106 8158
rect 17054 8082 17106 8094
rect 17278 8146 17330 8158
rect 17278 8082 17330 8094
rect 17950 8146 18002 8158
rect 17950 8082 18002 8094
rect 3054 8034 3106 8046
rect 3054 7970 3106 7982
rect 3502 8034 3554 8046
rect 3502 7970 3554 7982
rect 4286 8034 4338 8046
rect 4286 7970 4338 7982
rect 4734 8034 4786 8046
rect 4734 7970 4786 7982
rect 5966 8034 6018 8046
rect 5966 7970 6018 7982
rect 6302 8034 6354 8046
rect 6302 7970 6354 7982
rect 6974 8034 7026 8046
rect 6974 7970 7026 7982
rect 17614 8034 17666 8046
rect 17614 7970 17666 7982
rect 1344 7866 18752 7900
rect 1344 7814 5526 7866
rect 5578 7814 5630 7866
rect 5682 7814 5734 7866
rect 5786 7814 9838 7866
rect 9890 7814 9942 7866
rect 9994 7814 10046 7866
rect 10098 7814 14150 7866
rect 14202 7814 14254 7866
rect 14306 7814 14358 7866
rect 14410 7814 18462 7866
rect 18514 7814 18566 7866
rect 18618 7814 18670 7866
rect 18722 7814 18752 7866
rect 1344 7780 18752 7814
rect 2046 7698 2098 7710
rect 2046 7634 2098 7646
rect 2718 7698 2770 7710
rect 2718 7634 2770 7646
rect 3614 7698 3666 7710
rect 7634 7646 7646 7698
rect 7698 7646 7710 7698
rect 3614 7634 3666 7646
rect 1710 7586 1762 7598
rect 1710 7522 1762 7534
rect 3278 7586 3330 7598
rect 3278 7522 3330 7534
rect 4734 7586 4786 7598
rect 4734 7522 4786 7534
rect 6750 7586 6802 7598
rect 6750 7522 6802 7534
rect 9998 7586 10050 7598
rect 9998 7522 10050 7534
rect 10782 7586 10834 7598
rect 17390 7586 17442 7598
rect 12114 7534 12126 7586
rect 12178 7534 12190 7586
rect 10782 7522 10834 7534
rect 17390 7522 17442 7534
rect 17502 7586 17554 7598
rect 17602 7534 17614 7586
rect 17666 7534 17678 7586
rect 17502 7522 17554 7534
rect 8094 7474 8146 7486
rect 2482 7422 2494 7474
rect 2546 7422 2558 7474
rect 4050 7422 4062 7474
rect 4114 7422 4126 7474
rect 7858 7422 7870 7474
rect 7922 7422 7934 7474
rect 8094 7410 8146 7422
rect 8542 7474 8594 7486
rect 8542 7410 8594 7422
rect 8766 7474 8818 7486
rect 8766 7410 8818 7422
rect 9662 7474 9714 7486
rect 9662 7410 9714 7422
rect 10446 7474 10498 7486
rect 16706 7422 16718 7474
rect 16770 7422 16782 7474
rect 17938 7422 17950 7474
rect 18002 7422 18014 7474
rect 10446 7410 10498 7422
rect 8654 7362 8706 7374
rect 8654 7298 8706 7310
rect 11230 7362 11282 7374
rect 11230 7298 11282 7310
rect 17838 7250 17890 7262
rect 17838 7186 17890 7198
rect 1344 7082 18592 7116
rect 1344 7030 3370 7082
rect 3422 7030 3474 7082
rect 3526 7030 3578 7082
rect 3630 7030 7682 7082
rect 7734 7030 7786 7082
rect 7838 7030 7890 7082
rect 7942 7030 11994 7082
rect 12046 7030 12098 7082
rect 12150 7030 12202 7082
rect 12254 7030 16306 7082
rect 16358 7030 16410 7082
rect 16462 7030 16514 7082
rect 16566 7030 18592 7082
rect 1344 6996 18592 7030
rect 12574 6914 12626 6926
rect 12574 6850 12626 6862
rect 12910 6914 12962 6926
rect 12910 6850 12962 6862
rect 1822 6690 1874 6702
rect 1822 6626 1874 6638
rect 2494 6690 2546 6702
rect 2494 6626 2546 6638
rect 3054 6690 3106 6702
rect 4622 6690 4674 6702
rect 3938 6638 3950 6690
rect 4002 6638 4014 6690
rect 3054 6626 3106 6638
rect 4622 6626 4674 6638
rect 4846 6690 4898 6702
rect 4846 6626 4898 6638
rect 4958 6690 5010 6702
rect 13470 6690 13522 6702
rect 5730 6638 5742 6690
rect 5794 6638 5806 6690
rect 7634 6638 7646 6690
rect 7698 6638 7710 6690
rect 9650 6638 9662 6690
rect 9714 6638 9726 6690
rect 12114 6638 12126 6690
rect 12178 6638 12190 6690
rect 4958 6626 5010 6638
rect 13470 6626 13522 6638
rect 13806 6690 13858 6702
rect 13806 6626 13858 6638
rect 14030 6690 14082 6702
rect 14354 6638 14366 6690
rect 14418 6638 14430 6690
rect 18162 6638 18174 6690
rect 18226 6638 18238 6690
rect 14030 6626 14082 6638
rect 3390 6578 3442 6590
rect 5070 6578 5122 6590
rect 2146 6526 2158 6578
rect 2210 6526 2222 6578
rect 4162 6526 4174 6578
rect 4226 6526 4238 6578
rect 3390 6514 3442 6526
rect 5070 6514 5122 6526
rect 6414 6578 6466 6590
rect 6414 6514 6466 6526
rect 6526 6578 6578 6590
rect 6526 6514 6578 6526
rect 7086 6578 7138 6590
rect 7086 6514 7138 6526
rect 7198 6578 7250 6590
rect 7198 6514 7250 6526
rect 7422 6578 7474 6590
rect 15038 6578 15090 6590
rect 17054 6578 17106 6590
rect 7746 6526 7758 6578
rect 7810 6526 7822 6578
rect 11442 6526 11454 6578
rect 11506 6526 11518 6578
rect 16258 6526 16270 6578
rect 16322 6526 16334 6578
rect 7422 6514 7474 6526
rect 15038 6514 15090 6526
rect 17054 6514 17106 6526
rect 3502 6466 3554 6478
rect 3502 6402 3554 6414
rect 5966 6466 6018 6478
rect 5966 6402 6018 6414
rect 6190 6466 6242 6478
rect 11902 6466 11954 6478
rect 8642 6414 8654 6466
rect 8706 6414 8718 6466
rect 6190 6402 6242 6414
rect 11902 6402 11954 6414
rect 12798 6466 12850 6478
rect 12798 6402 12850 6414
rect 13694 6466 13746 6478
rect 13694 6402 13746 6414
rect 1344 6298 18752 6332
rect 1344 6246 5526 6298
rect 5578 6246 5630 6298
rect 5682 6246 5734 6298
rect 5786 6246 9838 6298
rect 9890 6246 9942 6298
rect 9994 6246 10046 6298
rect 10098 6246 14150 6298
rect 14202 6246 14254 6298
rect 14306 6246 14358 6298
rect 14410 6246 18462 6298
rect 18514 6246 18566 6298
rect 18618 6246 18670 6298
rect 18722 6246 18752 6298
rect 1344 6212 18752 6246
rect 1822 6130 1874 6142
rect 3502 6130 3554 6142
rect 2818 6078 2830 6130
rect 2882 6078 2894 6130
rect 1822 6066 1874 6078
rect 3502 6066 3554 6078
rect 17390 6130 17442 6142
rect 17390 6066 17442 6078
rect 17502 6130 17554 6142
rect 17502 6066 17554 6078
rect 17614 6130 17666 6142
rect 17614 6066 17666 6078
rect 3838 6018 3890 6030
rect 2146 5966 2158 6018
rect 2210 5966 2222 6018
rect 3838 5954 3890 5966
rect 4174 6018 4226 6030
rect 4174 5954 4226 5966
rect 4846 6018 4898 6030
rect 4846 5954 4898 5966
rect 5854 6018 5906 6030
rect 5854 5954 5906 5966
rect 7870 6018 7922 6030
rect 7870 5954 7922 5966
rect 9886 6018 9938 6030
rect 9886 5954 9938 5966
rect 10222 6018 10274 6030
rect 10222 5954 10274 5966
rect 11230 6018 11282 6030
rect 16146 5966 16158 6018
rect 16210 5966 16222 6018
rect 11230 5954 11282 5966
rect 4510 5906 4562 5918
rect 2594 5854 2606 5906
rect 2658 5854 2670 5906
rect 3266 5854 3278 5906
rect 3330 5854 3342 5906
rect 4510 5842 4562 5854
rect 5294 5906 5346 5918
rect 5294 5842 5346 5854
rect 7310 5906 7362 5918
rect 10994 5854 11006 5906
rect 11058 5854 11070 5906
rect 12338 5854 12350 5906
rect 12402 5854 12414 5906
rect 17938 5854 17950 5906
rect 18002 5854 18014 5906
rect 7310 5842 7362 5854
rect 6738 5742 6750 5794
rect 6802 5742 6814 5794
rect 1344 5514 18592 5548
rect 1344 5462 3370 5514
rect 3422 5462 3474 5514
rect 3526 5462 3578 5514
rect 3630 5462 7682 5514
rect 7734 5462 7786 5514
rect 7838 5462 7890 5514
rect 7942 5462 11994 5514
rect 12046 5462 12098 5514
rect 12150 5462 12202 5514
rect 12254 5462 16306 5514
rect 16358 5462 16410 5514
rect 16462 5462 16514 5514
rect 16566 5462 18592 5514
rect 1344 5428 18592 5462
rect 8754 5182 8766 5234
rect 8818 5182 8830 5234
rect 1822 5122 1874 5134
rect 4734 5122 4786 5134
rect 2818 5070 2830 5122
rect 2882 5070 2894 5122
rect 3490 5070 3502 5122
rect 3554 5070 3566 5122
rect 5954 5082 5966 5134
rect 6018 5082 6030 5134
rect 15598 5122 15650 5134
rect 9090 5070 9102 5122
rect 9154 5070 9166 5122
rect 11330 5070 11342 5122
rect 11394 5070 11406 5122
rect 13458 5070 13470 5122
rect 13522 5070 13534 5122
rect 1822 5058 1874 5070
rect 4734 5058 4786 5070
rect 15598 5058 15650 5070
rect 17950 5122 18002 5134
rect 17950 5058 18002 5070
rect 3054 5010 3106 5022
rect 2146 4958 2158 5010
rect 2210 4958 2222 5010
rect 3054 4946 3106 4958
rect 3726 5010 3778 5022
rect 3726 4946 3778 4958
rect 4062 5010 4114 5022
rect 4062 4946 4114 4958
rect 4398 5010 4450 5022
rect 4398 4946 4450 4958
rect 5070 5010 5122 5022
rect 9774 5010 9826 5022
rect 6626 4958 6638 5010
rect 6690 4958 6702 5010
rect 5070 4946 5122 4958
rect 9774 4946 9826 4958
rect 12350 5010 12402 5022
rect 12350 4946 12402 4958
rect 14142 5010 14194 5022
rect 14142 4946 14194 4958
rect 16718 5010 16770 5022
rect 16718 4946 16770 4958
rect 17614 5010 17666 5022
rect 17614 4946 17666 4958
rect 11330 4846 11342 4898
rect 11394 4846 11406 4898
rect 15810 4846 15822 4898
rect 15874 4846 15886 4898
rect 1344 4730 18752 4764
rect 1344 4678 5526 4730
rect 5578 4678 5630 4730
rect 5682 4678 5734 4730
rect 5786 4678 9838 4730
rect 9890 4678 9942 4730
rect 9994 4678 10046 4730
rect 10098 4678 14150 4730
rect 14202 4678 14254 4730
rect 14306 4678 14358 4730
rect 14410 4678 18462 4730
rect 18514 4678 18566 4730
rect 18618 4678 18670 4730
rect 18722 4678 18752 4730
rect 1344 4644 18752 4678
rect 2942 4562 2994 4574
rect 2942 4498 2994 4510
rect 4958 4562 5010 4574
rect 4958 4498 5010 4510
rect 9662 4562 9714 4574
rect 17390 4562 17442 4574
rect 14914 4510 14926 4562
rect 14978 4510 14990 4562
rect 9662 4498 9714 4510
rect 17390 4498 17442 4510
rect 18174 4562 18226 4574
rect 18174 4498 18226 4510
rect 5742 4450 5794 4462
rect 5742 4386 5794 4398
rect 8318 4450 8370 4462
rect 8318 4386 8370 4398
rect 9550 4450 9602 4462
rect 9550 4386 9602 4398
rect 10110 4450 10162 4462
rect 10110 4386 10162 4398
rect 10670 4450 10722 4462
rect 10670 4386 10722 4398
rect 10894 4450 10946 4462
rect 10894 4386 10946 4398
rect 11790 4450 11842 4462
rect 11790 4386 11842 4398
rect 13806 4450 13858 4462
rect 15362 4398 15374 4450
rect 15426 4398 15438 4450
rect 15586 4398 15598 4450
rect 15650 4398 15662 4450
rect 13806 4386 13858 4398
rect 9774 4338 9826 4350
rect 13358 4338 13410 4350
rect 3714 4286 3726 4338
rect 3778 4286 3790 4338
rect 3938 4286 3950 4338
rect 4002 4286 4014 4338
rect 4274 4286 4286 4338
rect 4338 4286 4350 4338
rect 5170 4286 5182 4338
rect 5234 4286 5246 4338
rect 8978 4286 8990 4338
rect 9042 4286 9054 4338
rect 11218 4286 11230 4338
rect 11282 4286 11294 4338
rect 15810 4286 15822 4338
rect 15874 4286 15886 4338
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 9774 4274 9826 4286
rect 13358 4274 13410 4286
rect 1934 4226 1986 4238
rect 8530 4174 8542 4226
rect 8594 4174 8606 4226
rect 10546 4174 10558 4226
rect 10610 4174 10622 4226
rect 1934 4162 1986 4174
rect 2158 4114 2210 4126
rect 2158 4050 2210 4062
rect 1344 3946 18592 3980
rect 1344 3894 3370 3946
rect 3422 3894 3474 3946
rect 3526 3894 3578 3946
rect 3630 3894 7682 3946
rect 7734 3894 7786 3946
rect 7838 3894 7890 3946
rect 7942 3894 11994 3946
rect 12046 3894 12098 3946
rect 12150 3894 12202 3946
rect 12254 3894 16306 3946
rect 16358 3894 16410 3946
rect 16462 3894 16514 3946
rect 16566 3894 18592 3946
rect 1344 3860 18592 3894
rect 7534 3778 7586 3790
rect 7534 3714 7586 3726
rect 12238 3778 12290 3790
rect 12238 3714 12290 3726
rect 12574 3778 12626 3790
rect 12574 3714 12626 3726
rect 4510 3666 4562 3678
rect 17838 3666 17890 3678
rect 3378 3614 3390 3666
rect 3442 3614 3454 3666
rect 11554 3614 11566 3666
rect 11618 3614 11630 3666
rect 13906 3614 13918 3666
rect 13970 3614 13982 3666
rect 18162 3614 18174 3666
rect 18226 3614 18238 3666
rect 18834 3614 18846 3666
rect 18898 3663 18910 3666
rect 19394 3663 19406 3666
rect 18898 3617 19406 3663
rect 18898 3614 18910 3617
rect 19394 3614 19406 3617
rect 19458 3614 19470 3666
rect 4510 3602 4562 3614
rect 17838 3602 17890 3614
rect 4062 3554 4114 3566
rect 2818 3502 2830 3554
rect 2882 3502 2894 3554
rect 4062 3490 4114 3502
rect 4398 3554 4450 3566
rect 4398 3490 4450 3502
rect 5070 3554 5122 3566
rect 5070 3490 5122 3502
rect 6638 3554 6690 3566
rect 6638 3490 6690 3502
rect 7310 3554 7362 3566
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 8754 3502 8766 3554
rect 8818 3502 8830 3554
rect 9314 3502 9326 3554
rect 9378 3502 9390 3554
rect 11330 3502 11342 3554
rect 11394 3502 11406 3554
rect 14802 3502 14814 3554
rect 14866 3502 14878 3554
rect 15922 3502 15934 3554
rect 15986 3502 15998 3554
rect 17154 3502 17166 3554
rect 17218 3502 17230 3554
rect 7310 3490 7362 3502
rect 4622 3442 4674 3454
rect 16942 3442 16994 3454
rect 5842 3390 5854 3442
rect 5906 3390 5918 3442
rect 6402 3390 6414 3442
rect 6466 3390 6478 3442
rect 7522 3390 7534 3442
rect 7586 3390 7598 3442
rect 10210 3390 10222 3442
rect 10274 3390 10286 3442
rect 14578 3390 14590 3442
rect 14642 3390 14654 3442
rect 15698 3390 15710 3442
rect 15762 3390 15774 3442
rect 4622 3378 4674 3390
rect 16942 3378 16994 3390
rect 1934 3330 1986 3342
rect 1934 3266 1986 3278
rect 2158 3330 2210 3342
rect 12350 3330 12402 3342
rect 6514 3278 6526 3330
rect 6578 3278 6590 3330
rect 2158 3266 2210 3278
rect 12350 3266 12402 3278
rect 1344 3162 18752 3196
rect 1344 3110 5526 3162
rect 5578 3110 5630 3162
rect 5682 3110 5734 3162
rect 5786 3110 9838 3162
rect 9890 3110 9942 3162
rect 9994 3110 10046 3162
rect 10098 3110 14150 3162
rect 14202 3110 14254 3162
rect 14306 3110 14358 3162
rect 14410 3110 18462 3162
rect 18514 3110 18566 3162
rect 18618 3110 18670 3162
rect 18722 3110 18752 3162
rect 1344 3076 18752 3110
rect 3938 2942 3950 2994
rect 4002 2991 4014 2994
rect 8082 2991 8094 2994
rect 4002 2945 8094 2991
rect 4002 2942 4014 2945
rect 8082 2942 8094 2945
rect 8146 2942 8158 2994
rect 14690 2942 14702 2994
rect 14754 2991 14766 2994
rect 19170 2991 19182 2994
rect 14754 2945 19182 2991
rect 14754 2942 14766 2945
rect 19170 2942 19182 2945
rect 19234 2942 19246 2994
rect 1922 2718 1934 2770
rect 1986 2767 1998 2770
rect 2930 2767 2942 2770
rect 1986 2721 2942 2767
rect 1986 2718 1998 2721
rect 2930 2718 2942 2721
rect 2994 2767 3006 2770
rect 6626 2767 6638 2770
rect 2994 2721 6638 2767
rect 2994 2718 3006 2721
rect 6626 2718 6638 2721
rect 6690 2718 6702 2770
<< via1 >>
rect 2494 12686 2546 12738
rect 3054 12686 3106 12738
rect 17166 12686 17218 12738
rect 19182 12686 19234 12738
rect 5526 12518 5578 12570
rect 5630 12518 5682 12570
rect 5734 12518 5786 12570
rect 9838 12518 9890 12570
rect 9942 12518 9994 12570
rect 10046 12518 10098 12570
rect 14150 12518 14202 12570
rect 14254 12518 14306 12570
rect 14358 12518 14410 12570
rect 18462 12518 18514 12570
rect 18566 12518 18618 12570
rect 18670 12518 18722 12570
rect 4286 12350 4338 12402
rect 4734 12350 4786 12402
rect 7646 12350 7698 12402
rect 16382 12350 16434 12402
rect 1710 12238 1762 12290
rect 2158 12238 2210 12290
rect 3054 12238 3106 12290
rect 15822 12238 15874 12290
rect 17166 12238 17218 12290
rect 17838 12238 17890 12290
rect 3950 12126 4002 12178
rect 13246 12126 13298 12178
rect 14926 12126 14978 12178
rect 17502 12126 17554 12178
rect 18062 12126 18114 12178
rect 5630 12014 5682 12066
rect 6078 12014 6130 12066
rect 6638 12014 6690 12066
rect 12238 12014 12290 12066
rect 12686 12014 12738 12066
rect 13582 12014 13634 12066
rect 14478 12014 14530 12066
rect 15374 12014 15426 12066
rect 3370 11734 3422 11786
rect 3474 11734 3526 11786
rect 3578 11734 3630 11786
rect 7682 11734 7734 11786
rect 7786 11734 7838 11786
rect 7890 11734 7942 11786
rect 11994 11734 12046 11786
rect 12098 11734 12150 11786
rect 12202 11734 12254 11786
rect 16306 11734 16358 11786
rect 16410 11734 16462 11786
rect 16514 11734 16566 11786
rect 16830 11454 16882 11506
rect 14814 11342 14866 11394
rect 16942 11342 16994 11394
rect 2158 11230 2210 11282
rect 2606 11230 2658 11282
rect 3054 11230 3106 11282
rect 3502 11230 3554 11282
rect 13694 11230 13746 11282
rect 16046 11230 16098 11282
rect 16382 11230 16434 11282
rect 17726 11230 17778 11282
rect 18062 11230 18114 11282
rect 1710 11118 1762 11170
rect 4510 11118 4562 11170
rect 4958 11118 5010 11170
rect 5854 11118 5906 11170
rect 6302 11118 6354 11170
rect 6638 11118 6690 11170
rect 7086 11118 7138 11170
rect 7534 11118 7586 11170
rect 11678 11118 11730 11170
rect 12126 11118 12178 11170
rect 12574 11118 12626 11170
rect 13022 11118 13074 11170
rect 14142 11118 14194 11170
rect 15150 11118 15202 11170
rect 15710 11118 15762 11170
rect 5526 10950 5578 11002
rect 5630 10950 5682 11002
rect 5734 10950 5786 11002
rect 9838 10950 9890 11002
rect 9942 10950 9994 11002
rect 10046 10950 10098 11002
rect 14150 10950 14202 11002
rect 14254 10950 14306 11002
rect 14358 10950 14410 11002
rect 18462 10950 18514 11002
rect 18566 10950 18618 11002
rect 18670 10950 18722 11002
rect 2158 10782 2210 10834
rect 13694 10782 13746 10834
rect 17390 10782 17442 10834
rect 1710 10670 1762 10722
rect 2606 10670 2658 10722
rect 3054 10670 3106 10722
rect 3502 10670 3554 10722
rect 8990 10670 9042 10722
rect 10670 10670 10722 10722
rect 14702 10670 14754 10722
rect 15374 10670 15426 10722
rect 16158 10670 16210 10722
rect 16830 10670 16882 10722
rect 6862 10558 6914 10610
rect 8206 10558 8258 10610
rect 11678 10558 11730 10610
rect 13134 10558 13186 10610
rect 13582 10558 13634 10610
rect 13806 10558 13858 10610
rect 14366 10558 14418 10610
rect 15038 10558 15090 10610
rect 15822 10558 15874 10610
rect 16606 10558 16658 10610
rect 17726 10558 17778 10610
rect 3950 10446 4002 10498
rect 6078 10446 6130 10498
rect 7310 10446 7362 10498
rect 7758 10446 7810 10498
rect 11230 10446 11282 10498
rect 12126 10446 12178 10498
rect 12574 10446 12626 10498
rect 13022 10446 13074 10498
rect 18174 10446 18226 10498
rect 3370 10166 3422 10218
rect 3474 10166 3526 10218
rect 3578 10166 3630 10218
rect 7682 10166 7734 10218
rect 7786 10166 7838 10218
rect 7890 10166 7942 10218
rect 11994 10166 12046 10218
rect 12098 10166 12150 10218
rect 12202 10166 12254 10218
rect 16306 10166 16358 10218
rect 16410 10166 16462 10218
rect 16514 10166 16566 10218
rect 11454 9998 11506 10050
rect 10222 9886 10274 9938
rect 18174 9886 18226 9938
rect 9886 9774 9938 9826
rect 12126 9774 12178 9826
rect 13694 9774 13746 9826
rect 13806 9774 13858 9826
rect 14030 9774 14082 9826
rect 14702 9774 14754 9826
rect 15374 9774 15426 9826
rect 1710 9662 1762 9714
rect 10558 9662 10610 9714
rect 10670 9662 10722 9714
rect 11342 9662 11394 9714
rect 12462 9662 12514 9714
rect 14254 9662 14306 9714
rect 16046 9662 16098 9714
rect 2158 9550 2210 9602
rect 2606 9550 2658 9602
rect 3054 9550 3106 9602
rect 3502 9550 3554 9602
rect 3950 9550 4002 9602
rect 4398 9550 4450 9602
rect 5070 9550 5122 9602
rect 5742 9550 5794 9602
rect 6302 9550 6354 9602
rect 6750 9550 6802 9602
rect 7198 9550 7250 9602
rect 7534 9550 7586 9602
rect 7982 9550 8034 9602
rect 8430 9550 8482 9602
rect 8878 9550 8930 9602
rect 9438 9550 9490 9602
rect 10894 9550 10946 9602
rect 11454 9550 11506 9602
rect 11790 9550 11842 9602
rect 12014 9550 12066 9602
rect 12574 9550 12626 9602
rect 12798 9550 12850 9602
rect 13806 9550 13858 9602
rect 14926 9550 14978 9602
rect 5526 9382 5578 9434
rect 5630 9382 5682 9434
rect 5734 9382 5786 9434
rect 9838 9382 9890 9434
rect 9942 9382 9994 9434
rect 10046 9382 10098 9434
rect 14150 9382 14202 9434
rect 14254 9382 14306 9434
rect 14358 9382 14410 9434
rect 18462 9382 18514 9434
rect 18566 9382 18618 9434
rect 18670 9382 18722 9434
rect 1710 9102 1762 9154
rect 2158 9102 2210 9154
rect 2606 9102 2658 9154
rect 3054 9102 3106 9154
rect 3502 9102 3554 9154
rect 3950 9102 4002 9154
rect 4398 9102 4450 9154
rect 5294 9102 5346 9154
rect 8318 9102 8370 9154
rect 10110 9102 10162 9154
rect 13246 9102 13298 9154
rect 17390 9102 17442 9154
rect 5182 8990 5234 9042
rect 7198 8990 7250 9042
rect 9550 8990 9602 9042
rect 11566 8990 11618 9042
rect 16718 8990 16770 9042
rect 17614 8990 17666 9042
rect 8206 8878 8258 8930
rect 12910 8878 12962 8930
rect 13918 8878 13970 8930
rect 16046 8878 16098 8930
rect 18174 8878 18226 8930
rect 17950 8766 18002 8818
rect 18286 8766 18338 8818
rect 3370 8598 3422 8650
rect 3474 8598 3526 8650
rect 3578 8598 3630 8650
rect 7682 8598 7734 8650
rect 7786 8598 7838 8650
rect 7890 8598 7942 8650
rect 11994 8598 12046 8650
rect 12098 8598 12150 8650
rect 12202 8598 12254 8650
rect 16306 8598 16358 8650
rect 16410 8598 16462 8650
rect 16514 8598 16566 8650
rect 13470 8318 13522 8370
rect 16830 8318 16882 8370
rect 2158 8206 2210 8258
rect 7198 8206 7250 8258
rect 12126 8206 12178 8258
rect 16270 8206 16322 8258
rect 2382 8094 2434 8146
rect 4174 8094 4226 8146
rect 4622 8094 4674 8146
rect 5630 8094 5682 8146
rect 7870 8094 7922 8146
rect 15598 8094 15650 8146
rect 16718 8094 16770 8146
rect 17054 8094 17106 8146
rect 17278 8094 17330 8146
rect 17950 8094 18002 8146
rect 3054 7982 3106 8034
rect 3502 7982 3554 8034
rect 4286 7982 4338 8034
rect 4734 7982 4786 8034
rect 5966 7982 6018 8034
rect 6302 7982 6354 8034
rect 6974 7982 7026 8034
rect 17614 7982 17666 8034
rect 5526 7814 5578 7866
rect 5630 7814 5682 7866
rect 5734 7814 5786 7866
rect 9838 7814 9890 7866
rect 9942 7814 9994 7866
rect 10046 7814 10098 7866
rect 14150 7814 14202 7866
rect 14254 7814 14306 7866
rect 14358 7814 14410 7866
rect 18462 7814 18514 7866
rect 18566 7814 18618 7866
rect 18670 7814 18722 7866
rect 2046 7646 2098 7698
rect 2718 7646 2770 7698
rect 3614 7646 3666 7698
rect 7646 7646 7698 7698
rect 1710 7534 1762 7586
rect 3278 7534 3330 7586
rect 4734 7534 4786 7586
rect 6750 7534 6802 7586
rect 9998 7534 10050 7586
rect 10782 7534 10834 7586
rect 12126 7534 12178 7586
rect 17390 7534 17442 7586
rect 17502 7534 17554 7586
rect 17614 7534 17666 7586
rect 2494 7422 2546 7474
rect 4062 7422 4114 7474
rect 7870 7422 7922 7474
rect 8094 7422 8146 7474
rect 8542 7422 8594 7474
rect 8766 7422 8818 7474
rect 9662 7422 9714 7474
rect 10446 7422 10498 7474
rect 16718 7422 16770 7474
rect 17950 7422 18002 7474
rect 8654 7310 8706 7362
rect 11230 7310 11282 7362
rect 17838 7198 17890 7250
rect 3370 7030 3422 7082
rect 3474 7030 3526 7082
rect 3578 7030 3630 7082
rect 7682 7030 7734 7082
rect 7786 7030 7838 7082
rect 7890 7030 7942 7082
rect 11994 7030 12046 7082
rect 12098 7030 12150 7082
rect 12202 7030 12254 7082
rect 16306 7030 16358 7082
rect 16410 7030 16462 7082
rect 16514 7030 16566 7082
rect 12574 6862 12626 6914
rect 12910 6862 12962 6914
rect 1822 6638 1874 6690
rect 2494 6638 2546 6690
rect 3054 6638 3106 6690
rect 3950 6638 4002 6690
rect 4622 6638 4674 6690
rect 4846 6638 4898 6690
rect 4958 6638 5010 6690
rect 5742 6638 5794 6690
rect 7646 6638 7698 6690
rect 9662 6638 9714 6690
rect 12126 6638 12178 6690
rect 13470 6638 13522 6690
rect 13806 6638 13858 6690
rect 14030 6638 14082 6690
rect 14366 6638 14418 6690
rect 18174 6638 18226 6690
rect 2158 6526 2210 6578
rect 3390 6526 3442 6578
rect 4174 6526 4226 6578
rect 5070 6526 5122 6578
rect 6414 6526 6466 6578
rect 6526 6526 6578 6578
rect 7086 6526 7138 6578
rect 7198 6526 7250 6578
rect 7422 6526 7474 6578
rect 7758 6526 7810 6578
rect 11454 6526 11506 6578
rect 15038 6526 15090 6578
rect 16270 6526 16322 6578
rect 17054 6526 17106 6578
rect 3502 6414 3554 6466
rect 5966 6414 6018 6466
rect 6190 6414 6242 6466
rect 8654 6414 8706 6466
rect 11902 6414 11954 6466
rect 12798 6414 12850 6466
rect 13694 6414 13746 6466
rect 5526 6246 5578 6298
rect 5630 6246 5682 6298
rect 5734 6246 5786 6298
rect 9838 6246 9890 6298
rect 9942 6246 9994 6298
rect 10046 6246 10098 6298
rect 14150 6246 14202 6298
rect 14254 6246 14306 6298
rect 14358 6246 14410 6298
rect 18462 6246 18514 6298
rect 18566 6246 18618 6298
rect 18670 6246 18722 6298
rect 1822 6078 1874 6130
rect 2830 6078 2882 6130
rect 3502 6078 3554 6130
rect 17390 6078 17442 6130
rect 17502 6078 17554 6130
rect 17614 6078 17666 6130
rect 2158 5966 2210 6018
rect 3838 5966 3890 6018
rect 4174 5966 4226 6018
rect 4846 5966 4898 6018
rect 5854 5966 5906 6018
rect 7870 5966 7922 6018
rect 9886 5966 9938 6018
rect 10222 5966 10274 6018
rect 11230 5966 11282 6018
rect 16158 5966 16210 6018
rect 2606 5854 2658 5906
rect 3278 5854 3330 5906
rect 4510 5854 4562 5906
rect 5294 5854 5346 5906
rect 7310 5854 7362 5906
rect 11006 5854 11058 5906
rect 12350 5854 12402 5906
rect 17950 5854 18002 5906
rect 6750 5742 6802 5794
rect 3370 5462 3422 5514
rect 3474 5462 3526 5514
rect 3578 5462 3630 5514
rect 7682 5462 7734 5514
rect 7786 5462 7838 5514
rect 7890 5462 7942 5514
rect 11994 5462 12046 5514
rect 12098 5462 12150 5514
rect 12202 5462 12254 5514
rect 16306 5462 16358 5514
rect 16410 5462 16462 5514
rect 16514 5462 16566 5514
rect 8766 5182 8818 5234
rect 1822 5070 1874 5122
rect 2830 5070 2882 5122
rect 3502 5070 3554 5122
rect 4734 5070 4786 5122
rect 5966 5082 6018 5134
rect 9102 5070 9154 5122
rect 11342 5070 11394 5122
rect 13470 5070 13522 5122
rect 15598 5070 15650 5122
rect 17950 5070 18002 5122
rect 2158 4958 2210 5010
rect 3054 4958 3106 5010
rect 3726 4958 3778 5010
rect 4062 4958 4114 5010
rect 4398 4958 4450 5010
rect 5070 4958 5122 5010
rect 6638 4958 6690 5010
rect 9774 4958 9826 5010
rect 12350 4958 12402 5010
rect 14142 4958 14194 5010
rect 16718 4958 16770 5010
rect 17614 4958 17666 5010
rect 11342 4846 11394 4898
rect 15822 4846 15874 4898
rect 5526 4678 5578 4730
rect 5630 4678 5682 4730
rect 5734 4678 5786 4730
rect 9838 4678 9890 4730
rect 9942 4678 9994 4730
rect 10046 4678 10098 4730
rect 14150 4678 14202 4730
rect 14254 4678 14306 4730
rect 14358 4678 14410 4730
rect 18462 4678 18514 4730
rect 18566 4678 18618 4730
rect 18670 4678 18722 4730
rect 2942 4510 2994 4562
rect 4958 4510 5010 4562
rect 9662 4510 9714 4562
rect 14926 4510 14978 4562
rect 17390 4510 17442 4562
rect 18174 4510 18226 4562
rect 5742 4398 5794 4450
rect 8318 4398 8370 4450
rect 9550 4398 9602 4450
rect 10110 4398 10162 4450
rect 10670 4398 10722 4450
rect 10894 4398 10946 4450
rect 11790 4398 11842 4450
rect 13806 4398 13858 4450
rect 15374 4398 15426 4450
rect 15598 4398 15650 4450
rect 3726 4286 3778 4338
rect 3950 4286 4002 4338
rect 4286 4286 4338 4338
rect 5182 4286 5234 4338
rect 8990 4286 9042 4338
rect 9774 4286 9826 4338
rect 11230 4286 11282 4338
rect 13358 4286 13410 4338
rect 15822 4286 15874 4338
rect 17614 4286 17666 4338
rect 1934 4174 1986 4226
rect 8542 4174 8594 4226
rect 10558 4174 10610 4226
rect 2158 4062 2210 4114
rect 3370 3894 3422 3946
rect 3474 3894 3526 3946
rect 3578 3894 3630 3946
rect 7682 3894 7734 3946
rect 7786 3894 7838 3946
rect 7890 3894 7942 3946
rect 11994 3894 12046 3946
rect 12098 3894 12150 3946
rect 12202 3894 12254 3946
rect 16306 3894 16358 3946
rect 16410 3894 16462 3946
rect 16514 3894 16566 3946
rect 7534 3726 7586 3778
rect 12238 3726 12290 3778
rect 12574 3726 12626 3778
rect 3390 3614 3442 3666
rect 4510 3614 4562 3666
rect 11566 3614 11618 3666
rect 13918 3614 13970 3666
rect 17838 3614 17890 3666
rect 18174 3614 18226 3666
rect 18846 3614 18898 3666
rect 19406 3614 19458 3666
rect 2830 3502 2882 3554
rect 4062 3502 4114 3554
rect 4398 3502 4450 3554
rect 5070 3502 5122 3554
rect 6638 3502 6690 3554
rect 7310 3502 7362 3554
rect 7870 3502 7922 3554
rect 8766 3502 8818 3554
rect 9326 3502 9378 3554
rect 11342 3502 11394 3554
rect 14814 3502 14866 3554
rect 15934 3502 15986 3554
rect 17166 3502 17218 3554
rect 4622 3390 4674 3442
rect 5854 3390 5906 3442
rect 6414 3390 6466 3442
rect 7534 3390 7586 3442
rect 10222 3390 10274 3442
rect 14590 3390 14642 3442
rect 15710 3390 15762 3442
rect 16942 3390 16994 3442
rect 1934 3278 1986 3330
rect 2158 3278 2210 3330
rect 6526 3278 6578 3330
rect 12350 3278 12402 3330
rect 5526 3110 5578 3162
rect 5630 3110 5682 3162
rect 5734 3110 5786 3162
rect 9838 3110 9890 3162
rect 9942 3110 9994 3162
rect 10046 3110 10098 3162
rect 14150 3110 14202 3162
rect 14254 3110 14306 3162
rect 14358 3110 14410 3162
rect 18462 3110 18514 3162
rect 18566 3110 18618 3162
rect 18670 3110 18722 3162
rect 3950 2942 4002 2994
rect 8094 2942 8146 2994
rect 14702 2942 14754 2994
rect 19182 2942 19234 2994
rect 1934 2718 1986 2770
rect 2942 2718 2994 2770
rect 6638 2718 6690 2770
<< metal2 >>
rect 1708 15316 1764 15326
rect 1764 15260 1876 15316
rect 1708 15250 1764 15260
rect 1708 12290 1764 12302
rect 1708 12238 1710 12290
rect 1762 12238 1764 12290
rect 1708 11956 1764 12238
rect 1708 11890 1764 11900
rect 1708 11172 1764 11182
rect 1708 11078 1764 11116
rect 1708 10722 1764 10734
rect 1708 10670 1710 10722
rect 1762 10670 1764 10722
rect 1372 10612 1428 10622
rect 1260 8372 1316 8382
rect 1260 7588 1316 8316
rect 1260 3388 1316 7532
rect 1372 3556 1428 10556
rect 1708 10388 1764 10670
rect 1708 10322 1764 10332
rect 1708 9716 1764 9726
rect 1820 9716 1876 15260
rect 2464 15200 2576 16000
rect 7392 15200 7504 16000
rect 12320 15200 12432 16000
rect 17248 15200 17360 16000
rect 1932 13076 1988 13086
rect 1988 13020 2100 13076
rect 1932 13010 1988 13020
rect 1932 12068 1988 12078
rect 1932 10612 1988 12012
rect 2044 10836 2100 13020
rect 2492 12738 2548 15200
rect 4732 14868 4788 14878
rect 4284 14420 4340 14430
rect 3500 13972 3556 13982
rect 2828 13524 2884 13534
rect 2884 13468 2996 13524
rect 2828 13458 2884 13468
rect 2492 12686 2494 12738
rect 2546 12686 2548 12738
rect 2492 12674 2548 12686
rect 2604 12628 2660 12638
rect 2156 12292 2212 12302
rect 2156 12198 2212 12236
rect 2156 11284 2212 11294
rect 2156 11190 2212 11228
rect 2604 11282 2660 12572
rect 2604 11230 2606 11282
rect 2658 11230 2660 11282
rect 2604 11218 2660 11230
rect 2940 11284 2996 13468
rect 3052 12738 3108 12750
rect 3052 12686 3054 12738
rect 3106 12686 3108 12738
rect 3052 12290 3108 12686
rect 3052 12238 3054 12290
rect 3106 12238 3108 12290
rect 3052 12226 3108 12238
rect 3500 11956 3556 13916
rect 4284 12402 4340 14364
rect 4284 12350 4286 12402
rect 4338 12350 4340 12402
rect 4284 12338 4340 12350
rect 4732 12402 4788 14812
rect 5524 12572 5788 12582
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5524 12506 5788 12516
rect 4732 12350 4734 12402
rect 4786 12350 4788 12402
rect 4732 12338 4788 12350
rect 7420 12404 7476 15200
rect 9836 12572 10100 12582
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 9836 12506 10100 12516
rect 7644 12404 7700 12414
rect 7420 12402 7700 12404
rect 7420 12350 7646 12402
rect 7698 12350 7700 12402
rect 7420 12348 7700 12350
rect 7644 12338 7700 12348
rect 12348 12404 12404 15200
rect 17164 12738 17220 12750
rect 17164 12686 17166 12738
rect 17218 12686 17220 12738
rect 14148 12572 14412 12582
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14148 12506 14412 12516
rect 12348 12338 12404 12348
rect 13580 12404 13636 12414
rect 3948 12178 4004 12190
rect 3948 12126 3950 12178
rect 4002 12126 4004 12178
rect 3500 11900 3780 11956
rect 3368 11788 3632 11798
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3368 11722 3632 11732
rect 3052 11284 3108 11294
rect 2940 11282 3108 11284
rect 2940 11230 3054 11282
rect 3106 11230 3108 11282
rect 2940 11228 3108 11230
rect 3052 11218 3108 11228
rect 3500 11284 3556 11294
rect 3724 11284 3780 11900
rect 3500 11282 3780 11284
rect 3500 11230 3502 11282
rect 3554 11230 3780 11282
rect 3500 11228 3780 11230
rect 3500 11218 3556 11228
rect 2156 10836 2212 10846
rect 2044 10834 2212 10836
rect 2044 10782 2158 10834
rect 2210 10782 2212 10834
rect 2044 10780 2212 10782
rect 2156 10770 2212 10780
rect 2604 10722 2660 10734
rect 3052 10724 3108 10734
rect 2604 10670 2606 10722
rect 2658 10670 2660 10722
rect 1932 10556 2100 10612
rect 1708 9714 1876 9716
rect 1708 9662 1710 9714
rect 1762 9662 1876 9714
rect 1708 9660 1876 9662
rect 1932 10388 1988 10398
rect 1708 9650 1764 9660
rect 1708 9154 1764 9166
rect 1708 9102 1710 9154
rect 1762 9102 1764 9154
rect 1708 7924 1764 9102
rect 1596 7868 1764 7924
rect 1820 8820 1876 8830
rect 1484 7812 1540 7822
rect 1484 4564 1540 7756
rect 1596 6692 1652 7868
rect 1708 7588 1764 7598
rect 1708 7494 1764 7532
rect 1820 7028 1876 8764
rect 1596 6626 1652 6636
rect 1708 6972 1876 7028
rect 1484 4498 1540 4508
rect 1372 3490 1428 3500
rect 1260 3332 1428 3388
rect 1372 800 1428 3332
rect 1708 2772 1764 6972
rect 1820 6692 1876 6702
rect 1820 6598 1876 6636
rect 1932 6244 1988 10332
rect 2044 9716 2100 10556
rect 2604 9940 2660 10670
rect 2604 9874 2660 9884
rect 2828 10722 3108 10724
rect 2828 10670 3054 10722
rect 3106 10670 3108 10722
rect 2828 10668 3108 10670
rect 2044 9650 2100 9660
rect 2156 9604 2212 9614
rect 2604 9604 2660 9614
rect 2156 9510 2212 9548
rect 2492 9602 2660 9604
rect 2492 9550 2606 9602
rect 2658 9550 2660 9602
rect 2492 9548 2660 9550
rect 2156 9154 2212 9166
rect 2156 9102 2158 9154
rect 2210 9102 2212 9154
rect 2156 8596 2212 9102
rect 2156 8530 2212 8540
rect 2268 9156 2324 9166
rect 2156 8258 2212 8270
rect 2156 8206 2158 8258
rect 2210 8206 2212 8258
rect 2156 8148 2212 8206
rect 2156 8082 2212 8092
rect 2044 8036 2100 8046
rect 2044 7698 2100 7980
rect 2044 7646 2046 7698
rect 2098 7646 2100 7698
rect 2044 7634 2100 7646
rect 2156 6916 2212 6926
rect 1820 6188 1988 6244
rect 2044 6692 2100 6702
rect 1820 6130 1876 6188
rect 1820 6078 1822 6130
rect 1874 6078 1876 6130
rect 1820 5348 1876 6078
rect 1820 5292 1988 5348
rect 1820 5124 1876 5134
rect 1820 5030 1876 5068
rect 1932 4452 1988 5292
rect 2044 4452 2100 6636
rect 2156 6578 2212 6860
rect 2156 6526 2158 6578
rect 2210 6526 2212 6578
rect 2156 6514 2212 6526
rect 2156 6020 2212 6030
rect 2156 5926 2212 5964
rect 2156 5236 2212 5246
rect 2156 5010 2212 5180
rect 2156 4958 2158 5010
rect 2210 4958 2212 5010
rect 2156 4946 2212 4958
rect 2268 4676 2324 9100
rect 2380 8932 2436 8942
rect 2380 8146 2436 8876
rect 2380 8094 2382 8146
rect 2434 8094 2436 8146
rect 2380 8082 2436 8094
rect 2492 7700 2548 9548
rect 2604 9538 2660 9548
rect 2268 4610 2324 4620
rect 2380 7644 2548 7700
rect 2604 9154 2660 9166
rect 2604 9102 2606 9154
rect 2658 9102 2660 9154
rect 2044 4396 2324 4452
rect 1932 4386 1988 4396
rect 1932 4226 1988 4238
rect 1932 4174 1934 4226
rect 1986 4174 1988 4226
rect 1708 2706 1764 2716
rect 1820 4004 1876 4014
rect 1820 800 1876 3948
rect 1932 3780 1988 4174
rect 2156 4116 2212 4126
rect 1932 3714 1988 3724
rect 2044 4114 2212 4116
rect 2044 4062 2158 4114
rect 2210 4062 2212 4114
rect 2044 4060 2212 4062
rect 1932 3330 1988 3342
rect 1932 3278 1934 3330
rect 1986 3278 1988 3330
rect 1932 2770 1988 3278
rect 1932 2718 1934 2770
rect 1986 2718 1988 2770
rect 1932 2706 1988 2718
rect 2044 1876 2100 4060
rect 2156 4050 2212 4060
rect 2044 1810 2100 1820
rect 2156 3330 2212 3342
rect 2156 3278 2158 3330
rect 2210 3278 2212 3330
rect 2156 1540 2212 3278
rect 2156 1474 2212 1484
rect 2268 800 2324 4396
rect 2380 3668 2436 7644
rect 2492 7476 2548 7486
rect 2492 7382 2548 7420
rect 2492 6692 2548 6702
rect 2492 6598 2548 6636
rect 2604 6132 2660 9102
rect 2828 8820 2884 10668
rect 3052 10658 3108 10668
rect 3500 10724 3556 10734
rect 3500 10722 3780 10724
rect 3500 10670 3502 10722
rect 3554 10670 3780 10722
rect 3500 10668 3780 10670
rect 3500 10658 3556 10668
rect 3368 10220 3632 10230
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3368 10154 3632 10164
rect 3052 9604 3108 9614
rect 2828 8754 2884 8764
rect 2940 9602 3108 9604
rect 2940 9550 3054 9602
rect 3106 9550 3108 9602
rect 2940 9548 3108 9550
rect 2828 8484 2884 8494
rect 2716 8148 2772 8158
rect 2716 7698 2772 8092
rect 2716 7646 2718 7698
rect 2770 7646 2772 7698
rect 2716 7634 2772 7646
rect 2492 6076 2660 6132
rect 2716 7476 2772 7486
rect 2492 5012 2548 6076
rect 2604 5908 2660 5918
rect 2604 5814 2660 5852
rect 2716 5460 2772 7420
rect 2828 6692 2884 8428
rect 2828 6626 2884 6636
rect 2716 5394 2772 5404
rect 2828 6132 2884 6142
rect 2828 5348 2884 6076
rect 2828 5282 2884 5292
rect 2828 5124 2884 5134
rect 2828 5030 2884 5068
rect 2492 4946 2548 4956
rect 2940 4900 2996 9548
rect 3052 9538 3108 9548
rect 3500 9604 3556 9614
rect 3500 9510 3556 9548
rect 3164 9380 3220 9390
rect 3052 9156 3108 9166
rect 3052 9062 3108 9100
rect 3164 8372 3220 9324
rect 3276 9156 3332 9166
rect 3276 8820 3332 9100
rect 3500 9156 3556 9166
rect 3500 9062 3556 9100
rect 3276 8754 3332 8764
rect 3368 8652 3632 8662
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3368 8586 3632 8596
rect 3164 8306 3220 8316
rect 3612 8372 3668 8382
rect 3052 8036 3108 8046
rect 3052 8034 3220 8036
rect 3052 7982 3054 8034
rect 3106 7982 3220 8034
rect 3052 7980 3220 7982
rect 3052 7970 3108 7980
rect 3052 6690 3108 6702
rect 3052 6638 3054 6690
rect 3106 6638 3108 6690
rect 3052 6580 3108 6638
rect 3052 6514 3108 6524
rect 3164 6244 3220 7980
rect 3500 8034 3556 8046
rect 3500 7982 3502 8034
rect 3554 7982 3556 8034
rect 3276 7924 3332 7934
rect 3276 7586 3332 7868
rect 3276 7534 3278 7586
rect 3330 7534 3332 7586
rect 3276 7522 3332 7534
rect 3500 7588 3556 7982
rect 3612 7698 3668 8316
rect 3612 7646 3614 7698
rect 3666 7646 3668 7698
rect 3612 7634 3668 7646
rect 3724 7700 3780 10668
rect 3948 10498 4004 12126
rect 13244 12178 13300 12190
rect 13244 12126 13246 12178
rect 13298 12126 13300 12178
rect 5628 12068 5684 12078
rect 6076 12068 6132 12078
rect 6636 12068 6692 12078
rect 5628 11974 5684 12012
rect 5964 12066 6132 12068
rect 5964 12014 6078 12066
rect 6130 12014 6132 12066
rect 5964 12012 6132 12014
rect 3948 10446 3950 10498
rect 4002 10446 4004 10498
rect 3948 9828 4004 10446
rect 3948 9762 4004 9772
rect 4508 11170 4564 11182
rect 4508 11118 4510 11170
rect 4562 11118 4564 11170
rect 3948 9604 4004 9614
rect 4396 9604 4452 9614
rect 3948 9510 4004 9548
rect 4284 9602 4452 9604
rect 4284 9550 4398 9602
rect 4450 9550 4452 9602
rect 4284 9548 4452 9550
rect 3724 7634 3780 7644
rect 3948 9154 4004 9166
rect 3948 9102 3950 9154
rect 4002 9102 4004 9154
rect 3500 7522 3556 7532
rect 3724 7476 3780 7486
rect 3368 7084 3632 7094
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3368 7018 3632 7028
rect 3388 6578 3444 6590
rect 3388 6526 3390 6578
rect 3442 6526 3444 6578
rect 3164 6178 3220 6188
rect 3276 6468 3332 6478
rect 3276 5906 3332 6412
rect 3388 6132 3444 6526
rect 3500 6468 3556 6478
rect 3500 6466 3668 6468
rect 3500 6414 3502 6466
rect 3554 6414 3668 6466
rect 3500 6412 3668 6414
rect 3500 6402 3556 6412
rect 3500 6132 3556 6142
rect 3388 6130 3556 6132
rect 3388 6078 3502 6130
rect 3554 6078 3556 6130
rect 3388 6076 3556 6078
rect 3500 6066 3556 6076
rect 3276 5854 3278 5906
rect 3330 5854 3332 5906
rect 3276 5684 3332 5854
rect 3612 5684 3668 6412
rect 3724 5796 3780 7420
rect 3948 7252 4004 9102
rect 4284 8260 4340 9548
rect 4396 9538 4452 9548
rect 4396 9156 4452 9166
rect 4396 9062 4452 9100
rect 4284 8194 4340 8204
rect 4396 8484 4452 8494
rect 4172 8146 4228 8158
rect 4172 8094 4174 8146
rect 4226 8094 4228 8146
rect 4060 8036 4116 8046
rect 4060 7700 4116 7980
rect 4060 7634 4116 7644
rect 4060 7476 4116 7486
rect 4060 7382 4116 7420
rect 3948 7186 4004 7196
rect 3948 7028 4004 7038
rect 3948 6690 4004 6972
rect 3948 6638 3950 6690
rect 4002 6638 4004 6690
rect 3836 6244 3892 6254
rect 3836 6018 3892 6188
rect 3836 5966 3838 6018
rect 3890 5966 3892 6018
rect 3836 5954 3892 5966
rect 3948 5908 4004 6638
rect 4172 6916 4228 8094
rect 4284 8036 4340 8046
rect 4284 7942 4340 7980
rect 4172 6578 4228 6860
rect 4172 6526 4174 6578
rect 4226 6526 4228 6578
rect 4172 6514 4228 6526
rect 4284 6244 4340 6254
rect 4172 6020 4228 6058
rect 4172 5954 4228 5964
rect 4284 5908 4340 6188
rect 3948 5852 4116 5908
rect 4060 5796 4116 5852
rect 3724 5740 4004 5796
rect 4060 5740 4228 5796
rect 3612 5628 3892 5684
rect 3276 5618 3332 5628
rect 3368 5516 3632 5526
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3368 5450 3632 5460
rect 3724 5460 3780 5470
rect 3612 5348 3668 5358
rect 3388 5236 3444 5246
rect 3052 5180 3388 5236
rect 3052 5010 3108 5180
rect 3388 5170 3444 5180
rect 3052 4958 3054 5010
rect 3106 4958 3108 5010
rect 3052 4946 3108 4958
rect 3500 5122 3556 5134
rect 3500 5070 3502 5122
rect 3554 5070 3556 5122
rect 3500 5012 3556 5070
rect 3500 4946 3556 4956
rect 2380 3602 2436 3612
rect 2604 4844 2996 4900
rect 2604 3220 2660 4844
rect 2940 4564 2996 4574
rect 2940 4470 2996 4508
rect 3500 4452 3556 4462
rect 3500 4228 3556 4396
rect 3612 4340 3668 5292
rect 3724 5010 3780 5404
rect 3724 4958 3726 5010
rect 3778 4958 3780 5010
rect 3724 4946 3780 4958
rect 3836 4676 3892 5628
rect 3836 4610 3892 4620
rect 3948 5124 4004 5740
rect 3724 4340 3780 4350
rect 3612 4338 3780 4340
rect 3612 4286 3726 4338
rect 3778 4286 3780 4338
rect 3612 4284 3780 4286
rect 3724 4274 3780 4284
rect 3948 4338 4004 5068
rect 3948 4286 3950 4338
rect 4002 4286 4004 4338
rect 3948 4274 4004 4286
rect 4060 5348 4116 5358
rect 4060 5010 4116 5292
rect 4060 4958 4062 5010
rect 4114 4958 4116 5010
rect 3500 4172 3668 4228
rect 3612 4116 3668 4172
rect 4060 4116 4116 4958
rect 3612 4060 3780 4116
rect 3052 4004 3108 4014
rect 3108 3948 3220 4004
rect 3052 3938 3108 3948
rect 2604 3154 2660 3164
rect 2716 3892 2772 3902
rect 2716 800 2772 3836
rect 2828 3556 2884 3566
rect 2828 3462 2884 3500
rect 2940 2772 2996 2782
rect 2940 2678 2996 2716
rect 3164 800 3220 3948
rect 3368 3948 3632 3958
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3368 3882 3632 3892
rect 3724 3780 3780 4060
rect 3612 3724 3780 3780
rect 3948 4060 4116 4116
rect 3388 3666 3444 3678
rect 3388 3614 3390 3666
rect 3442 3614 3444 3666
rect 3388 868 3444 3614
rect 3388 802 3444 812
rect 3612 800 3668 3724
rect 3948 2994 4004 4060
rect 4060 3556 4116 3566
rect 4060 3462 4116 3500
rect 4172 3388 4228 5740
rect 4284 4338 4340 5852
rect 4396 5010 4452 8428
rect 4508 7700 4564 11118
rect 4956 11172 5012 11182
rect 4956 11078 5012 11116
rect 5852 11170 5908 11182
rect 5852 11118 5854 11170
rect 5906 11118 5908 11170
rect 5524 11004 5788 11014
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5524 10938 5788 10948
rect 5852 10724 5908 11118
rect 5852 10658 5908 10668
rect 4956 10164 5012 10174
rect 4620 8148 4676 8158
rect 4620 8054 4676 8092
rect 4732 8036 4788 8046
rect 4732 8034 4900 8036
rect 4732 7982 4734 8034
rect 4786 7982 4900 8034
rect 4732 7980 4900 7982
rect 4732 7970 4788 7980
rect 4508 7644 4676 7700
rect 4508 7476 4564 7486
rect 4508 6132 4564 7420
rect 4620 7028 4676 7644
rect 4620 6962 4676 6972
rect 4732 7586 4788 7598
rect 4732 7534 4734 7586
rect 4786 7534 4788 7586
rect 4508 6066 4564 6076
rect 4620 6690 4676 6702
rect 4620 6638 4622 6690
rect 4674 6638 4676 6690
rect 4508 5908 4564 5946
rect 4508 5842 4564 5852
rect 4396 4958 4398 5010
rect 4450 4958 4452 5010
rect 4396 4946 4452 4958
rect 4508 5684 4564 5694
rect 4508 4788 4564 5628
rect 4284 4286 4286 4338
rect 4338 4286 4340 4338
rect 4284 4274 4340 4286
rect 4396 4732 4564 4788
rect 4396 3554 4452 4732
rect 4508 3668 4564 3678
rect 4620 3668 4676 6638
rect 4732 6244 4788 7534
rect 4844 6690 4900 7980
rect 4844 6638 4846 6690
rect 4898 6638 4900 6690
rect 4844 6626 4900 6638
rect 4956 6690 5012 10108
rect 5068 9602 5124 9614
rect 5068 9550 5070 9602
rect 5122 9550 5124 9602
rect 5068 7924 5124 9550
rect 5740 9604 5796 9614
rect 5740 9602 5908 9604
rect 5740 9550 5742 9602
rect 5794 9550 5908 9602
rect 5740 9548 5908 9550
rect 5740 9538 5796 9548
rect 5524 9436 5788 9446
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 5524 9370 5788 9380
rect 5292 9154 5348 9166
rect 5292 9102 5294 9154
rect 5346 9102 5348 9154
rect 5180 9044 5236 9054
rect 5180 8950 5236 8988
rect 5292 8484 5348 9102
rect 5292 8418 5348 8428
rect 5628 8148 5684 8158
rect 5852 8148 5908 9548
rect 5964 8260 6020 12012
rect 6076 12002 6132 12012
rect 6524 12066 6692 12068
rect 6524 12014 6638 12066
rect 6690 12014 6692 12066
rect 6524 12012 6692 12014
rect 6300 11170 6356 11182
rect 6300 11118 6302 11170
rect 6354 11118 6356 11170
rect 6076 10498 6132 10510
rect 6076 10446 6078 10498
rect 6130 10446 6132 10498
rect 6076 10164 6132 10446
rect 6300 10500 6356 11118
rect 6300 10434 6356 10444
rect 6076 10098 6132 10108
rect 6300 9604 6356 9614
rect 5964 8194 6020 8204
rect 6188 9602 6356 9604
rect 6188 9550 6302 9602
rect 6354 9550 6356 9602
rect 6188 9548 6356 9550
rect 5628 8146 5908 8148
rect 5628 8094 5630 8146
rect 5682 8094 5908 8146
rect 5628 8092 5908 8094
rect 6076 8148 6132 8158
rect 5628 8036 5684 8092
rect 5068 7140 5124 7868
rect 5068 7074 5124 7084
rect 5180 7980 5684 8036
rect 5964 8034 6020 8046
rect 5964 7982 5966 8034
rect 6018 7982 6020 8034
rect 4956 6638 4958 6690
rect 5010 6638 5012 6690
rect 4956 6626 5012 6638
rect 4732 6178 4788 6188
rect 5068 6578 5124 6590
rect 5068 6526 5070 6578
rect 5122 6526 5124 6578
rect 4844 6076 5012 6132
rect 4844 6018 4900 6076
rect 4844 5966 4846 6018
rect 4898 5966 4900 6018
rect 4844 5954 4900 5966
rect 4956 6020 5012 6076
rect 4956 5954 5012 5964
rect 4956 5796 5012 5806
rect 4732 5348 4788 5358
rect 4732 5122 4788 5292
rect 4732 5070 4734 5122
rect 4786 5070 4788 5122
rect 4732 5058 4788 5070
rect 4732 4900 4788 4910
rect 4732 4340 4788 4844
rect 4956 4562 5012 5740
rect 5068 5684 5124 6526
rect 5180 5684 5236 7980
rect 5524 7868 5788 7878
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5524 7802 5788 7812
rect 5964 7028 6020 7982
rect 5404 6972 6020 7028
rect 5404 6244 5460 6972
rect 5740 6692 5796 6702
rect 5852 6692 5908 6702
rect 5740 6690 5852 6692
rect 5740 6638 5742 6690
rect 5794 6638 5852 6690
rect 5740 6636 5852 6638
rect 5740 6626 5796 6636
rect 5292 6188 5460 6244
rect 5524 6300 5788 6310
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5524 6234 5788 6244
rect 5852 6244 5908 6636
rect 5964 6468 6020 6478
rect 5964 6374 6020 6412
rect 5852 6188 6020 6244
rect 5292 5906 5348 6188
rect 5292 5854 5294 5906
rect 5346 5854 5348 5906
rect 5292 5842 5348 5854
rect 5852 6018 5908 6030
rect 5852 5966 5854 6018
rect 5906 5966 5908 6018
rect 5180 5628 5460 5684
rect 5068 5618 5124 5628
rect 5068 5124 5124 5134
rect 5068 5010 5124 5068
rect 5068 4958 5070 5010
rect 5122 4958 5124 5010
rect 5068 4946 5124 4958
rect 5180 4900 5236 4910
rect 4956 4510 4958 4562
rect 5010 4510 5012 4562
rect 4956 4498 5012 4510
rect 5068 4788 5124 4798
rect 5068 4452 5124 4732
rect 5068 4386 5124 4396
rect 4732 4284 5012 4340
rect 4508 3666 4676 3668
rect 4508 3614 4510 3666
rect 4562 3614 4676 3666
rect 4508 3612 4676 3614
rect 4508 3602 4564 3612
rect 4396 3502 4398 3554
rect 4450 3502 4452 3554
rect 4396 3490 4452 3502
rect 4620 3444 4676 3482
rect 3948 2942 3950 2994
rect 4002 2942 4004 2994
rect 3948 2930 4004 2942
rect 4060 3332 4116 3342
rect 4172 3332 4564 3388
rect 4620 3378 4676 3388
rect 4060 800 4116 3276
rect 4508 800 4564 3332
rect 4956 800 5012 4284
rect 5180 4338 5236 4844
rect 5180 4286 5182 4338
rect 5234 4286 5236 4338
rect 5180 4274 5236 4286
rect 5068 4004 5124 4014
rect 5068 3554 5124 3948
rect 5068 3502 5070 3554
rect 5122 3502 5124 3554
rect 5068 3490 5124 3502
rect 5404 800 5460 5628
rect 5852 5236 5908 5966
rect 5964 5908 6020 6188
rect 5964 5842 6020 5852
rect 6076 5684 6132 8092
rect 6188 6692 6244 9548
rect 6300 9538 6356 9548
rect 6300 8034 6356 8046
rect 6300 7982 6302 8034
rect 6354 7982 6356 8034
rect 6300 7252 6356 7982
rect 6300 7186 6356 7196
rect 6412 8036 6468 8046
rect 6188 6626 6244 6636
rect 6412 6578 6468 7980
rect 6524 7028 6580 12012
rect 6636 12002 6692 12012
rect 12236 12066 12292 12078
rect 12236 12014 12238 12066
rect 12290 12014 12292 12066
rect 12236 11956 12292 12014
rect 11788 11900 12292 11956
rect 12684 12066 12740 12078
rect 12684 12014 12686 12066
rect 12738 12014 12740 12066
rect 7680 11788 7944 11798
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 7680 11722 7944 11732
rect 6636 11170 6692 11182
rect 7084 11172 7140 11182
rect 6636 11118 6638 11170
rect 6690 11118 6692 11170
rect 6636 9604 6692 11118
rect 6972 11170 7140 11172
rect 6972 11118 7086 11170
rect 7138 11118 7140 11170
rect 6972 11116 7140 11118
rect 6972 10724 7028 11116
rect 7084 11106 7140 11116
rect 7532 11170 7588 11182
rect 7532 11118 7534 11170
rect 7586 11118 7588 11170
rect 6860 10610 6916 10622
rect 6860 10558 6862 10610
rect 6914 10558 6916 10610
rect 6636 9538 6692 9548
rect 6748 9602 6804 9614
rect 6748 9550 6750 9602
rect 6802 9550 6804 9602
rect 6524 6962 6580 6972
rect 6636 9380 6692 9390
rect 6636 7588 6692 9324
rect 6748 7812 6804 9550
rect 6860 8148 6916 10558
rect 6972 8260 7028 10668
rect 7308 10498 7364 10510
rect 7308 10446 7310 10498
rect 7362 10446 7364 10498
rect 7308 10276 7364 10446
rect 7308 10210 7364 10220
rect 7532 10052 7588 11118
rect 11676 11172 11732 11182
rect 11676 11078 11732 11116
rect 9836 11004 10100 11014
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 9836 10938 10100 10948
rect 8988 10724 9044 10734
rect 8988 10630 9044 10668
rect 10220 10724 10276 10734
rect 8204 10612 8260 10622
rect 8204 10518 8260 10556
rect 7756 10498 7812 10510
rect 7756 10446 7758 10498
rect 7810 10446 7812 10498
rect 7756 10388 7812 10446
rect 7756 10322 7812 10332
rect 7680 10220 7944 10230
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7680 10154 7944 10164
rect 7532 9986 7588 9996
rect 10220 10052 10276 10668
rect 10668 10724 10724 10734
rect 10668 10630 10724 10668
rect 11676 10612 11732 10622
rect 11452 10610 11732 10612
rect 11452 10558 11678 10610
rect 11730 10558 11732 10610
rect 11452 10556 11732 10558
rect 11228 10498 11284 10510
rect 11228 10446 11230 10498
rect 11282 10446 11284 10498
rect 11228 10276 11284 10446
rect 11452 10388 11508 10556
rect 11676 10546 11732 10556
rect 11788 10612 11844 11900
rect 11992 11788 12256 11798
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 11992 11722 12256 11732
rect 12684 11396 12740 12014
rect 12684 11330 12740 11340
rect 13132 11732 13188 11742
rect 12124 11172 12180 11182
rect 12124 11078 12180 11116
rect 12572 11172 12628 11182
rect 13020 11172 13076 11182
rect 12572 11170 12964 11172
rect 12572 11118 12574 11170
rect 12626 11118 12964 11170
rect 12572 11116 12964 11118
rect 12572 11106 12628 11116
rect 11788 10546 11844 10556
rect 12124 10500 12180 10510
rect 12572 10500 12628 10510
rect 12124 10498 12404 10500
rect 12124 10446 12126 10498
rect 12178 10446 12404 10498
rect 12124 10444 12404 10446
rect 12124 10434 12180 10444
rect 11452 10332 11732 10388
rect 11228 10210 11284 10220
rect 11452 10052 11508 10062
rect 10220 9938 10276 9996
rect 11228 10050 11508 10052
rect 11228 9998 11454 10050
rect 11506 9998 11508 10050
rect 11228 9996 11508 9998
rect 10220 9886 10222 9938
rect 10274 9886 10276 9938
rect 10220 9874 10276 9886
rect 10668 9940 10724 9950
rect 9884 9828 9940 9838
rect 9324 9826 9940 9828
rect 9324 9774 9886 9826
rect 9938 9774 9940 9826
rect 9324 9772 9940 9774
rect 7196 9604 7252 9614
rect 7196 9602 7364 9604
rect 7196 9550 7198 9602
rect 7250 9550 7364 9602
rect 7196 9548 7364 9550
rect 7196 9538 7252 9548
rect 7196 9042 7252 9054
rect 7196 8990 7198 9042
rect 7250 8990 7252 9042
rect 7196 8596 7252 8990
rect 7196 8530 7252 8540
rect 6972 8204 7140 8260
rect 6860 8082 6916 8092
rect 6972 8034 7028 8046
rect 6972 7982 6974 8034
rect 7026 7982 7028 8034
rect 6748 7756 6916 7812
rect 6412 6526 6414 6578
rect 6466 6526 6468 6578
rect 6412 6514 6468 6526
rect 6524 6580 6580 6590
rect 5852 5170 5908 5180
rect 5964 5628 6132 5684
rect 6188 6466 6244 6478
rect 6188 6414 6190 6466
rect 6242 6414 6244 6466
rect 5964 5134 6020 5628
rect 5964 5082 5966 5134
rect 6018 5082 6020 5134
rect 5964 5070 6020 5082
rect 6188 5012 6244 6414
rect 6524 5796 6580 6524
rect 6524 5730 6580 5740
rect 6636 5572 6692 7532
rect 6748 7586 6804 7598
rect 6748 7534 6750 7586
rect 6802 7534 6804 7586
rect 6748 6804 6804 7534
rect 6748 6738 6804 6748
rect 6860 7028 6916 7756
rect 6412 5516 6692 5572
rect 6748 5794 6804 5806
rect 6748 5742 6750 5794
rect 6802 5742 6804 5794
rect 5852 4956 6244 5012
rect 6300 5460 6356 5470
rect 5524 4732 5788 4742
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5524 4666 5788 4676
rect 5740 4452 5796 4462
rect 5852 4452 5908 4956
rect 5740 4450 5908 4452
rect 5740 4398 5742 4450
rect 5794 4398 5908 4450
rect 5740 4396 5908 4398
rect 5964 4788 6020 4798
rect 5964 4452 6020 4732
rect 5740 4386 5796 4396
rect 5852 3444 5908 3454
rect 5852 3350 5908 3388
rect 5524 3164 5788 3174
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5524 3098 5788 3108
rect 5964 1764 6020 4396
rect 5852 1708 6020 1764
rect 5852 800 5908 1708
rect 6300 800 6356 5404
rect 6412 3442 6468 5516
rect 6636 5236 6692 5246
rect 6524 5180 6636 5236
rect 6524 4340 6580 5180
rect 6636 5170 6692 5180
rect 6636 5010 6692 5022
rect 6636 4958 6638 5010
rect 6690 4958 6692 5010
rect 6636 4564 6692 4958
rect 6636 4498 6692 4508
rect 6524 4284 6692 4340
rect 6412 3390 6414 3442
rect 6466 3390 6468 3442
rect 6412 3378 6468 3390
rect 6524 3556 6580 3566
rect 6524 3330 6580 3500
rect 6524 3278 6526 3330
rect 6578 3278 6580 3330
rect 6524 3266 6580 3278
rect 6636 3554 6692 4284
rect 6636 3502 6638 3554
rect 6690 3502 6692 3554
rect 6636 2770 6692 3502
rect 6748 3556 6804 5742
rect 6748 3490 6804 3500
rect 6860 3388 6916 6972
rect 6972 5908 7028 7982
rect 7084 7476 7140 8204
rect 7084 7410 7140 7420
rect 7196 8258 7252 8270
rect 7196 8206 7198 8258
rect 7250 8206 7252 8258
rect 7196 7028 7252 8206
rect 7196 6962 7252 6972
rect 7196 6804 7252 6814
rect 7084 6580 7140 6590
rect 7084 6486 7140 6524
rect 7196 6578 7252 6748
rect 7196 6526 7198 6578
rect 7250 6526 7252 6578
rect 7196 6514 7252 6526
rect 7308 6356 7364 9548
rect 7532 9602 7588 9614
rect 7532 9550 7534 9602
rect 7586 9550 7588 9602
rect 7532 8708 7588 9550
rect 7980 9602 8036 9614
rect 7980 9550 7982 9602
rect 8034 9550 8036 9602
rect 7980 8820 8036 9550
rect 8428 9602 8484 9614
rect 8428 9550 8430 9602
rect 8482 9550 8484 9602
rect 8316 9154 8372 9166
rect 8316 9102 8318 9154
rect 8370 9102 8372 9154
rect 7980 8754 8036 8764
rect 8204 8930 8260 8942
rect 8204 8878 8206 8930
rect 8258 8878 8260 8930
rect 7532 8642 7588 8652
rect 7680 8652 7944 8662
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7680 8586 7944 8596
rect 7868 8148 7924 8158
rect 7868 8054 7924 8092
rect 7644 8036 7700 8046
rect 7644 7698 7700 7980
rect 7644 7646 7646 7698
rect 7698 7646 7700 7698
rect 7644 7634 7700 7646
rect 7868 7812 7924 7822
rect 7868 7474 7924 7756
rect 7868 7422 7870 7474
rect 7922 7422 7924 7474
rect 7868 7410 7924 7422
rect 8092 7476 8148 7486
rect 8092 7382 8148 7420
rect 7680 7084 7944 7094
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7680 7018 7944 7028
rect 7644 6692 7700 6702
rect 7532 6690 7700 6692
rect 7532 6638 7646 6690
rect 7698 6638 7700 6690
rect 7532 6636 7700 6638
rect 7420 6580 7476 6590
rect 7420 6486 7476 6524
rect 7308 6300 7476 6356
rect 7308 5908 7364 5918
rect 6972 5906 7364 5908
rect 6972 5854 7310 5906
rect 7362 5854 7364 5906
rect 6972 5852 7364 5854
rect 7308 5842 7364 5852
rect 7308 5348 7364 5358
rect 7420 5348 7476 6300
rect 7364 5292 7476 5348
rect 7308 5282 7364 5292
rect 7532 5012 7588 6636
rect 7644 6626 7700 6636
rect 7756 6578 7812 6590
rect 7756 6526 7758 6578
rect 7810 6526 7812 6578
rect 7756 6244 7812 6526
rect 7756 6178 7812 6188
rect 7868 6132 7924 6142
rect 7868 6018 7924 6076
rect 7868 5966 7870 6018
rect 7922 5966 7924 6018
rect 7868 5954 7924 5966
rect 7680 5516 7944 5526
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7680 5450 7944 5460
rect 7420 4956 7588 5012
rect 7420 3780 7476 4956
rect 7680 3948 7944 3958
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7680 3882 7944 3892
rect 7532 3780 7588 3790
rect 8204 3780 8260 8878
rect 8316 6020 8372 9102
rect 8428 8372 8484 9550
rect 8876 9602 8932 9614
rect 8876 9550 8878 9602
rect 8930 9550 8932 9602
rect 8876 9268 8932 9550
rect 8876 9202 8932 9212
rect 8428 8306 8484 8316
rect 8988 8820 9044 8830
rect 8316 5954 8372 5964
rect 8540 7588 8596 7598
rect 8540 7474 8596 7532
rect 8540 7422 8542 7474
rect 8594 7422 8596 7474
rect 8540 5236 8596 7422
rect 8764 7474 8820 7486
rect 8764 7422 8766 7474
rect 8818 7422 8820 7474
rect 8652 7362 8708 7374
rect 8652 7310 8654 7362
rect 8706 7310 8708 7362
rect 8652 6692 8708 7310
rect 8652 6626 8708 6636
rect 8652 6468 8708 6478
rect 8764 6468 8820 7422
rect 8652 6466 8820 6468
rect 8652 6414 8654 6466
rect 8706 6414 8820 6466
rect 8652 6412 8820 6414
rect 8652 5796 8708 6412
rect 8652 5730 8708 5740
rect 8876 5348 8932 5358
rect 8764 5236 8820 5246
rect 8540 5234 8820 5236
rect 8540 5182 8766 5234
rect 8818 5182 8820 5234
rect 8540 5180 8820 5182
rect 8764 5170 8820 5180
rect 8428 5012 8484 5022
rect 8316 4450 8372 4462
rect 8316 4398 8318 4450
rect 8370 4398 8372 4450
rect 8316 4340 8372 4398
rect 8316 4274 8372 4284
rect 7420 3778 7588 3780
rect 7420 3726 7534 3778
rect 7586 3726 7588 3778
rect 7420 3724 7588 3726
rect 7532 3714 7588 3724
rect 7868 3724 8260 3780
rect 6636 2718 6638 2770
rect 6690 2718 6692 2770
rect 6636 2706 6692 2718
rect 6748 3332 6916 3388
rect 7308 3554 7364 3566
rect 7308 3502 7310 3554
rect 7362 3502 7364 3554
rect 7308 3444 7364 3502
rect 7308 3378 7364 3388
rect 7532 3556 7588 3566
rect 7532 3442 7588 3500
rect 7868 3554 7924 3724
rect 8204 3668 8260 3724
rect 8204 3602 8260 3612
rect 7868 3502 7870 3554
rect 7922 3502 7924 3554
rect 7868 3490 7924 3502
rect 8428 3556 8484 4956
rect 8540 4226 8596 4238
rect 8540 4174 8542 4226
rect 8594 4174 8596 4226
rect 8540 4004 8596 4174
rect 8876 4004 8932 5292
rect 8988 5012 9044 8764
rect 9324 6020 9380 9772
rect 9884 9762 9940 9772
rect 10556 9716 10612 9726
rect 10332 9660 10556 9716
rect 9436 9602 9492 9614
rect 9436 9550 9438 9602
rect 9490 9550 9492 9602
rect 9436 7476 9492 9550
rect 9836 9436 10100 9446
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 9836 9370 10100 9380
rect 10108 9156 10164 9166
rect 10108 9154 10276 9156
rect 10108 9102 10110 9154
rect 10162 9102 10276 9154
rect 10108 9100 10276 9102
rect 10108 9090 10164 9100
rect 9548 9042 9604 9054
rect 9548 8990 9550 9042
rect 9602 8990 9604 9042
rect 9548 7700 9604 8990
rect 9836 7868 10100 7878
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 9836 7802 10100 7812
rect 9548 7644 9828 7700
rect 9660 7476 9716 7486
rect 9436 7420 9660 7476
rect 9660 7382 9716 7420
rect 9660 6692 9716 6702
rect 9772 6692 9828 7644
rect 9548 6690 9828 6692
rect 9548 6638 9662 6690
rect 9714 6638 9828 6690
rect 9548 6636 9828 6638
rect 9996 7586 10052 7598
rect 9996 7534 9998 7586
rect 10050 7534 10052 7586
rect 9548 6020 9604 6636
rect 9660 6626 9716 6636
rect 9996 6468 10052 7534
rect 10220 6804 10276 9100
rect 10332 6916 10388 9660
rect 10556 9622 10612 9660
rect 10668 9714 10724 9884
rect 10668 9662 10670 9714
rect 10722 9662 10724 9714
rect 10668 9650 10724 9662
rect 10892 9602 10948 9614
rect 10892 9550 10894 9602
rect 10946 9550 10948 9602
rect 10556 8932 10612 8942
rect 10332 6850 10388 6860
rect 10444 7474 10500 7486
rect 10444 7422 10446 7474
rect 10498 7422 10500 7474
rect 10444 7364 10500 7422
rect 10108 6748 10276 6804
rect 10108 6580 10164 6748
rect 10108 6514 10164 6524
rect 10332 6692 10388 6702
rect 9660 6412 10052 6468
rect 9660 6132 9716 6412
rect 9836 6300 10100 6310
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 9836 6234 10100 6244
rect 9660 6076 9828 6132
rect 9548 5964 9716 6020
rect 9324 5954 9380 5964
rect 9548 5684 9604 5694
rect 9100 5124 9156 5134
rect 9100 5030 9156 5068
rect 8988 4946 9044 4956
rect 9548 4450 9604 5628
rect 9660 4900 9716 5964
rect 9772 5010 9828 6076
rect 9772 4958 9774 5010
rect 9826 4958 9828 5010
rect 9772 4946 9828 4958
rect 9884 6020 9940 6030
rect 9660 4834 9716 4844
rect 9884 4900 9940 5964
rect 10220 6018 10276 6030
rect 10220 5966 10222 6018
rect 10274 5966 10276 6018
rect 10108 5908 10164 5918
rect 10108 5348 10164 5852
rect 10108 5282 10164 5292
rect 10220 5124 10276 5966
rect 10220 5058 10276 5068
rect 9996 5012 10052 5022
rect 9996 4900 10052 4956
rect 9996 4844 10276 4900
rect 9884 4834 9940 4844
rect 10220 4788 10276 4844
rect 9836 4732 10100 4742
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10220 4722 10276 4732
rect 9836 4666 10100 4676
rect 9660 4564 9716 4574
rect 10332 4564 10388 6636
rect 9660 4470 9716 4508
rect 10108 4508 10388 4564
rect 9548 4398 9550 4450
rect 9602 4398 9604 4450
rect 9548 4386 9604 4398
rect 9772 4452 9828 4462
rect 8988 4338 9044 4350
rect 8988 4286 8990 4338
rect 9042 4286 9044 4338
rect 8988 4228 9044 4286
rect 9772 4338 9828 4396
rect 10108 4450 10164 4508
rect 10108 4398 10110 4450
rect 10162 4398 10164 4450
rect 10108 4386 10164 4398
rect 10444 4340 10500 7308
rect 9772 4286 9774 4338
rect 9826 4286 9828 4338
rect 9772 4274 9828 4286
rect 10332 4284 10500 4340
rect 8988 4162 9044 4172
rect 8876 3948 9044 4004
rect 8540 3938 8596 3948
rect 8428 3490 8484 3500
rect 8764 3556 8820 3566
rect 8764 3462 8820 3500
rect 7532 3390 7534 3442
rect 7586 3390 7588 3442
rect 7532 3378 7588 3390
rect 6748 800 6804 3332
rect 8092 2994 8148 3006
rect 8092 2942 8094 2994
rect 8146 2942 8148 2994
rect 7196 2772 7252 2782
rect 7196 800 7252 2716
rect 7644 2660 7700 2670
rect 7644 800 7700 2604
rect 8092 800 8148 2942
rect 8540 2996 8596 3006
rect 8540 800 8596 2940
rect 8988 800 9044 3948
rect 9324 3668 9380 3678
rect 9324 3554 9380 3612
rect 9324 3502 9326 3554
rect 9378 3502 9380 3554
rect 9324 3490 9380 3502
rect 10220 3444 10276 3482
rect 10220 3378 10276 3388
rect 9836 3164 10100 3174
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 9836 3098 10100 3108
rect 9884 2884 9940 2894
rect 9436 1092 9492 1102
rect 9436 800 9492 1036
rect 9884 800 9940 2828
rect 10332 800 10388 4284
rect 10556 4226 10612 8876
rect 10892 8148 10948 9550
rect 11116 8484 11172 8494
rect 10892 8082 10948 8092
rect 11004 8428 11116 8484
rect 10780 7586 10836 7598
rect 10780 7534 10782 7586
rect 10834 7534 10836 7586
rect 10668 6916 10724 6926
rect 10668 4676 10724 6860
rect 10780 5124 10836 7534
rect 11004 6804 11060 8428
rect 11116 8418 11172 8428
rect 11228 8036 11284 9996
rect 11452 9986 11508 9996
rect 11452 9828 11508 9838
rect 11340 9716 11396 9726
rect 11340 9622 11396 9660
rect 11228 7970 11284 7980
rect 11452 9602 11508 9772
rect 11452 9550 11454 9602
rect 11506 9550 11508 9602
rect 11452 7588 11508 9550
rect 11452 7522 11508 7532
rect 11564 9042 11620 9054
rect 11564 8990 11566 9042
rect 11618 8990 11620 9042
rect 11228 7364 11284 7374
rect 11228 7270 11284 7308
rect 10780 5058 10836 5068
rect 10892 6748 11060 6804
rect 10780 4676 10836 4686
rect 10668 4620 10780 4676
rect 10780 4610 10836 4620
rect 10556 4174 10558 4226
rect 10610 4174 10612 4226
rect 10556 4162 10612 4174
rect 10668 4450 10724 4462
rect 10668 4398 10670 4450
rect 10722 4398 10724 4450
rect 10668 3780 10724 4398
rect 10780 4452 10836 4462
rect 10780 4228 10836 4396
rect 10892 4450 10948 6748
rect 11452 6580 11508 6590
rect 11564 6580 11620 8990
rect 11452 6578 11620 6580
rect 11452 6526 11454 6578
rect 11506 6526 11620 6578
rect 11452 6524 11620 6526
rect 11676 6692 11732 10332
rect 11992 10220 12256 10230
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 11992 10154 12256 10164
rect 12348 10164 12404 10444
rect 12572 10498 12740 10500
rect 12572 10446 12574 10498
rect 12626 10446 12740 10498
rect 12572 10444 12740 10446
rect 12572 10434 12628 10444
rect 12348 10108 12628 10164
rect 12124 10052 12180 10062
rect 12124 9826 12180 9996
rect 12572 9940 12628 10108
rect 12124 9774 12126 9826
rect 12178 9774 12180 9826
rect 12124 9762 12180 9774
rect 12348 9884 12628 9940
rect 12012 9716 12068 9726
rect 11788 9602 11844 9614
rect 11788 9550 11790 9602
rect 11842 9550 11844 9602
rect 11788 8484 11844 9550
rect 12012 9602 12068 9660
rect 12012 9550 12014 9602
rect 12066 9550 12068 9602
rect 12012 9044 12068 9550
rect 12012 8978 12068 8988
rect 11992 8652 12256 8662
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 11992 8586 12256 8596
rect 11788 8418 11844 8428
rect 12124 8258 12180 8270
rect 12124 8206 12126 8258
rect 12178 8206 12180 8258
rect 12124 7588 12180 8206
rect 12348 7700 12404 9884
rect 12460 9716 12516 9726
rect 12460 9622 12516 9660
rect 12572 9604 12628 9614
rect 12572 9510 12628 9548
rect 12348 7644 12516 7700
rect 12124 7586 12404 7588
rect 12124 7534 12126 7586
rect 12178 7534 12404 7586
rect 12124 7532 12404 7534
rect 12124 7522 12180 7532
rect 11992 7084 12256 7094
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 11992 7018 12256 7028
rect 12124 6692 12180 6702
rect 11676 6690 12180 6692
rect 11676 6638 12126 6690
rect 12178 6638 12180 6690
rect 11676 6636 12180 6638
rect 11004 6020 11060 6030
rect 11228 6020 11284 6030
rect 11004 5906 11060 5964
rect 11004 5854 11006 5906
rect 11058 5854 11060 5906
rect 11004 5842 11060 5854
rect 11116 6018 11284 6020
rect 11116 5966 11230 6018
rect 11282 5966 11284 6018
rect 11116 5964 11284 5966
rect 10892 4398 10894 4450
rect 10946 4398 10948 4450
rect 10892 4386 10948 4398
rect 11116 4340 11172 5964
rect 11228 5954 11284 5964
rect 11452 5796 11508 6524
rect 11228 5740 11508 5796
rect 11228 4564 11284 5740
rect 11340 5124 11396 5162
rect 11340 5058 11396 5068
rect 11228 4498 11284 4508
rect 11340 4898 11396 4910
rect 11340 4846 11342 4898
rect 11394 4846 11396 4898
rect 11228 4340 11284 4350
rect 11116 4338 11284 4340
rect 11116 4286 11230 4338
rect 11282 4286 11284 4338
rect 11116 4284 11284 4286
rect 11228 4274 11284 4284
rect 10780 4162 10836 4172
rect 10668 3714 10724 3724
rect 10780 3892 10836 3902
rect 10780 800 10836 3836
rect 11340 3556 11396 4846
rect 11340 3462 11396 3500
rect 11452 4900 11508 4910
rect 11452 3388 11508 4844
rect 11564 4788 11620 4798
rect 11564 4340 11620 4732
rect 11564 3666 11620 4284
rect 11564 3614 11566 3666
rect 11618 3614 11620 3666
rect 11564 3602 11620 3614
rect 11228 3332 11508 3388
rect 11228 800 11284 3332
rect 11676 800 11732 6636
rect 12124 6626 12180 6636
rect 11900 6468 11956 6478
rect 11788 6466 11956 6468
rect 11788 6414 11902 6466
rect 11954 6414 11956 6466
rect 11788 6412 11956 6414
rect 11788 5348 11844 6412
rect 11900 6402 11956 6412
rect 12348 5906 12404 7532
rect 12348 5854 12350 5906
rect 12402 5854 12404 5906
rect 12348 5842 12404 5854
rect 12460 6020 12516 7644
rect 12684 7476 12740 10444
rect 12908 9940 12964 11116
rect 13020 11078 13076 11116
rect 13132 10610 13188 11676
rect 13132 10558 13134 10610
rect 13186 10558 13188 10610
rect 13020 10500 13076 10510
rect 13020 10406 13076 10444
rect 13132 10388 13188 10558
rect 13132 10322 13188 10332
rect 13132 10164 13188 10174
rect 12908 9884 13076 9940
rect 12684 7410 12740 7420
rect 12796 9604 12852 9614
rect 12572 7252 12628 7262
rect 12796 7252 12852 9548
rect 12628 7196 12852 7252
rect 12908 9492 12964 9502
rect 12908 8930 12964 9436
rect 12908 8878 12910 8930
rect 12962 8878 12964 8930
rect 12572 6914 12628 7196
rect 12908 7140 12964 8878
rect 12572 6862 12574 6914
rect 12626 6862 12628 6914
rect 12572 6850 12628 6862
rect 12684 7084 12964 7140
rect 11992 5516 12256 5526
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 11992 5450 12256 5460
rect 11788 5292 11956 5348
rect 11788 4452 11844 4462
rect 11900 4452 11956 5292
rect 11788 4450 11956 4452
rect 11788 4398 11790 4450
rect 11842 4398 11956 4450
rect 11788 4396 11956 4398
rect 12348 5010 12404 5022
rect 12348 4958 12350 5010
rect 12402 4958 12404 5010
rect 11788 4386 11844 4396
rect 12348 4116 12404 4958
rect 12348 4050 12404 4060
rect 11788 4004 11844 4014
rect 11788 3556 11844 3948
rect 11992 3948 12256 3958
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 11992 3882 12256 3892
rect 12236 3780 12292 3790
rect 12236 3686 12292 3724
rect 12460 3556 12516 5964
rect 12572 3780 12628 3790
rect 12684 3780 12740 7084
rect 12908 6916 12964 6926
rect 12908 6822 12964 6860
rect 12796 6468 12852 6478
rect 12796 5236 12852 6412
rect 12796 5170 12852 5180
rect 13020 4340 13076 9884
rect 13020 4274 13076 4284
rect 12572 3778 12740 3780
rect 12572 3726 12574 3778
rect 12626 3726 12740 3778
rect 12572 3724 12740 3726
rect 12572 3714 12628 3724
rect 11788 3490 11844 3500
rect 12124 3500 12516 3556
rect 12572 3556 12628 3566
rect 12124 800 12180 3500
rect 12572 3388 12628 3500
rect 12348 3332 12628 3388
rect 12348 3330 12404 3332
rect 12348 3278 12350 3330
rect 12402 3278 12404 3330
rect 12348 3266 12404 3278
rect 12572 3220 12628 3230
rect 12572 800 12628 3164
rect 13132 1988 13188 10108
rect 13244 9828 13300 12126
rect 13580 12066 13636 12348
rect 16380 12404 16436 12414
rect 16380 12310 16436 12348
rect 15820 12292 15876 12302
rect 15820 12198 15876 12236
rect 17164 12290 17220 12686
rect 17276 12404 17332 15200
rect 19180 12738 19236 12750
rect 19180 12686 19182 12738
rect 19234 12686 19236 12738
rect 18460 12572 18724 12582
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18460 12506 18724 12516
rect 17276 12338 17332 12348
rect 17164 12238 17166 12290
rect 17218 12238 17220 12290
rect 17164 12226 17220 12238
rect 17836 12290 17892 12302
rect 17836 12238 17838 12290
rect 17890 12238 17892 12290
rect 14924 12180 14980 12190
rect 14924 12086 14980 12124
rect 17500 12178 17556 12190
rect 17500 12126 17502 12178
rect 17554 12126 17556 12178
rect 13580 12014 13582 12066
rect 13634 12014 13636 12066
rect 13580 12002 13636 12014
rect 14476 12066 14532 12078
rect 14476 12014 14478 12066
rect 14530 12014 14532 12066
rect 14476 11732 14532 12014
rect 15372 12066 15428 12078
rect 15372 12014 15374 12066
rect 15426 12014 15428 12066
rect 15372 11956 15428 12014
rect 15372 11890 15428 11900
rect 16716 11844 16772 11854
rect 16304 11788 16568 11798
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16304 11722 16568 11732
rect 14476 11666 14532 11676
rect 14588 11508 14644 11518
rect 14476 11452 14588 11508
rect 13692 11284 13748 11294
rect 13692 11190 13748 11228
rect 13244 9762 13300 9772
rect 13356 11172 13412 11182
rect 13244 9154 13300 9166
rect 13244 9102 13246 9154
rect 13298 9102 13300 9154
rect 13244 4788 13300 9102
rect 13356 5124 13412 11116
rect 14140 11172 14196 11210
rect 14140 11106 14196 11116
rect 14148 11004 14412 11014
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14148 10938 14412 10948
rect 13692 10836 13748 10846
rect 14364 10836 14420 10846
rect 13692 10834 13972 10836
rect 13692 10782 13694 10834
rect 13746 10782 13972 10834
rect 13692 10780 13972 10782
rect 13692 10770 13748 10780
rect 13580 10612 13636 10622
rect 13468 10610 13636 10612
rect 13468 10558 13582 10610
rect 13634 10558 13636 10610
rect 13468 10556 13636 10558
rect 13468 8372 13524 10556
rect 13580 10546 13636 10556
rect 13804 10610 13860 10622
rect 13804 10558 13806 10610
rect 13858 10558 13860 10610
rect 13804 10164 13860 10558
rect 13468 8306 13524 8316
rect 13580 10108 13860 10164
rect 13468 8148 13524 8158
rect 13468 6690 13524 8092
rect 13580 6916 13636 10108
rect 13692 9826 13748 9838
rect 13692 9774 13694 9826
rect 13746 9774 13748 9826
rect 13692 9380 13748 9774
rect 13804 9828 13860 9866
rect 13804 9762 13860 9772
rect 13692 8708 13748 9324
rect 13692 8642 13748 8652
rect 13804 9602 13860 9614
rect 13804 9550 13806 9602
rect 13858 9550 13860 9602
rect 13804 8596 13860 9550
rect 13916 9156 13972 10780
rect 14364 10610 14420 10780
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14364 10164 14420 10558
rect 14364 10098 14420 10108
rect 14476 9940 14532 11452
rect 14588 11442 14644 11452
rect 14812 11396 14868 11406
rect 16044 11396 16100 11406
rect 14812 11394 14980 11396
rect 14812 11342 14814 11394
rect 14866 11342 14980 11394
rect 14812 11340 14980 11342
rect 14812 11330 14868 11340
rect 14812 11172 14868 11182
rect 14700 10724 14756 10734
rect 14140 9884 14532 9940
rect 14588 10722 14756 10724
rect 14588 10670 14702 10722
rect 14754 10670 14756 10722
rect 14588 10668 14756 10670
rect 14028 9828 14084 9838
rect 14140 9828 14196 9884
rect 14028 9826 14196 9828
rect 14028 9774 14030 9826
rect 14082 9774 14196 9826
rect 14028 9772 14196 9774
rect 14028 9762 14084 9772
rect 14252 9714 14308 9726
rect 14252 9662 14254 9714
rect 14306 9662 14308 9714
rect 14252 9604 14308 9662
rect 14252 9538 14308 9548
rect 14148 9436 14412 9446
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14148 9370 14412 9380
rect 13916 9100 14084 9156
rect 13916 8930 13972 8942
rect 13916 8878 13918 8930
rect 13970 8878 13972 8930
rect 13916 8820 13972 8878
rect 13916 8754 13972 8764
rect 13804 8530 13860 8540
rect 13804 8260 13860 8270
rect 13580 6850 13636 6860
rect 13692 8148 13748 8158
rect 13468 6638 13470 6690
rect 13522 6638 13524 6690
rect 13468 6626 13524 6638
rect 13692 6466 13748 8092
rect 13804 6690 13860 8204
rect 13804 6638 13806 6690
rect 13858 6638 13860 6690
rect 13804 6626 13860 6638
rect 14028 6690 14084 9100
rect 14148 7868 14412 7878
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14148 7802 14412 7812
rect 14028 6638 14030 6690
rect 14082 6638 14084 6690
rect 14028 6626 14084 6638
rect 14364 6692 14420 6702
rect 14364 6598 14420 6636
rect 13692 6414 13694 6466
rect 13746 6414 13748 6466
rect 13692 6402 13748 6414
rect 14148 6300 14412 6310
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14148 6234 14412 6244
rect 14588 6132 14644 10668
rect 14700 10658 14756 10668
rect 14812 10500 14868 11116
rect 14924 10612 14980 11340
rect 16044 11282 16100 11340
rect 16044 11230 16046 11282
rect 16098 11230 16100 11282
rect 15148 11172 15204 11182
rect 15708 11172 15764 11182
rect 15148 11078 15204 11116
rect 15484 11170 15764 11172
rect 15484 11118 15710 11170
rect 15762 11118 15764 11170
rect 15484 11116 15764 11118
rect 16044 11172 16100 11230
rect 16380 11282 16436 11294
rect 16380 11230 16382 11282
rect 16434 11230 16436 11282
rect 16156 11172 16212 11182
rect 16044 11116 16156 11172
rect 15372 10724 15428 10734
rect 15260 10722 15428 10724
rect 15260 10670 15374 10722
rect 15426 10670 15428 10722
rect 15260 10668 15428 10670
rect 15036 10612 15092 10622
rect 14924 10610 15092 10612
rect 14924 10558 15038 10610
rect 15090 10558 15092 10610
rect 14924 10556 15092 10558
rect 14140 6076 14644 6132
rect 14700 10444 14868 10500
rect 14700 9826 14756 10444
rect 15036 9828 15092 10556
rect 14700 9774 14702 9826
rect 14754 9774 14756 9826
rect 13356 5058 13412 5068
rect 13468 5122 13524 5134
rect 13468 5070 13470 5122
rect 13522 5070 13524 5122
rect 13244 4722 13300 4732
rect 13468 4452 13524 5070
rect 13804 5012 13860 5022
rect 13468 4396 13636 4452
rect 13356 4340 13412 4350
rect 13356 4338 13524 4340
rect 13356 4286 13358 4338
rect 13410 4286 13524 4338
rect 13356 4284 13524 4286
rect 13356 4274 13412 4284
rect 13468 3332 13524 4284
rect 13580 3444 13636 4396
rect 13804 4450 13860 4956
rect 14140 5010 14196 6076
rect 14700 6020 14756 9774
rect 14812 9772 15092 9828
rect 14812 6356 14868 9772
rect 14924 9602 14980 9614
rect 14924 9550 14926 9602
rect 14978 9550 14980 9602
rect 14924 7364 14980 9550
rect 14924 7298 14980 7308
rect 15036 6580 15092 6590
rect 15260 6580 15316 10668
rect 15372 10658 15428 10668
rect 15372 9826 15428 9838
rect 15372 9774 15374 9826
rect 15426 9774 15428 9826
rect 15372 9044 15428 9774
rect 15372 8978 15428 8988
rect 15036 6578 15316 6580
rect 15036 6526 15038 6578
rect 15090 6526 15316 6578
rect 15036 6524 15316 6526
rect 15036 6514 15092 6524
rect 14812 6300 15092 6356
rect 14140 4958 14142 5010
rect 14194 4958 14196 5010
rect 14140 4946 14196 4958
rect 14476 5964 14756 6020
rect 14148 4732 14412 4742
rect 13804 4398 13806 4450
rect 13858 4398 13860 4450
rect 13804 4386 13860 4398
rect 13916 4676 13972 4686
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14148 4666 14412 4676
rect 13580 3378 13636 3388
rect 13692 3668 13748 3678
rect 13468 3266 13524 3276
rect 13020 1932 13188 1988
rect 13020 800 13076 1932
rect 13692 1764 13748 3612
rect 13916 3666 13972 4620
rect 13916 3614 13918 3666
rect 13970 3614 13972 3666
rect 13916 3602 13972 3614
rect 14476 3388 14532 5964
rect 14924 4564 14980 4574
rect 14924 4470 14980 4508
rect 14812 3556 14868 3594
rect 14812 3490 14868 3500
rect 13468 1708 13748 1764
rect 13916 3332 14532 3388
rect 14588 3444 14644 3454
rect 14588 3442 14756 3444
rect 14588 3390 14590 3442
rect 14642 3390 14756 3442
rect 14588 3388 14756 3390
rect 14588 3378 14644 3388
rect 13468 800 13524 1708
rect 13916 800 13972 3332
rect 14148 3164 14412 3174
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14148 3098 14412 3108
rect 14364 2996 14420 3006
rect 14364 800 14420 2940
rect 14700 2994 14756 3388
rect 15036 3332 15092 6300
rect 15372 4452 15428 4462
rect 15372 4358 15428 4396
rect 14700 2942 14702 2994
rect 14754 2942 14756 2994
rect 14700 2930 14756 2942
rect 14812 3276 15092 3332
rect 15260 4340 15316 4350
rect 14812 800 14868 3276
rect 15260 800 15316 4284
rect 15484 3556 15540 11116
rect 15708 11106 15764 11116
rect 16156 11106 16212 11116
rect 16380 10948 16436 11230
rect 15932 10892 16436 10948
rect 15820 10612 15876 10622
rect 15820 10518 15876 10556
rect 15932 10388 15988 10892
rect 15820 10332 15988 10388
rect 16156 10722 16212 10734
rect 16156 10670 16158 10722
rect 16210 10670 16212 10722
rect 15596 8148 15652 8158
rect 15820 8148 15876 10332
rect 16044 9716 16100 9726
rect 15932 9714 16100 9716
rect 15932 9662 16046 9714
rect 16098 9662 16100 9714
rect 15932 9660 16100 9662
rect 15932 8372 15988 9660
rect 16044 9650 16100 9660
rect 16156 9156 16212 10670
rect 16604 10610 16660 10622
rect 16604 10558 16606 10610
rect 16658 10558 16660 10610
rect 16604 10388 16660 10558
rect 16604 10322 16660 10332
rect 16304 10220 16568 10230
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16304 10154 16568 10164
rect 16716 10052 16772 11788
rect 17500 11844 17556 12126
rect 17500 11778 17556 11788
rect 16828 11506 16884 11518
rect 16828 11454 16830 11506
rect 16882 11454 16884 11506
rect 16828 10948 16884 11454
rect 17836 11508 17892 12238
rect 17836 11442 17892 11452
rect 17948 12292 18004 12302
rect 16940 11396 16996 11406
rect 16940 11394 17220 11396
rect 16940 11342 16942 11394
rect 16994 11342 17220 11394
rect 16940 11340 17220 11342
rect 16940 11330 16996 11340
rect 17164 11284 17220 11340
rect 17724 11284 17780 11294
rect 17164 11282 17780 11284
rect 17164 11230 17726 11282
rect 17778 11230 17780 11282
rect 17164 11228 17780 11230
rect 17948 11284 18004 12236
rect 18060 12180 18116 12190
rect 18060 12086 18116 12124
rect 18060 11284 18116 11294
rect 17948 11282 18116 11284
rect 17948 11230 18062 11282
rect 18114 11230 18116 11282
rect 17948 11228 18116 11230
rect 17724 11218 17780 11228
rect 16828 10892 17444 10948
rect 17388 10834 17444 10892
rect 17388 10782 17390 10834
rect 17442 10782 17444 10834
rect 17388 10770 17444 10782
rect 16828 10724 16884 10734
rect 17948 10724 18004 10734
rect 16828 10722 16996 10724
rect 16828 10670 16830 10722
rect 16882 10670 16996 10722
rect 16828 10668 16996 10670
rect 16828 10658 16884 10668
rect 16156 9090 16212 9100
rect 16604 9996 16772 10052
rect 16044 8932 16100 8942
rect 16604 8932 16660 9996
rect 16044 8838 16100 8876
rect 16156 8876 16660 8932
rect 16716 9044 16772 9054
rect 16156 8708 16212 8876
rect 15932 8306 15988 8316
rect 16044 8652 16212 8708
rect 16304 8652 16568 8662
rect 15820 8092 15988 8148
rect 15596 8054 15652 8092
rect 15596 7364 15652 7374
rect 15596 5122 15652 7308
rect 15596 5070 15598 5122
rect 15650 5070 15652 5122
rect 15596 5058 15652 5070
rect 15708 4900 15764 4910
rect 15596 4452 15652 4462
rect 15596 4358 15652 4396
rect 15484 3490 15540 3500
rect 15708 3442 15764 4844
rect 15820 4898 15876 4910
rect 15820 4846 15822 4898
rect 15874 4846 15876 4898
rect 15820 4338 15876 4846
rect 15820 4286 15822 4338
rect 15874 4286 15876 4338
rect 15820 4274 15876 4286
rect 15932 3554 15988 8092
rect 15932 3502 15934 3554
rect 15986 3502 15988 3554
rect 15932 3490 15988 3502
rect 15708 3390 15710 3442
rect 15762 3390 15764 3442
rect 15708 3378 15764 3390
rect 16044 3388 16100 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16304 8586 16568 8596
rect 16716 8484 16772 8988
rect 16268 8428 16772 8484
rect 16268 8260 16324 8428
rect 16828 8372 16884 8382
rect 16828 8278 16884 8316
rect 16156 8258 16324 8260
rect 16156 8206 16270 8258
rect 16322 8206 16324 8258
rect 16156 8204 16324 8206
rect 16156 6018 16212 8204
rect 16268 8194 16324 8204
rect 16716 8148 16772 8158
rect 16716 8054 16772 8092
rect 16828 7924 16884 7934
rect 16716 7476 16772 7486
rect 16716 7140 16772 7420
rect 16304 7084 16568 7094
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16716 7074 16772 7084
rect 16304 7018 16568 7028
rect 16828 6916 16884 7868
rect 16604 6860 16884 6916
rect 16156 5966 16158 6018
rect 16210 5966 16212 6018
rect 16156 5954 16212 5966
rect 16268 6578 16324 6590
rect 16268 6526 16270 6578
rect 16322 6526 16324 6578
rect 16268 5684 16324 6526
rect 16604 6468 16660 6860
rect 16604 6412 16772 6468
rect 16156 5628 16324 5684
rect 16156 4900 16212 5628
rect 16304 5516 16568 5526
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16304 5450 16568 5460
rect 16716 5010 16772 6412
rect 16716 4958 16718 5010
rect 16770 4958 16772 5010
rect 16716 4946 16772 4958
rect 16828 6244 16884 6254
rect 16156 4834 16212 4844
rect 16304 3948 16568 3958
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16304 3882 16568 3892
rect 16044 3332 16660 3388
rect 16156 3220 16212 3230
rect 15708 980 15764 990
rect 15708 800 15764 924
rect 16156 800 16212 3164
rect 16604 800 16660 3332
rect 16828 1764 16884 6188
rect 16940 4004 16996 10668
rect 18060 10724 18116 11228
rect 18460 11004 18724 11014
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18460 10938 18724 10948
rect 18060 10668 19124 10724
rect 17724 10610 17780 10622
rect 17724 10558 17726 10610
rect 17778 10558 17780 10610
rect 17052 9604 17108 9614
rect 17108 9548 17220 9604
rect 17052 9538 17108 9548
rect 17052 8146 17108 8158
rect 17052 8094 17054 8146
rect 17106 8094 17108 8146
rect 17052 7588 17108 8094
rect 17164 7924 17220 9548
rect 17388 9154 17444 9166
rect 17388 9102 17390 9154
rect 17442 9102 17444 9154
rect 17388 8596 17444 9102
rect 17612 9044 17668 9054
rect 17612 8950 17668 8988
rect 17724 8820 17780 10558
rect 17948 10052 18004 10668
rect 18172 10500 18228 10510
rect 18172 10406 18228 10444
rect 18844 10500 18900 10510
rect 17948 9996 18228 10052
rect 17948 8820 18004 8830
rect 17724 8818 18004 8820
rect 17724 8766 17950 8818
rect 18002 8766 18004 8818
rect 17724 8764 18004 8766
rect 17948 8754 18004 8764
rect 17388 8540 17780 8596
rect 17724 8372 17780 8540
rect 18060 8484 18116 9996
rect 18172 9938 18228 9996
rect 18172 9886 18174 9938
rect 18226 9886 18228 9938
rect 18172 9874 18228 9886
rect 18460 9436 18724 9446
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18460 9370 18724 9380
rect 18172 8932 18228 8942
rect 18172 8930 18340 8932
rect 18172 8878 18174 8930
rect 18226 8878 18340 8930
rect 18172 8876 18340 8878
rect 18172 8866 18228 8876
rect 18284 8818 18340 8876
rect 18284 8766 18286 8818
rect 18338 8766 18340 8818
rect 18060 8428 18228 8484
rect 17724 8316 18116 8372
rect 17276 8148 17332 8158
rect 17276 8054 17332 8092
rect 17724 8148 17780 8158
rect 17612 8036 17668 8046
rect 17612 7942 17668 7980
rect 17164 7868 17444 7924
rect 17052 7522 17108 7532
rect 17388 7586 17444 7868
rect 17612 7812 17668 7822
rect 17388 7534 17390 7586
rect 17442 7534 17444 7586
rect 17388 7522 17444 7534
rect 17500 7588 17556 7598
rect 17500 7494 17556 7532
rect 17612 7586 17668 7756
rect 17612 7534 17614 7586
rect 17666 7534 17668 7586
rect 17612 7522 17668 7534
rect 17276 6916 17332 6926
rect 17724 6916 17780 8092
rect 17948 8148 18004 8158
rect 17948 8054 18004 8092
rect 17948 7474 18004 7486
rect 17948 7422 17950 7474
rect 18002 7422 18004 7474
rect 17836 7252 17892 7262
rect 17836 7158 17892 7196
rect 17052 6578 17108 6590
rect 17052 6526 17054 6578
rect 17106 6526 17108 6578
rect 17052 4676 17108 6526
rect 17276 6132 17332 6860
rect 17500 6860 17780 6916
rect 17836 7028 17892 7038
rect 17388 6132 17444 6142
rect 17276 6130 17444 6132
rect 17276 6078 17390 6130
rect 17442 6078 17444 6130
rect 17276 6076 17444 6078
rect 17388 6066 17444 6076
rect 17500 6130 17556 6860
rect 17612 6692 17668 6702
rect 17668 6636 17780 6692
rect 17612 6626 17668 6636
rect 17500 6078 17502 6130
rect 17554 6078 17556 6130
rect 17500 6066 17556 6078
rect 17612 6356 17668 6366
rect 17612 6130 17668 6300
rect 17612 6078 17614 6130
rect 17666 6078 17668 6130
rect 17612 6066 17668 6078
rect 17724 5124 17780 6636
rect 17612 5068 17780 5124
rect 17612 5010 17668 5068
rect 17612 4958 17614 5010
rect 17666 4958 17668 5010
rect 17612 4946 17668 4958
rect 17836 4900 17892 6972
rect 17948 6468 18004 7422
rect 18060 6692 18116 8316
rect 18172 6916 18228 8428
rect 18172 6850 18228 6860
rect 18172 6692 18228 6702
rect 18060 6690 18228 6692
rect 18060 6638 18174 6690
rect 18226 6638 18228 6690
rect 18060 6636 18228 6638
rect 18172 6626 18228 6636
rect 17948 6132 18004 6412
rect 18172 6244 18228 6254
rect 18284 6244 18340 8766
rect 18460 7868 18724 7878
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18460 7802 18724 7812
rect 18228 6188 18340 6244
rect 18460 6300 18724 6310
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18460 6234 18724 6244
rect 18172 6178 18228 6188
rect 17948 6076 18116 6132
rect 17948 5908 18004 5918
rect 17948 5814 18004 5852
rect 17948 5124 18004 5134
rect 17948 5030 18004 5068
rect 17836 4844 18004 4900
rect 17052 4620 17444 4676
rect 17388 4562 17444 4620
rect 17388 4510 17390 4562
rect 17442 4510 17444 4562
rect 17388 4498 17444 4510
rect 17612 4340 17668 4350
rect 17612 4246 17668 4284
rect 16940 3948 17892 4004
rect 17836 3666 17892 3948
rect 17836 3614 17838 3666
rect 17890 3614 17892 3666
rect 17836 3602 17892 3614
rect 17164 3554 17220 3566
rect 17164 3502 17166 3554
rect 17218 3502 17220 3554
rect 16940 3444 16996 3482
rect 16940 3378 16996 3388
rect 17164 3332 17220 3502
rect 17164 3266 17220 3276
rect 17500 3444 17556 3454
rect 16828 1708 17108 1764
rect 17052 800 17108 1708
rect 17500 800 17556 3388
rect 17948 800 18004 4844
rect 18060 4564 18116 6076
rect 18172 5908 18228 5918
rect 18228 5852 18340 5908
rect 18172 5842 18228 5852
rect 18172 4564 18228 4574
rect 18060 4562 18228 4564
rect 18060 4510 18174 4562
rect 18226 4510 18228 4562
rect 18060 4508 18228 4510
rect 18172 4498 18228 4508
rect 18172 3668 18228 3678
rect 18284 3668 18340 5852
rect 18460 4732 18724 4742
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18460 4666 18724 4676
rect 18844 3892 18900 10444
rect 18956 8148 19012 8158
rect 18956 4116 19012 8092
rect 18956 4050 19012 4060
rect 18844 3826 18900 3836
rect 18172 3666 18340 3668
rect 18172 3614 18174 3666
rect 18226 3614 18340 3666
rect 18172 3612 18340 3614
rect 18844 3666 18900 3678
rect 18844 3614 18846 3666
rect 18898 3614 18900 3666
rect 18172 3602 18228 3612
rect 18460 3164 18724 3174
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18460 3098 18724 3108
rect 18844 1764 18900 3614
rect 18956 3444 19012 3454
rect 19068 3444 19124 10668
rect 19012 3388 19124 3444
rect 18956 3378 19012 3388
rect 19180 2994 19236 12686
rect 19404 10388 19460 10398
rect 19292 9940 19348 9950
rect 19292 5908 19348 9884
rect 19292 5842 19348 5852
rect 19404 3666 19460 10332
rect 19404 3614 19406 3666
rect 19458 3614 19460 3666
rect 19404 3602 19460 3614
rect 19180 2942 19182 2994
rect 19234 2942 19236 2994
rect 19180 2930 19236 2942
rect 18396 1708 18900 1764
rect 18396 800 18452 1708
rect 1344 0 1456 800
rect 1792 0 1904 800
rect 2240 0 2352 800
rect 2688 0 2800 800
rect 3136 0 3248 800
rect 3584 0 3696 800
rect 4032 0 4144 800
rect 4480 0 4592 800
rect 4928 0 5040 800
rect 5376 0 5488 800
rect 5824 0 5936 800
rect 6272 0 6384 800
rect 6720 0 6832 800
rect 7168 0 7280 800
rect 7616 0 7728 800
rect 8064 0 8176 800
rect 8512 0 8624 800
rect 8960 0 9072 800
rect 9408 0 9520 800
rect 9856 0 9968 800
rect 10304 0 10416 800
rect 10752 0 10864 800
rect 11200 0 11312 800
rect 11648 0 11760 800
rect 12096 0 12208 800
rect 12544 0 12656 800
rect 12992 0 13104 800
rect 13440 0 13552 800
rect 13888 0 14000 800
rect 14336 0 14448 800
rect 14784 0 14896 800
rect 15232 0 15344 800
rect 15680 0 15792 800
rect 16128 0 16240 800
rect 16576 0 16688 800
rect 17024 0 17136 800
rect 17472 0 17584 800
rect 17920 0 18032 800
rect 18368 0 18480 800
<< via2 >>
rect 1708 15260 1764 15316
rect 1708 11900 1764 11956
rect 1708 11170 1764 11172
rect 1708 11118 1710 11170
rect 1710 11118 1762 11170
rect 1762 11118 1764 11170
rect 1708 11116 1764 11118
rect 1372 10556 1428 10612
rect 1260 8316 1316 8372
rect 1260 7532 1316 7588
rect 1708 10332 1764 10388
rect 1932 13020 1988 13076
rect 1932 12012 1988 12068
rect 4732 14812 4788 14868
rect 4284 14364 4340 14420
rect 3500 13916 3556 13972
rect 2828 13468 2884 13524
rect 2604 12572 2660 12628
rect 2156 12290 2212 12292
rect 2156 12238 2158 12290
rect 2158 12238 2210 12290
rect 2210 12238 2212 12290
rect 2156 12236 2212 12238
rect 2156 11282 2212 11284
rect 2156 11230 2158 11282
rect 2158 11230 2210 11282
rect 2210 11230 2212 11282
rect 2156 11228 2212 11230
rect 5524 12570 5580 12572
rect 5524 12518 5526 12570
rect 5526 12518 5578 12570
rect 5578 12518 5580 12570
rect 5524 12516 5580 12518
rect 5628 12570 5684 12572
rect 5628 12518 5630 12570
rect 5630 12518 5682 12570
rect 5682 12518 5684 12570
rect 5628 12516 5684 12518
rect 5732 12570 5788 12572
rect 5732 12518 5734 12570
rect 5734 12518 5786 12570
rect 5786 12518 5788 12570
rect 5732 12516 5788 12518
rect 9836 12570 9892 12572
rect 9836 12518 9838 12570
rect 9838 12518 9890 12570
rect 9890 12518 9892 12570
rect 9836 12516 9892 12518
rect 9940 12570 9996 12572
rect 9940 12518 9942 12570
rect 9942 12518 9994 12570
rect 9994 12518 9996 12570
rect 9940 12516 9996 12518
rect 10044 12570 10100 12572
rect 10044 12518 10046 12570
rect 10046 12518 10098 12570
rect 10098 12518 10100 12570
rect 10044 12516 10100 12518
rect 14148 12570 14204 12572
rect 14148 12518 14150 12570
rect 14150 12518 14202 12570
rect 14202 12518 14204 12570
rect 14148 12516 14204 12518
rect 14252 12570 14308 12572
rect 14252 12518 14254 12570
rect 14254 12518 14306 12570
rect 14306 12518 14308 12570
rect 14252 12516 14308 12518
rect 14356 12570 14412 12572
rect 14356 12518 14358 12570
rect 14358 12518 14410 12570
rect 14410 12518 14412 12570
rect 14356 12516 14412 12518
rect 12348 12348 12404 12404
rect 13580 12348 13636 12404
rect 3368 11786 3424 11788
rect 3368 11734 3370 11786
rect 3370 11734 3422 11786
rect 3422 11734 3424 11786
rect 3368 11732 3424 11734
rect 3472 11786 3528 11788
rect 3472 11734 3474 11786
rect 3474 11734 3526 11786
rect 3526 11734 3528 11786
rect 3472 11732 3528 11734
rect 3576 11786 3632 11788
rect 3576 11734 3578 11786
rect 3578 11734 3630 11786
rect 3630 11734 3632 11786
rect 3576 11732 3632 11734
rect 1932 10332 1988 10388
rect 1820 8764 1876 8820
rect 1484 7756 1540 7812
rect 1708 7586 1764 7588
rect 1708 7534 1710 7586
rect 1710 7534 1762 7586
rect 1762 7534 1764 7586
rect 1708 7532 1764 7534
rect 1596 6636 1652 6692
rect 1484 4508 1540 4564
rect 1372 3500 1428 3556
rect 1820 6690 1876 6692
rect 1820 6638 1822 6690
rect 1822 6638 1874 6690
rect 1874 6638 1876 6690
rect 1820 6636 1876 6638
rect 2604 9884 2660 9940
rect 2044 9660 2100 9716
rect 2156 9602 2212 9604
rect 2156 9550 2158 9602
rect 2158 9550 2210 9602
rect 2210 9550 2212 9602
rect 2156 9548 2212 9550
rect 2156 8540 2212 8596
rect 2268 9100 2324 9156
rect 2156 8092 2212 8148
rect 2044 7980 2100 8036
rect 2156 6860 2212 6916
rect 2044 6636 2100 6692
rect 1820 5122 1876 5124
rect 1820 5070 1822 5122
rect 1822 5070 1874 5122
rect 1874 5070 1876 5122
rect 1820 5068 1876 5070
rect 1932 4396 1988 4452
rect 2156 6018 2212 6020
rect 2156 5966 2158 6018
rect 2158 5966 2210 6018
rect 2210 5966 2212 6018
rect 2156 5964 2212 5966
rect 2156 5180 2212 5236
rect 2380 8876 2436 8932
rect 2268 4620 2324 4676
rect 1708 2716 1764 2772
rect 1820 3948 1876 4004
rect 1932 3724 1988 3780
rect 2044 1820 2100 1876
rect 2156 1484 2212 1540
rect 2492 7474 2548 7476
rect 2492 7422 2494 7474
rect 2494 7422 2546 7474
rect 2546 7422 2548 7474
rect 2492 7420 2548 7422
rect 2492 6690 2548 6692
rect 2492 6638 2494 6690
rect 2494 6638 2546 6690
rect 2546 6638 2548 6690
rect 2492 6636 2548 6638
rect 3368 10218 3424 10220
rect 3368 10166 3370 10218
rect 3370 10166 3422 10218
rect 3422 10166 3424 10218
rect 3368 10164 3424 10166
rect 3472 10218 3528 10220
rect 3472 10166 3474 10218
rect 3474 10166 3526 10218
rect 3526 10166 3528 10218
rect 3472 10164 3528 10166
rect 3576 10218 3632 10220
rect 3576 10166 3578 10218
rect 3578 10166 3630 10218
rect 3630 10166 3632 10218
rect 3576 10164 3632 10166
rect 2828 8764 2884 8820
rect 2828 8428 2884 8484
rect 2716 8092 2772 8148
rect 2716 7420 2772 7476
rect 2604 5906 2660 5908
rect 2604 5854 2606 5906
rect 2606 5854 2658 5906
rect 2658 5854 2660 5906
rect 2604 5852 2660 5854
rect 2828 6636 2884 6692
rect 2716 5404 2772 5460
rect 2828 6130 2884 6132
rect 2828 6078 2830 6130
rect 2830 6078 2882 6130
rect 2882 6078 2884 6130
rect 2828 6076 2884 6078
rect 2828 5292 2884 5348
rect 2828 5122 2884 5124
rect 2828 5070 2830 5122
rect 2830 5070 2882 5122
rect 2882 5070 2884 5122
rect 2828 5068 2884 5070
rect 2492 4956 2548 5012
rect 3500 9602 3556 9604
rect 3500 9550 3502 9602
rect 3502 9550 3554 9602
rect 3554 9550 3556 9602
rect 3500 9548 3556 9550
rect 3164 9324 3220 9380
rect 3052 9154 3108 9156
rect 3052 9102 3054 9154
rect 3054 9102 3106 9154
rect 3106 9102 3108 9154
rect 3052 9100 3108 9102
rect 3276 9100 3332 9156
rect 3500 9154 3556 9156
rect 3500 9102 3502 9154
rect 3502 9102 3554 9154
rect 3554 9102 3556 9154
rect 3500 9100 3556 9102
rect 3276 8764 3332 8820
rect 3368 8650 3424 8652
rect 3368 8598 3370 8650
rect 3370 8598 3422 8650
rect 3422 8598 3424 8650
rect 3368 8596 3424 8598
rect 3472 8650 3528 8652
rect 3472 8598 3474 8650
rect 3474 8598 3526 8650
rect 3526 8598 3528 8650
rect 3472 8596 3528 8598
rect 3576 8650 3632 8652
rect 3576 8598 3578 8650
rect 3578 8598 3630 8650
rect 3630 8598 3632 8650
rect 3576 8596 3632 8598
rect 3164 8316 3220 8372
rect 3612 8316 3668 8372
rect 3052 6524 3108 6580
rect 3276 7868 3332 7924
rect 5628 12066 5684 12068
rect 5628 12014 5630 12066
rect 5630 12014 5682 12066
rect 5682 12014 5684 12066
rect 5628 12012 5684 12014
rect 3948 9772 4004 9828
rect 3948 9602 4004 9604
rect 3948 9550 3950 9602
rect 3950 9550 4002 9602
rect 4002 9550 4004 9602
rect 3948 9548 4004 9550
rect 3724 7644 3780 7700
rect 3500 7532 3556 7588
rect 3724 7420 3780 7476
rect 3368 7082 3424 7084
rect 3368 7030 3370 7082
rect 3370 7030 3422 7082
rect 3422 7030 3424 7082
rect 3368 7028 3424 7030
rect 3472 7082 3528 7084
rect 3472 7030 3474 7082
rect 3474 7030 3526 7082
rect 3526 7030 3528 7082
rect 3472 7028 3528 7030
rect 3576 7082 3632 7084
rect 3576 7030 3578 7082
rect 3578 7030 3630 7082
rect 3630 7030 3632 7082
rect 3576 7028 3632 7030
rect 3164 6188 3220 6244
rect 3276 6412 3332 6468
rect 3276 5628 3332 5684
rect 4396 9154 4452 9156
rect 4396 9102 4398 9154
rect 4398 9102 4450 9154
rect 4450 9102 4452 9154
rect 4396 9100 4452 9102
rect 4284 8204 4340 8260
rect 4396 8428 4452 8484
rect 4060 7980 4116 8036
rect 4060 7644 4116 7700
rect 4060 7474 4116 7476
rect 4060 7422 4062 7474
rect 4062 7422 4114 7474
rect 4114 7422 4116 7474
rect 4060 7420 4116 7422
rect 3948 7196 4004 7252
rect 3948 6972 4004 7028
rect 3836 6188 3892 6244
rect 4284 8034 4340 8036
rect 4284 7982 4286 8034
rect 4286 7982 4338 8034
rect 4338 7982 4340 8034
rect 4284 7980 4340 7982
rect 4172 6860 4228 6916
rect 4284 6188 4340 6244
rect 4172 6018 4228 6020
rect 4172 5966 4174 6018
rect 4174 5966 4226 6018
rect 4226 5966 4228 6018
rect 4172 5964 4228 5966
rect 4284 5852 4340 5908
rect 3368 5514 3424 5516
rect 3368 5462 3370 5514
rect 3370 5462 3422 5514
rect 3422 5462 3424 5514
rect 3368 5460 3424 5462
rect 3472 5514 3528 5516
rect 3472 5462 3474 5514
rect 3474 5462 3526 5514
rect 3526 5462 3528 5514
rect 3472 5460 3528 5462
rect 3576 5514 3632 5516
rect 3576 5462 3578 5514
rect 3578 5462 3630 5514
rect 3630 5462 3632 5514
rect 3576 5460 3632 5462
rect 3724 5404 3780 5460
rect 3612 5292 3668 5348
rect 3388 5180 3444 5236
rect 3500 4956 3556 5012
rect 2380 3612 2436 3668
rect 2940 4562 2996 4564
rect 2940 4510 2942 4562
rect 2942 4510 2994 4562
rect 2994 4510 2996 4562
rect 2940 4508 2996 4510
rect 3500 4396 3556 4452
rect 3836 4620 3892 4676
rect 3948 5068 4004 5124
rect 4060 5292 4116 5348
rect 3052 3948 3108 4004
rect 2604 3164 2660 3220
rect 2716 3836 2772 3892
rect 2828 3554 2884 3556
rect 2828 3502 2830 3554
rect 2830 3502 2882 3554
rect 2882 3502 2884 3554
rect 2828 3500 2884 3502
rect 2940 2770 2996 2772
rect 2940 2718 2942 2770
rect 2942 2718 2994 2770
rect 2994 2718 2996 2770
rect 2940 2716 2996 2718
rect 3368 3946 3424 3948
rect 3368 3894 3370 3946
rect 3370 3894 3422 3946
rect 3422 3894 3424 3946
rect 3368 3892 3424 3894
rect 3472 3946 3528 3948
rect 3472 3894 3474 3946
rect 3474 3894 3526 3946
rect 3526 3894 3528 3946
rect 3472 3892 3528 3894
rect 3576 3946 3632 3948
rect 3576 3894 3578 3946
rect 3578 3894 3630 3946
rect 3630 3894 3632 3946
rect 3576 3892 3632 3894
rect 3388 812 3444 868
rect 4060 3554 4116 3556
rect 4060 3502 4062 3554
rect 4062 3502 4114 3554
rect 4114 3502 4116 3554
rect 4060 3500 4116 3502
rect 4956 11170 5012 11172
rect 4956 11118 4958 11170
rect 4958 11118 5010 11170
rect 5010 11118 5012 11170
rect 4956 11116 5012 11118
rect 5524 11002 5580 11004
rect 5524 10950 5526 11002
rect 5526 10950 5578 11002
rect 5578 10950 5580 11002
rect 5524 10948 5580 10950
rect 5628 11002 5684 11004
rect 5628 10950 5630 11002
rect 5630 10950 5682 11002
rect 5682 10950 5684 11002
rect 5628 10948 5684 10950
rect 5732 11002 5788 11004
rect 5732 10950 5734 11002
rect 5734 10950 5786 11002
rect 5786 10950 5788 11002
rect 5732 10948 5788 10950
rect 5852 10668 5908 10724
rect 4956 10108 5012 10164
rect 4620 8146 4676 8148
rect 4620 8094 4622 8146
rect 4622 8094 4674 8146
rect 4674 8094 4676 8146
rect 4620 8092 4676 8094
rect 4508 7420 4564 7476
rect 4620 6972 4676 7028
rect 4508 6076 4564 6132
rect 4508 5906 4564 5908
rect 4508 5854 4510 5906
rect 4510 5854 4562 5906
rect 4562 5854 4564 5906
rect 4508 5852 4564 5854
rect 4508 5628 4564 5684
rect 5524 9434 5580 9436
rect 5524 9382 5526 9434
rect 5526 9382 5578 9434
rect 5578 9382 5580 9434
rect 5524 9380 5580 9382
rect 5628 9434 5684 9436
rect 5628 9382 5630 9434
rect 5630 9382 5682 9434
rect 5682 9382 5684 9434
rect 5628 9380 5684 9382
rect 5732 9434 5788 9436
rect 5732 9382 5734 9434
rect 5734 9382 5786 9434
rect 5786 9382 5788 9434
rect 5732 9380 5788 9382
rect 5180 9042 5236 9044
rect 5180 8990 5182 9042
rect 5182 8990 5234 9042
rect 5234 8990 5236 9042
rect 5180 8988 5236 8990
rect 5292 8428 5348 8484
rect 6300 10444 6356 10500
rect 6076 10108 6132 10164
rect 5964 8204 6020 8260
rect 6076 8092 6132 8148
rect 5068 7868 5124 7924
rect 5068 7084 5124 7140
rect 4732 6188 4788 6244
rect 4956 5964 5012 6020
rect 4956 5740 5012 5796
rect 4732 5292 4788 5348
rect 4732 4844 4788 4900
rect 5068 5628 5124 5684
rect 5524 7866 5580 7868
rect 5524 7814 5526 7866
rect 5526 7814 5578 7866
rect 5578 7814 5580 7866
rect 5524 7812 5580 7814
rect 5628 7866 5684 7868
rect 5628 7814 5630 7866
rect 5630 7814 5682 7866
rect 5682 7814 5684 7866
rect 5628 7812 5684 7814
rect 5732 7866 5788 7868
rect 5732 7814 5734 7866
rect 5734 7814 5786 7866
rect 5786 7814 5788 7866
rect 5732 7812 5788 7814
rect 5852 6636 5908 6692
rect 5524 6298 5580 6300
rect 5524 6246 5526 6298
rect 5526 6246 5578 6298
rect 5578 6246 5580 6298
rect 5524 6244 5580 6246
rect 5628 6298 5684 6300
rect 5628 6246 5630 6298
rect 5630 6246 5682 6298
rect 5682 6246 5684 6298
rect 5628 6244 5684 6246
rect 5732 6298 5788 6300
rect 5732 6246 5734 6298
rect 5734 6246 5786 6298
rect 5786 6246 5788 6298
rect 5732 6244 5788 6246
rect 5964 6466 6020 6468
rect 5964 6414 5966 6466
rect 5966 6414 6018 6466
rect 6018 6414 6020 6466
rect 5964 6412 6020 6414
rect 5068 5068 5124 5124
rect 5180 4844 5236 4900
rect 5068 4732 5124 4788
rect 5068 4396 5124 4452
rect 4620 3442 4676 3444
rect 4620 3390 4622 3442
rect 4622 3390 4674 3442
rect 4674 3390 4676 3442
rect 4620 3388 4676 3390
rect 4060 3276 4116 3332
rect 5068 3948 5124 4004
rect 5964 5852 6020 5908
rect 6300 7196 6356 7252
rect 6412 7980 6468 8036
rect 6188 6636 6244 6692
rect 7680 11786 7736 11788
rect 7680 11734 7682 11786
rect 7682 11734 7734 11786
rect 7734 11734 7736 11786
rect 7680 11732 7736 11734
rect 7784 11786 7840 11788
rect 7784 11734 7786 11786
rect 7786 11734 7838 11786
rect 7838 11734 7840 11786
rect 7784 11732 7840 11734
rect 7888 11786 7944 11788
rect 7888 11734 7890 11786
rect 7890 11734 7942 11786
rect 7942 11734 7944 11786
rect 7888 11732 7944 11734
rect 6972 10668 7028 10724
rect 6636 9548 6692 9604
rect 6524 6972 6580 7028
rect 6636 9324 6692 9380
rect 7308 10220 7364 10276
rect 11676 11170 11732 11172
rect 11676 11118 11678 11170
rect 11678 11118 11730 11170
rect 11730 11118 11732 11170
rect 11676 11116 11732 11118
rect 9836 11002 9892 11004
rect 9836 10950 9838 11002
rect 9838 10950 9890 11002
rect 9890 10950 9892 11002
rect 9836 10948 9892 10950
rect 9940 11002 9996 11004
rect 9940 10950 9942 11002
rect 9942 10950 9994 11002
rect 9994 10950 9996 11002
rect 9940 10948 9996 10950
rect 10044 11002 10100 11004
rect 10044 10950 10046 11002
rect 10046 10950 10098 11002
rect 10098 10950 10100 11002
rect 10044 10948 10100 10950
rect 8988 10722 9044 10724
rect 8988 10670 8990 10722
rect 8990 10670 9042 10722
rect 9042 10670 9044 10722
rect 8988 10668 9044 10670
rect 10220 10668 10276 10724
rect 8204 10610 8260 10612
rect 8204 10558 8206 10610
rect 8206 10558 8258 10610
rect 8258 10558 8260 10610
rect 8204 10556 8260 10558
rect 7756 10332 7812 10388
rect 7680 10218 7736 10220
rect 7680 10166 7682 10218
rect 7682 10166 7734 10218
rect 7734 10166 7736 10218
rect 7680 10164 7736 10166
rect 7784 10218 7840 10220
rect 7784 10166 7786 10218
rect 7786 10166 7838 10218
rect 7838 10166 7840 10218
rect 7784 10164 7840 10166
rect 7888 10218 7944 10220
rect 7888 10166 7890 10218
rect 7890 10166 7942 10218
rect 7942 10166 7944 10218
rect 7888 10164 7944 10166
rect 7532 9996 7588 10052
rect 10668 10722 10724 10724
rect 10668 10670 10670 10722
rect 10670 10670 10722 10722
rect 10722 10670 10724 10722
rect 10668 10668 10724 10670
rect 11992 11786 12048 11788
rect 11992 11734 11994 11786
rect 11994 11734 12046 11786
rect 12046 11734 12048 11786
rect 11992 11732 12048 11734
rect 12096 11786 12152 11788
rect 12096 11734 12098 11786
rect 12098 11734 12150 11786
rect 12150 11734 12152 11786
rect 12096 11732 12152 11734
rect 12200 11786 12256 11788
rect 12200 11734 12202 11786
rect 12202 11734 12254 11786
rect 12254 11734 12256 11786
rect 12200 11732 12256 11734
rect 12684 11340 12740 11396
rect 13132 11676 13188 11732
rect 12124 11170 12180 11172
rect 12124 11118 12126 11170
rect 12126 11118 12178 11170
rect 12178 11118 12180 11170
rect 12124 11116 12180 11118
rect 11788 10556 11844 10612
rect 11228 10220 11284 10276
rect 10220 9996 10276 10052
rect 10668 9884 10724 9940
rect 7196 8540 7252 8596
rect 6860 8092 6916 8148
rect 6636 7532 6692 7588
rect 6524 6578 6580 6580
rect 6524 6526 6526 6578
rect 6526 6526 6578 6578
rect 6578 6526 6580 6578
rect 6524 6524 6580 6526
rect 5852 5180 5908 5236
rect 6524 5740 6580 5796
rect 6748 6748 6804 6804
rect 6860 6972 6916 7028
rect 6300 5404 6356 5460
rect 5524 4730 5580 4732
rect 5524 4678 5526 4730
rect 5526 4678 5578 4730
rect 5578 4678 5580 4730
rect 5524 4676 5580 4678
rect 5628 4730 5684 4732
rect 5628 4678 5630 4730
rect 5630 4678 5682 4730
rect 5682 4678 5684 4730
rect 5628 4676 5684 4678
rect 5732 4730 5788 4732
rect 5732 4678 5734 4730
rect 5734 4678 5786 4730
rect 5786 4678 5788 4730
rect 5732 4676 5788 4678
rect 5964 4732 6020 4788
rect 5964 4396 6020 4452
rect 5852 3442 5908 3444
rect 5852 3390 5854 3442
rect 5854 3390 5906 3442
rect 5906 3390 5908 3442
rect 5852 3388 5908 3390
rect 5524 3162 5580 3164
rect 5524 3110 5526 3162
rect 5526 3110 5578 3162
rect 5578 3110 5580 3162
rect 5524 3108 5580 3110
rect 5628 3162 5684 3164
rect 5628 3110 5630 3162
rect 5630 3110 5682 3162
rect 5682 3110 5684 3162
rect 5628 3108 5684 3110
rect 5732 3162 5788 3164
rect 5732 3110 5734 3162
rect 5734 3110 5786 3162
rect 5786 3110 5788 3162
rect 5732 3108 5788 3110
rect 6636 5180 6692 5236
rect 6636 4508 6692 4564
rect 6524 3500 6580 3556
rect 6748 3500 6804 3556
rect 7084 7420 7140 7476
rect 7196 6972 7252 7028
rect 7196 6748 7252 6804
rect 7084 6578 7140 6580
rect 7084 6526 7086 6578
rect 7086 6526 7138 6578
rect 7138 6526 7140 6578
rect 7084 6524 7140 6526
rect 7980 8764 8036 8820
rect 7532 8652 7588 8708
rect 7680 8650 7736 8652
rect 7680 8598 7682 8650
rect 7682 8598 7734 8650
rect 7734 8598 7736 8650
rect 7680 8596 7736 8598
rect 7784 8650 7840 8652
rect 7784 8598 7786 8650
rect 7786 8598 7838 8650
rect 7838 8598 7840 8650
rect 7784 8596 7840 8598
rect 7888 8650 7944 8652
rect 7888 8598 7890 8650
rect 7890 8598 7942 8650
rect 7942 8598 7944 8650
rect 7888 8596 7944 8598
rect 7868 8146 7924 8148
rect 7868 8094 7870 8146
rect 7870 8094 7922 8146
rect 7922 8094 7924 8146
rect 7868 8092 7924 8094
rect 7644 7980 7700 8036
rect 7868 7756 7924 7812
rect 8092 7474 8148 7476
rect 8092 7422 8094 7474
rect 8094 7422 8146 7474
rect 8146 7422 8148 7474
rect 8092 7420 8148 7422
rect 7680 7082 7736 7084
rect 7680 7030 7682 7082
rect 7682 7030 7734 7082
rect 7734 7030 7736 7082
rect 7680 7028 7736 7030
rect 7784 7082 7840 7084
rect 7784 7030 7786 7082
rect 7786 7030 7838 7082
rect 7838 7030 7840 7082
rect 7784 7028 7840 7030
rect 7888 7082 7944 7084
rect 7888 7030 7890 7082
rect 7890 7030 7942 7082
rect 7942 7030 7944 7082
rect 7888 7028 7944 7030
rect 7420 6578 7476 6580
rect 7420 6526 7422 6578
rect 7422 6526 7474 6578
rect 7474 6526 7476 6578
rect 7420 6524 7476 6526
rect 7308 5292 7364 5348
rect 7756 6188 7812 6244
rect 7868 6076 7924 6132
rect 7680 5514 7736 5516
rect 7680 5462 7682 5514
rect 7682 5462 7734 5514
rect 7734 5462 7736 5514
rect 7680 5460 7736 5462
rect 7784 5514 7840 5516
rect 7784 5462 7786 5514
rect 7786 5462 7838 5514
rect 7838 5462 7840 5514
rect 7784 5460 7840 5462
rect 7888 5514 7944 5516
rect 7888 5462 7890 5514
rect 7890 5462 7942 5514
rect 7942 5462 7944 5514
rect 7888 5460 7944 5462
rect 7680 3946 7736 3948
rect 7680 3894 7682 3946
rect 7682 3894 7734 3946
rect 7734 3894 7736 3946
rect 7680 3892 7736 3894
rect 7784 3946 7840 3948
rect 7784 3894 7786 3946
rect 7786 3894 7838 3946
rect 7838 3894 7840 3946
rect 7784 3892 7840 3894
rect 7888 3946 7944 3948
rect 7888 3894 7890 3946
rect 7890 3894 7942 3946
rect 7942 3894 7944 3946
rect 7888 3892 7944 3894
rect 8876 9212 8932 9268
rect 8428 8316 8484 8372
rect 8988 8764 9044 8820
rect 8316 5964 8372 6020
rect 8540 7532 8596 7588
rect 8652 6636 8708 6692
rect 8652 5740 8708 5796
rect 8876 5292 8932 5348
rect 8428 4956 8484 5012
rect 8316 4284 8372 4340
rect 7308 3388 7364 3444
rect 7532 3500 7588 3556
rect 8204 3612 8260 3668
rect 8540 3948 8596 4004
rect 10556 9714 10612 9716
rect 10556 9662 10558 9714
rect 10558 9662 10610 9714
rect 10610 9662 10612 9714
rect 10556 9660 10612 9662
rect 9836 9434 9892 9436
rect 9836 9382 9838 9434
rect 9838 9382 9890 9434
rect 9890 9382 9892 9434
rect 9836 9380 9892 9382
rect 9940 9434 9996 9436
rect 9940 9382 9942 9434
rect 9942 9382 9994 9434
rect 9994 9382 9996 9434
rect 9940 9380 9996 9382
rect 10044 9434 10100 9436
rect 10044 9382 10046 9434
rect 10046 9382 10098 9434
rect 10098 9382 10100 9434
rect 10044 9380 10100 9382
rect 9836 7866 9892 7868
rect 9836 7814 9838 7866
rect 9838 7814 9890 7866
rect 9890 7814 9892 7866
rect 9836 7812 9892 7814
rect 9940 7866 9996 7868
rect 9940 7814 9942 7866
rect 9942 7814 9994 7866
rect 9994 7814 9996 7866
rect 9940 7812 9996 7814
rect 10044 7866 10100 7868
rect 10044 7814 10046 7866
rect 10046 7814 10098 7866
rect 10098 7814 10100 7866
rect 10044 7812 10100 7814
rect 9660 7474 9716 7476
rect 9660 7422 9662 7474
rect 9662 7422 9714 7474
rect 9714 7422 9716 7474
rect 9660 7420 9716 7422
rect 9324 5964 9380 6020
rect 10556 8876 10612 8932
rect 10332 6860 10388 6916
rect 10444 7308 10500 7364
rect 10108 6524 10164 6580
rect 10332 6636 10388 6692
rect 9836 6298 9892 6300
rect 9836 6246 9838 6298
rect 9838 6246 9890 6298
rect 9890 6246 9892 6298
rect 9836 6244 9892 6246
rect 9940 6298 9996 6300
rect 9940 6246 9942 6298
rect 9942 6246 9994 6298
rect 9994 6246 9996 6298
rect 9940 6244 9996 6246
rect 10044 6298 10100 6300
rect 10044 6246 10046 6298
rect 10046 6246 10098 6298
rect 10098 6246 10100 6298
rect 10044 6244 10100 6246
rect 9548 5628 9604 5684
rect 9100 5122 9156 5124
rect 9100 5070 9102 5122
rect 9102 5070 9154 5122
rect 9154 5070 9156 5122
rect 9100 5068 9156 5070
rect 8988 4956 9044 5012
rect 9884 6018 9940 6020
rect 9884 5966 9886 6018
rect 9886 5966 9938 6018
rect 9938 5966 9940 6018
rect 9884 5964 9940 5966
rect 9660 4844 9716 4900
rect 10108 5852 10164 5908
rect 10108 5292 10164 5348
rect 10220 5068 10276 5124
rect 9884 4844 9940 4900
rect 9996 4956 10052 5012
rect 9836 4730 9892 4732
rect 9836 4678 9838 4730
rect 9838 4678 9890 4730
rect 9890 4678 9892 4730
rect 9836 4676 9892 4678
rect 9940 4730 9996 4732
rect 9940 4678 9942 4730
rect 9942 4678 9994 4730
rect 9994 4678 9996 4730
rect 9940 4676 9996 4678
rect 10044 4730 10100 4732
rect 10044 4678 10046 4730
rect 10046 4678 10098 4730
rect 10098 4678 10100 4730
rect 10220 4732 10276 4788
rect 10044 4676 10100 4678
rect 9660 4562 9716 4564
rect 9660 4510 9662 4562
rect 9662 4510 9714 4562
rect 9714 4510 9716 4562
rect 9660 4508 9716 4510
rect 9772 4396 9828 4452
rect 8988 4172 9044 4228
rect 8428 3500 8484 3556
rect 8764 3554 8820 3556
rect 8764 3502 8766 3554
rect 8766 3502 8818 3554
rect 8818 3502 8820 3554
rect 8764 3500 8820 3502
rect 7196 2716 7252 2772
rect 7644 2604 7700 2660
rect 8540 2940 8596 2996
rect 9324 3612 9380 3668
rect 10220 3442 10276 3444
rect 10220 3390 10222 3442
rect 10222 3390 10274 3442
rect 10274 3390 10276 3442
rect 10220 3388 10276 3390
rect 9836 3162 9892 3164
rect 9836 3110 9838 3162
rect 9838 3110 9890 3162
rect 9890 3110 9892 3162
rect 9836 3108 9892 3110
rect 9940 3162 9996 3164
rect 9940 3110 9942 3162
rect 9942 3110 9994 3162
rect 9994 3110 9996 3162
rect 9940 3108 9996 3110
rect 10044 3162 10100 3164
rect 10044 3110 10046 3162
rect 10046 3110 10098 3162
rect 10098 3110 10100 3162
rect 10044 3108 10100 3110
rect 9884 2828 9940 2884
rect 9436 1036 9492 1092
rect 10892 8092 10948 8148
rect 11116 8428 11172 8484
rect 10668 6860 10724 6916
rect 11452 9772 11508 9828
rect 11340 9714 11396 9716
rect 11340 9662 11342 9714
rect 11342 9662 11394 9714
rect 11394 9662 11396 9714
rect 11340 9660 11396 9662
rect 11228 7980 11284 8036
rect 11452 7532 11508 7588
rect 11228 7362 11284 7364
rect 11228 7310 11230 7362
rect 11230 7310 11282 7362
rect 11282 7310 11284 7362
rect 11228 7308 11284 7310
rect 10780 5068 10836 5124
rect 10780 4620 10836 4676
rect 10780 4396 10836 4452
rect 11992 10218 12048 10220
rect 11992 10166 11994 10218
rect 11994 10166 12046 10218
rect 12046 10166 12048 10218
rect 11992 10164 12048 10166
rect 12096 10218 12152 10220
rect 12096 10166 12098 10218
rect 12098 10166 12150 10218
rect 12150 10166 12152 10218
rect 12096 10164 12152 10166
rect 12200 10218 12256 10220
rect 12200 10166 12202 10218
rect 12202 10166 12254 10218
rect 12254 10166 12256 10218
rect 12200 10164 12256 10166
rect 12124 9996 12180 10052
rect 12012 9660 12068 9716
rect 12012 8988 12068 9044
rect 11992 8650 12048 8652
rect 11992 8598 11994 8650
rect 11994 8598 12046 8650
rect 12046 8598 12048 8650
rect 11992 8596 12048 8598
rect 12096 8650 12152 8652
rect 12096 8598 12098 8650
rect 12098 8598 12150 8650
rect 12150 8598 12152 8650
rect 12096 8596 12152 8598
rect 12200 8650 12256 8652
rect 12200 8598 12202 8650
rect 12202 8598 12254 8650
rect 12254 8598 12256 8650
rect 12200 8596 12256 8598
rect 11788 8428 11844 8484
rect 12460 9714 12516 9716
rect 12460 9662 12462 9714
rect 12462 9662 12514 9714
rect 12514 9662 12516 9714
rect 12460 9660 12516 9662
rect 12572 9602 12628 9604
rect 12572 9550 12574 9602
rect 12574 9550 12626 9602
rect 12626 9550 12628 9602
rect 12572 9548 12628 9550
rect 11992 7082 12048 7084
rect 11992 7030 11994 7082
rect 11994 7030 12046 7082
rect 12046 7030 12048 7082
rect 11992 7028 12048 7030
rect 12096 7082 12152 7084
rect 12096 7030 12098 7082
rect 12098 7030 12150 7082
rect 12150 7030 12152 7082
rect 12096 7028 12152 7030
rect 12200 7082 12256 7084
rect 12200 7030 12202 7082
rect 12202 7030 12254 7082
rect 12254 7030 12256 7082
rect 12200 7028 12256 7030
rect 11004 5964 11060 6020
rect 11340 5122 11396 5124
rect 11340 5070 11342 5122
rect 11342 5070 11394 5122
rect 11394 5070 11396 5122
rect 11340 5068 11396 5070
rect 11228 4508 11284 4564
rect 10780 4172 10836 4228
rect 10668 3724 10724 3780
rect 10780 3836 10836 3892
rect 11340 3554 11396 3556
rect 11340 3502 11342 3554
rect 11342 3502 11394 3554
rect 11394 3502 11396 3554
rect 11340 3500 11396 3502
rect 11452 4844 11508 4900
rect 11564 4732 11620 4788
rect 11564 4284 11620 4340
rect 13020 11170 13076 11172
rect 13020 11118 13022 11170
rect 13022 11118 13074 11170
rect 13074 11118 13076 11170
rect 13020 11116 13076 11118
rect 13020 10498 13076 10500
rect 13020 10446 13022 10498
rect 13022 10446 13074 10498
rect 13074 10446 13076 10498
rect 13020 10444 13076 10446
rect 13132 10332 13188 10388
rect 13132 10108 13188 10164
rect 12684 7420 12740 7476
rect 12796 9602 12852 9604
rect 12796 9550 12798 9602
rect 12798 9550 12850 9602
rect 12850 9550 12852 9602
rect 12796 9548 12852 9550
rect 12572 7196 12628 7252
rect 12908 9436 12964 9492
rect 12460 5964 12516 6020
rect 11992 5514 12048 5516
rect 11992 5462 11994 5514
rect 11994 5462 12046 5514
rect 12046 5462 12048 5514
rect 11992 5460 12048 5462
rect 12096 5514 12152 5516
rect 12096 5462 12098 5514
rect 12098 5462 12150 5514
rect 12150 5462 12152 5514
rect 12096 5460 12152 5462
rect 12200 5514 12256 5516
rect 12200 5462 12202 5514
rect 12202 5462 12254 5514
rect 12254 5462 12256 5514
rect 12200 5460 12256 5462
rect 12348 4060 12404 4116
rect 11788 3948 11844 4004
rect 11992 3946 12048 3948
rect 11992 3894 11994 3946
rect 11994 3894 12046 3946
rect 12046 3894 12048 3946
rect 11992 3892 12048 3894
rect 12096 3946 12152 3948
rect 12096 3894 12098 3946
rect 12098 3894 12150 3946
rect 12150 3894 12152 3946
rect 12096 3892 12152 3894
rect 12200 3946 12256 3948
rect 12200 3894 12202 3946
rect 12202 3894 12254 3946
rect 12254 3894 12256 3946
rect 12200 3892 12256 3894
rect 12236 3778 12292 3780
rect 12236 3726 12238 3778
rect 12238 3726 12290 3778
rect 12290 3726 12292 3778
rect 12236 3724 12292 3726
rect 12908 6914 12964 6916
rect 12908 6862 12910 6914
rect 12910 6862 12962 6914
rect 12962 6862 12964 6914
rect 12908 6860 12964 6862
rect 12796 6466 12852 6468
rect 12796 6414 12798 6466
rect 12798 6414 12850 6466
rect 12850 6414 12852 6466
rect 12796 6412 12852 6414
rect 12796 5180 12852 5236
rect 13020 4284 13076 4340
rect 11788 3500 11844 3556
rect 12572 3500 12628 3556
rect 12572 3164 12628 3220
rect 16380 12402 16436 12404
rect 16380 12350 16382 12402
rect 16382 12350 16434 12402
rect 16434 12350 16436 12402
rect 16380 12348 16436 12350
rect 15820 12290 15876 12292
rect 15820 12238 15822 12290
rect 15822 12238 15874 12290
rect 15874 12238 15876 12290
rect 15820 12236 15876 12238
rect 18460 12570 18516 12572
rect 18460 12518 18462 12570
rect 18462 12518 18514 12570
rect 18514 12518 18516 12570
rect 18460 12516 18516 12518
rect 18564 12570 18620 12572
rect 18564 12518 18566 12570
rect 18566 12518 18618 12570
rect 18618 12518 18620 12570
rect 18564 12516 18620 12518
rect 18668 12570 18724 12572
rect 18668 12518 18670 12570
rect 18670 12518 18722 12570
rect 18722 12518 18724 12570
rect 18668 12516 18724 12518
rect 17276 12348 17332 12404
rect 14924 12178 14980 12180
rect 14924 12126 14926 12178
rect 14926 12126 14978 12178
rect 14978 12126 14980 12178
rect 14924 12124 14980 12126
rect 15372 11900 15428 11956
rect 14476 11676 14532 11732
rect 16304 11786 16360 11788
rect 16304 11734 16306 11786
rect 16306 11734 16358 11786
rect 16358 11734 16360 11786
rect 16304 11732 16360 11734
rect 16408 11786 16464 11788
rect 16408 11734 16410 11786
rect 16410 11734 16462 11786
rect 16462 11734 16464 11786
rect 16408 11732 16464 11734
rect 16512 11786 16568 11788
rect 16512 11734 16514 11786
rect 16514 11734 16566 11786
rect 16566 11734 16568 11786
rect 16512 11732 16568 11734
rect 16716 11788 16772 11844
rect 14588 11452 14644 11508
rect 13692 11282 13748 11284
rect 13692 11230 13694 11282
rect 13694 11230 13746 11282
rect 13746 11230 13748 11282
rect 13692 11228 13748 11230
rect 13244 9772 13300 9828
rect 13356 11116 13412 11172
rect 14140 11170 14196 11172
rect 14140 11118 14142 11170
rect 14142 11118 14194 11170
rect 14194 11118 14196 11170
rect 14140 11116 14196 11118
rect 14148 11002 14204 11004
rect 14148 10950 14150 11002
rect 14150 10950 14202 11002
rect 14202 10950 14204 11002
rect 14148 10948 14204 10950
rect 14252 11002 14308 11004
rect 14252 10950 14254 11002
rect 14254 10950 14306 11002
rect 14306 10950 14308 11002
rect 14252 10948 14308 10950
rect 14356 11002 14412 11004
rect 14356 10950 14358 11002
rect 14358 10950 14410 11002
rect 14410 10950 14412 11002
rect 14356 10948 14412 10950
rect 13468 8370 13524 8372
rect 13468 8318 13470 8370
rect 13470 8318 13522 8370
rect 13522 8318 13524 8370
rect 13468 8316 13524 8318
rect 13468 8092 13524 8148
rect 13804 9826 13860 9828
rect 13804 9774 13806 9826
rect 13806 9774 13858 9826
rect 13858 9774 13860 9826
rect 13804 9772 13860 9774
rect 13692 9324 13748 9380
rect 13692 8652 13748 8708
rect 14364 10780 14420 10836
rect 14364 10108 14420 10164
rect 14812 11116 14868 11172
rect 14252 9548 14308 9604
rect 14148 9434 14204 9436
rect 14148 9382 14150 9434
rect 14150 9382 14202 9434
rect 14202 9382 14204 9434
rect 14148 9380 14204 9382
rect 14252 9434 14308 9436
rect 14252 9382 14254 9434
rect 14254 9382 14306 9434
rect 14306 9382 14308 9434
rect 14252 9380 14308 9382
rect 14356 9434 14412 9436
rect 14356 9382 14358 9434
rect 14358 9382 14410 9434
rect 14410 9382 14412 9434
rect 14356 9380 14412 9382
rect 13916 8764 13972 8820
rect 13804 8540 13860 8596
rect 13804 8204 13860 8260
rect 13580 6860 13636 6916
rect 13692 8092 13748 8148
rect 14148 7866 14204 7868
rect 14148 7814 14150 7866
rect 14150 7814 14202 7866
rect 14202 7814 14204 7866
rect 14148 7812 14204 7814
rect 14252 7866 14308 7868
rect 14252 7814 14254 7866
rect 14254 7814 14306 7866
rect 14306 7814 14308 7866
rect 14252 7812 14308 7814
rect 14356 7866 14412 7868
rect 14356 7814 14358 7866
rect 14358 7814 14410 7866
rect 14410 7814 14412 7866
rect 14356 7812 14412 7814
rect 14364 6690 14420 6692
rect 14364 6638 14366 6690
rect 14366 6638 14418 6690
rect 14418 6638 14420 6690
rect 14364 6636 14420 6638
rect 14148 6298 14204 6300
rect 14148 6246 14150 6298
rect 14150 6246 14202 6298
rect 14202 6246 14204 6298
rect 14148 6244 14204 6246
rect 14252 6298 14308 6300
rect 14252 6246 14254 6298
rect 14254 6246 14306 6298
rect 14306 6246 14308 6298
rect 14252 6244 14308 6246
rect 14356 6298 14412 6300
rect 14356 6246 14358 6298
rect 14358 6246 14410 6298
rect 14410 6246 14412 6298
rect 14356 6244 14412 6246
rect 16044 11340 16100 11396
rect 15148 11170 15204 11172
rect 15148 11118 15150 11170
rect 15150 11118 15202 11170
rect 15202 11118 15204 11170
rect 15148 11116 15204 11118
rect 16156 11116 16212 11172
rect 13356 5068 13412 5124
rect 13244 4732 13300 4788
rect 13804 4956 13860 5012
rect 14924 7308 14980 7364
rect 15372 8988 15428 9044
rect 14148 4730 14204 4732
rect 13916 4620 13972 4676
rect 14148 4678 14150 4730
rect 14150 4678 14202 4730
rect 14202 4678 14204 4730
rect 14148 4676 14204 4678
rect 14252 4730 14308 4732
rect 14252 4678 14254 4730
rect 14254 4678 14306 4730
rect 14306 4678 14308 4730
rect 14252 4676 14308 4678
rect 14356 4730 14412 4732
rect 14356 4678 14358 4730
rect 14358 4678 14410 4730
rect 14410 4678 14412 4730
rect 14356 4676 14412 4678
rect 13580 3388 13636 3444
rect 13692 3612 13748 3668
rect 13468 3276 13524 3332
rect 14924 4562 14980 4564
rect 14924 4510 14926 4562
rect 14926 4510 14978 4562
rect 14978 4510 14980 4562
rect 14924 4508 14980 4510
rect 14812 3554 14868 3556
rect 14812 3502 14814 3554
rect 14814 3502 14866 3554
rect 14866 3502 14868 3554
rect 14812 3500 14868 3502
rect 14148 3162 14204 3164
rect 14148 3110 14150 3162
rect 14150 3110 14202 3162
rect 14202 3110 14204 3162
rect 14148 3108 14204 3110
rect 14252 3162 14308 3164
rect 14252 3110 14254 3162
rect 14254 3110 14306 3162
rect 14306 3110 14308 3162
rect 14252 3108 14308 3110
rect 14356 3162 14412 3164
rect 14356 3110 14358 3162
rect 14358 3110 14410 3162
rect 14410 3110 14412 3162
rect 14356 3108 14412 3110
rect 14364 2940 14420 2996
rect 15372 4450 15428 4452
rect 15372 4398 15374 4450
rect 15374 4398 15426 4450
rect 15426 4398 15428 4450
rect 15372 4396 15428 4398
rect 15260 4284 15316 4340
rect 15820 10610 15876 10612
rect 15820 10558 15822 10610
rect 15822 10558 15874 10610
rect 15874 10558 15876 10610
rect 15820 10556 15876 10558
rect 15596 8146 15652 8148
rect 15596 8094 15598 8146
rect 15598 8094 15650 8146
rect 15650 8094 15652 8146
rect 15596 8092 15652 8094
rect 16604 10332 16660 10388
rect 16304 10218 16360 10220
rect 16304 10166 16306 10218
rect 16306 10166 16358 10218
rect 16358 10166 16360 10218
rect 16304 10164 16360 10166
rect 16408 10218 16464 10220
rect 16408 10166 16410 10218
rect 16410 10166 16462 10218
rect 16462 10166 16464 10218
rect 16408 10164 16464 10166
rect 16512 10218 16568 10220
rect 16512 10166 16514 10218
rect 16514 10166 16566 10218
rect 16566 10166 16568 10218
rect 16512 10164 16568 10166
rect 17500 11788 17556 11844
rect 17836 11452 17892 11508
rect 17948 12236 18004 12292
rect 18060 12178 18116 12180
rect 18060 12126 18062 12178
rect 18062 12126 18114 12178
rect 18114 12126 18116 12178
rect 18060 12124 18116 12126
rect 16156 9100 16212 9156
rect 16044 8930 16100 8932
rect 16044 8878 16046 8930
rect 16046 8878 16098 8930
rect 16098 8878 16100 8930
rect 16044 8876 16100 8878
rect 16716 9042 16772 9044
rect 16716 8990 16718 9042
rect 16718 8990 16770 9042
rect 16770 8990 16772 9042
rect 16716 8988 16772 8990
rect 15932 8316 15988 8372
rect 15596 7308 15652 7364
rect 15708 4844 15764 4900
rect 15596 4450 15652 4452
rect 15596 4398 15598 4450
rect 15598 4398 15650 4450
rect 15650 4398 15652 4450
rect 15596 4396 15652 4398
rect 15484 3500 15540 3556
rect 16304 8650 16360 8652
rect 16304 8598 16306 8650
rect 16306 8598 16358 8650
rect 16358 8598 16360 8650
rect 16304 8596 16360 8598
rect 16408 8650 16464 8652
rect 16408 8598 16410 8650
rect 16410 8598 16462 8650
rect 16462 8598 16464 8650
rect 16408 8596 16464 8598
rect 16512 8650 16568 8652
rect 16512 8598 16514 8650
rect 16514 8598 16566 8650
rect 16566 8598 16568 8650
rect 16512 8596 16568 8598
rect 16828 8370 16884 8372
rect 16828 8318 16830 8370
rect 16830 8318 16882 8370
rect 16882 8318 16884 8370
rect 16828 8316 16884 8318
rect 16716 8146 16772 8148
rect 16716 8094 16718 8146
rect 16718 8094 16770 8146
rect 16770 8094 16772 8146
rect 16716 8092 16772 8094
rect 16828 7868 16884 7924
rect 16716 7474 16772 7476
rect 16716 7422 16718 7474
rect 16718 7422 16770 7474
rect 16770 7422 16772 7474
rect 16716 7420 16772 7422
rect 16304 7082 16360 7084
rect 16304 7030 16306 7082
rect 16306 7030 16358 7082
rect 16358 7030 16360 7082
rect 16304 7028 16360 7030
rect 16408 7082 16464 7084
rect 16408 7030 16410 7082
rect 16410 7030 16462 7082
rect 16462 7030 16464 7082
rect 16408 7028 16464 7030
rect 16512 7082 16568 7084
rect 16512 7030 16514 7082
rect 16514 7030 16566 7082
rect 16566 7030 16568 7082
rect 16716 7084 16772 7140
rect 16512 7028 16568 7030
rect 16304 5514 16360 5516
rect 16304 5462 16306 5514
rect 16306 5462 16358 5514
rect 16358 5462 16360 5514
rect 16304 5460 16360 5462
rect 16408 5514 16464 5516
rect 16408 5462 16410 5514
rect 16410 5462 16462 5514
rect 16462 5462 16464 5514
rect 16408 5460 16464 5462
rect 16512 5514 16568 5516
rect 16512 5462 16514 5514
rect 16514 5462 16566 5514
rect 16566 5462 16568 5514
rect 16512 5460 16568 5462
rect 16828 6188 16884 6244
rect 16156 4844 16212 4900
rect 16304 3946 16360 3948
rect 16304 3894 16306 3946
rect 16306 3894 16358 3946
rect 16358 3894 16360 3946
rect 16304 3892 16360 3894
rect 16408 3946 16464 3948
rect 16408 3894 16410 3946
rect 16410 3894 16462 3946
rect 16462 3894 16464 3946
rect 16408 3892 16464 3894
rect 16512 3946 16568 3948
rect 16512 3894 16514 3946
rect 16514 3894 16566 3946
rect 16566 3894 16568 3946
rect 16512 3892 16568 3894
rect 16156 3164 16212 3220
rect 15708 924 15764 980
rect 17948 10668 18004 10724
rect 18460 11002 18516 11004
rect 18460 10950 18462 11002
rect 18462 10950 18514 11002
rect 18514 10950 18516 11002
rect 18460 10948 18516 10950
rect 18564 11002 18620 11004
rect 18564 10950 18566 11002
rect 18566 10950 18618 11002
rect 18618 10950 18620 11002
rect 18564 10948 18620 10950
rect 18668 11002 18724 11004
rect 18668 10950 18670 11002
rect 18670 10950 18722 11002
rect 18722 10950 18724 11002
rect 18668 10948 18724 10950
rect 17052 9548 17108 9604
rect 17612 9042 17668 9044
rect 17612 8990 17614 9042
rect 17614 8990 17666 9042
rect 17666 8990 17668 9042
rect 17612 8988 17668 8990
rect 18172 10498 18228 10500
rect 18172 10446 18174 10498
rect 18174 10446 18226 10498
rect 18226 10446 18228 10498
rect 18172 10444 18228 10446
rect 18844 10444 18900 10500
rect 18460 9434 18516 9436
rect 18460 9382 18462 9434
rect 18462 9382 18514 9434
rect 18514 9382 18516 9434
rect 18460 9380 18516 9382
rect 18564 9434 18620 9436
rect 18564 9382 18566 9434
rect 18566 9382 18618 9434
rect 18618 9382 18620 9434
rect 18564 9380 18620 9382
rect 18668 9434 18724 9436
rect 18668 9382 18670 9434
rect 18670 9382 18722 9434
rect 18722 9382 18724 9434
rect 18668 9380 18724 9382
rect 17276 8146 17332 8148
rect 17276 8094 17278 8146
rect 17278 8094 17330 8146
rect 17330 8094 17332 8146
rect 17276 8092 17332 8094
rect 17724 8092 17780 8148
rect 17612 8034 17668 8036
rect 17612 7982 17614 8034
rect 17614 7982 17666 8034
rect 17666 7982 17668 8034
rect 17612 7980 17668 7982
rect 17052 7532 17108 7588
rect 17612 7756 17668 7812
rect 17500 7586 17556 7588
rect 17500 7534 17502 7586
rect 17502 7534 17554 7586
rect 17554 7534 17556 7586
rect 17500 7532 17556 7534
rect 17948 8146 18004 8148
rect 17948 8094 17950 8146
rect 17950 8094 18002 8146
rect 18002 8094 18004 8146
rect 17948 8092 18004 8094
rect 17836 7250 17892 7252
rect 17836 7198 17838 7250
rect 17838 7198 17890 7250
rect 17890 7198 17892 7250
rect 17836 7196 17892 7198
rect 17276 6860 17332 6916
rect 17836 6972 17892 7028
rect 17612 6636 17668 6692
rect 17612 6300 17668 6356
rect 18172 6860 18228 6916
rect 17948 6412 18004 6468
rect 18460 7866 18516 7868
rect 18460 7814 18462 7866
rect 18462 7814 18514 7866
rect 18514 7814 18516 7866
rect 18460 7812 18516 7814
rect 18564 7866 18620 7868
rect 18564 7814 18566 7866
rect 18566 7814 18618 7866
rect 18618 7814 18620 7866
rect 18564 7812 18620 7814
rect 18668 7866 18724 7868
rect 18668 7814 18670 7866
rect 18670 7814 18722 7866
rect 18722 7814 18724 7866
rect 18668 7812 18724 7814
rect 18172 6188 18228 6244
rect 18460 6298 18516 6300
rect 18460 6246 18462 6298
rect 18462 6246 18514 6298
rect 18514 6246 18516 6298
rect 18460 6244 18516 6246
rect 18564 6298 18620 6300
rect 18564 6246 18566 6298
rect 18566 6246 18618 6298
rect 18618 6246 18620 6298
rect 18564 6244 18620 6246
rect 18668 6298 18724 6300
rect 18668 6246 18670 6298
rect 18670 6246 18722 6298
rect 18722 6246 18724 6298
rect 18668 6244 18724 6246
rect 17948 5906 18004 5908
rect 17948 5854 17950 5906
rect 17950 5854 18002 5906
rect 18002 5854 18004 5906
rect 17948 5852 18004 5854
rect 17948 5122 18004 5124
rect 17948 5070 17950 5122
rect 17950 5070 18002 5122
rect 18002 5070 18004 5122
rect 17948 5068 18004 5070
rect 17612 4338 17668 4340
rect 17612 4286 17614 4338
rect 17614 4286 17666 4338
rect 17666 4286 17668 4338
rect 17612 4284 17668 4286
rect 16940 3442 16996 3444
rect 16940 3390 16942 3442
rect 16942 3390 16994 3442
rect 16994 3390 16996 3442
rect 16940 3388 16996 3390
rect 17164 3276 17220 3332
rect 17500 3388 17556 3444
rect 18172 5852 18228 5908
rect 18460 4730 18516 4732
rect 18460 4678 18462 4730
rect 18462 4678 18514 4730
rect 18514 4678 18516 4730
rect 18460 4676 18516 4678
rect 18564 4730 18620 4732
rect 18564 4678 18566 4730
rect 18566 4678 18618 4730
rect 18618 4678 18620 4730
rect 18564 4676 18620 4678
rect 18668 4730 18724 4732
rect 18668 4678 18670 4730
rect 18670 4678 18722 4730
rect 18722 4678 18724 4730
rect 18668 4676 18724 4678
rect 18956 8092 19012 8148
rect 18956 4060 19012 4116
rect 18844 3836 18900 3892
rect 18460 3162 18516 3164
rect 18460 3110 18462 3162
rect 18462 3110 18514 3162
rect 18514 3110 18516 3162
rect 18460 3108 18516 3110
rect 18564 3162 18620 3164
rect 18564 3110 18566 3162
rect 18566 3110 18618 3162
rect 18618 3110 18620 3162
rect 18564 3108 18620 3110
rect 18668 3162 18724 3164
rect 18668 3110 18670 3162
rect 18670 3110 18722 3162
rect 18722 3110 18724 3162
rect 18668 3108 18724 3110
rect 18956 3388 19012 3444
rect 19404 10332 19460 10388
rect 19292 9884 19348 9940
rect 19292 5852 19348 5908
<< metal3 >>
rect 0 15316 800 15344
rect 0 15260 1708 15316
rect 1764 15260 1774 15316
rect 0 15232 800 15260
rect 0 14868 800 14896
rect 0 14812 4732 14868
rect 4788 14812 4798 14868
rect 0 14784 800 14812
rect 0 14420 800 14448
rect 0 14364 4284 14420
rect 4340 14364 4350 14420
rect 0 14336 800 14364
rect 0 13972 800 14000
rect 0 13916 3500 13972
rect 3556 13916 3566 13972
rect 0 13888 800 13916
rect 0 13524 800 13552
rect 0 13468 2828 13524
rect 2884 13468 2894 13524
rect 0 13440 800 13468
rect 0 13076 800 13104
rect 0 13020 1932 13076
rect 1988 13020 1998 13076
rect 0 12992 800 13020
rect 0 12628 800 12656
rect 0 12572 2604 12628
rect 2660 12572 2670 12628
rect 0 12544 800 12572
rect 5514 12516 5524 12572
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5788 12516 5798 12572
rect 9826 12516 9836 12572
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 10100 12516 10110 12572
rect 14138 12516 14148 12572
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14412 12516 14422 12572
rect 18450 12516 18460 12572
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18724 12516 18734 12572
rect 12338 12348 12348 12404
rect 12404 12348 13580 12404
rect 13636 12348 13646 12404
rect 16370 12348 16380 12404
rect 16436 12348 17276 12404
rect 17332 12348 17342 12404
rect 2146 12236 2156 12292
rect 2212 12236 2222 12292
rect 15810 12236 15820 12292
rect 15876 12236 17948 12292
rect 18004 12236 18014 12292
rect 0 12180 800 12208
rect 2156 12180 2212 12236
rect 0 12124 2212 12180
rect 14914 12124 14924 12180
rect 14980 12124 18060 12180
rect 18116 12124 18126 12180
rect 0 12096 800 12124
rect 1922 12012 1932 12068
rect 1988 12012 5628 12068
rect 5684 12012 5694 12068
rect 18060 11956 18116 12124
rect 19200 11956 20000 11984
rect 1698 11900 1708 11956
rect 1764 11900 1774 11956
rect 15362 11900 15372 11956
rect 15428 11900 16772 11956
rect 18060 11900 20000 11956
rect 0 11732 800 11760
rect 1708 11732 1764 11900
rect 16716 11844 16772 11900
rect 19200 11872 20000 11900
rect 16706 11788 16716 11844
rect 16772 11788 17500 11844
rect 17556 11788 17566 11844
rect 3358 11732 3368 11788
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3632 11732 3642 11788
rect 7670 11732 7680 11788
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 7944 11732 7954 11788
rect 11982 11732 11992 11788
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 12256 11732 12266 11788
rect 16294 11732 16304 11788
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16568 11732 16578 11788
rect 0 11676 1764 11732
rect 13122 11676 13132 11732
rect 13188 11676 14476 11732
rect 14532 11676 14542 11732
rect 0 11648 800 11676
rect 14578 11452 14588 11508
rect 14644 11452 17836 11508
rect 17892 11452 17902 11508
rect 12674 11340 12684 11396
rect 12740 11340 16044 11396
rect 16100 11340 16110 11396
rect 0 11284 800 11312
rect 0 11228 2156 11284
rect 2212 11228 2222 11284
rect 13682 11228 13692 11284
rect 13748 11228 17612 11284
rect 17668 11228 17678 11284
rect 0 11200 800 11228
rect 1698 11116 1708 11172
rect 1764 11116 1774 11172
rect 2146 11116 2156 11172
rect 2212 11116 4956 11172
rect 5012 11116 5022 11172
rect 11638 11116 11676 11172
rect 11732 11116 12124 11172
rect 12180 11116 12190 11172
rect 13010 11116 13020 11172
rect 13076 11116 13356 11172
rect 13412 11116 13422 11172
rect 14130 11116 14140 11172
rect 14196 11116 14644 11172
rect 14802 11116 14812 11172
rect 14868 11116 15148 11172
rect 15204 11116 15214 11172
rect 16118 11116 16156 11172
rect 16212 11116 16222 11172
rect 0 10836 800 10864
rect 1708 10836 1764 11116
rect 5514 10948 5524 11004
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5788 10948 5798 11004
rect 9826 10948 9836 11004
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 10100 10948 10110 11004
rect 14138 10948 14148 11004
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14412 10948 14422 11004
rect 14588 10836 14644 11116
rect 18450 10948 18460 11004
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18724 10948 18734 11004
rect 0 10780 1764 10836
rect 14354 10780 14364 10836
rect 14420 10780 14644 10836
rect 0 10752 800 10780
rect 4162 10668 4172 10724
rect 4228 10668 5852 10724
rect 5908 10668 5918 10724
rect 6962 10668 6972 10724
rect 7028 10668 8988 10724
rect 9044 10668 10220 10724
rect 10276 10668 10668 10724
rect 10724 10668 10734 10724
rect 15092 10668 17948 10724
rect 18004 10668 18014 10724
rect 15092 10612 15148 10668
rect 1362 10556 1372 10612
rect 1428 10556 8204 10612
rect 8260 10556 11788 10612
rect 11844 10556 15148 10612
rect 15810 10556 15820 10612
rect 15876 10556 18228 10612
rect 18172 10500 18228 10556
rect 4386 10444 4396 10500
rect 4452 10444 6300 10500
rect 6356 10444 6366 10500
rect 13010 10444 13020 10500
rect 13076 10444 15148 10500
rect 18162 10444 18172 10500
rect 18228 10444 18844 10500
rect 18900 10444 18910 10500
rect 0 10388 800 10416
rect 15092 10388 15148 10444
rect 0 10332 1708 10388
rect 1764 10332 1774 10388
rect 1922 10332 1932 10388
rect 1988 10332 7756 10388
rect 7812 10332 7822 10388
rect 12908 10332 13132 10388
rect 13188 10332 13198 10388
rect 15092 10332 16604 10388
rect 16660 10332 19404 10388
rect 19460 10332 19470 10388
rect 0 10304 800 10332
rect 4722 10220 4732 10276
rect 4788 10220 7308 10276
rect 7364 10220 7374 10276
rect 11218 10220 11228 10276
rect 11284 10220 11788 10276
rect 11844 10220 11854 10276
rect 3358 10164 3368 10220
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3632 10164 3642 10220
rect 7670 10164 7680 10220
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7944 10164 7954 10220
rect 11982 10164 11992 10220
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 12256 10164 12266 10220
rect 4946 10108 4956 10164
rect 5012 10108 6076 10164
rect 6132 10108 6142 10164
rect 12908 10052 12964 10332
rect 16294 10164 16304 10220
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16568 10164 16578 10220
rect 13122 10108 13132 10164
rect 13188 10108 14364 10164
rect 14420 10108 14430 10164
rect 2482 9996 2492 10052
rect 2548 9996 7532 10052
rect 7588 9996 7598 10052
rect 10210 9996 10220 10052
rect 10276 9996 12124 10052
rect 12180 9996 12964 10052
rect 0 9940 800 9968
rect 12908 9940 12964 9996
rect 0 9884 2604 9940
rect 2660 9884 2670 9940
rect 4620 9884 10668 9940
rect 10724 9884 10734 9940
rect 12908 9884 19292 9940
rect 19348 9884 19358 9940
rect 0 9856 800 9884
rect 4620 9828 4676 9884
rect 3938 9772 3948 9828
rect 4004 9772 4620 9828
rect 4676 9772 4686 9828
rect 11442 9772 11452 9828
rect 11508 9772 13244 9828
rect 13300 9772 13310 9828
rect 13794 9772 13804 9828
rect 13860 9772 13870 9828
rect 1810 9660 1820 9716
rect 1876 9660 2044 9716
rect 2100 9660 2110 9716
rect 10546 9660 10556 9716
rect 10612 9660 11340 9716
rect 11396 9660 11406 9716
rect 12002 9660 12012 9716
rect 12068 9660 12460 9716
rect 12516 9660 12526 9716
rect 13804 9604 13860 9772
rect 2146 9548 2156 9604
rect 2212 9548 2222 9604
rect 3490 9548 3500 9604
rect 3556 9548 3724 9604
rect 3780 9548 3790 9604
rect 3910 9548 3948 9604
rect 4004 9548 4014 9604
rect 5068 9548 6636 9604
rect 6692 9548 6702 9604
rect 6860 9548 12572 9604
rect 12628 9548 12638 9604
rect 12786 9548 12796 9604
rect 12852 9548 13860 9604
rect 13916 9548 14252 9604
rect 14308 9548 17052 9604
rect 17108 9548 17118 9604
rect 0 9492 800 9520
rect 2156 9492 2212 9548
rect 0 9436 2212 9492
rect 0 9408 800 9436
rect 5068 9380 5124 9548
rect 5514 9380 5524 9436
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 5788 9380 5798 9436
rect 6860 9380 6916 9548
rect 13916 9492 13972 9548
rect 11666 9436 11676 9492
rect 11732 9436 11956 9492
rect 12898 9436 12908 9492
rect 12964 9436 13972 9492
rect 9826 9380 9836 9436
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 10100 9380 10110 9436
rect 11900 9380 11956 9436
rect 14138 9380 14148 9436
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14412 9380 14422 9436
rect 18450 9380 18460 9436
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18724 9380 18734 9436
rect 3154 9324 3164 9380
rect 3220 9324 5124 9380
rect 6626 9324 6636 9380
rect 6692 9324 6916 9380
rect 11900 9324 13692 9380
rect 13748 9324 13758 9380
rect 1922 9212 1932 9268
rect 1988 9212 8876 9268
rect 8932 9212 8942 9268
rect 2258 9100 2268 9156
rect 2324 9100 3052 9156
rect 3108 9100 3118 9156
rect 3266 9100 3276 9156
rect 3332 9100 3500 9156
rect 3556 9100 3566 9156
rect 4386 9100 4396 9156
rect 4452 9100 4462 9156
rect 16146 9100 16156 9156
rect 16212 9100 16940 9156
rect 16996 9100 17006 9156
rect 0 9044 800 9072
rect 4396 9044 4452 9100
rect 0 8988 4452 9044
rect 5170 8988 5180 9044
rect 5236 8988 5246 9044
rect 6402 8988 6412 9044
rect 6468 8988 12012 9044
rect 12068 8988 12078 9044
rect 15362 8988 15372 9044
rect 15428 8988 16716 9044
rect 16772 8988 16782 9044
rect 17574 8988 17612 9044
rect 17668 8988 17678 9044
rect 0 8960 800 8988
rect 5180 8932 5236 8988
rect 2370 8876 2380 8932
rect 2436 8876 5236 8932
rect 10546 8876 10556 8932
rect 10612 8876 16044 8932
rect 16100 8876 16110 8932
rect 1810 8764 1820 8820
rect 1876 8764 2828 8820
rect 2884 8764 2894 8820
rect 3154 8764 3164 8820
rect 3220 8764 3276 8820
rect 3332 8764 3342 8820
rect 4274 8764 4284 8820
rect 4340 8764 7980 8820
rect 8036 8764 8046 8820
rect 8978 8764 8988 8820
rect 9044 8764 13916 8820
rect 13972 8764 13982 8820
rect 4050 8652 4060 8708
rect 4116 8652 7532 8708
rect 7588 8652 7598 8708
rect 13654 8652 13692 8708
rect 13748 8652 13758 8708
rect 0 8596 800 8624
rect 3358 8596 3368 8652
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3632 8596 3642 8652
rect 7670 8596 7680 8652
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7944 8596 7954 8652
rect 11982 8596 11992 8652
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 12256 8596 12266 8652
rect 16294 8596 16304 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16568 8596 16578 8652
rect 0 8540 2156 8596
rect 2212 8540 2222 8596
rect 4498 8540 4508 8596
rect 4564 8540 7196 8596
rect 7252 8540 7262 8596
rect 13794 8540 13804 8596
rect 13860 8540 13870 8596
rect 0 8512 800 8540
rect 2818 8428 2828 8484
rect 2884 8428 4116 8484
rect 4386 8428 4396 8484
rect 4452 8428 5292 8484
rect 5348 8428 5358 8484
rect 11106 8428 11116 8484
rect 11172 8428 11788 8484
rect 11844 8428 11854 8484
rect 4060 8372 4116 8428
rect 1250 8316 1260 8372
rect 1316 8316 3164 8372
rect 3220 8316 3230 8372
rect 3602 8316 3612 8372
rect 3668 8316 3836 8372
rect 3892 8316 3902 8372
rect 4060 8316 8428 8372
rect 8484 8316 8494 8372
rect 13458 8316 13468 8372
rect 13524 8316 13534 8372
rect 13468 8260 13524 8316
rect 13804 8260 13860 8540
rect 15922 8316 15932 8372
rect 15988 8316 16828 8372
rect 16884 8316 16894 8372
rect 1708 8204 4284 8260
rect 4340 8204 4350 8260
rect 5954 8204 5964 8260
rect 6020 8204 6076 8260
rect 6132 8204 6142 8260
rect 10220 8204 13524 8260
rect 13794 8204 13804 8260
rect 13860 8204 13870 8260
rect 0 8148 800 8176
rect 1708 8148 1764 8204
rect 0 8092 1764 8148
rect 2118 8092 2156 8148
rect 2212 8092 2222 8148
rect 2706 8092 2716 8148
rect 2772 8092 4620 8148
rect 4676 8092 4686 8148
rect 6066 8092 6076 8148
rect 6132 8092 6860 8148
rect 6916 8092 7868 8148
rect 7924 8092 7934 8148
rect 0 8064 800 8092
rect 2034 7980 2044 8036
rect 2100 7980 4060 8036
rect 4116 7980 4126 8036
rect 4274 7980 4284 8036
rect 4340 7980 6412 8036
rect 6468 7980 6478 8036
rect 7186 7980 7196 8036
rect 7252 7980 7644 8036
rect 7700 7980 7710 8036
rect 3266 7868 3276 7924
rect 3332 7868 5068 7924
rect 5124 7868 5134 7924
rect 5514 7812 5524 7868
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5788 7812 5798 7868
rect 9826 7812 9836 7868
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 10100 7812 10110 7868
rect 1474 7756 1484 7812
rect 1540 7756 5348 7812
rect 5954 7756 5964 7812
rect 6020 7756 7868 7812
rect 7924 7756 7934 7812
rect 0 7700 800 7728
rect 5292 7700 5348 7756
rect 10220 7700 10276 8204
rect 10882 8092 10892 8148
rect 10948 8092 13468 8148
rect 13524 8092 13534 8148
rect 13682 8092 13692 8148
rect 13748 8092 15596 8148
rect 15652 8092 15662 8148
rect 16706 8092 16716 8148
rect 16772 8092 16782 8148
rect 17266 8092 17276 8148
rect 17332 8092 17724 8148
rect 17780 8092 17790 8148
rect 17938 8092 17948 8148
rect 18004 8092 18956 8148
rect 19012 8092 19022 8148
rect 16716 8036 16772 8092
rect 11218 7980 11228 8036
rect 11284 7980 16772 8036
rect 17602 7980 17612 8036
rect 17668 7980 17678 8036
rect 17612 7924 17668 7980
rect 16818 7868 16828 7924
rect 16884 7868 17668 7924
rect 14138 7812 14148 7868
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14412 7812 14422 7868
rect 18450 7812 18460 7868
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18724 7812 18734 7868
rect 16930 7756 16940 7812
rect 16996 7756 17612 7812
rect 17668 7756 17678 7812
rect 0 7644 3724 7700
rect 3780 7644 3790 7700
rect 4050 7644 4060 7700
rect 4116 7644 5236 7700
rect 5292 7644 10276 7700
rect 0 7616 800 7644
rect 5180 7588 5236 7644
rect 1250 7532 1260 7588
rect 1316 7532 1708 7588
rect 1764 7532 1774 7588
rect 3490 7532 3500 7588
rect 3556 7532 3566 7588
rect 3826 7532 3836 7588
rect 3892 7532 4956 7588
rect 5012 7532 5022 7588
rect 5180 7532 6636 7588
rect 6692 7532 6702 7588
rect 8530 7532 8540 7588
rect 8596 7532 11452 7588
rect 11508 7532 11518 7588
rect 17042 7532 17052 7588
rect 17108 7532 17500 7588
rect 17556 7532 17566 7588
rect 3500 7476 3556 7532
rect 2454 7420 2492 7476
rect 2548 7420 2558 7476
rect 2706 7420 2716 7476
rect 2772 7420 3556 7476
rect 3714 7420 3724 7476
rect 3780 7420 4060 7476
rect 4116 7420 4126 7476
rect 4498 7420 4508 7476
rect 4564 7420 5964 7476
rect 6020 7420 6030 7476
rect 7074 7420 7084 7476
rect 7140 7420 7532 7476
rect 7588 7420 8092 7476
rect 8148 7420 8158 7476
rect 9426 7420 9436 7476
rect 9492 7420 9660 7476
rect 9716 7420 9726 7476
rect 12674 7420 12684 7476
rect 12740 7420 16716 7476
rect 16772 7420 16782 7476
rect 2930 7308 2940 7364
rect 2996 7308 4228 7364
rect 10434 7308 10444 7364
rect 10500 7308 11228 7364
rect 11284 7308 11294 7364
rect 14914 7308 14924 7364
rect 14980 7308 15596 7364
rect 15652 7308 15662 7364
rect 0 7252 800 7280
rect 4172 7252 4228 7308
rect 0 7196 3948 7252
rect 4004 7196 4014 7252
rect 4172 7196 6300 7252
rect 6356 7196 6366 7252
rect 12562 7196 12572 7252
rect 12628 7196 17836 7252
rect 17892 7196 17902 7252
rect 0 7168 800 7196
rect 5030 7084 5068 7140
rect 5124 7084 5134 7140
rect 16706 7084 16716 7140
rect 16772 7084 17892 7140
rect 3358 7028 3368 7084
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3632 7028 3642 7084
rect 7670 7028 7680 7084
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7944 7028 7954 7084
rect 11982 7028 11992 7084
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 12256 7028 12266 7084
rect 16294 7028 16304 7084
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16568 7028 16578 7084
rect 17836 7028 17892 7084
rect 3938 6972 3948 7028
rect 4004 6972 4620 7028
rect 4676 6972 4686 7028
rect 5170 6972 5180 7028
rect 5236 6972 6524 7028
rect 6580 6972 6590 7028
rect 6850 6972 6860 7028
rect 6916 6972 7196 7028
rect 7252 6972 7262 7028
rect 17826 6972 17836 7028
rect 17892 6972 17902 7028
rect 2146 6860 2156 6916
rect 2212 6860 3556 6916
rect 4162 6860 4172 6916
rect 4228 6860 6804 6916
rect 10322 6860 10332 6916
rect 10388 6860 10668 6916
rect 10724 6860 10734 6916
rect 12898 6860 12908 6916
rect 12964 6860 13580 6916
rect 13636 6860 17276 6916
rect 17332 6860 17342 6916
rect 18162 6860 18172 6916
rect 18228 6860 18238 6916
rect 0 6804 800 6832
rect 3500 6804 3556 6860
rect 6748 6804 6804 6860
rect 0 6748 2940 6804
rect 2996 6748 3006 6804
rect 3500 6748 6468 6804
rect 6738 6748 6748 6804
rect 6804 6748 7196 6804
rect 7252 6748 7262 6804
rect 0 6720 800 6748
rect 6412 6692 6468 6748
rect 1586 6636 1596 6692
rect 1652 6636 1662 6692
rect 1810 6636 1820 6692
rect 1876 6636 1914 6692
rect 2034 6636 2044 6692
rect 2100 6636 2492 6692
rect 2548 6636 2828 6692
rect 2884 6636 2894 6692
rect 5842 6636 5852 6692
rect 5908 6636 6188 6692
rect 6244 6636 6254 6692
rect 6402 6636 6412 6692
rect 6468 6636 6478 6692
rect 8642 6636 8652 6692
rect 8708 6636 10332 6692
rect 10388 6636 10398 6692
rect 14354 6636 14364 6692
rect 14420 6636 17612 6692
rect 17668 6636 17678 6692
rect 0 6356 800 6384
rect 1596 6356 1652 6636
rect 3042 6524 3052 6580
rect 3108 6524 3118 6580
rect 6514 6524 6524 6580
rect 6580 6524 7084 6580
rect 7140 6524 7150 6580
rect 7410 6524 7420 6580
rect 7476 6524 10108 6580
rect 10164 6524 10174 6580
rect 3052 6468 3108 6524
rect 2930 6412 2940 6468
rect 2996 6412 3108 6468
rect 3266 6412 3276 6468
rect 3332 6412 4284 6468
rect 4340 6412 4350 6468
rect 5926 6412 5964 6468
rect 6020 6412 6030 6468
rect 12786 6412 12796 6468
rect 12852 6412 13692 6468
rect 13748 6412 17948 6468
rect 18004 6412 18014 6468
rect 18172 6356 18228 6860
rect 0 6300 1652 6356
rect 17602 6300 17612 6356
rect 17668 6300 18228 6356
rect 0 6272 800 6300
rect 5514 6244 5524 6300
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5788 6244 5798 6300
rect 9826 6244 9836 6300
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 10100 6244 10110 6300
rect 14138 6244 14148 6300
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14412 6244 14422 6300
rect 18450 6244 18460 6300
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18724 6244 18734 6300
rect 1596 6188 3164 6244
rect 3220 6188 3230 6244
rect 3826 6188 3836 6244
rect 3892 6188 4060 6244
rect 4116 6188 4126 6244
rect 4274 6188 4284 6244
rect 4340 6188 4732 6244
rect 4788 6188 4798 6244
rect 6514 6188 6524 6244
rect 6580 6188 7756 6244
rect 7812 6188 7822 6244
rect 16818 6188 16828 6244
rect 16884 6188 18172 6244
rect 18228 6188 18238 6244
rect 0 5908 800 5936
rect 1596 5908 1652 6188
rect 2818 6076 2828 6132
rect 2884 6076 4508 6132
rect 4564 6076 4574 6132
rect 4732 6076 7868 6132
rect 7924 6076 7934 6132
rect 4732 6020 4788 6076
rect 2146 5964 2156 6020
rect 2212 5964 4004 6020
rect 4162 5964 4172 6020
rect 4228 5964 4788 6020
rect 4946 5964 4956 6020
rect 5012 5964 8316 6020
rect 8372 5964 8382 6020
rect 9314 5964 9324 6020
rect 9380 5964 9884 6020
rect 9940 5964 9950 6020
rect 10994 5964 11004 6020
rect 11060 5964 12460 6020
rect 12516 5964 12526 6020
rect 3948 5908 4004 5964
rect 0 5852 1652 5908
rect 2594 5852 2604 5908
rect 2660 5852 3388 5908
rect 3948 5852 4284 5908
rect 4340 5852 4350 5908
rect 4498 5852 4508 5908
rect 4564 5852 5180 5908
rect 5236 5852 5246 5908
rect 5954 5852 5964 5908
rect 6020 5852 10108 5908
rect 10164 5852 10174 5908
rect 17938 5852 17948 5908
rect 18004 5852 18172 5908
rect 18228 5852 19292 5908
rect 19348 5852 19358 5908
rect 0 5824 800 5852
rect 3332 5796 3388 5852
rect 3332 5740 4732 5796
rect 4788 5740 4798 5796
rect 4946 5740 4956 5796
rect 5012 5740 6524 5796
rect 6580 5740 6590 5796
rect 7308 5740 8652 5796
rect 8708 5740 8718 5796
rect 7308 5684 7364 5740
rect 3042 5628 3052 5684
rect 3108 5628 3276 5684
rect 3332 5628 3342 5684
rect 4498 5628 4508 5684
rect 4564 5628 5068 5684
rect 5124 5628 7364 5684
rect 8652 5684 8708 5740
rect 8652 5628 9548 5684
rect 9604 5628 9614 5684
rect 3724 5516 4508 5572
rect 4564 5516 4574 5572
rect 0 5460 800 5488
rect 3358 5460 3368 5516
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3632 5460 3642 5516
rect 3724 5460 3780 5516
rect 7670 5460 7680 5516
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7944 5460 7954 5516
rect 11982 5460 11992 5516
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 12256 5460 12266 5516
rect 16294 5460 16304 5516
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16568 5460 16578 5516
rect 0 5404 2716 5460
rect 2772 5404 2782 5460
rect 3714 5404 3724 5460
rect 3780 5404 3790 5460
rect 4050 5404 4060 5460
rect 4116 5404 6300 5460
rect 6356 5404 6366 5460
rect 0 5376 800 5404
rect 2818 5292 2828 5348
rect 2884 5292 3612 5348
rect 3668 5292 3678 5348
rect 4050 5292 4060 5348
rect 4116 5292 4172 5348
rect 4228 5292 4238 5348
rect 4722 5292 4732 5348
rect 4788 5292 7308 5348
rect 7364 5292 8876 5348
rect 8932 5292 8942 5348
rect 10098 5292 10108 5348
rect 10164 5292 10668 5348
rect 10724 5292 10734 5348
rect 2146 5180 2156 5236
rect 2212 5180 3108 5236
rect 3378 5180 3388 5236
rect 3444 5180 5852 5236
rect 5908 5180 5918 5236
rect 6626 5180 6636 5236
rect 6692 5180 12796 5236
rect 12852 5180 12862 5236
rect 3052 5124 3108 5180
rect 1810 5068 1820 5124
rect 1876 5068 1932 5124
rect 1988 5068 1998 5124
rect 2818 5068 2828 5124
rect 2884 5068 2996 5124
rect 3052 5068 3948 5124
rect 4004 5068 4014 5124
rect 5058 5068 5068 5124
rect 5124 5068 9100 5124
rect 9156 5068 9166 5124
rect 10210 5068 10220 5124
rect 10276 5068 10286 5124
rect 10770 5068 10780 5124
rect 10836 5068 11340 5124
rect 11396 5068 11406 5124
rect 13346 5068 13356 5124
rect 13412 5068 14588 5124
rect 14644 5068 17948 5124
rect 18004 5068 18014 5124
rect 0 5012 800 5040
rect 0 4956 2492 5012
rect 2548 4956 2558 5012
rect 0 4928 800 4956
rect 2940 4900 2996 5068
rect 10220 5012 10276 5068
rect 3490 4956 3500 5012
rect 3556 4956 4508 5012
rect 4564 4956 4574 5012
rect 8418 4956 8428 5012
rect 8484 4956 8988 5012
rect 9044 4956 9054 5012
rect 9660 4956 9996 5012
rect 10052 4956 10062 5012
rect 10220 4956 13804 5012
rect 13860 4956 13870 5012
rect 9660 4900 9716 4956
rect 2940 4844 3388 4900
rect 4694 4844 4732 4900
rect 4788 4844 4798 4900
rect 5170 4844 5180 4900
rect 5236 4844 9660 4900
rect 9716 4844 9726 4900
rect 9874 4844 9884 4900
rect 9940 4844 11452 4900
rect 11508 4844 11518 4900
rect 15698 4844 15708 4900
rect 15764 4844 16156 4900
rect 16212 4844 16222 4900
rect 3332 4788 3388 4844
rect 3332 4732 5068 4788
rect 5124 4732 5134 4788
rect 5954 4732 5964 4788
rect 6020 4732 6076 4788
rect 6132 4732 6142 4788
rect 10210 4732 10220 4788
rect 10276 4732 11060 4788
rect 11554 4732 11564 4788
rect 11620 4732 13244 4788
rect 13300 4732 13310 4788
rect 5514 4676 5524 4732
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5788 4676 5798 4732
rect 9826 4676 9836 4732
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10100 4676 10110 4732
rect 11004 4676 11060 4732
rect 14138 4676 14148 4732
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14412 4676 14422 4732
rect 18450 4676 18460 4732
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18724 4676 18734 4732
rect 1260 4620 2268 4676
rect 2324 4620 2334 4676
rect 3826 4620 3836 4676
rect 3892 4620 3902 4676
rect 10742 4620 10780 4676
rect 10836 4620 10846 4676
rect 11004 4620 13916 4676
rect 13972 4620 13982 4676
rect 0 4564 800 4592
rect 1260 4564 1316 4620
rect 3836 4564 3892 4620
rect 0 4508 1316 4564
rect 1474 4508 1484 4564
rect 1540 4508 2940 4564
rect 2996 4508 3006 4564
rect 3836 4508 6468 4564
rect 6626 4508 6636 4564
rect 6692 4508 9660 4564
rect 9716 4508 9726 4564
rect 11218 4508 11228 4564
rect 11284 4508 11294 4564
rect 14914 4508 14924 4564
rect 14980 4508 15652 4564
rect 0 4480 800 4508
rect 6412 4452 6468 4508
rect 11228 4452 11284 4508
rect 15596 4452 15652 4508
rect 1922 4396 1932 4452
rect 1988 4396 3500 4452
rect 3556 4396 3566 4452
rect 5058 4396 5068 4452
rect 5124 4396 5964 4452
rect 6020 4396 6030 4452
rect 6412 4396 9772 4452
rect 9828 4396 9838 4452
rect 10770 4396 10780 4452
rect 10836 4396 15372 4452
rect 15428 4396 15438 4452
rect 15586 4396 15596 4452
rect 15652 4396 15662 4452
rect 3154 4284 3164 4340
rect 3220 4284 3230 4340
rect 8306 4284 8316 4340
rect 8372 4284 11564 4340
rect 11620 4284 11630 4340
rect 13010 4284 13020 4340
rect 13076 4284 15260 4340
rect 15316 4284 17612 4340
rect 17668 4284 17678 4340
rect 0 4116 800 4144
rect 3164 4116 3220 4284
rect 8978 4172 8988 4228
rect 9044 4172 10780 4228
rect 10836 4172 10846 4228
rect 0 4060 3220 4116
rect 4946 4060 4956 4116
rect 5012 4060 12348 4116
rect 12404 4060 12414 4116
rect 13692 4060 18956 4116
rect 19012 4060 19022 4116
rect 0 4032 800 4060
rect 1782 3948 1820 4004
rect 1876 3948 1886 4004
rect 3014 3948 3052 4004
rect 3108 3948 3118 4004
rect 5058 3948 5068 4004
rect 5124 3948 7532 4004
rect 7588 3948 7598 4004
rect 8530 3948 8540 4004
rect 8596 3948 10780 4004
rect 10836 3948 11788 4004
rect 11844 3948 11854 4004
rect 3358 3892 3368 3948
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3632 3892 3642 3948
rect 7670 3892 7680 3948
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7944 3892 7954 3948
rect 11982 3892 11992 3948
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 12256 3892 12266 3948
rect 1922 3836 1932 3892
rect 1988 3836 2716 3892
rect 2772 3836 2782 3892
rect 10658 3836 10668 3892
rect 10724 3836 10780 3892
rect 10836 3836 10846 3892
rect 1922 3724 1932 3780
rect 1988 3724 10500 3780
rect 10658 3724 10668 3780
rect 10724 3724 12236 3780
rect 12292 3724 12302 3780
rect 0 3668 800 3696
rect 10444 3668 10500 3724
rect 13692 3668 13748 4060
rect 16294 3892 16304 3948
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16568 3892 16578 3948
rect 19200 3892 20000 3920
rect 18834 3836 18844 3892
rect 18900 3836 20000 3892
rect 19200 3808 20000 3836
rect 0 3612 2380 3668
rect 2436 3612 2446 3668
rect 4060 3612 8036 3668
rect 8194 3612 8204 3668
rect 8260 3612 9324 3668
rect 9380 3612 9390 3668
rect 10444 3612 13692 3668
rect 13748 3612 13758 3668
rect 0 3584 800 3612
rect 4060 3556 4116 3612
rect 7980 3556 8036 3612
rect 1362 3500 1372 3556
rect 1428 3500 2828 3556
rect 2884 3500 2894 3556
rect 4050 3500 4060 3556
rect 4116 3500 4126 3556
rect 6486 3500 6524 3556
rect 6580 3500 6590 3556
rect 6738 3500 6748 3556
rect 6804 3500 7532 3556
rect 7588 3500 7598 3556
rect 7980 3500 8428 3556
rect 8484 3500 8494 3556
rect 8754 3500 8764 3556
rect 8820 3500 11340 3556
rect 11396 3500 11406 3556
rect 11778 3500 11788 3556
rect 11844 3500 12572 3556
rect 12628 3500 12638 3556
rect 14802 3500 14812 3556
rect 14868 3500 15484 3556
rect 15540 3500 15550 3556
rect 7532 3444 7588 3500
rect 4582 3388 4620 3444
rect 4676 3388 4686 3444
rect 5842 3388 5852 3444
rect 5908 3388 6412 3444
rect 6468 3388 6478 3444
rect 7186 3388 7196 3444
rect 7252 3388 7308 3444
rect 7364 3388 7374 3444
rect 7532 3388 10220 3444
rect 10276 3388 10286 3444
rect 13570 3388 13580 3444
rect 13636 3388 16940 3444
rect 16996 3388 17006 3444
rect 17490 3388 17500 3444
rect 17556 3388 18956 3444
rect 19012 3388 19022 3444
rect 2482 3276 2492 3332
rect 2548 3276 4060 3332
rect 4116 3276 4126 3332
rect 5954 3276 5964 3332
rect 6020 3276 13468 3332
rect 13524 3276 13534 3332
rect 13916 3276 17164 3332
rect 17220 3276 17230 3332
rect 0 3220 800 3248
rect 13916 3220 13972 3276
rect 0 3164 2604 3220
rect 2660 3164 2670 3220
rect 11778 3164 11788 3220
rect 11844 3164 12572 3220
rect 12628 3164 13972 3220
rect 16118 3164 16156 3220
rect 16212 3164 16222 3220
rect 0 3136 800 3164
rect 5514 3108 5524 3164
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5788 3108 5798 3164
rect 9826 3108 9836 3164
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 10100 3108 10110 3164
rect 14138 3108 14148 3164
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14412 3108 14422 3164
rect 18450 3108 18460 3164
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18724 3108 18734 3164
rect 2146 2940 2156 2996
rect 2212 2940 8540 2996
rect 8596 2940 8606 2996
rect 14354 2940 14364 2996
rect 14420 2940 14588 2996
rect 14644 2940 14654 2996
rect 5058 2828 5068 2884
rect 5124 2828 9884 2884
rect 9940 2828 9950 2884
rect 0 2772 800 2800
rect 0 2716 1708 2772
rect 1764 2716 1774 2772
rect 2902 2716 2940 2772
rect 2996 2716 3006 2772
rect 4498 2716 4508 2772
rect 4564 2716 7196 2772
rect 7252 2716 7262 2772
rect 0 2688 800 2716
rect 5170 2604 5180 2660
rect 5236 2604 7644 2660
rect 7700 2604 7710 2660
rect 0 2324 800 2352
rect 0 2268 3836 2324
rect 3892 2268 3902 2324
rect 0 2240 800 2268
rect 0 1876 800 1904
rect 0 1820 2044 1876
rect 2100 1820 2110 1876
rect 0 1792 800 1820
rect 2146 1484 2156 1540
rect 2212 1484 2222 1540
rect 0 1428 800 1456
rect 2156 1428 2212 1484
rect 0 1372 2212 1428
rect 0 1344 800 1372
rect 9398 1036 9436 1092
rect 9492 1036 9502 1092
rect 0 980 800 1008
rect 0 924 4060 980
rect 4116 924 4126 980
rect 15698 924 15708 980
rect 15764 924 17612 980
rect 17668 924 17678 980
rect 0 896 800 924
rect 0 532 800 560
rect 3332 532 3388 868
rect 3444 812 3454 868
rect 0 476 3388 532
rect 0 448 800 476
<< via3 >>
rect 5524 12516 5580 12572
rect 5628 12516 5684 12572
rect 5732 12516 5788 12572
rect 9836 12516 9892 12572
rect 9940 12516 9996 12572
rect 10044 12516 10100 12572
rect 14148 12516 14204 12572
rect 14252 12516 14308 12572
rect 14356 12516 14412 12572
rect 18460 12516 18516 12572
rect 18564 12516 18620 12572
rect 18668 12516 18724 12572
rect 3368 11732 3424 11788
rect 3472 11732 3528 11788
rect 3576 11732 3632 11788
rect 7680 11732 7736 11788
rect 7784 11732 7840 11788
rect 7888 11732 7944 11788
rect 11992 11732 12048 11788
rect 12096 11732 12152 11788
rect 12200 11732 12256 11788
rect 16304 11732 16360 11788
rect 16408 11732 16464 11788
rect 16512 11732 16568 11788
rect 17612 11228 17668 11284
rect 2156 11116 2212 11172
rect 11676 11116 11732 11172
rect 16156 11116 16212 11172
rect 5524 10948 5580 11004
rect 5628 10948 5684 11004
rect 5732 10948 5788 11004
rect 9836 10948 9892 11004
rect 9940 10948 9996 11004
rect 10044 10948 10100 11004
rect 14148 10948 14204 11004
rect 14252 10948 14308 11004
rect 14356 10948 14412 11004
rect 18460 10948 18516 11004
rect 18564 10948 18620 11004
rect 18668 10948 18724 11004
rect 4172 10668 4228 10724
rect 4396 10444 4452 10500
rect 4732 10220 4788 10276
rect 11788 10220 11844 10276
rect 3368 10164 3424 10220
rect 3472 10164 3528 10220
rect 3576 10164 3632 10220
rect 7680 10164 7736 10220
rect 7784 10164 7840 10220
rect 7888 10164 7944 10220
rect 11992 10164 12048 10220
rect 12096 10164 12152 10220
rect 12200 10164 12256 10220
rect 16304 10164 16360 10220
rect 16408 10164 16464 10220
rect 16512 10164 16568 10220
rect 2492 9996 2548 10052
rect 4620 9772 4676 9828
rect 1820 9660 1876 9716
rect 3724 9548 3780 9604
rect 3948 9548 4004 9604
rect 5524 9380 5580 9436
rect 5628 9380 5684 9436
rect 5732 9380 5788 9436
rect 11676 9436 11732 9492
rect 9836 9380 9892 9436
rect 9940 9380 9996 9436
rect 10044 9380 10100 9436
rect 14148 9380 14204 9436
rect 14252 9380 14308 9436
rect 14356 9380 14412 9436
rect 18460 9380 18516 9436
rect 18564 9380 18620 9436
rect 18668 9380 18724 9436
rect 1932 9212 1988 9268
rect 16940 9100 16996 9156
rect 6412 8988 6468 9044
rect 17612 8988 17668 9044
rect 3164 8764 3220 8820
rect 4284 8764 4340 8820
rect 4060 8652 4116 8708
rect 13692 8652 13748 8708
rect 3368 8596 3424 8652
rect 3472 8596 3528 8652
rect 3576 8596 3632 8652
rect 7680 8596 7736 8652
rect 7784 8596 7840 8652
rect 7888 8596 7944 8652
rect 11992 8596 12048 8652
rect 12096 8596 12152 8652
rect 12200 8596 12256 8652
rect 16304 8596 16360 8652
rect 16408 8596 16464 8652
rect 16512 8596 16568 8652
rect 4508 8540 4564 8596
rect 3836 8316 3892 8372
rect 6076 8204 6132 8260
rect 2156 8092 2212 8148
rect 7196 7980 7252 8036
rect 5524 7812 5580 7868
rect 5628 7812 5684 7868
rect 5732 7812 5788 7868
rect 9836 7812 9892 7868
rect 9940 7812 9996 7868
rect 10044 7812 10100 7868
rect 5964 7756 6020 7812
rect 14148 7812 14204 7868
rect 14252 7812 14308 7868
rect 14356 7812 14412 7868
rect 18460 7812 18516 7868
rect 18564 7812 18620 7868
rect 18668 7812 18724 7868
rect 16940 7756 16996 7812
rect 3836 7532 3892 7588
rect 4956 7532 5012 7588
rect 2492 7420 2548 7476
rect 5964 7420 6020 7476
rect 7532 7420 7588 7476
rect 9436 7420 9492 7476
rect 2940 7308 2996 7364
rect 5068 7084 5124 7140
rect 3368 7028 3424 7084
rect 3472 7028 3528 7084
rect 3576 7028 3632 7084
rect 7680 7028 7736 7084
rect 7784 7028 7840 7084
rect 7888 7028 7944 7084
rect 11992 7028 12048 7084
rect 12096 7028 12152 7084
rect 12200 7028 12256 7084
rect 16304 7028 16360 7084
rect 16408 7028 16464 7084
rect 16512 7028 16568 7084
rect 5180 6972 5236 7028
rect 2940 6748 2996 6804
rect 1820 6636 1876 6692
rect 6412 6636 6468 6692
rect 2940 6412 2996 6468
rect 4284 6412 4340 6468
rect 5964 6412 6020 6468
rect 13692 6412 13748 6468
rect 5524 6244 5580 6300
rect 5628 6244 5684 6300
rect 5732 6244 5788 6300
rect 9836 6244 9892 6300
rect 9940 6244 9996 6300
rect 10044 6244 10100 6300
rect 14148 6244 14204 6300
rect 14252 6244 14308 6300
rect 14356 6244 14412 6300
rect 18460 6244 18516 6300
rect 18564 6244 18620 6300
rect 18668 6244 18724 6300
rect 4060 6188 4116 6244
rect 6524 6188 6580 6244
rect 5180 5852 5236 5908
rect 4732 5740 4788 5796
rect 3052 5628 3108 5684
rect 4508 5516 4564 5572
rect 3368 5460 3424 5516
rect 3472 5460 3528 5516
rect 3576 5460 3632 5516
rect 7680 5460 7736 5516
rect 7784 5460 7840 5516
rect 7888 5460 7944 5516
rect 11992 5460 12048 5516
rect 12096 5460 12152 5516
rect 12200 5460 12256 5516
rect 16304 5460 16360 5516
rect 16408 5460 16464 5516
rect 16512 5460 16568 5516
rect 4060 5404 4116 5460
rect 4172 5292 4228 5348
rect 10668 5292 10724 5348
rect 1932 5068 1988 5124
rect 14588 5068 14644 5124
rect 4508 4956 4564 5012
rect 4732 4844 4788 4900
rect 6076 4732 6132 4788
rect 5524 4676 5580 4732
rect 5628 4676 5684 4732
rect 5732 4676 5788 4732
rect 9836 4676 9892 4732
rect 9940 4676 9996 4732
rect 10044 4676 10100 4732
rect 14148 4676 14204 4732
rect 14252 4676 14308 4732
rect 14356 4676 14412 4732
rect 18460 4676 18516 4732
rect 18564 4676 18620 4732
rect 18668 4676 18724 4732
rect 10780 4620 10836 4676
rect 3164 4284 3220 4340
rect 4956 4060 5012 4116
rect 1820 3948 1876 4004
rect 3052 3948 3108 4004
rect 7532 3948 7588 4004
rect 10780 3948 10836 4004
rect 3368 3892 3424 3948
rect 3472 3892 3528 3948
rect 3576 3892 3632 3948
rect 7680 3892 7736 3948
rect 7784 3892 7840 3948
rect 7888 3892 7944 3948
rect 11992 3892 12048 3948
rect 12096 3892 12152 3948
rect 12200 3892 12256 3948
rect 1932 3836 1988 3892
rect 10668 3836 10724 3892
rect 16304 3892 16360 3948
rect 16408 3892 16464 3948
rect 16512 3892 16568 3948
rect 6524 3500 6580 3556
rect 4620 3388 4676 3444
rect 6412 3388 6468 3444
rect 7196 3388 7252 3444
rect 2492 3276 2548 3332
rect 5964 3276 6020 3332
rect 11788 3164 11844 3220
rect 16156 3164 16212 3220
rect 5524 3108 5580 3164
rect 5628 3108 5684 3164
rect 5732 3108 5788 3164
rect 9836 3108 9892 3164
rect 9940 3108 9996 3164
rect 10044 3108 10100 3164
rect 14148 3108 14204 3164
rect 14252 3108 14308 3164
rect 14356 3108 14412 3164
rect 18460 3108 18516 3164
rect 18564 3108 18620 3164
rect 18668 3108 18724 3164
rect 2156 2940 2212 2996
rect 14588 2940 14644 2996
rect 5068 2828 5124 2884
rect 2940 2716 2996 2772
rect 4508 2716 4564 2772
rect 5180 2604 5236 2660
rect 3836 2268 3892 2324
rect 9436 1036 9492 1092
rect 4060 924 4116 980
rect 17612 924 17668 980
<< metal4 >>
rect 3340 11788 3660 12604
rect 3340 11732 3368 11788
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3632 11732 3660 11788
rect 2156 11172 2212 11182
rect 1820 9716 1876 9726
rect 1820 6692 1876 9660
rect 1820 4004 1876 6636
rect 1820 3938 1876 3948
rect 1932 9268 1988 9278
rect 1932 5124 1988 9212
rect 1932 3892 1988 5068
rect 1932 3826 1988 3836
rect 2156 8148 2212 11116
rect 3340 10220 3660 11732
rect 5496 12572 5816 12604
rect 5496 12516 5524 12572
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5788 12516 5816 12572
rect 5496 11004 5816 12516
rect 5496 10948 5524 11004
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5788 10948 5816 11004
rect 3340 10164 3368 10220
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3632 10164 3660 10220
rect 2156 2996 2212 8092
rect 2492 10052 2548 10062
rect 2492 7476 2548 9996
rect 2492 3332 2548 7420
rect 3164 8820 3220 8830
rect 2940 7364 2996 7374
rect 2940 6804 2996 7308
rect 2940 6738 2996 6748
rect 2492 3266 2548 3276
rect 2940 6468 2996 6478
rect 2156 2930 2212 2940
rect 2940 2772 2996 6412
rect 3052 5684 3108 5694
rect 3052 4004 3108 5628
rect 3164 4340 3220 8764
rect 3164 4274 3220 4284
rect 3340 8652 3660 10164
rect 4172 10724 4228 10734
rect 3340 8596 3368 8652
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3632 8596 3660 8652
rect 3340 7084 3660 8596
rect 3340 7028 3368 7084
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3632 7028 3660 7084
rect 3340 5516 3660 7028
rect 3340 5460 3368 5516
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3632 5460 3660 5516
rect 3052 3938 3108 3948
rect 3340 3948 3660 5460
rect 3340 3892 3368 3948
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3632 3892 3660 3948
rect 3340 3076 3660 3892
rect 3724 9604 3780 9614
rect 3724 3388 3780 9548
rect 3948 9604 4004 9614
rect 3836 8372 3892 8382
rect 3836 7588 3892 8316
rect 3836 7522 3892 7532
rect 3948 3388 4004 9548
rect 4060 8708 4116 8718
rect 4060 6244 4116 8652
rect 4060 5460 4116 6188
rect 4060 5394 4116 5404
rect 4172 5348 4228 10668
rect 4396 10500 4452 10510
rect 4284 8820 4340 8830
rect 4284 6468 4340 8764
rect 4284 6402 4340 6412
rect 4396 5348 4452 10444
rect 4732 10276 4788 10286
rect 4620 9828 4676 9838
rect 4508 8596 4564 8606
rect 4508 5572 4564 8540
rect 4508 5506 4564 5516
rect 4396 5292 4564 5348
rect 4172 5282 4228 5292
rect 4508 5012 4564 5292
rect 3724 3332 3892 3388
rect 3948 3332 4116 3388
rect 2940 2706 2996 2716
rect 3836 2324 3892 3332
rect 3836 2258 3892 2268
rect 4060 980 4116 3332
rect 4508 2772 4564 4956
rect 4620 3444 4676 9772
rect 4732 5796 4788 10220
rect 5496 9436 5816 10948
rect 5496 9380 5524 9436
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 5788 9380 5816 9436
rect 5496 7868 5816 9380
rect 7652 11788 7972 12604
rect 7652 11732 7680 11788
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 7944 11732 7972 11788
rect 7652 10220 7972 11732
rect 7652 10164 7680 10220
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7944 10164 7972 10220
rect 6412 9044 6468 9054
rect 5496 7812 5524 7868
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5788 7812 5816 7868
rect 6076 8260 6132 8270
rect 4732 4900 4788 5740
rect 4732 4834 4788 4844
rect 4956 7588 5012 7598
rect 4956 4116 5012 7532
rect 4956 4050 5012 4060
rect 5068 7140 5124 7150
rect 4620 3378 4676 3388
rect 5068 2884 5124 7084
rect 5068 2818 5124 2828
rect 5180 7028 5236 7038
rect 5180 5908 5236 6972
rect 4508 2706 4564 2716
rect 5180 2660 5236 5852
rect 5496 6300 5816 7812
rect 5964 7812 6020 7822
rect 5964 7476 6020 7756
rect 5964 7410 6020 7420
rect 5496 6244 5524 6300
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5788 6244 5816 6300
rect 5496 4732 5816 6244
rect 5496 4676 5524 4732
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5788 4676 5816 4732
rect 5496 3164 5816 4676
rect 5964 6468 6020 6478
rect 5964 3332 6020 6412
rect 6076 4788 6132 8204
rect 6076 4722 6132 4732
rect 6412 6692 6468 8988
rect 7652 8652 7972 10164
rect 7652 8596 7680 8652
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7944 8596 7972 8652
rect 6412 3444 6468 6636
rect 7196 8036 7252 8046
rect 6524 6244 6580 6254
rect 6524 3556 6580 6188
rect 6524 3490 6580 3500
rect 6412 3378 6468 3388
rect 7196 3444 7252 7980
rect 7532 7476 7588 7486
rect 7532 4004 7588 7420
rect 7532 3938 7588 3948
rect 7652 7084 7972 8596
rect 9808 12572 10128 12604
rect 9808 12516 9836 12572
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 10100 12516 10128 12572
rect 9808 11004 10128 12516
rect 11964 11788 12284 12604
rect 11964 11732 11992 11788
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 12256 11732 12284 11788
rect 9808 10948 9836 11004
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 10100 10948 10128 11004
rect 9808 9436 10128 10948
rect 9808 9380 9836 9436
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 10100 9380 10128 9436
rect 11676 11172 11732 11182
rect 11676 9492 11732 11116
rect 11676 9426 11732 9436
rect 11788 10276 11844 10286
rect 9808 7868 10128 9380
rect 9808 7812 9836 7868
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 10100 7812 10128 7868
rect 7652 7028 7680 7084
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7944 7028 7972 7084
rect 7652 5516 7972 7028
rect 7652 5460 7680 5516
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7944 5460 7972 5516
rect 7652 3948 7972 5460
rect 7196 3378 7252 3388
rect 7652 3892 7680 3948
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7944 3892 7972 3948
rect 5964 3266 6020 3276
rect 5496 3108 5524 3164
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5788 3108 5816 3164
rect 5496 3076 5816 3108
rect 7652 3076 7972 3892
rect 9436 7476 9492 7486
rect 5180 2594 5236 2604
rect 9436 1092 9492 7420
rect 9808 6300 10128 7812
rect 9808 6244 9836 6300
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 10100 6244 10128 6300
rect 9808 4732 10128 6244
rect 9808 4676 9836 4732
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10100 4676 10128 4732
rect 9808 3164 10128 4676
rect 10668 5348 10724 5358
rect 10668 3892 10724 5292
rect 10780 4676 10836 4686
rect 10780 4004 10836 4620
rect 10780 3938 10836 3948
rect 10668 3826 10724 3836
rect 9808 3108 9836 3164
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 10100 3108 10128 3164
rect 11788 3220 11844 10220
rect 11788 3154 11844 3164
rect 11964 10220 12284 11732
rect 11964 10164 11992 10220
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 12256 10164 12284 10220
rect 11964 8652 12284 10164
rect 14120 12572 14440 12604
rect 14120 12516 14148 12572
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14412 12516 14440 12572
rect 14120 11004 14440 12516
rect 16276 11788 16596 12604
rect 16276 11732 16304 11788
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16568 11732 16596 11788
rect 14120 10948 14148 11004
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14412 10948 14440 11004
rect 14120 9436 14440 10948
rect 14120 9380 14148 9436
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14412 9380 14440 9436
rect 11964 8596 11992 8652
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 12256 8596 12284 8652
rect 11964 7084 12284 8596
rect 11964 7028 11992 7084
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 12256 7028 12284 7084
rect 11964 5516 12284 7028
rect 13692 8708 13748 8718
rect 13692 6468 13748 8652
rect 13692 6402 13748 6412
rect 14120 7868 14440 9380
rect 14120 7812 14148 7868
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14412 7812 14440 7868
rect 11964 5460 11992 5516
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 12256 5460 12284 5516
rect 11964 3948 12284 5460
rect 11964 3892 11992 3948
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 12256 3892 12284 3948
rect 9808 3076 10128 3108
rect 11964 3076 12284 3892
rect 14120 6300 14440 7812
rect 14120 6244 14148 6300
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14412 6244 14440 6300
rect 14120 4732 14440 6244
rect 16156 11172 16212 11182
rect 14120 4676 14148 4732
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14412 4676 14440 4732
rect 14120 3164 14440 4676
rect 14120 3108 14148 3164
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14412 3108 14440 3164
rect 14120 3076 14440 3108
rect 14588 5124 14644 5134
rect 14588 2996 14644 5068
rect 16156 3220 16212 11116
rect 16156 3154 16212 3164
rect 16276 10220 16596 11732
rect 18432 12572 18752 12604
rect 18432 12516 18460 12572
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18724 12516 18752 12572
rect 16276 10164 16304 10220
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16568 10164 16596 10220
rect 16276 8652 16596 10164
rect 17612 11284 17668 11294
rect 16276 8596 16304 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16568 8596 16596 8652
rect 16276 7084 16596 8596
rect 16940 9156 16996 9166
rect 16940 7812 16996 9100
rect 16940 7746 16996 7756
rect 17612 9044 17668 11228
rect 16276 7028 16304 7084
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16568 7028 16596 7084
rect 16276 5516 16596 7028
rect 16276 5460 16304 5516
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16568 5460 16596 5516
rect 16276 3948 16596 5460
rect 16276 3892 16304 3948
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16568 3892 16596 3948
rect 16276 3076 16596 3892
rect 14588 2930 14644 2940
rect 9436 1026 9492 1036
rect 4060 914 4116 924
rect 17612 980 17668 8988
rect 18432 11004 18752 12516
rect 18432 10948 18460 11004
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18724 10948 18752 11004
rect 18432 9436 18752 10948
rect 18432 9380 18460 9436
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18724 9380 18752 9436
rect 18432 7868 18752 9380
rect 18432 7812 18460 7868
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18724 7812 18752 7868
rect 18432 6300 18752 7812
rect 18432 6244 18460 6300
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18724 6244 18752 6300
rect 18432 4732 18752 6244
rect 18432 4676 18460 4732
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18724 4676 18752 4732
rect 18432 3164 18752 4676
rect 18432 3108 18460 3164
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18724 3108 18752 3164
rect 18432 3076 18752 3108
rect 17612 914 17668 924
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _040_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _041_
timestamp 1698431365
transform 1 0 3248 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _042_
timestamp 1698431365
transform 1 0 4032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _043_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _044_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _045_
timestamp 1698431365
transform 1 0 5040 0 -1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _046_
timestamp 1698431365
transform -1 0 9184 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _047_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _048_
timestamp 1698431365
transform -1 0 17472 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _049_
timestamp 1698431365
transform 1 0 11088 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _050_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _051_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17360 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _052_
timestamp 1698431365
transform -1 0 18368 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _053_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _054_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5040 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _055_
timestamp 1698431365
transform -1 0 8064 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _056_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6720 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _057_
timestamp 1698431365
transform 1 0 5040 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _058_
timestamp 1698431365
transform 1 0 6944 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _059_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _060_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _061_
timestamp 1698431365
transform -1 0 12320 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _062_
timestamp 1698431365
transform -1 0 11088 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _063_
timestamp 1698431365
transform 1 0 12320 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _064_
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _065_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _066_
timestamp 1698431365
transform 1 0 11200 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _067_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _068_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _069_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16576 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _070_
timestamp 1698431365
transform -1 0 14448 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _071_
timestamp 1698431365
transform 1 0 10416 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _072_
timestamp 1698431365
transform -1 0 14000 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _073_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _074_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6832 0 1 3136
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _075_
timestamp 1698431365
transform 1 0 7504 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _076_
timestamp 1698431365
transform -1 0 8960 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _077_
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _078_
timestamp 1698431365
transform 1 0 4256 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _079_
timestamp 1698431365
transform -1 0 5264 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _080_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _081_
timestamp 1698431365
transform 1 0 15120 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _082_
timestamp 1698431365
transform -1 0 16576 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _083_
timestamp 1698431365
transform 1 0 5712 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _084_
timestamp 1698431365
transform -1 0 7056 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__A2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__A1
timestamp 1698431365
transform -1 0 11760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__C
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__A1
timestamp 1698431365
transform -1 0 12320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__B
timestamp 1698431365
transform 1 0 10640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__C
timestamp 1698431365
transform -1 0 12208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__B
timestamp 1698431365
transform -1 0 14560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__A3
timestamp 1698431365
transform -1 0 2016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__B
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__B
timestamp 1698431365
transform 1 0 7056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 12656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 8848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 5936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 7280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 9520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 5152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 11200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 9968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 11760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 12208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 7728 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 11312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 14224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 2016 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 14896 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 12768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 15456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 4592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 15904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 7280 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 7504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 6832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 6384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 6720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 6608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 7504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform 1 0 5600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 13104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output44_I
timestamp 1698431365
transform 1 0 8176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 11424 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_49
timestamp 1698431365
transform 1 0 6832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_51 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7056 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_144
timestamp 1698431365
transform 1 0 17472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_16
timestamp 1698431365
transform 1 0 3136 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_80
timestamp 1698431365
transform 1 0 10304 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_9
timestamp 1698431365
transform 1 0 2352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_150
timestamp 1698431365
transform 1 0 18144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_74
timestamp 1698431365
transform 1 0 9632 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_81
timestamp 1698431365
transform 1 0 10416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_83
timestamp 1698431365
transform 1 0 10640 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_48
timestamp 1698431365
transform 1 0 6720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_92
timestamp 1698431365
transform 1 0 11648 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_14
timestamp 1698431365
transform 1 0 2912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_22
timestamp 1698431365
transform 1 0 3808 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_79
timestamp 1698431365
transform 1 0 10192 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_86
timestamp 1698431365
transform 1 0 10976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_4
timestamp 1698431365
transform 1 0 1792 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_11
timestamp 1698431365
transform 1 0 2576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_13
timestamp 1698431365
transform 1 0 2800 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_22
timestamp 1698431365
transform 1 0 3808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_47
timestamp 1698431365
transform 1 0 6608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_150
timestamp 1698431365
transform 1 0 18144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_30
timestamp 1698431365
transform 1 0 4704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_32
timestamp 1698431365
transform 1 0 4928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_109
timestamp 1698431365
transform 1 0 13552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_148
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_30
timestamp 1698431365
transform 1 0 4704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_41
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_49
timestamp 1698431365
transform 1 0 6832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_57
timestamp 1698431365
transform 1 0 7728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_65
timestamp 1698431365
transform 1 0 8624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_73
timestamp 1698431365
transform 1 0 9520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_77
timestamp 1698431365
transform 1 0 9968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_86
timestamp 1698431365
transform 1 0 10976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698431365
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_51
timestamp 1698431365
transform 1 0 7056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_55
timestamp 1698431365
transform 1 0 7504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_59
timestamp 1698431365
transform 1 0 7952 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_63 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_82
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_85
timestamp 1698431365
transform 1 0 10864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_89
timestamp 1698431365
transform 1 0 11312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_93
timestamp 1698431365
transform 1 0 11760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_97
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_101
timestamp 1698431365
transform 1 0 12656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_113
timestamp 1698431365
transform 1 0 14000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_127
timestamp 1698431365
transform 1 0 15568 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_148
timestamp 1698431365
transform 1 0 17920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_22
timestamp 1698431365
transform 1 0 3808 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_29
timestamp 1698431365
transform 1 0 4592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_33
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_49
timestamp 1698431365
transform 1 0 6832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_57 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7728 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_89
timestamp 1698431365
transform 1 0 11312 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_93
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_97
timestamp 1698431365
transform 1 0 12208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_115
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_121
timestamp 1698431365
transform 1 0 14896 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_125
timestamp 1698431365
transform 1 0 15344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_143
timestamp 1698431365
transform 1 0 17360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_151
timestamp 1698431365
transform 1 0 18256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_33
timestamp 1698431365
transform 1 0 5040 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_36
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_40
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_44
timestamp 1698431365
transform 1 0 6272 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_48
timestamp 1698431365
transform 1 0 6720 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_52
timestamp 1698431365
transform 1 0 7168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_54
timestamp 1698431365
transform 1 0 7392 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_59
timestamp 1698431365
transform 1 0 7952 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_67
timestamp 1698431365
transform 1 0 8848 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_70 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_86
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_94
timestamp 1698431365
transform 1 0 11872 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_98
timestamp 1698431365
transform 1 0 12320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_114
timestamp 1698431365
transform 1 0 14112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_118
timestamp 1698431365
transform 1 0 14560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_126
timestamp 1698431365
transform 1 0 15456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_130
timestamp 1698431365
transform 1 0 15904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 18368 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1680 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 3920 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 1904 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 4592 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 9520 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 3136 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 9744 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 12432 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 10752 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1698431365
transform 1 0 1680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 17472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 14224 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 18144 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 14448 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 18144 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 14896 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 17920 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 17920 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698431365
transform -1 0 16240 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input24
timestamp 1698431365
transform -1 0 17696 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698431365
transform 1 0 3696 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 17920 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 18256 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input28
timestamp 1698431365
transform 1 0 2352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 2576 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 3696 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 7504 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 3248 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 4368 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 3024 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input38
timestamp 1698431365
transform 1 0 1680 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input39 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2352 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 16352 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output41 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output42 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4144 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43
timestamp 1698431365
transform -1 0 4256 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform -1 0 3136 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output45
timestamp 1698431365
transform -1 0 3136 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_12 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_13
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_14
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 18592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_15
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 18592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_16
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 18592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_17
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_18
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 18592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_19
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 18592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_20
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 18592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_21
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 18592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_22
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 18592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_23
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 18592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_24 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_25
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_26
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_27
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_28
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_29
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_30
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_31
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_32
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_33
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_34
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_35
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_36
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_37
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_38
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_39
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_40
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_41
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_42
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_43
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_44
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_45
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_46
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_47
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_48
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_49
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_50
timestamp 1698431365
transform 1 0 12768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_51
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_46 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_47
timestamp 1698431365
transform -1 0 7952 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_48
timestamp 1698431365
transform -1 0 3808 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_49
timestamp 1698431365
transform -1 0 3360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_50
timestamp 1698431365
transform -1 0 3360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_51
timestamp 1698431365
transform -1 0 2912 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_52
timestamp 1698431365
transform -1 0 3808 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_53
timestamp 1698431365
transform -1 0 3360 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_54
timestamp 1698431365
transform -1 0 2912 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_55
timestamp 1698431365
transform -1 0 3808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_56
timestamp 1698431365
transform -1 0 3360 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_57
timestamp 1698431365
transform -1 0 2016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_58
timestamp 1698431365
transform -1 0 6608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_59
timestamp 1698431365
transform -1 0 4256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_60
timestamp 1698431365
transform -1 0 3808 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_61
timestamp 1698431365
transform -1 0 4704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_62
timestamp 1698431365
transform -1 0 2464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_63
timestamp 1698431365
transform -1 0 4704 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_64
timestamp 1698431365
transform -1 0 2464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_65
timestamp 1698431365
transform -1 0 2912 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_66
timestamp 1698431365
transform -1 0 2016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_67
timestamp 1698431365
transform -1 0 2016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_68
timestamp 1698431365
transform -1 0 2464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_69
timestamp 1698431365
transform -1 0 2016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_70
timestamp 1698431365
transform -1 0 2464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_71
timestamp 1698431365
transform -1 0 2912 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_72
timestamp 1698431365
transform -1 0 2464 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_73
timestamp 1698431365
transform -1 0 3360 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_74
timestamp 1698431365
transform -1 0 3808 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_75
timestamp 1698431365
transform -1 0 4592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_76
timestamp 1698431365
transform -1 0 5040 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_77
timestamp 1698431365
transform -1 0 2016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wb_buttons_leds_78
timestamp 1698431365
transform -1 0 4256 0 1 9408
box -86 -86 534 870
<< labels >>
flabel metal4 s 3340 3076 3660 12604 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 7652 3076 7972 12604 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 11964 3076 12284 12604 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 16276 3076 16596 12604 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 5496 3076 5816 12604 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 9808 3076 10128 12604 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 14120 3076 14440 12604 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 18432 3076 18752 12604 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 s 19200 3808 20000 3920 0 FreeSans 448 0 0 0 buttons[0]
port 2 nsew signal input
flabel metal3 s 19200 11872 20000 11984 0 FreeSans 448 0 0 0 buttons[1]
port 3 nsew signal input
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 clk
port 4 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 i_wb_addr[0]
port 5 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 i_wb_addr[10]
port 6 nsew signal input
flabel metal2 s 8512 0 8624 800 0 FreeSans 448 90 0 0 i_wb_addr[11]
port 7 nsew signal input
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 i_wb_addr[12]
port 8 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 i_wb_addr[13]
port 9 nsew signal input
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 i_wb_addr[14]
port 10 nsew signal input
flabel metal2 s 10304 0 10416 800 0 FreeSans 448 90 0 0 i_wb_addr[15]
port 11 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 i_wb_addr[16]
port 12 nsew signal input
flabel metal2 s 11200 0 11312 800 0 FreeSans 448 90 0 0 i_wb_addr[17]
port 13 nsew signal input
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 i_wb_addr[18]
port 14 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 i_wb_addr[19]
port 15 nsew signal input
flabel metal2 s 3584 0 3696 800 0 FreeSans 448 90 0 0 i_wb_addr[1]
port 16 nsew signal input
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 i_wb_addr[20]
port 17 nsew signal input
flabel metal2 s 12992 0 13104 800 0 FreeSans 448 90 0 0 i_wb_addr[21]
port 18 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 i_wb_addr[22]
port 19 nsew signal input
flabel metal2 s 13888 0 14000 800 0 FreeSans 448 90 0 0 i_wb_addr[23]
port 20 nsew signal input
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 i_wb_addr[24]
port 21 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 i_wb_addr[25]
port 22 nsew signal input
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 i_wb_addr[26]
port 23 nsew signal input
flabel metal2 s 15680 0 15792 800 0 FreeSans 448 90 0 0 i_wb_addr[27]
port 24 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 i_wb_addr[28]
port 25 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 i_wb_addr[29]
port 26 nsew signal input
flabel metal2 s 4480 0 4592 800 0 FreeSans 448 90 0 0 i_wb_addr[2]
port 27 nsew signal input
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 i_wb_addr[30]
port 28 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 i_wb_addr[31]
port 29 nsew signal input
flabel metal2 s 4928 0 5040 800 0 FreeSans 448 90 0 0 i_wb_addr[3]
port 30 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 i_wb_addr[4]
port 31 nsew signal input
flabel metal2 s 5824 0 5936 800 0 FreeSans 448 90 0 0 i_wb_addr[5]
port 32 nsew signal input
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 i_wb_addr[6]
port 33 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 i_wb_addr[7]
port 34 nsew signal input
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 i_wb_addr[8]
port 35 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 i_wb_addr[9]
port 36 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 i_wb_cyc
port 37 nsew signal input
flabel metal2 s 3136 0 3248 800 0 FreeSans 448 90 0 0 i_wb_data[0]
port 38 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 i_wb_data[1]
port 39 nsew signal input
flabel metal2 s 1792 0 1904 800 0 FreeSans 448 90 0 0 i_wb_stb
port 40 nsew signal input
flabel metal2 s 2240 0 2352 800 0 FreeSans 448 90 0 0 i_wb_we
port 41 nsew signal input
flabel metal2 s 17248 15200 17360 16000 0 FreeSans 448 90 0 0 led_enb[0]
port 42 nsew signal tristate
flabel metal2 s 7392 15200 7504 16000 0 FreeSans 448 90 0 0 led_enb[1]
port 43 nsew signal tristate
flabel metal2 s 12320 15200 12432 16000 0 FreeSans 448 90 0 0 leds[0]
port 44 nsew signal tristate
flabel metal2 s 2464 15200 2576 16000 0 FreeSans 448 90 0 0 leds[1]
port 45 nsew signal tristate
flabel metal3 s 0 448 800 560 0 FreeSans 448 0 0 0 o_wb_ack
port 46 nsew signal tristate
flabel metal3 s 0 1344 800 1456 0 FreeSans 448 0 0 0 o_wb_data[0]
port 47 nsew signal tristate
flabel metal3 s 0 5824 800 5936 0 FreeSans 448 0 0 0 o_wb_data[10]
port 48 nsew signal tristate
flabel metal3 s 0 6272 800 6384 0 FreeSans 448 0 0 0 o_wb_data[11]
port 49 nsew signal tristate
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 o_wb_data[12]
port 50 nsew signal tristate
flabel metal3 s 0 7168 800 7280 0 FreeSans 448 0 0 0 o_wb_data[13]
port 51 nsew signal tristate
flabel metal3 s 0 7616 800 7728 0 FreeSans 448 0 0 0 o_wb_data[14]
port 52 nsew signal tristate
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 o_wb_data[15]
port 53 nsew signal tristate
flabel metal3 s 0 8512 800 8624 0 FreeSans 448 0 0 0 o_wb_data[16]
port 54 nsew signal tristate
flabel metal3 s 0 8960 800 9072 0 FreeSans 448 0 0 0 o_wb_data[17]
port 55 nsew signal tristate
flabel metal3 s 0 9408 800 9520 0 FreeSans 448 0 0 0 o_wb_data[18]
port 56 nsew signal tristate
flabel metal3 s 0 9856 800 9968 0 FreeSans 448 0 0 0 o_wb_data[19]
port 57 nsew signal tristate
flabel metal3 s 0 1792 800 1904 0 FreeSans 448 0 0 0 o_wb_data[1]
port 58 nsew signal tristate
flabel metal3 s 0 10304 800 10416 0 FreeSans 448 0 0 0 o_wb_data[20]
port 59 nsew signal tristate
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 o_wb_data[21]
port 60 nsew signal tristate
flabel metal3 s 0 11200 800 11312 0 FreeSans 448 0 0 0 o_wb_data[22]
port 61 nsew signal tristate
flabel metal3 s 0 11648 800 11760 0 FreeSans 448 0 0 0 o_wb_data[23]
port 62 nsew signal tristate
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 o_wb_data[24]
port 63 nsew signal tristate
flabel metal3 s 0 12544 800 12656 0 FreeSans 448 0 0 0 o_wb_data[25]
port 64 nsew signal tristate
flabel metal3 s 0 12992 800 13104 0 FreeSans 448 0 0 0 o_wb_data[26]
port 65 nsew signal tristate
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 o_wb_data[27]
port 66 nsew signal tristate
flabel metal3 s 0 13888 800 14000 0 FreeSans 448 0 0 0 o_wb_data[28]
port 67 nsew signal tristate
flabel metal3 s 0 14336 800 14448 0 FreeSans 448 0 0 0 o_wb_data[29]
port 68 nsew signal tristate
flabel metal3 s 0 2240 800 2352 0 FreeSans 448 0 0 0 o_wb_data[2]
port 69 nsew signal tristate
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 o_wb_data[30]
port 70 nsew signal tristate
flabel metal3 s 0 15232 800 15344 0 FreeSans 448 0 0 0 o_wb_data[31]
port 71 nsew signal tristate
flabel metal3 s 0 2688 800 2800 0 FreeSans 448 0 0 0 o_wb_data[3]
port 72 nsew signal tristate
flabel metal3 s 0 3136 800 3248 0 FreeSans 448 0 0 0 o_wb_data[4]
port 73 nsew signal tristate
flabel metal3 s 0 3584 800 3696 0 FreeSans 448 0 0 0 o_wb_data[5]
port 74 nsew signal tristate
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 o_wb_data[6]
port 75 nsew signal tristate
flabel metal3 s 0 4480 800 4592 0 FreeSans 448 0 0 0 o_wb_data[7]
port 76 nsew signal tristate
flabel metal3 s 0 4928 800 5040 0 FreeSans 448 0 0 0 o_wb_data[8]
port 77 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 o_wb_data[9]
port 78 nsew signal tristate
flabel metal3 s 0 896 800 1008 0 FreeSans 448 0 0 0 o_wb_stall
port 79 nsew signal tristate
flabel metal2 s 18368 0 18480 800 0 FreeSans 448 90 0 0 reset
port 80 nsew signal input
rlabel metal1 9968 11760 9968 11760 0 VDD
rlabel via1 10048 12544 10048 12544 0 VSS
rlabel metal2 10584 6552 10584 6552 0 _000_
rlabel metal3 16408 8344 16408 8344 0 _001_
rlabel metal2 13720 7280 13720 7280 0 _002_
rlabel metal3 8176 4536 8176 4536 0 _003_
rlabel metal2 4984 8400 4984 8400 0 _004_
rlabel metal2 4872 7336 4872 7336 0 _005_
rlabel metal2 9800 4368 9800 4368 0 _006_
rlabel metal2 6440 7280 6440 7280 0 _007_
rlabel metal3 18648 5880 18648 5880 0 _008_
rlabel metal2 11368 4200 11368 4200 0 _009_
rlabel metal2 7896 3640 7896 3640 0 _010_
rlabel metal2 7560 3472 7560 3472 0 _011_
rlabel metal2 11592 4200 11592 4200 0 _012_
rlabel metal2 15848 4592 15848 4592 0 _013_
rlabel metal3 15624 4480 15624 4480 0 _014_
rlabel metal2 11480 6160 11480 6160 0 _015_
rlabel metal2 16408 11088 16408 11088 0 _016_
rlabel metal2 15736 4144 15736 4144 0 _017_
rlabel metal2 13944 4144 13944 4144 0 _018_
rlabel metal2 6552 6160 6552 6160 0 _019_
rlabel metal2 7336 3472 7336 3472 0 _020_
rlabel metal2 5824 4424 5824 4424 0 _021_
rlabel metal2 12376 3332 12376 3332 0 _022_
rlabel metal3 8792 6552 8792 6552 0 _023_
rlabel metal2 17416 7728 17416 7728 0 _024_
rlabel metal3 11480 3752 11480 3752 0 _025_
rlabel metal2 10920 5600 10920 5600 0 _026_
rlabel metal2 12600 7056 12600 7056 0 _027_
rlabel metal2 17360 6104 17360 6104 0 _028_
rlabel metal2 17080 7840 17080 7840 0 _029_
rlabel metal3 16744 8064 16744 8064 0 _030_
rlabel metal2 7504 3752 7504 3752 0 _031_
rlabel metal2 17528 6496 17528 6496 0 _032_
rlabel metal2 13832 7448 13832 7448 0 _033_
rlabel metal2 13496 7392 13496 7392 0 _034_
rlabel metal2 14056 7896 14056 7896 0 _035_
rlabel metal2 6552 3416 6552 3416 0 _036_
rlabel metal2 5096 6104 5096 6104 0 _037_
rlabel metal2 10136 4480 10136 4480 0 _038_
rlabel metal2 4592 3640 4592 3640 0 _039_
rlabel metal3 18536 10472 18536 10472 0 buttons[0]
rlabel metal3 18690 11928 18690 11928 0 buttons[1]
rlabel metal2 16744 7280 16744 7280 0 clk
rlabel metal2 12152 7896 12152 7896 0 clknet_0_clk
rlabel metal3 7000 8120 7000 8120 0 clknet_1_0__leaf_clk
rlabel metal2 16240 8232 16240 8232 0 clknet_1_1__leaf_clk
rlabel metal3 1904 5096 1904 5096 0 i_wb_addr[0]
rlabel metal2 4088 4536 4088 4536 0 i_wb_addr[10]
rlabel metal2 2184 8176 2184 8176 0 i_wb_addr[11]
rlabel metal2 4760 5208 4760 5208 0 i_wb_addr[12]
rlabel metal3 9576 7448 9576 7448 0 i_wb_addr[13]
rlabel metal2 5096 8344 5096 8344 0 i_wb_addr[14]
rlabel metal2 10472 5880 10472 5880 0 i_wb_addr[15]
rlabel metal2 5824 6664 5824 6664 0 i_wb_addr[16]
rlabel metal2 11256 2058 11256 2058 0 i_wb_addr[17]
rlabel metal2 11704 3710 11704 3710 0 i_wb_addr[18]
rlabel metal2 12320 3528 12320 3528 0 i_wb_addr[19]
rlabel metal2 1848 6160 1848 6160 0 i_wb_addr[1]
rlabel metal2 11256 10360 11256 10360 0 i_wb_addr[20]
rlabel metal2 14392 10360 14392 10360 0 i_wb_addr[21]
rlabel metal2 1960 3976 1960 3976 0 i_wb_addr[22]
rlabel metal2 13944 2058 13944 2058 0 i_wb_addr[23]
rlabel metal3 15680 5096 15680 5096 0 i_wb_addr[24]
rlabel metal2 15064 10192 15064 10192 0 i_wb_addr[25]
rlabel metal2 15288 2534 15288 2534 0 i_wb_addr[26]
rlabel metal4 17640 4984 17640 4984 0 i_wb_addr[27]
rlabel metal2 16072 11200 16072 11200 0 i_wb_addr[28]
rlabel metal2 16632 2058 16632 2058 0 i_wb_addr[29]
rlabel metal2 3976 6272 3976 6272 0 i_wb_addr[2]
rlabel metal2 17080 1246 17080 1246 0 i_wb_addr[30]
rlabel metal2 18088 10976 18088 10976 0 i_wb_addr[31]
rlabel metal3 2996 5880 2996 5880 0 i_wb_addr[3]
rlabel metal2 5656 8064 5656 8064 0 i_wb_addr[4]
rlabel metal3 2968 4984 2968 4984 0 i_wb_addr[5]
rlabel metal2 3864 6104 3864 6104 0 i_wb_addr[6]
rlabel metal2 7224 7616 7224 7616 0 i_wb_addr[7]
rlabel metal2 3528 5040 3528 5040 0 i_wb_addr[8]
rlabel metal2 6608 12040 6608 12040 0 i_wb_addr[9]
rlabel metal2 1400 2058 1400 2058 0 i_wb_cyc
rlabel metal2 3304 6160 3304 6160 0 i_wb_data[0]
rlabel metal4 2520 8736 2520 8736 0 i_wb_data[1]
rlabel metal4 1848 8176 1848 8176 0 i_wb_stb
rlabel metal3 2688 6664 2688 6664 0 i_wb_we
rlabel metal2 13608 12208 13608 12208 0 leds[0]
rlabel metal2 3080 12488 3080 12488 0 leds[1]
rlabel metal2 17640 7672 17640 7672 0 net1
rlabel metal3 9744 3304 9744 3304 0 net10
rlabel metal2 10248 5544 10248 5544 0 net11
rlabel metal2 11872 6440 11872 6440 0 net12
rlabel metal2 11200 4312 11200 4312 0 net13
rlabel metal3 3976 5936 3976 5936 0 net14
rlabel metal2 13496 4760 13496 4760 0 net15
rlabel metal2 14168 5544 14168 5544 0 net16
rlabel metal2 16744 5712 16744 5712 0 net17
rlabel metal2 14952 8456 14952 8456 0 net18
rlabel metal2 17640 5040 17640 5040 0 net19
rlabel metal2 17864 11872 17864 11872 0 net2
rlabel metal2 15344 10696 15344 10696 0 net20
rlabel metal2 17416 4592 17416 4592 0 net21
rlabel metal2 17416 8848 17416 8848 0 net22
rlabel metal3 15176 3528 15176 3528 0 net23
rlabel metal1 18200 12712 18200 12712 0 net24
rlabel metal2 7224 6664 7224 6664 0 net25
rlabel metal2 17416 10864 17416 10864 0 net26
rlabel metal2 17080 11368 17080 11368 0 net27
rlabel metal2 2856 5712 2856 5712 0 net28
rlabel metal2 5992 7504 5992 7504 0 net29
rlabel metal2 3976 5040 3976 5040 0 net3
rlabel metal2 3080 5096 3080 5096 0 net30
rlabel metal3 4480 5992 4480 5992 0 net31
rlabel metal2 7000 6944 7000 6944 0 net32
rlabel metal2 3752 5208 3752 5208 0 net33
rlabel metal2 4872 6048 4872 6048 0 net34
rlabel metal2 6440 4480 6440 4480 0 net35
rlabel metal2 3472 6104 3472 6104 0 net36
rlabel metal2 2744 7896 2744 7896 0 net37
rlabel metal2 12040 9296 12040 9296 0 net38
rlabel metal2 17976 6776 17976 6776 0 net39
rlabel metal2 4424 6720 4424 6720 0 net4
rlabel metal2 17864 3808 17864 3808 0 net40
rlabel metal2 13272 10976 13272 10976 0 net41
rlabel metal2 3976 10136 3976 10136 0 net42
rlabel metal2 13944 8848 13944 8848 0 net43
rlabel metal3 2128 3528 2128 3528 0 net44
rlabel metal2 1512 6160 1512 6160 0 net45
rlabel metal3 16856 12376 16856 12376 0 net46
rlabel metal2 7560 12376 7560 12376 0 net47
rlabel metal3 2310 2296 2310 2296 0 net48
rlabel metal3 1246 2744 1246 2744 0 net49
rlabel metal2 2408 8512 2408 8512 0 net5
rlabel metal3 1694 3192 1694 3192 0 net50
rlabel metal3 1582 3640 1582 3640 0 net51
rlabel metal3 1974 4088 1974 4088 0 net52
rlabel metal3 1022 4536 1022 4536 0 net53
rlabel metal3 1638 4984 1638 4984 0 net54
rlabel metal3 1750 5432 1750 5432 0 net55
rlabel metal3 1190 5880 1190 5880 0 net56
rlabel metal3 1190 6328 1190 6328 0 net57
rlabel metal3 1862 6776 1862 6776 0 net58
rlabel metal2 3976 8176 3976 8176 0 net59
rlabel metal2 5096 5040 5096 5040 0 net6
rlabel metal2 3752 9184 3752 9184 0 net60
rlabel metal3 1246 8120 1246 8120 0 net61
rlabel metal3 1470 8568 1470 8568 0 net62
rlabel metal3 4424 9072 4424 9072 0 net63
rlabel metal3 1470 9464 1470 9464 0 net64
rlabel metal3 1694 9912 1694 9912 0 net65
rlabel metal3 1246 10360 1246 10360 0 net66
rlabel metal3 1246 10808 1246 10808 0 net67
rlabel metal3 1470 11256 1470 11256 0 net68
rlabel metal3 1246 11704 1246 11704 0 net69
rlabel metal2 10024 7000 10024 7000 0 net7
rlabel metal3 1470 12152 1470 12152 0 net70
rlabel metal2 2632 11928 2632 11928 0 net71
rlabel metal2 2128 10808 2128 10808 0 net72
rlabel metal2 3024 11256 3024 11256 0 net73
rlabel metal2 3640 11256 3640 11256 0 net74
rlabel metal2 4312 13384 4312 13384 0 net75
rlabel metal2 4760 13608 4760 13608 0 net76
rlabel metal2 1792 9688 1792 9688 0 net77
rlabel metal3 2422 952 2422 952 0 net78
rlabel metal2 3640 8008 3640 8008 0 net8
rlabel metal2 10808 6328 10808 6328 0 net9
rlabel metal3 2058 504 2058 504 0 o_wb_ack
rlabel metal3 1470 1400 1470 1400 0 o_wb_data[0]
rlabel metal3 1414 1848 1414 1848 0 o_wb_data[1]
rlabel metal2 18424 1246 18424 1246 0 reset
<< properties >>
string FIXED_BBOX 0 0 20000 16000
<< end >>
