VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pinmux_top
  CLASS BLOCK ;
  FOREIGN pinmux_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 1000.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
  END VSS
  PIN digital_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 937.440 4.000 938.000 ;
    END
  END digital_io_in[21]
  PIN digital_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 880.320 4.000 880.880 ;
    END
  END digital_io_in[22]
  PIN digital_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 823.200 4.000 823.760 ;
    END
  END digital_io_in[23]
  PIN digital_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 804.160 4.000 804.720 ;
    END
  END digital_io_in[24]
  PIN digital_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 747.040 4.000 747.600 ;
    END
  END digital_io_in[25]
  PIN digital_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 689.920 4.000 690.480 ;
    END
  END digital_io_in[26]
  PIN digital_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 632.800 4.000 633.360 ;
    END
  END digital_io_in[27]
  PIN digital_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 575.680 4.000 576.240 ;
    END
  END digital_io_in[28]
  PIN digital_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 518.560 4.000 519.120 ;
    END
  END digital_io_in[29]
  PIN digital_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 461.440 4.000 462.000 ;
    END
  END digital_io_in[30]
  PIN digital_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 404.320 4.000 404.880 ;
    END
  END digital_io_in[31]
  PIN digital_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.200 4.000 347.760 ;
    END
  END digital_io_in[32]
  PIN digital_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 290.080 4.000 290.640 ;
    END
  END digital_io_in[33]
  PIN digital_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.960 4.000 233.520 ;
    END
  END digital_io_in[34]
  PIN digital_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 175.840 4.000 176.400 ;
    END
  END digital_io_in[35]
  PIN digital_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END digital_io_in[36]
  PIN digital_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 4.000 62.160 ;
    END
  END digital_io_in[37]
  PIN digital_io_oen[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 975.520 4.000 976.080 ;
    END
  END digital_io_oen[21]
  PIN digital_io_oen[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 918.400 4.000 918.960 ;
    END
  END digital_io_oen[22]
  PIN digital_io_oen[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 861.280 4.000 861.840 ;
    END
  END digital_io_oen[23]
  PIN digital_io_oen[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 766.080 4.000 766.640 ;
    END
  END digital_io_oen[24]
  PIN digital_io_oen[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 708.960 4.000 709.520 ;
    END
  END digital_io_oen[25]
  PIN digital_io_oen[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 651.840 4.000 652.400 ;
    END
  END digital_io_oen[26]
  PIN digital_io_oen[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 594.720 4.000 595.280 ;
    END
  END digital_io_oen[27]
  PIN digital_io_oen[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END digital_io_oen[28]
  PIN digital_io_oen[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 480.480 4.000 481.040 ;
    END
  END digital_io_oen[29]
  PIN digital_io_oen[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 423.360 4.000 423.920 ;
    END
  END digital_io_oen[30]
  PIN digital_io_oen[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 366.240 4.000 366.800 ;
    END
  END digital_io_oen[31]
  PIN digital_io_oen[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.120 4.000 309.680 ;
    END
  END digital_io_oen[32]
  PIN digital_io_oen[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END digital_io_oen[33]
  PIN digital_io_oen[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END digital_io_oen[34]
  PIN digital_io_oen[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END digital_io_oen[35]
  PIN digital_io_oen[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END digital_io_oen[36]
  PIN digital_io_oen[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END digital_io_oen[37]
  PIN digital_io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 956.480 4.000 957.040 ;
    END
  END digital_io_out[21]
  PIN digital_io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 899.360 4.000 899.920 ;
    END
  END digital_io_out[22]
  PIN digital_io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 842.240 4.000 842.800 ;
    END
  END digital_io_out[23]
  PIN digital_io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 785.120 4.000 785.680 ;
    END
  END digital_io_out[24]
  PIN digital_io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 728.000 4.000 728.560 ;
    END
  END digital_io_out[25]
  PIN digital_io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 670.880 4.000 671.440 ;
    END
  END digital_io_out[26]
  PIN digital_io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 613.760 4.000 614.320 ;
    END
  END digital_io_out[27]
  PIN digital_io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 556.640 4.000 557.200 ;
    END
  END digital_io_out[28]
  PIN digital_io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 499.520 4.000 500.080 ;
    END
  END digital_io_out[29]
  PIN digital_io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.400 4.000 442.960 ;
    END
  END digital_io_out[30]
  PIN digital_io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 385.280 4.000 385.840 ;
    END
  END digital_io_out[31]
  PIN digital_io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.160 4.000 328.720 ;
    END
  END digital_io_out[32]
  PIN digital_io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.040 4.000 271.600 ;
    END
  END digital_io_out[33]
  PIN digital_io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.920 4.000 214.480 ;
    END
  END digital_io_out[34]
  PIN digital_io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 156.800 4.000 157.360 ;
    END
  END digital_io_out[35]
  PIN digital_io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 4.000 100.240 ;
    END
  END digital_io_out[36]
  PIN digital_io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 4.000 43.120 ;
    END
  END digital_io_out[37]
  PIN e_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 4.000 ;
    END
  END e_reset_n
  PIN i2cm_clk_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 996.000 485.520 1000.000 ;
    END
  END i2cm_clk_i
  PIN i2cm_clk_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 996.000 449.680 1000.000 ;
    END
  END i2cm_clk_o
  PIN i2cm_clk_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 996.000 521.360 1000.000 ;
    END
  END i2cm_clk_oen
  PIN i2cm_data_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 996.000 628.880 1000.000 ;
    END
  END i2cm_data_i
  PIN i2cm_data_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 996.000 593.040 1000.000 ;
    END
  END i2cm_data_o
  PIN i2cm_data_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 556.640 996.000 557.200 1000.000 ;
    END
  END i2cm_data_oen
  PIN i2cm_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 996.000 342.160 1000.000 ;
    END
  END i2cm_intr
  PIN i2cm_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 996.000 127.120 1000.000 ;
    END
  END i2cm_rst_n
  PIN mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END mclk
  PIN p_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 4.000 ;
    END
  END p_reset_n
  PIN pulse1m_mclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 996.000 413.840 1000.000 ;
    END
  END pulse1m_mclk
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 825.440 0.000 826.000 4.000 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END reg_addr[10]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 0.000 189.840 4.000 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 0.000 180.880 4.000 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 4.000 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 4.000 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 0.000 136.080 4.000 ;
    END
  END reg_addr[8]
  PIN reg_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END reg_addr[9]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 0.000 243.600 4.000 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 4.000 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 0.000 216.720 4.000 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 4.000 ;
    END
  END reg_cs
  PIN reg_peri_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 953.120 900.000 953.680 ;
    END
  END reg_peri_ack
  PIN reg_peri_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 257.600 900.000 258.160 ;
    END
  END reg_peri_addr[0]
  PIN reg_peri_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 156.800 900.000 157.360 ;
    END
  END reg_peri_addr[10]
  PIN reg_peri_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 247.520 900.000 248.080 ;
    END
  END reg_peri_addr[1]
  PIN reg_peri_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 237.440 900.000 238.000 ;
    END
  END reg_peri_addr[2]
  PIN reg_peri_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 227.360 900.000 227.920 ;
    END
  END reg_peri_addr[3]
  PIN reg_peri_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 217.280 900.000 217.840 ;
    END
  END reg_peri_addr[4]
  PIN reg_peri_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 207.200 900.000 207.760 ;
    END
  END reg_peri_addr[5]
  PIN reg_peri_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 197.120 900.000 197.680 ;
    END
  END reg_peri_addr[6]
  PIN reg_peri_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 187.040 900.000 187.600 ;
    END
  END reg_peri_addr[7]
  PIN reg_peri_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 176.960 900.000 177.520 ;
    END
  END reg_peri_addr[8]
  PIN reg_peri_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 166.880 900.000 167.440 ;
    END
  END reg_peri_addr[9]
  PIN reg_peri_be[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 297.920 900.000 298.480 ;
    END
  END reg_peri_be[0]
  PIN reg_peri_be[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 287.840 900.000 288.400 ;
    END
  END reg_peri_be[1]
  PIN reg_peri_be[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 277.760 900.000 278.320 ;
    END
  END reg_peri_be[2]
  PIN reg_peri_be[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 267.680 900.000 268.240 ;
    END
  END reg_peri_be[3]
  PIN reg_peri_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 136.640 900.000 137.200 ;
    END
  END reg_peri_cs
  PIN reg_peri_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 943.040 900.000 943.600 ;
    END
  END reg_peri_rdata[0]
  PIN reg_peri_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 842.240 900.000 842.800 ;
    END
  END reg_peri_rdata[10]
  PIN reg_peri_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 832.160 900.000 832.720 ;
    END
  END reg_peri_rdata[11]
  PIN reg_peri_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 822.080 900.000 822.640 ;
    END
  END reg_peri_rdata[12]
  PIN reg_peri_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 812.000 900.000 812.560 ;
    END
  END reg_peri_rdata[13]
  PIN reg_peri_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 801.920 900.000 802.480 ;
    END
  END reg_peri_rdata[14]
  PIN reg_peri_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 791.840 900.000 792.400 ;
    END
  END reg_peri_rdata[15]
  PIN reg_peri_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 781.760 900.000 782.320 ;
    END
  END reg_peri_rdata[16]
  PIN reg_peri_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 771.680 900.000 772.240 ;
    END
  END reg_peri_rdata[17]
  PIN reg_peri_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 761.600 900.000 762.160 ;
    END
  END reg_peri_rdata[18]
  PIN reg_peri_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 751.520 900.000 752.080 ;
    END
  END reg_peri_rdata[19]
  PIN reg_peri_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 932.960 900.000 933.520 ;
    END
  END reg_peri_rdata[1]
  PIN reg_peri_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 741.440 900.000 742.000 ;
    END
  END reg_peri_rdata[20]
  PIN reg_peri_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 731.360 900.000 731.920 ;
    END
  END reg_peri_rdata[21]
  PIN reg_peri_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 721.280 900.000 721.840 ;
    END
  END reg_peri_rdata[22]
  PIN reg_peri_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 711.200 900.000 711.760 ;
    END
  END reg_peri_rdata[23]
  PIN reg_peri_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 701.120 900.000 701.680 ;
    END
  END reg_peri_rdata[24]
  PIN reg_peri_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 691.040 900.000 691.600 ;
    END
  END reg_peri_rdata[25]
  PIN reg_peri_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 680.960 900.000 681.520 ;
    END
  END reg_peri_rdata[26]
  PIN reg_peri_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 670.880 900.000 671.440 ;
    END
  END reg_peri_rdata[27]
  PIN reg_peri_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 660.800 900.000 661.360 ;
    END
  END reg_peri_rdata[28]
  PIN reg_peri_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 650.720 900.000 651.280 ;
    END
  END reg_peri_rdata[29]
  PIN reg_peri_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 922.880 900.000 923.440 ;
    END
  END reg_peri_rdata[2]
  PIN reg_peri_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 640.640 900.000 641.200 ;
    END
  END reg_peri_rdata[30]
  PIN reg_peri_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 630.560 900.000 631.120 ;
    END
  END reg_peri_rdata[31]
  PIN reg_peri_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 912.800 900.000 913.360 ;
    END
  END reg_peri_rdata[3]
  PIN reg_peri_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 902.720 900.000 903.280 ;
    END
  END reg_peri_rdata[4]
  PIN reg_peri_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 892.640 900.000 893.200 ;
    END
  END reg_peri_rdata[5]
  PIN reg_peri_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 882.560 900.000 883.120 ;
    END
  END reg_peri_rdata[6]
  PIN reg_peri_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 872.480 900.000 873.040 ;
    END
  END reg_peri_rdata[7]
  PIN reg_peri_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 862.400 900.000 862.960 ;
    END
  END reg_peri_rdata[8]
  PIN reg_peri_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 852.320 900.000 852.880 ;
    END
  END reg_peri_rdata[9]
  PIN reg_peri_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 620.480 900.000 621.040 ;
    END
  END reg_peri_wdata[0]
  PIN reg_peri_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 519.680 900.000 520.240 ;
    END
  END reg_peri_wdata[10]
  PIN reg_peri_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 509.600 900.000 510.160 ;
    END
  END reg_peri_wdata[11]
  PIN reg_peri_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 499.520 900.000 500.080 ;
    END
  END reg_peri_wdata[12]
  PIN reg_peri_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 489.440 900.000 490.000 ;
    END
  END reg_peri_wdata[13]
  PIN reg_peri_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 479.360 900.000 479.920 ;
    END
  END reg_peri_wdata[14]
  PIN reg_peri_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 469.280 900.000 469.840 ;
    END
  END reg_peri_wdata[15]
  PIN reg_peri_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 459.200 900.000 459.760 ;
    END
  END reg_peri_wdata[16]
  PIN reg_peri_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 449.120 900.000 449.680 ;
    END
  END reg_peri_wdata[17]
  PIN reg_peri_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 439.040 900.000 439.600 ;
    END
  END reg_peri_wdata[18]
  PIN reg_peri_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 428.960 900.000 429.520 ;
    END
  END reg_peri_wdata[19]
  PIN reg_peri_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 610.400 900.000 610.960 ;
    END
  END reg_peri_wdata[1]
  PIN reg_peri_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 418.880 900.000 419.440 ;
    END
  END reg_peri_wdata[20]
  PIN reg_peri_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 408.800 900.000 409.360 ;
    END
  END reg_peri_wdata[21]
  PIN reg_peri_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 398.720 900.000 399.280 ;
    END
  END reg_peri_wdata[22]
  PIN reg_peri_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 388.640 900.000 389.200 ;
    END
  END reg_peri_wdata[23]
  PIN reg_peri_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 378.560 900.000 379.120 ;
    END
  END reg_peri_wdata[24]
  PIN reg_peri_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 368.480 900.000 369.040 ;
    END
  END reg_peri_wdata[25]
  PIN reg_peri_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 358.400 900.000 358.960 ;
    END
  END reg_peri_wdata[26]
  PIN reg_peri_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 348.320 900.000 348.880 ;
    END
  END reg_peri_wdata[27]
  PIN reg_peri_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 338.240 900.000 338.800 ;
    END
  END reg_peri_wdata[28]
  PIN reg_peri_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 328.160 900.000 328.720 ;
    END
  END reg_peri_wdata[29]
  PIN reg_peri_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 600.320 900.000 600.880 ;
    END
  END reg_peri_wdata[2]
  PIN reg_peri_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 318.080 900.000 318.640 ;
    END
  END reg_peri_wdata[30]
  PIN reg_peri_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 308.000 900.000 308.560 ;
    END
  END reg_peri_wdata[31]
  PIN reg_peri_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 590.240 900.000 590.800 ;
    END
  END reg_peri_wdata[3]
  PIN reg_peri_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 580.160 900.000 580.720 ;
    END
  END reg_peri_wdata[4]
  PIN reg_peri_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 570.080 900.000 570.640 ;
    END
  END reg_peri_wdata[5]
  PIN reg_peri_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 560.000 900.000 560.560 ;
    END
  END reg_peri_wdata[6]
  PIN reg_peri_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 549.920 900.000 550.480 ;
    END
  END reg_peri_wdata[7]
  PIN reg_peri_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 539.840 900.000 540.400 ;
    END
  END reg_peri_wdata[8]
  PIN reg_peri_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 529.760 900.000 530.320 ;
    END
  END reg_peri_wdata[9]
  PIN reg_peri_wr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 146.720 900.000 147.280 ;
    END
  END reg_peri_wr
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 0.000 817.040 4.000 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 726.880 0.000 727.440 4.000 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 717.920 0.000 718.480 4.000 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 0.000 709.520 4.000 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 700.000 0.000 700.560 4.000 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 691.040 0.000 691.600 4.000 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 0.000 682.640 4.000 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 673.120 0.000 673.680 4.000 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 664.160 0.000 664.720 4.000 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 0.000 655.760 4.000 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 0.000 646.800 4.000 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 807.520 0.000 808.080 4.000 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 637.280 0.000 637.840 4.000 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 0.000 628.880 4.000 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 619.360 0.000 619.920 4.000 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 610.400 0.000 610.960 4.000 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 0.000 602.000 4.000 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 0.000 593.040 4.000 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 583.520 0.000 584.080 4.000 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 0.000 566.160 4.000 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 556.640 0.000 557.200 4.000 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 798.560 0.000 799.120 4.000 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 0.000 548.240 4.000 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 0.000 539.280 4.000 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 0.000 790.160 4.000 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 780.640 0.000 781.200 4.000 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 0.000 772.240 4.000 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 0.000 763.280 4.000 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 753.760 0.000 754.320 4.000 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 744.800 0.000 745.360 4.000 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 0.000 736.400 4.000 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 0.000 530.320 4.000 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 0.000 440.720 4.000 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 0.000 431.760 4.000 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 0.000 422.800 4.000 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 0.000 413.840 4.000 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 404.320 0.000 404.880 4.000 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 395.360 0.000 395.920 4.000 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 0.000 378.000 4.000 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 0.000 369.040 4.000 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 0.000 360.080 4.000 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 0.000 521.360 4.000 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 350.560 0.000 351.120 4.000 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 0.000 342.160 4.000 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 0.000 324.240 4.000 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 314.720 0.000 315.280 4.000 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 0.000 288.400 4.000 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 4.000 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 511.840 0.000 512.400 4.000 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 4.000 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 4.000 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 0.000 503.440 4.000 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 0.000 494.480 4.000 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 0.000 485.520 4.000 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 476.000 0.000 476.560 4.000 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 0.000 467.600 4.000 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 4.000 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 0.000 449.680 4.000 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 4.000 ;
    END
  END reg_wr
  PIN rtc_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 996.000 270.480 1000.000 ;
    END
  END rtc_clk
  PIN rtc_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 996.000 306.320 1000.000 ;
    END
  END rtc_intr
  PIN s_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END s_reset_n
  PIN spim_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 996.000 843.920 1000.000 ;
    END
  END spim_miso
  PIN spim_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 879.200 996.000 879.760 1000.000 ;
    END
  END spim_mosi
  PIN spim_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 664.160 996.000 664.720 1000.000 ;
    END
  END spim_sck
  PIN spim_ssn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 807.520 996.000 808.080 1000.000 ;
    END
  END spim_ssn[0]
  PIN spim_ssn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 996.000 772.240 1000.000 ;
    END
  END spim_ssn[1]
  PIN spim_ssn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 996.000 736.400 1000.000 ;
    END
  END spim_ssn[2]
  PIN spim_ssn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 700.000 996.000 700.560 1000.000 ;
    END
  END spim_ssn[3]
  PIN sspim_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 996.000 19.600 1000.000 ;
    END
  END sspim_rst_n
  PIN uart_rst_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 996.000 91.280 1000.000 ;
    END
  END uart_rst_n[0]
  PIN uart_rst_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 996.000 55.440 1000.000 ;
    END
  END uart_rst_n[1]
  PIN uart_rxd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 126.560 900.000 127.120 ;
    END
  END uart_rxd[0]
  PIN uart_rxd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 106.400 900.000 106.960 ;
    END
  END uart_rxd[1]
  PIN uart_txd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 116.480 900.000 117.040 ;
    END
  END uart_txd[0]
  PIN uart_txd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 96.320 900.000 96.880 ;
    END
  END uart_txd[1]
  PIN usb_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 996.000 234.640 1000.000 ;
    END
  END usb_clk
  PIN usb_dn_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 86.240 900.000 86.800 ;
    END
  END usb_dn_i
  PIN usb_dn_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 56.000 900.000 56.560 ;
    END
  END usb_dn_o
  PIN usb_dp_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 76.160 900.000 76.720 ;
    END
  END usb_dp_i
  PIN usb_dp_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 45.920 900.000 46.480 ;
    END
  END usb_dp_o
  PIN usb_intr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 996.000 378.000 1000.000 ;
    END
  END usb_intr
  PIN usb_oen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 66.080 900.000 66.640 ;
    END
  END usb_oen
  PIN usb_rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 996.000 162.960 1000.000 ;
    END
  END usb_rst_n
  PIN user_clock1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 0.000 55.440 4.000 ;
    END
  END user_clock1
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 834.400 0.000 834.960 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 0.000 843.920 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 0.000 852.880 4.000 ;
    END
  END user_irq[2]
  PIN xtal_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 996.000 198.800 1000.000 ;
    END
  END xtal_clk
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 893.200 984.220 ;
      LAYER Metal2 ;
        RECT 8.540 995.700 18.740 996.660 ;
        RECT 19.900 995.700 54.580 996.660 ;
        RECT 55.740 995.700 90.420 996.660 ;
        RECT 91.580 995.700 126.260 996.660 ;
        RECT 127.420 995.700 162.100 996.660 ;
        RECT 163.260 995.700 197.940 996.660 ;
        RECT 199.100 995.700 233.780 996.660 ;
        RECT 234.940 995.700 269.620 996.660 ;
        RECT 270.780 995.700 305.460 996.660 ;
        RECT 306.620 995.700 341.300 996.660 ;
        RECT 342.460 995.700 377.140 996.660 ;
        RECT 378.300 995.700 412.980 996.660 ;
        RECT 414.140 995.700 448.820 996.660 ;
        RECT 449.980 995.700 484.660 996.660 ;
        RECT 485.820 995.700 520.500 996.660 ;
        RECT 521.660 995.700 556.340 996.660 ;
        RECT 557.500 995.700 592.180 996.660 ;
        RECT 593.340 995.700 628.020 996.660 ;
        RECT 629.180 995.700 663.860 996.660 ;
        RECT 665.020 995.700 699.700 996.660 ;
        RECT 700.860 995.700 735.540 996.660 ;
        RECT 736.700 995.700 771.380 996.660 ;
        RECT 772.540 995.700 807.220 996.660 ;
        RECT 808.380 995.700 843.060 996.660 ;
        RECT 844.220 995.700 878.900 996.660 ;
        RECT 880.060 995.700 894.180 996.660 ;
        RECT 8.540 4.300 894.180 995.700 ;
        RECT 8.540 3.500 45.620 4.300 ;
        RECT 46.780 3.500 54.580 4.300 ;
        RECT 55.740 3.500 63.540 4.300 ;
        RECT 64.700 3.500 72.500 4.300 ;
        RECT 73.660 3.500 81.460 4.300 ;
        RECT 82.620 3.500 90.420 4.300 ;
        RECT 91.580 3.500 99.380 4.300 ;
        RECT 100.540 3.500 108.340 4.300 ;
        RECT 109.500 3.500 117.300 4.300 ;
        RECT 118.460 3.500 126.260 4.300 ;
        RECT 127.420 3.500 135.220 4.300 ;
        RECT 136.380 3.500 144.180 4.300 ;
        RECT 145.340 3.500 153.140 4.300 ;
        RECT 154.300 3.500 162.100 4.300 ;
        RECT 163.260 3.500 171.060 4.300 ;
        RECT 172.220 3.500 180.020 4.300 ;
        RECT 181.180 3.500 188.980 4.300 ;
        RECT 190.140 3.500 197.940 4.300 ;
        RECT 199.100 3.500 206.900 4.300 ;
        RECT 208.060 3.500 215.860 4.300 ;
        RECT 217.020 3.500 224.820 4.300 ;
        RECT 225.980 3.500 233.780 4.300 ;
        RECT 234.940 3.500 242.740 4.300 ;
        RECT 243.900 3.500 251.700 4.300 ;
        RECT 252.860 3.500 260.660 4.300 ;
        RECT 261.820 3.500 269.620 4.300 ;
        RECT 270.780 3.500 278.580 4.300 ;
        RECT 279.740 3.500 287.540 4.300 ;
        RECT 288.700 3.500 296.500 4.300 ;
        RECT 297.660 3.500 305.460 4.300 ;
        RECT 306.620 3.500 314.420 4.300 ;
        RECT 315.580 3.500 323.380 4.300 ;
        RECT 324.540 3.500 332.340 4.300 ;
        RECT 333.500 3.500 341.300 4.300 ;
        RECT 342.460 3.500 350.260 4.300 ;
        RECT 351.420 3.500 359.220 4.300 ;
        RECT 360.380 3.500 368.180 4.300 ;
        RECT 369.340 3.500 377.140 4.300 ;
        RECT 378.300 3.500 386.100 4.300 ;
        RECT 387.260 3.500 395.060 4.300 ;
        RECT 396.220 3.500 404.020 4.300 ;
        RECT 405.180 3.500 412.980 4.300 ;
        RECT 414.140 3.500 421.940 4.300 ;
        RECT 423.100 3.500 430.900 4.300 ;
        RECT 432.060 3.500 439.860 4.300 ;
        RECT 441.020 3.500 448.820 4.300 ;
        RECT 449.980 3.500 457.780 4.300 ;
        RECT 458.940 3.500 466.740 4.300 ;
        RECT 467.900 3.500 475.700 4.300 ;
        RECT 476.860 3.500 484.660 4.300 ;
        RECT 485.820 3.500 493.620 4.300 ;
        RECT 494.780 3.500 502.580 4.300 ;
        RECT 503.740 3.500 511.540 4.300 ;
        RECT 512.700 3.500 520.500 4.300 ;
        RECT 521.660 3.500 529.460 4.300 ;
        RECT 530.620 3.500 538.420 4.300 ;
        RECT 539.580 3.500 547.380 4.300 ;
        RECT 548.540 3.500 556.340 4.300 ;
        RECT 557.500 3.500 565.300 4.300 ;
        RECT 566.460 3.500 574.260 4.300 ;
        RECT 575.420 3.500 583.220 4.300 ;
        RECT 584.380 3.500 592.180 4.300 ;
        RECT 593.340 3.500 601.140 4.300 ;
        RECT 602.300 3.500 610.100 4.300 ;
        RECT 611.260 3.500 619.060 4.300 ;
        RECT 620.220 3.500 628.020 4.300 ;
        RECT 629.180 3.500 636.980 4.300 ;
        RECT 638.140 3.500 645.940 4.300 ;
        RECT 647.100 3.500 654.900 4.300 ;
        RECT 656.060 3.500 663.860 4.300 ;
        RECT 665.020 3.500 672.820 4.300 ;
        RECT 673.980 3.500 681.780 4.300 ;
        RECT 682.940 3.500 690.740 4.300 ;
        RECT 691.900 3.500 699.700 4.300 ;
        RECT 700.860 3.500 708.660 4.300 ;
        RECT 709.820 3.500 717.620 4.300 ;
        RECT 718.780 3.500 726.580 4.300 ;
        RECT 727.740 3.500 735.540 4.300 ;
        RECT 736.700 3.500 744.500 4.300 ;
        RECT 745.660 3.500 753.460 4.300 ;
        RECT 754.620 3.500 762.420 4.300 ;
        RECT 763.580 3.500 771.380 4.300 ;
        RECT 772.540 3.500 780.340 4.300 ;
        RECT 781.500 3.500 789.300 4.300 ;
        RECT 790.460 3.500 798.260 4.300 ;
        RECT 799.420 3.500 807.220 4.300 ;
        RECT 808.380 3.500 816.180 4.300 ;
        RECT 817.340 3.500 825.140 4.300 ;
        RECT 826.300 3.500 834.100 4.300 ;
        RECT 835.260 3.500 843.060 4.300 ;
        RECT 844.220 3.500 852.020 4.300 ;
        RECT 853.180 3.500 894.180 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 976.380 896.000 984.060 ;
        RECT 4.300 975.220 896.000 976.380 ;
        RECT 4.000 957.340 896.000 975.220 ;
        RECT 4.300 956.180 896.000 957.340 ;
        RECT 4.000 953.980 896.000 956.180 ;
        RECT 4.000 952.820 895.700 953.980 ;
        RECT 4.000 943.900 896.000 952.820 ;
        RECT 4.000 942.740 895.700 943.900 ;
        RECT 4.000 938.300 896.000 942.740 ;
        RECT 4.300 937.140 896.000 938.300 ;
        RECT 4.000 933.820 896.000 937.140 ;
        RECT 4.000 932.660 895.700 933.820 ;
        RECT 4.000 923.740 896.000 932.660 ;
        RECT 4.000 922.580 895.700 923.740 ;
        RECT 4.000 919.260 896.000 922.580 ;
        RECT 4.300 918.100 896.000 919.260 ;
        RECT 4.000 913.660 896.000 918.100 ;
        RECT 4.000 912.500 895.700 913.660 ;
        RECT 4.000 903.580 896.000 912.500 ;
        RECT 4.000 902.420 895.700 903.580 ;
        RECT 4.000 900.220 896.000 902.420 ;
        RECT 4.300 899.060 896.000 900.220 ;
        RECT 4.000 893.500 896.000 899.060 ;
        RECT 4.000 892.340 895.700 893.500 ;
        RECT 4.000 883.420 896.000 892.340 ;
        RECT 4.000 882.260 895.700 883.420 ;
        RECT 4.000 881.180 896.000 882.260 ;
        RECT 4.300 880.020 896.000 881.180 ;
        RECT 4.000 873.340 896.000 880.020 ;
        RECT 4.000 872.180 895.700 873.340 ;
        RECT 4.000 863.260 896.000 872.180 ;
        RECT 4.000 862.140 895.700 863.260 ;
        RECT 4.300 862.100 895.700 862.140 ;
        RECT 4.300 860.980 896.000 862.100 ;
        RECT 4.000 853.180 896.000 860.980 ;
        RECT 4.000 852.020 895.700 853.180 ;
        RECT 4.000 843.100 896.000 852.020 ;
        RECT 4.300 841.940 895.700 843.100 ;
        RECT 4.000 833.020 896.000 841.940 ;
        RECT 4.000 831.860 895.700 833.020 ;
        RECT 4.000 824.060 896.000 831.860 ;
        RECT 4.300 822.940 896.000 824.060 ;
        RECT 4.300 822.900 895.700 822.940 ;
        RECT 4.000 821.780 895.700 822.900 ;
        RECT 4.000 812.860 896.000 821.780 ;
        RECT 4.000 811.700 895.700 812.860 ;
        RECT 4.000 805.020 896.000 811.700 ;
        RECT 4.300 803.860 896.000 805.020 ;
        RECT 4.000 802.780 896.000 803.860 ;
        RECT 4.000 801.620 895.700 802.780 ;
        RECT 4.000 792.700 896.000 801.620 ;
        RECT 4.000 791.540 895.700 792.700 ;
        RECT 4.000 785.980 896.000 791.540 ;
        RECT 4.300 784.820 896.000 785.980 ;
        RECT 4.000 782.620 896.000 784.820 ;
        RECT 4.000 781.460 895.700 782.620 ;
        RECT 4.000 772.540 896.000 781.460 ;
        RECT 4.000 771.380 895.700 772.540 ;
        RECT 4.000 766.940 896.000 771.380 ;
        RECT 4.300 765.780 896.000 766.940 ;
        RECT 4.000 762.460 896.000 765.780 ;
        RECT 4.000 761.300 895.700 762.460 ;
        RECT 4.000 752.380 896.000 761.300 ;
        RECT 4.000 751.220 895.700 752.380 ;
        RECT 4.000 747.900 896.000 751.220 ;
        RECT 4.300 746.740 896.000 747.900 ;
        RECT 4.000 742.300 896.000 746.740 ;
        RECT 4.000 741.140 895.700 742.300 ;
        RECT 4.000 732.220 896.000 741.140 ;
        RECT 4.000 731.060 895.700 732.220 ;
        RECT 4.000 728.860 896.000 731.060 ;
        RECT 4.300 727.700 896.000 728.860 ;
        RECT 4.000 722.140 896.000 727.700 ;
        RECT 4.000 720.980 895.700 722.140 ;
        RECT 4.000 712.060 896.000 720.980 ;
        RECT 4.000 710.900 895.700 712.060 ;
        RECT 4.000 709.820 896.000 710.900 ;
        RECT 4.300 708.660 896.000 709.820 ;
        RECT 4.000 701.980 896.000 708.660 ;
        RECT 4.000 700.820 895.700 701.980 ;
        RECT 4.000 691.900 896.000 700.820 ;
        RECT 4.000 690.780 895.700 691.900 ;
        RECT 4.300 690.740 895.700 690.780 ;
        RECT 4.300 689.620 896.000 690.740 ;
        RECT 4.000 681.820 896.000 689.620 ;
        RECT 4.000 680.660 895.700 681.820 ;
        RECT 4.000 671.740 896.000 680.660 ;
        RECT 4.300 670.580 895.700 671.740 ;
        RECT 4.000 661.660 896.000 670.580 ;
        RECT 4.000 660.500 895.700 661.660 ;
        RECT 4.000 652.700 896.000 660.500 ;
        RECT 4.300 651.580 896.000 652.700 ;
        RECT 4.300 651.540 895.700 651.580 ;
        RECT 4.000 650.420 895.700 651.540 ;
        RECT 4.000 641.500 896.000 650.420 ;
        RECT 4.000 640.340 895.700 641.500 ;
        RECT 4.000 633.660 896.000 640.340 ;
        RECT 4.300 632.500 896.000 633.660 ;
        RECT 4.000 631.420 896.000 632.500 ;
        RECT 4.000 630.260 895.700 631.420 ;
        RECT 4.000 621.340 896.000 630.260 ;
        RECT 4.000 620.180 895.700 621.340 ;
        RECT 4.000 614.620 896.000 620.180 ;
        RECT 4.300 613.460 896.000 614.620 ;
        RECT 4.000 611.260 896.000 613.460 ;
        RECT 4.000 610.100 895.700 611.260 ;
        RECT 4.000 601.180 896.000 610.100 ;
        RECT 4.000 600.020 895.700 601.180 ;
        RECT 4.000 595.580 896.000 600.020 ;
        RECT 4.300 594.420 896.000 595.580 ;
        RECT 4.000 591.100 896.000 594.420 ;
        RECT 4.000 589.940 895.700 591.100 ;
        RECT 4.000 581.020 896.000 589.940 ;
        RECT 4.000 579.860 895.700 581.020 ;
        RECT 4.000 576.540 896.000 579.860 ;
        RECT 4.300 575.380 896.000 576.540 ;
        RECT 4.000 570.940 896.000 575.380 ;
        RECT 4.000 569.780 895.700 570.940 ;
        RECT 4.000 560.860 896.000 569.780 ;
        RECT 4.000 559.700 895.700 560.860 ;
        RECT 4.000 557.500 896.000 559.700 ;
        RECT 4.300 556.340 896.000 557.500 ;
        RECT 4.000 550.780 896.000 556.340 ;
        RECT 4.000 549.620 895.700 550.780 ;
        RECT 4.000 540.700 896.000 549.620 ;
        RECT 4.000 539.540 895.700 540.700 ;
        RECT 4.000 538.460 896.000 539.540 ;
        RECT 4.300 537.300 896.000 538.460 ;
        RECT 4.000 530.620 896.000 537.300 ;
        RECT 4.000 529.460 895.700 530.620 ;
        RECT 4.000 520.540 896.000 529.460 ;
        RECT 4.000 519.420 895.700 520.540 ;
        RECT 4.300 519.380 895.700 519.420 ;
        RECT 4.300 518.260 896.000 519.380 ;
        RECT 4.000 510.460 896.000 518.260 ;
        RECT 4.000 509.300 895.700 510.460 ;
        RECT 4.000 500.380 896.000 509.300 ;
        RECT 4.300 499.220 895.700 500.380 ;
        RECT 4.000 490.300 896.000 499.220 ;
        RECT 4.000 489.140 895.700 490.300 ;
        RECT 4.000 481.340 896.000 489.140 ;
        RECT 4.300 480.220 896.000 481.340 ;
        RECT 4.300 480.180 895.700 480.220 ;
        RECT 4.000 479.060 895.700 480.180 ;
        RECT 4.000 470.140 896.000 479.060 ;
        RECT 4.000 468.980 895.700 470.140 ;
        RECT 4.000 462.300 896.000 468.980 ;
        RECT 4.300 461.140 896.000 462.300 ;
        RECT 4.000 460.060 896.000 461.140 ;
        RECT 4.000 458.900 895.700 460.060 ;
        RECT 4.000 449.980 896.000 458.900 ;
        RECT 4.000 448.820 895.700 449.980 ;
        RECT 4.000 443.260 896.000 448.820 ;
        RECT 4.300 442.100 896.000 443.260 ;
        RECT 4.000 439.900 896.000 442.100 ;
        RECT 4.000 438.740 895.700 439.900 ;
        RECT 4.000 429.820 896.000 438.740 ;
        RECT 4.000 428.660 895.700 429.820 ;
        RECT 4.000 424.220 896.000 428.660 ;
        RECT 4.300 423.060 896.000 424.220 ;
        RECT 4.000 419.740 896.000 423.060 ;
        RECT 4.000 418.580 895.700 419.740 ;
        RECT 4.000 409.660 896.000 418.580 ;
        RECT 4.000 408.500 895.700 409.660 ;
        RECT 4.000 405.180 896.000 408.500 ;
        RECT 4.300 404.020 896.000 405.180 ;
        RECT 4.000 399.580 896.000 404.020 ;
        RECT 4.000 398.420 895.700 399.580 ;
        RECT 4.000 389.500 896.000 398.420 ;
        RECT 4.000 388.340 895.700 389.500 ;
        RECT 4.000 386.140 896.000 388.340 ;
        RECT 4.300 384.980 896.000 386.140 ;
        RECT 4.000 379.420 896.000 384.980 ;
        RECT 4.000 378.260 895.700 379.420 ;
        RECT 4.000 369.340 896.000 378.260 ;
        RECT 4.000 368.180 895.700 369.340 ;
        RECT 4.000 367.100 896.000 368.180 ;
        RECT 4.300 365.940 896.000 367.100 ;
        RECT 4.000 359.260 896.000 365.940 ;
        RECT 4.000 358.100 895.700 359.260 ;
        RECT 4.000 349.180 896.000 358.100 ;
        RECT 4.000 348.060 895.700 349.180 ;
        RECT 4.300 348.020 895.700 348.060 ;
        RECT 4.300 346.900 896.000 348.020 ;
        RECT 4.000 339.100 896.000 346.900 ;
        RECT 4.000 337.940 895.700 339.100 ;
        RECT 4.000 329.020 896.000 337.940 ;
        RECT 4.300 327.860 895.700 329.020 ;
        RECT 4.000 318.940 896.000 327.860 ;
        RECT 4.000 317.780 895.700 318.940 ;
        RECT 4.000 309.980 896.000 317.780 ;
        RECT 4.300 308.860 896.000 309.980 ;
        RECT 4.300 308.820 895.700 308.860 ;
        RECT 4.000 307.700 895.700 308.820 ;
        RECT 4.000 298.780 896.000 307.700 ;
        RECT 4.000 297.620 895.700 298.780 ;
        RECT 4.000 290.940 896.000 297.620 ;
        RECT 4.300 289.780 896.000 290.940 ;
        RECT 4.000 288.700 896.000 289.780 ;
        RECT 4.000 287.540 895.700 288.700 ;
        RECT 4.000 278.620 896.000 287.540 ;
        RECT 4.000 277.460 895.700 278.620 ;
        RECT 4.000 271.900 896.000 277.460 ;
        RECT 4.300 270.740 896.000 271.900 ;
        RECT 4.000 268.540 896.000 270.740 ;
        RECT 4.000 267.380 895.700 268.540 ;
        RECT 4.000 258.460 896.000 267.380 ;
        RECT 4.000 257.300 895.700 258.460 ;
        RECT 4.000 252.860 896.000 257.300 ;
        RECT 4.300 251.700 896.000 252.860 ;
        RECT 4.000 248.380 896.000 251.700 ;
        RECT 4.000 247.220 895.700 248.380 ;
        RECT 4.000 238.300 896.000 247.220 ;
        RECT 4.000 237.140 895.700 238.300 ;
        RECT 4.000 233.820 896.000 237.140 ;
        RECT 4.300 232.660 896.000 233.820 ;
        RECT 4.000 228.220 896.000 232.660 ;
        RECT 4.000 227.060 895.700 228.220 ;
        RECT 4.000 218.140 896.000 227.060 ;
        RECT 4.000 216.980 895.700 218.140 ;
        RECT 4.000 214.780 896.000 216.980 ;
        RECT 4.300 213.620 896.000 214.780 ;
        RECT 4.000 208.060 896.000 213.620 ;
        RECT 4.000 206.900 895.700 208.060 ;
        RECT 4.000 197.980 896.000 206.900 ;
        RECT 4.000 196.820 895.700 197.980 ;
        RECT 4.000 195.740 896.000 196.820 ;
        RECT 4.300 194.580 896.000 195.740 ;
        RECT 4.000 187.900 896.000 194.580 ;
        RECT 4.000 186.740 895.700 187.900 ;
        RECT 4.000 177.820 896.000 186.740 ;
        RECT 4.000 176.700 895.700 177.820 ;
        RECT 4.300 176.660 895.700 176.700 ;
        RECT 4.300 175.540 896.000 176.660 ;
        RECT 4.000 167.740 896.000 175.540 ;
        RECT 4.000 166.580 895.700 167.740 ;
        RECT 4.000 157.660 896.000 166.580 ;
        RECT 4.300 156.500 895.700 157.660 ;
        RECT 4.000 147.580 896.000 156.500 ;
        RECT 4.000 146.420 895.700 147.580 ;
        RECT 4.000 138.620 896.000 146.420 ;
        RECT 4.300 137.500 896.000 138.620 ;
        RECT 4.300 137.460 895.700 137.500 ;
        RECT 4.000 136.340 895.700 137.460 ;
        RECT 4.000 127.420 896.000 136.340 ;
        RECT 4.000 126.260 895.700 127.420 ;
        RECT 4.000 119.580 896.000 126.260 ;
        RECT 4.300 118.420 896.000 119.580 ;
        RECT 4.000 117.340 896.000 118.420 ;
        RECT 4.000 116.180 895.700 117.340 ;
        RECT 4.000 107.260 896.000 116.180 ;
        RECT 4.000 106.100 895.700 107.260 ;
        RECT 4.000 100.540 896.000 106.100 ;
        RECT 4.300 99.380 896.000 100.540 ;
        RECT 4.000 97.180 896.000 99.380 ;
        RECT 4.000 96.020 895.700 97.180 ;
        RECT 4.000 87.100 896.000 96.020 ;
        RECT 4.000 85.940 895.700 87.100 ;
        RECT 4.000 81.500 896.000 85.940 ;
        RECT 4.300 80.340 896.000 81.500 ;
        RECT 4.000 77.020 896.000 80.340 ;
        RECT 4.000 75.860 895.700 77.020 ;
        RECT 4.000 66.940 896.000 75.860 ;
        RECT 4.000 65.780 895.700 66.940 ;
        RECT 4.000 62.460 896.000 65.780 ;
        RECT 4.300 61.300 896.000 62.460 ;
        RECT 4.000 56.860 896.000 61.300 ;
        RECT 4.000 55.700 895.700 56.860 ;
        RECT 4.000 46.780 896.000 55.700 ;
        RECT 4.000 45.620 895.700 46.780 ;
        RECT 4.000 43.420 896.000 45.620 ;
        RECT 4.300 42.260 896.000 43.420 ;
        RECT 4.000 24.380 896.000 42.260 ;
        RECT 4.300 23.220 896.000 24.380 ;
        RECT 4.000 15.540 896.000 23.220 ;
      LAYER Metal4 ;
        RECT 35.980 16.890 98.740 981.030 ;
        RECT 100.940 16.890 175.540 981.030 ;
        RECT 177.740 16.890 252.340 981.030 ;
        RECT 254.540 16.890 329.140 981.030 ;
        RECT 331.340 16.890 405.940 981.030 ;
        RECT 408.140 16.890 482.740 981.030 ;
        RECT 484.940 16.890 559.540 981.030 ;
        RECT 561.740 16.890 636.340 981.030 ;
        RECT 638.540 16.890 713.140 981.030 ;
        RECT 715.340 16.890 789.940 981.030 ;
        RECT 792.140 16.890 866.740 981.030 ;
        RECT 868.940 16.890 891.380 981.030 ;
      LAYER Metal5 ;
        RECT 119.340 17.330 883.060 763.870 ;
  END
END pinmux_top
END LIBRARY

