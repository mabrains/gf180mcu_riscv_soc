magic
tech gf180mcuD
magscale 1 10
timestamp 1700742297
<< metal1 >>
rect 8530 118750 8542 118802
rect 8594 118799 8606 118802
rect 9314 118799 9326 118802
rect 8594 118753 9326 118799
rect 8594 118750 8606 118753
rect 9314 118750 9326 118753
rect 9378 118750 9390 118802
rect 1344 118410 28560 118444
rect 1344 118358 4616 118410
rect 4668 118358 4720 118410
rect 4772 118358 4824 118410
rect 4876 118358 11420 118410
rect 11472 118358 11524 118410
rect 11576 118358 11628 118410
rect 11680 118358 18224 118410
rect 18276 118358 18328 118410
rect 18380 118358 18432 118410
rect 18484 118358 25028 118410
rect 25080 118358 25132 118410
rect 25184 118358 25236 118410
rect 25288 118358 28560 118410
rect 1344 118324 28560 118358
rect 13794 117966 13806 118018
rect 13858 117966 13870 118018
rect 14690 117966 14702 118018
rect 14754 117966 14766 118018
rect 19394 117966 19406 118018
rect 19458 117966 19470 118018
rect 20066 117966 20078 118018
rect 20130 117966 20142 118018
rect 1710 117906 1762 117918
rect 1710 117842 1762 117854
rect 3390 117906 3442 117918
rect 3390 117842 3442 117854
rect 5518 117906 5570 117918
rect 5518 117842 5570 117854
rect 6974 117906 7026 117918
rect 6974 117842 7026 117854
rect 9326 117906 9378 117918
rect 9326 117842 9378 117854
rect 10558 117906 10610 117918
rect 10558 117842 10610 117854
rect 12350 117906 12402 117918
rect 12350 117842 12402 117854
rect 13358 117906 13410 117918
rect 13358 117842 13410 117854
rect 16046 117794 16098 117806
rect 16046 117730 16098 117742
rect 16382 117794 16434 117806
rect 16382 117730 16434 117742
rect 17838 117794 17890 117806
rect 17838 117730 17890 117742
rect 20862 117794 20914 117806
rect 20862 117730 20914 117742
rect 1344 117626 28720 117660
rect 1344 117574 8018 117626
rect 8070 117574 8122 117626
rect 8174 117574 8226 117626
rect 8278 117574 14822 117626
rect 14874 117574 14926 117626
rect 14978 117574 15030 117626
rect 15082 117574 21626 117626
rect 21678 117574 21730 117626
rect 21782 117574 21834 117626
rect 21886 117574 28430 117626
rect 28482 117574 28534 117626
rect 28586 117574 28638 117626
rect 28690 117574 28720 117626
rect 1344 117540 28720 117574
rect 25678 117458 25730 117470
rect 25678 117394 25730 117406
rect 17390 117234 17442 117246
rect 25342 117234 25394 117246
rect 13794 117182 13806 117234
rect 13858 117182 13870 117234
rect 14690 117182 14702 117234
rect 14754 117182 14766 117234
rect 18386 117182 18398 117234
rect 18450 117182 18462 117234
rect 20066 117182 20078 117234
rect 20130 117182 20142 117234
rect 20738 117182 20750 117234
rect 20802 117182 20814 117234
rect 17390 117170 17442 117182
rect 25342 117170 25394 117182
rect 16046 117122 16098 117134
rect 16046 117058 16098 117070
rect 16382 117122 16434 117134
rect 16382 117058 16434 117070
rect 16830 117122 16882 117134
rect 16830 117058 16882 117070
rect 22318 117122 22370 117134
rect 22318 117058 22370 117070
rect 22654 117122 22706 117134
rect 22654 117058 22706 117070
rect 24670 117122 24722 117134
rect 24670 117058 24722 117070
rect 19518 117010 19570 117022
rect 19518 116946 19570 116958
rect 1344 116842 28560 116876
rect 1344 116790 4616 116842
rect 4668 116790 4720 116842
rect 4772 116790 4824 116842
rect 4876 116790 11420 116842
rect 11472 116790 11524 116842
rect 11576 116790 11628 116842
rect 11680 116790 18224 116842
rect 18276 116790 18328 116842
rect 18380 116790 18432 116842
rect 18484 116790 25028 116842
rect 25080 116790 25132 116842
rect 25184 116790 25236 116842
rect 25288 116790 28560 116842
rect 1344 116756 28560 116790
rect 16270 116562 16322 116574
rect 16270 116498 16322 116510
rect 18622 116562 18674 116574
rect 18622 116498 18674 116510
rect 19854 116562 19906 116574
rect 19854 116498 19906 116510
rect 13918 116450 13970 116462
rect 10770 116398 10782 116450
rect 10834 116398 10846 116450
rect 11442 116398 11454 116450
rect 11506 116398 11518 116450
rect 14914 116398 14926 116450
rect 14978 116398 14990 116450
rect 16706 116398 16718 116450
rect 16770 116398 16782 116450
rect 17714 116398 17726 116450
rect 17778 116398 17790 116450
rect 13918 116386 13970 116398
rect 13022 116226 13074 116238
rect 13022 116162 13074 116174
rect 13582 116226 13634 116238
rect 13582 116162 13634 116174
rect 20302 116226 20354 116238
rect 20302 116162 20354 116174
rect 20750 116226 20802 116238
rect 20750 116162 20802 116174
rect 1344 116058 28720 116092
rect 1344 116006 8018 116058
rect 8070 116006 8122 116058
rect 8174 116006 8226 116058
rect 8278 116006 14822 116058
rect 14874 116006 14926 116058
rect 14978 116006 15030 116058
rect 15082 116006 21626 116058
rect 21678 116006 21730 116058
rect 21782 116006 21834 116058
rect 21886 116006 28430 116058
rect 28482 116006 28534 116058
rect 28586 116006 28638 116058
rect 28690 116006 28720 116058
rect 1344 115972 28720 116006
rect 12686 115890 12738 115902
rect 12686 115826 12738 115838
rect 16158 115890 16210 115902
rect 16158 115826 16210 115838
rect 19742 115890 19794 115902
rect 19742 115826 19794 115838
rect 1710 115778 1762 115790
rect 1710 115714 1762 115726
rect 12238 115666 12290 115678
rect 11218 115614 11230 115666
rect 11282 115614 11294 115666
rect 12238 115602 12290 115614
rect 13470 115666 13522 115678
rect 14466 115614 14478 115666
rect 14530 115614 14542 115666
rect 17490 115614 17502 115666
rect 17554 115614 17566 115666
rect 18386 115614 18398 115666
rect 18450 115614 18462 115666
rect 20066 115614 20078 115666
rect 20130 115614 20142 115666
rect 20850 115614 20862 115666
rect 20914 115614 20926 115666
rect 13470 115602 13522 115614
rect 22318 115554 22370 115566
rect 22318 115490 22370 115502
rect 22654 115554 22706 115566
rect 22654 115490 22706 115502
rect 10110 115442 10162 115454
rect 10110 115378 10162 115390
rect 15598 115442 15650 115454
rect 15598 115378 15650 115390
rect 1344 115274 28560 115308
rect 1344 115222 4616 115274
rect 4668 115222 4720 115274
rect 4772 115222 4824 115274
rect 4876 115222 11420 115274
rect 11472 115222 11524 115274
rect 11576 115222 11628 115274
rect 11680 115222 18224 115274
rect 18276 115222 18328 115274
rect 18380 115222 18432 115274
rect 18484 115222 25028 115274
rect 25080 115222 25132 115274
rect 25184 115222 25236 115274
rect 25288 115222 28560 115274
rect 1344 115188 28560 115222
rect 15710 114994 15762 115006
rect 15710 114930 15762 114942
rect 19854 114994 19906 115006
rect 19854 114930 19906 114942
rect 18062 114882 18114 114894
rect 17266 114830 17278 114882
rect 17330 114830 17342 114882
rect 18062 114818 18114 114830
rect 21422 114882 21474 114894
rect 22418 114830 22430 114882
rect 22482 114830 22494 114882
rect 21422 114818 21474 114830
rect 18510 114658 18562 114670
rect 18510 114594 18562 114606
rect 23774 114658 23826 114670
rect 23774 114594 23826 114606
rect 24110 114658 24162 114670
rect 24110 114594 24162 114606
rect 1344 114490 28720 114524
rect 1344 114438 8018 114490
rect 8070 114438 8122 114490
rect 8174 114438 8226 114490
rect 8278 114438 14822 114490
rect 14874 114438 14926 114490
rect 14978 114438 15030 114490
rect 15082 114438 21626 114490
rect 21678 114438 21730 114490
rect 21782 114438 21834 114490
rect 21886 114438 28430 114490
rect 28482 114438 28534 114490
rect 28586 114438 28638 114490
rect 28690 114438 28720 114490
rect 1344 114404 28720 114438
rect 13582 114098 13634 114110
rect 11218 114046 11230 114098
rect 11282 114046 11294 114098
rect 12114 114046 12126 114098
rect 12178 114046 12190 114098
rect 14578 114046 14590 114098
rect 14642 114046 14654 114098
rect 17490 114046 17502 114098
rect 17554 114046 17566 114098
rect 18162 114046 18174 114098
rect 18226 114046 18238 114098
rect 20066 114046 20078 114098
rect 20130 114046 20142 114098
rect 20850 114046 20862 114098
rect 20914 114046 20926 114098
rect 13582 114034 13634 114046
rect 16270 113986 16322 113998
rect 16270 113922 16322 113934
rect 22654 113986 22706 113998
rect 22654 113922 22706 113934
rect 10110 113874 10162 113886
rect 10110 113810 10162 113822
rect 15710 113874 15762 113886
rect 15710 113810 15762 113822
rect 19518 113874 19570 113886
rect 19518 113810 19570 113822
rect 22094 113874 22146 113886
rect 22094 113810 22146 113822
rect 1344 113706 28560 113740
rect 1344 113654 4616 113706
rect 4668 113654 4720 113706
rect 4772 113654 4824 113706
rect 4876 113654 11420 113706
rect 11472 113654 11524 113706
rect 11576 113654 11628 113706
rect 11680 113654 18224 113706
rect 18276 113654 18328 113706
rect 18380 113654 18432 113706
rect 18484 113654 25028 113706
rect 25080 113654 25132 113706
rect 25184 113654 25236 113706
rect 25288 113654 28560 113706
rect 1344 113620 28560 113654
rect 22094 113538 22146 113550
rect 22094 113474 22146 113486
rect 16382 113426 16434 113438
rect 16382 113362 16434 113374
rect 25902 113314 25954 113326
rect 7970 113262 7982 113314
rect 8034 113262 8046 113314
rect 8866 113262 8878 113314
rect 8930 113262 8942 113314
rect 10546 113262 10558 113314
rect 10610 113262 10622 113314
rect 11218 113262 11230 113314
rect 11282 113262 11294 113314
rect 18610 113262 18622 113314
rect 18674 113262 18686 113314
rect 19282 113262 19294 113314
rect 19346 113262 19358 113314
rect 23426 113262 23438 113314
rect 23490 113262 23502 113314
rect 24098 113262 24110 113314
rect 24162 113262 24174 113314
rect 26674 113262 26686 113314
rect 26738 113262 26750 113314
rect 25902 113250 25954 113262
rect 10222 113090 10274 113102
rect 10222 113026 10274 113038
rect 12798 113090 12850 113102
rect 12798 113026 12850 113038
rect 13806 113090 13858 113102
rect 13806 113026 13858 113038
rect 20862 113090 20914 113102
rect 20862 113026 20914 113038
rect 21422 113090 21474 113102
rect 21422 113026 21474 113038
rect 28254 113090 28306 113102
rect 28254 113026 28306 113038
rect 1344 112922 28720 112956
rect 1344 112870 8018 112922
rect 8070 112870 8122 112922
rect 8174 112870 8226 112922
rect 8278 112870 14822 112922
rect 14874 112870 14926 112922
rect 14978 112870 15030 112922
rect 15082 112870 21626 112922
rect 21678 112870 21730 112922
rect 21782 112870 21834 112922
rect 21886 112870 28430 112922
rect 28482 112870 28534 112922
rect 28586 112870 28638 112922
rect 28690 112870 28720 112922
rect 1344 112836 28720 112870
rect 28254 112754 28306 112766
rect 28254 112690 28306 112702
rect 13918 112530 13970 112542
rect 16606 112530 16658 112542
rect 11442 112478 11454 112530
rect 11506 112478 11518 112530
rect 12114 112478 12126 112530
rect 12178 112478 12190 112530
rect 14690 112478 14702 112530
rect 14754 112478 14766 112530
rect 13918 112466 13970 112478
rect 16606 112466 16658 112478
rect 19182 112530 19234 112542
rect 24782 112530 24834 112542
rect 19954 112478 19966 112530
rect 20018 112478 20030 112530
rect 22530 112478 22542 112530
rect 22594 112478 22606 112530
rect 23426 112478 23438 112530
rect 23490 112478 23502 112530
rect 19182 112466 19234 112478
rect 24782 112466 24834 112478
rect 25902 112530 25954 112542
rect 26674 112478 26686 112530
rect 26738 112478 26750 112530
rect 25902 112466 25954 112478
rect 21534 112418 21586 112430
rect 21534 112354 21586 112366
rect 21870 112418 21922 112430
rect 21870 112354 21922 112366
rect 13470 112306 13522 112318
rect 13470 112242 13522 112254
rect 16046 112306 16098 112318
rect 16046 112242 16098 112254
rect 1344 112138 28560 112172
rect 1344 112086 4616 112138
rect 4668 112086 4720 112138
rect 4772 112086 4824 112138
rect 4876 112086 11420 112138
rect 11472 112086 11524 112138
rect 11576 112086 11628 112138
rect 11680 112086 18224 112138
rect 18276 112086 18328 112138
rect 18380 112086 18432 112138
rect 18484 112086 25028 112138
rect 25080 112086 25132 112138
rect 25184 112086 25236 112138
rect 25288 112086 28560 112138
rect 1344 112052 28560 112086
rect 11678 111970 11730 111982
rect 11678 111906 11730 111918
rect 16046 111970 16098 111982
rect 16046 111906 16098 111918
rect 25230 111970 25282 111982
rect 25230 111906 25282 111918
rect 28030 111858 28082 111870
rect 28030 111794 28082 111806
rect 9214 111746 9266 111758
rect 8306 111694 8318 111746
rect 8370 111694 8382 111746
rect 9214 111682 9266 111694
rect 9550 111746 9602 111758
rect 13918 111746 13970 111758
rect 18958 111746 19010 111758
rect 10322 111694 10334 111746
rect 10386 111694 10398 111746
rect 14690 111694 14702 111746
rect 14754 111694 14766 111746
rect 16706 111694 16718 111746
rect 16770 111694 16782 111746
rect 17378 111694 17390 111746
rect 17442 111694 17454 111746
rect 9550 111682 9602 111694
rect 13918 111682 13970 111694
rect 18958 111682 19010 111694
rect 19294 111746 19346 111758
rect 23202 111694 23214 111746
rect 23266 111694 23278 111746
rect 24098 111694 24110 111746
rect 24162 111694 24174 111746
rect 25778 111694 25790 111746
rect 25842 111694 25854 111746
rect 26674 111694 26686 111746
rect 26738 111694 26750 111746
rect 19294 111682 19346 111694
rect 6862 111522 6914 111534
rect 6862 111458 6914 111470
rect 12350 111522 12402 111534
rect 12350 111458 12402 111470
rect 13694 111522 13746 111534
rect 13694 111458 13746 111470
rect 1344 111354 28720 111388
rect 1344 111302 8018 111354
rect 8070 111302 8122 111354
rect 8174 111302 8226 111354
rect 8278 111302 14822 111354
rect 14874 111302 14926 111354
rect 14978 111302 15030 111354
rect 15082 111302 21626 111354
rect 21678 111302 21730 111354
rect 21782 111302 21834 111354
rect 21886 111302 28430 111354
rect 28482 111302 28534 111354
rect 28586 111302 28638 111354
rect 28690 111302 28720 111354
rect 1344 111268 28720 111302
rect 28254 111186 28306 111198
rect 28254 111122 28306 111134
rect 12686 111074 12738 111086
rect 12686 111010 12738 111022
rect 9550 110962 9602 110974
rect 12126 110962 12178 110974
rect 10322 110910 10334 110962
rect 10386 110910 10398 110962
rect 9550 110898 9602 110910
rect 12126 110898 12178 110910
rect 13918 110962 13970 110974
rect 25902 110962 25954 110974
rect 14690 110910 14702 110962
rect 14754 110910 14766 110962
rect 17490 110910 17502 110962
rect 17554 110910 17566 110962
rect 18162 110910 18174 110962
rect 18226 110910 18238 110962
rect 20066 110910 20078 110962
rect 20130 110910 20142 110962
rect 20738 110910 20750 110962
rect 20802 110910 20814 110962
rect 26674 110910 26686 110962
rect 26738 110910 26750 110962
rect 13918 110898 13970 110910
rect 25902 110898 25954 110910
rect 13134 110850 13186 110862
rect 13134 110786 13186 110798
rect 13582 110850 13634 110862
rect 13582 110786 13634 110798
rect 16606 110850 16658 110862
rect 16606 110786 16658 110798
rect 22318 110850 22370 110862
rect 22318 110786 22370 110798
rect 22654 110850 22706 110862
rect 22654 110786 22706 110798
rect 11678 110738 11730 110750
rect 11678 110674 11730 110686
rect 16046 110738 16098 110750
rect 16046 110674 16098 110686
rect 19518 110738 19570 110750
rect 19518 110674 19570 110686
rect 1344 110570 28560 110604
rect 1344 110518 4616 110570
rect 4668 110518 4720 110570
rect 4772 110518 4824 110570
rect 4876 110518 11420 110570
rect 11472 110518 11524 110570
rect 11576 110518 11628 110570
rect 11680 110518 18224 110570
rect 18276 110518 18328 110570
rect 18380 110518 18432 110570
rect 18484 110518 25028 110570
rect 25080 110518 25132 110570
rect 25184 110518 25236 110570
rect 25288 110518 28560 110570
rect 1344 110484 28560 110518
rect 11006 110402 11058 110414
rect 16046 110402 16098 110414
rect 12002 110350 12014 110402
rect 12066 110350 12078 110402
rect 11006 110338 11058 110350
rect 16046 110338 16098 110350
rect 11454 110290 11506 110302
rect 11454 110226 11506 110238
rect 16606 110290 16658 110302
rect 16606 110226 16658 110238
rect 19854 110290 19906 110302
rect 19854 110226 19906 110238
rect 28254 110290 28306 110302
rect 28254 110226 28306 110238
rect 8878 110178 8930 110190
rect 11678 110178 11730 110190
rect 9650 110126 9662 110178
rect 9714 110126 9726 110178
rect 8878 110114 8930 110126
rect 11678 110114 11730 110126
rect 12686 110178 12738 110190
rect 12686 110114 12738 110126
rect 12910 110178 12962 110190
rect 12910 110114 12962 110126
rect 13918 110178 13970 110190
rect 25902 110178 25954 110190
rect 14690 110126 14702 110178
rect 14754 110126 14766 110178
rect 21410 110126 21422 110178
rect 21474 110126 21486 110178
rect 22306 110126 22318 110178
rect 22370 110126 22382 110178
rect 26674 110126 26686 110178
rect 26738 110126 26750 110178
rect 13918 110114 13970 110126
rect 25902 110114 25954 110126
rect 13470 110066 13522 110078
rect 13470 110002 13522 110014
rect 23662 110066 23714 110078
rect 23662 110002 23714 110014
rect 13582 109954 13634 109966
rect 12338 109902 12350 109954
rect 12402 109902 12414 109954
rect 13582 109890 13634 109902
rect 19406 109954 19458 109966
rect 19406 109890 19458 109902
rect 20638 109954 20690 109966
rect 20638 109890 20690 109902
rect 23998 109954 24050 109966
rect 23998 109890 24050 109902
rect 1344 109786 28720 109820
rect 1344 109734 8018 109786
rect 8070 109734 8122 109786
rect 8174 109734 8226 109786
rect 8278 109734 14822 109786
rect 14874 109734 14926 109786
rect 14978 109734 15030 109786
rect 15082 109734 21626 109786
rect 21678 109734 21730 109786
rect 21782 109734 21834 109786
rect 21886 109734 28430 109786
rect 28482 109734 28534 109786
rect 28586 109734 28638 109786
rect 28690 109734 28720 109786
rect 1344 109700 28720 109734
rect 28254 109618 28306 109630
rect 21410 109566 21422 109618
rect 21474 109566 21486 109618
rect 28254 109554 28306 109566
rect 12114 109454 12126 109506
rect 12178 109454 12190 109506
rect 14242 109454 14254 109506
rect 14306 109454 14318 109506
rect 20514 109454 20526 109506
rect 20578 109454 20590 109506
rect 15374 109394 15426 109406
rect 10770 109342 10782 109394
rect 10834 109342 10846 109394
rect 11666 109342 11678 109394
rect 11730 109342 11742 109394
rect 12338 109342 12350 109394
rect 12402 109342 12414 109394
rect 13570 109342 13582 109394
rect 13634 109342 13646 109394
rect 15374 109330 15426 109342
rect 15822 109394 15874 109406
rect 15822 109330 15874 109342
rect 16718 109394 16770 109406
rect 16718 109330 16770 109342
rect 19518 109394 19570 109406
rect 25902 109394 25954 109406
rect 21298 109342 21310 109394
rect 21362 109342 21374 109394
rect 26674 109342 26686 109394
rect 26738 109342 26750 109394
rect 19518 109330 19570 109342
rect 25902 109330 25954 109342
rect 16158 109282 16210 109294
rect 13010 109230 13022 109282
rect 13074 109230 13086 109282
rect 16158 109218 16210 109230
rect 18174 109282 18226 109294
rect 18174 109218 18226 109230
rect 18958 109282 19010 109294
rect 18958 109218 19010 109230
rect 19966 109282 20018 109294
rect 19966 109218 20018 109230
rect 22430 109282 22482 109294
rect 22430 109218 22482 109230
rect 9662 109170 9714 109182
rect 9662 109106 9714 109118
rect 1344 109002 28560 109036
rect 1344 108950 4616 109002
rect 4668 108950 4720 109002
rect 4772 108950 4824 109002
rect 4876 108950 11420 109002
rect 11472 108950 11524 109002
rect 11576 108950 11628 109002
rect 11680 108950 18224 109002
rect 18276 108950 18328 109002
rect 18380 108950 18432 109002
rect 18484 108950 25028 109002
rect 25080 108950 25132 109002
rect 25184 108950 25236 109002
rect 25288 108950 28560 109002
rect 1344 108916 28560 108950
rect 9662 108834 9714 108846
rect 16942 108834 16994 108846
rect 12786 108782 12798 108834
rect 12850 108782 12862 108834
rect 14242 108782 14254 108834
rect 14306 108782 14318 108834
rect 9662 108770 9714 108782
rect 16942 108770 16994 108782
rect 21310 108834 21362 108846
rect 21310 108770 21362 108782
rect 15038 108722 15090 108734
rect 8978 108670 8990 108722
rect 9042 108670 9054 108722
rect 14018 108670 14030 108722
rect 14082 108670 14094 108722
rect 15038 108658 15090 108670
rect 17390 108722 17442 108734
rect 17390 108658 17442 108670
rect 18734 108722 18786 108734
rect 20402 108670 20414 108722
rect 20466 108670 20478 108722
rect 18734 108658 18786 108670
rect 12574 108610 12626 108622
rect 14926 108610 14978 108622
rect 18510 108610 18562 108622
rect 22318 108610 22370 108622
rect 24894 108610 24946 108622
rect 10770 108558 10782 108610
rect 10834 108558 10846 108610
rect 11666 108558 11678 108610
rect 11730 108558 11742 108610
rect 12786 108558 12798 108610
rect 12850 108558 12862 108610
rect 13682 108558 13694 108610
rect 13746 108558 13758 108610
rect 16930 108558 16942 108610
rect 16994 108558 17006 108610
rect 17826 108558 17838 108610
rect 17890 108558 17902 108610
rect 19842 108558 19854 108610
rect 19906 108558 19918 108610
rect 23090 108558 23102 108610
rect 23154 108558 23166 108610
rect 25666 108558 25678 108610
rect 25730 108558 25742 108610
rect 12574 108546 12626 108558
rect 14926 108546 14978 108558
rect 18510 108546 18562 108558
rect 22318 108546 22370 108558
rect 24894 108546 24946 108558
rect 9214 108498 9266 108510
rect 9214 108434 9266 108446
rect 16046 108498 16098 108510
rect 16046 108434 16098 108446
rect 16606 108498 16658 108510
rect 19182 108498 19234 108510
rect 18162 108446 18174 108498
rect 18226 108446 18238 108498
rect 16606 108434 16658 108446
rect 19182 108434 19234 108446
rect 20750 108498 20802 108510
rect 20750 108434 20802 108446
rect 21422 108498 21474 108510
rect 21422 108434 21474 108446
rect 15710 108386 15762 108398
rect 15710 108322 15762 108334
rect 17278 108386 17330 108398
rect 17278 108322 17330 108334
rect 17502 108386 17554 108398
rect 17502 108322 17554 108334
rect 19070 108386 19122 108398
rect 19070 108322 19122 108334
rect 21870 108386 21922 108398
rect 21870 108322 21922 108334
rect 24670 108386 24722 108398
rect 24670 108322 24722 108334
rect 27246 108386 27298 108398
rect 27246 108322 27298 108334
rect 1344 108218 28720 108252
rect 1344 108166 8018 108218
rect 8070 108166 8122 108218
rect 8174 108166 8226 108218
rect 8278 108166 14822 108218
rect 14874 108166 14926 108218
rect 14978 108166 15030 108218
rect 15082 108166 21626 108218
rect 21678 108166 21730 108218
rect 21782 108166 21834 108218
rect 21886 108166 28430 108218
rect 28482 108166 28534 108218
rect 28586 108166 28638 108218
rect 28690 108166 28720 108218
rect 1344 108132 28720 108166
rect 14478 108050 14530 108062
rect 14478 107986 14530 107998
rect 20526 108050 20578 108062
rect 20526 107986 20578 107998
rect 21086 108050 21138 108062
rect 21086 107986 21138 107998
rect 28254 108050 28306 108062
rect 28254 107986 28306 107998
rect 13134 107938 13186 107950
rect 13134 107874 13186 107886
rect 17390 107938 17442 107950
rect 17390 107874 17442 107886
rect 12126 107826 12178 107838
rect 10770 107774 10782 107826
rect 10834 107774 10846 107826
rect 11666 107774 11678 107826
rect 11730 107774 11742 107826
rect 12126 107762 12178 107774
rect 12350 107826 12402 107838
rect 17726 107826 17778 107838
rect 12674 107774 12686 107826
rect 12738 107774 12750 107826
rect 13570 107774 13582 107826
rect 13634 107774 13646 107826
rect 16034 107774 16046 107826
rect 16098 107774 16110 107826
rect 16706 107774 16718 107826
rect 16770 107774 16782 107826
rect 12350 107762 12402 107774
rect 17726 107762 17778 107774
rect 18174 107826 18226 107838
rect 20750 107826 20802 107838
rect 25902 107826 25954 107838
rect 19170 107774 19182 107826
rect 19234 107774 19246 107826
rect 22306 107774 22318 107826
rect 22370 107774 22382 107826
rect 23090 107774 23102 107826
rect 23154 107774 23166 107826
rect 26674 107774 26686 107826
rect 26738 107774 26750 107826
rect 18174 107762 18226 107774
rect 20750 107762 20802 107774
rect 25902 107762 25954 107774
rect 8990 107714 9042 107726
rect 8990 107650 9042 107662
rect 12238 107714 12290 107726
rect 21534 107714 21586 107726
rect 14018 107662 14030 107714
rect 14082 107662 14094 107714
rect 12238 107650 12290 107662
rect 21534 107650 21586 107662
rect 9662 107602 9714 107614
rect 9662 107538 9714 107550
rect 24334 107602 24386 107614
rect 24334 107538 24386 107550
rect 1344 107434 28560 107468
rect 1344 107382 4616 107434
rect 4668 107382 4720 107434
rect 4772 107382 4824 107434
rect 4876 107382 11420 107434
rect 11472 107382 11524 107434
rect 11576 107382 11628 107434
rect 11680 107382 18224 107434
rect 18276 107382 18328 107434
rect 18380 107382 18432 107434
rect 18484 107382 25028 107434
rect 25080 107382 25132 107434
rect 25184 107382 25236 107434
rect 25288 107382 28560 107434
rect 1344 107348 28560 107382
rect 21534 107266 21586 107278
rect 8530 107214 8542 107266
rect 8594 107263 8606 107266
rect 8978 107263 8990 107266
rect 8594 107217 8990 107263
rect 8594 107214 8606 107217
rect 8978 107214 8990 107217
rect 9042 107263 9054 107266
rect 9426 107263 9438 107266
rect 9042 107217 9438 107263
rect 9042 107214 9054 107217
rect 9426 107214 9438 107217
rect 9490 107263 9502 107266
rect 9874 107263 9886 107266
rect 9490 107217 9886 107263
rect 9490 107214 9502 107217
rect 9874 107214 9886 107217
rect 9938 107214 9950 107266
rect 14914 107214 14926 107266
rect 14978 107214 14990 107266
rect 21534 107202 21586 107214
rect 9438 107154 9490 107166
rect 9438 107090 9490 107102
rect 9886 107154 9938 107166
rect 20078 107154 20130 107166
rect 14242 107102 14254 107154
rect 14306 107102 14318 107154
rect 9886 107090 9938 107102
rect 20078 107090 20130 107102
rect 25006 107154 25058 107166
rect 25006 107090 25058 107102
rect 28254 107154 28306 107166
rect 28254 107090 28306 107102
rect 12462 107042 12514 107054
rect 11442 106990 11454 107042
rect 11506 106990 11518 107042
rect 12462 106978 12514 106990
rect 13582 107042 13634 107054
rect 21310 107042 21362 107054
rect 14578 106990 14590 107042
rect 14642 106990 14654 107042
rect 15474 106990 15486 107042
rect 15538 106990 15550 107042
rect 16146 106990 16158 107042
rect 16210 106990 16222 107042
rect 18162 106990 18174 107042
rect 18226 106990 18238 107042
rect 19170 106990 19182 107042
rect 19234 106990 19246 107042
rect 13582 106978 13634 106990
rect 21310 106978 21362 106990
rect 22318 107042 22370 107054
rect 25902 107042 25954 107054
rect 23090 106990 23102 107042
rect 23154 106990 23166 107042
rect 26674 106990 26686 107042
rect 26738 106990 26750 107042
rect 22318 106978 22370 106990
rect 25902 106978 25954 106990
rect 13470 106930 13522 106942
rect 13470 106866 13522 106878
rect 7534 106818 7586 106830
rect 7534 106754 7586 106766
rect 8094 106818 8146 106830
rect 8094 106754 8146 106766
rect 8542 106818 8594 106830
rect 8542 106754 8594 106766
rect 9102 106818 9154 106830
rect 9102 106754 9154 106766
rect 10110 106818 10162 106830
rect 10110 106754 10162 106766
rect 13022 106818 13074 106830
rect 13022 106754 13074 106766
rect 17726 106818 17778 106830
rect 24670 106818 24722 106830
rect 21858 106766 21870 106818
rect 21922 106766 21934 106818
rect 17726 106754 17778 106766
rect 24670 106754 24722 106766
rect 1344 106650 28720 106684
rect 1344 106598 8018 106650
rect 8070 106598 8122 106650
rect 8174 106598 8226 106650
rect 8278 106598 14822 106650
rect 14874 106598 14926 106650
rect 14978 106598 15030 106650
rect 15082 106598 21626 106650
rect 21678 106598 21730 106650
rect 21782 106598 21834 106650
rect 21886 106598 28430 106650
rect 28482 106598 28534 106650
rect 28586 106598 28638 106650
rect 28690 106598 28720 106650
rect 1344 106564 28720 106598
rect 9886 106482 9938 106494
rect 19854 106482 19906 106494
rect 16818 106430 16830 106482
rect 16882 106430 16894 106482
rect 9886 106418 9938 106430
rect 19854 106418 19906 106430
rect 21310 106482 21362 106494
rect 28254 106482 28306 106494
rect 22754 106430 22766 106482
rect 22818 106430 22830 106482
rect 21310 106418 21362 106430
rect 28254 106418 28306 106430
rect 3166 106370 3218 106382
rect 3166 106306 3218 106318
rect 9102 106370 9154 106382
rect 9102 106306 9154 106318
rect 9774 106370 9826 106382
rect 21858 106318 21870 106370
rect 21922 106318 21934 106370
rect 9774 106306 9826 106318
rect 8094 106258 8146 106270
rect 15934 106258 15986 106270
rect 6066 106206 6078 106258
rect 6130 106206 6142 106258
rect 15474 106206 15486 106258
rect 15538 106206 15550 106258
rect 8094 106194 8146 106206
rect 15934 106194 15986 106206
rect 17502 106258 17554 106270
rect 25342 106258 25394 106270
rect 18274 106206 18286 106258
rect 18338 106206 18350 106258
rect 22194 106206 22206 106258
rect 22258 106206 22270 106258
rect 17502 106194 17554 106206
rect 25342 106194 25394 106206
rect 25902 106258 25954 106270
rect 26674 106206 26686 106258
rect 26738 106206 26750 106258
rect 25902 106194 25954 106206
rect 3278 106146 3330 106158
rect 3278 106082 3330 106094
rect 3838 106146 3890 106158
rect 3838 106082 3890 106094
rect 4734 106146 4786 106158
rect 4734 106082 4786 106094
rect 5294 106146 5346 106158
rect 5294 106082 5346 106094
rect 5742 106146 5794 106158
rect 5742 106082 5794 106094
rect 6302 106146 6354 106158
rect 6302 106082 6354 106094
rect 7310 106146 7362 106158
rect 7310 106082 7362 106094
rect 7646 106146 7698 106158
rect 7646 106082 7698 106094
rect 8542 106146 8594 106158
rect 16270 106146 16322 106158
rect 11218 106094 11230 106146
rect 11282 106094 11294 106146
rect 8542 106082 8594 106094
rect 16270 106082 16322 106094
rect 20190 106146 20242 106158
rect 20190 106082 20242 106094
rect 23326 106146 23378 106158
rect 23326 106082 23378 106094
rect 23774 106146 23826 106158
rect 23774 106082 23826 106094
rect 3390 106034 3442 106046
rect 3390 105970 3442 105982
rect 6414 106034 6466 106046
rect 15822 106034 15874 106046
rect 7298 105982 7310 106034
rect 7362 106031 7374 106034
rect 8306 106031 8318 106034
rect 7362 105985 8318 106031
rect 7362 105982 7374 105985
rect 8306 105982 8318 105985
rect 8370 105982 8382 106034
rect 8530 105982 8542 106034
rect 8594 106031 8606 106034
rect 9090 106031 9102 106034
rect 8594 105985 9102 106031
rect 8594 105982 8606 105985
rect 9090 105982 9102 105985
rect 9154 105982 9166 106034
rect 6414 105970 6466 105982
rect 15822 105970 15874 105982
rect 16494 106034 16546 106046
rect 16494 105970 16546 105982
rect 23438 106034 23490 106046
rect 23438 105970 23490 105982
rect 23998 106034 24050 106046
rect 24322 105982 24334 106034
rect 24386 105982 24398 106034
rect 23998 105970 24050 105982
rect 1344 105866 28560 105900
rect 1344 105814 4616 105866
rect 4668 105814 4720 105866
rect 4772 105814 4824 105866
rect 4876 105814 11420 105866
rect 11472 105814 11524 105866
rect 11576 105814 11628 105866
rect 11680 105814 18224 105866
rect 18276 105814 18328 105866
rect 18380 105814 18432 105866
rect 18484 105814 25028 105866
rect 25080 105814 25132 105866
rect 25184 105814 25236 105866
rect 25288 105814 28560 105866
rect 1344 105780 28560 105814
rect 9662 105698 9714 105710
rect 22542 105698 22594 105710
rect 19954 105646 19966 105698
rect 20018 105646 20030 105698
rect 9662 105634 9714 105646
rect 22542 105634 22594 105646
rect 22206 105586 22258 105598
rect 1698 105534 1710 105586
rect 1762 105534 1774 105586
rect 3826 105534 3838 105586
rect 3890 105534 3902 105586
rect 5618 105534 5630 105586
rect 5682 105534 5694 105586
rect 7746 105534 7758 105586
rect 7810 105534 7822 105586
rect 16370 105534 16382 105586
rect 16434 105534 16446 105586
rect 22206 105522 22258 105534
rect 26238 105586 26290 105598
rect 26238 105522 26290 105534
rect 12686 105474 12738 105486
rect 4498 105422 4510 105474
rect 4562 105422 4574 105474
rect 8530 105422 8542 105474
rect 8594 105422 8606 105474
rect 10770 105422 10782 105474
rect 10834 105422 10846 105474
rect 11666 105422 11678 105474
rect 11730 105422 11742 105474
rect 12686 105410 12738 105422
rect 13806 105474 13858 105486
rect 13806 105410 13858 105422
rect 14030 105474 14082 105486
rect 20302 105474 20354 105486
rect 14578 105422 14590 105474
rect 14642 105422 14654 105474
rect 14030 105410 14082 105422
rect 20302 105410 20354 105422
rect 20526 105474 20578 105486
rect 25006 105474 25058 105486
rect 22530 105422 22542 105474
rect 22594 105422 22606 105474
rect 23202 105422 23214 105474
rect 23266 105422 23278 105474
rect 24434 105422 24446 105474
rect 24498 105422 24510 105474
rect 20526 105410 20578 105422
rect 25006 105410 25058 105422
rect 8878 105362 8930 105374
rect 8878 105298 8930 105310
rect 21310 105362 21362 105374
rect 21310 105298 21362 105310
rect 21534 105362 21586 105374
rect 21534 105298 21586 105310
rect 23886 105362 23938 105374
rect 23886 105298 23938 105310
rect 5182 105250 5234 105262
rect 5182 105186 5234 105198
rect 8990 105250 9042 105262
rect 8990 105186 9042 105198
rect 12462 105250 12514 105262
rect 12462 105186 12514 105198
rect 12798 105250 12850 105262
rect 12798 105186 12850 105198
rect 12910 105250 12962 105262
rect 21422 105250 21474 105262
rect 13458 105198 13470 105250
rect 13522 105198 13534 105250
rect 12910 105186 12962 105198
rect 21422 105186 21474 105198
rect 25342 105250 25394 105262
rect 25342 105186 25394 105198
rect 25678 105250 25730 105262
rect 25678 105186 25730 105198
rect 26686 105250 26738 105262
rect 26686 105186 26738 105198
rect 1344 105082 28720 105116
rect 1344 105030 8018 105082
rect 8070 105030 8122 105082
rect 8174 105030 8226 105082
rect 8278 105030 14822 105082
rect 14874 105030 14926 105082
rect 14978 105030 15030 105082
rect 15082 105030 21626 105082
rect 21678 105030 21730 105082
rect 21782 105030 21834 105082
rect 21886 105030 28430 105082
rect 28482 105030 28534 105082
rect 28586 105030 28638 105082
rect 28690 105030 28720 105082
rect 1344 104996 28720 105030
rect 3838 104914 3890 104926
rect 3838 104850 3890 104862
rect 3950 104914 4002 104926
rect 3950 104850 4002 104862
rect 4062 104914 4114 104926
rect 4062 104850 4114 104862
rect 6750 104914 6802 104926
rect 6750 104850 6802 104862
rect 7982 104914 8034 104926
rect 7982 104850 8034 104862
rect 8094 104914 8146 104926
rect 8094 104850 8146 104862
rect 28030 104914 28082 104926
rect 28030 104850 28082 104862
rect 4286 104802 4338 104814
rect 8318 104802 8370 104814
rect 10446 104802 10498 104814
rect 7298 104750 7310 104802
rect 7362 104799 7374 104802
rect 7522 104799 7534 104802
rect 7362 104753 7534 104799
rect 7362 104750 7374 104753
rect 7522 104750 7534 104753
rect 7586 104750 7598 104802
rect 8978 104750 8990 104802
rect 9042 104750 9054 104802
rect 4286 104738 4338 104750
rect 8318 104738 8370 104750
rect 10446 104738 10498 104750
rect 19070 104802 19122 104814
rect 19070 104738 19122 104750
rect 25230 104802 25282 104814
rect 25230 104738 25282 104750
rect 3726 104690 3778 104702
rect 3726 104626 3778 104638
rect 5182 104690 5234 104702
rect 5182 104626 5234 104638
rect 6526 104690 6578 104702
rect 6526 104626 6578 104638
rect 6638 104690 6690 104702
rect 6638 104626 6690 104638
rect 6862 104690 6914 104702
rect 7870 104690 7922 104702
rect 7074 104638 7086 104690
rect 7138 104638 7150 104690
rect 7634 104638 7646 104690
rect 7698 104638 7710 104690
rect 6862 104626 6914 104638
rect 7870 104626 7922 104638
rect 8654 104690 8706 104702
rect 25678 104690 25730 104702
rect 9650 104638 9662 104690
rect 9714 104638 9726 104690
rect 11218 104638 11230 104690
rect 11282 104638 11294 104690
rect 11778 104638 11790 104690
rect 11842 104638 11854 104690
rect 18162 104638 18174 104690
rect 18226 104638 18238 104690
rect 19394 104638 19406 104690
rect 19458 104638 19470 104690
rect 26674 104638 26686 104690
rect 26738 104638 26750 104690
rect 8654 104626 8706 104638
rect 25678 104626 25730 104638
rect 2830 104578 2882 104590
rect 2830 104514 2882 104526
rect 3278 104578 3330 104590
rect 3278 104514 3330 104526
rect 4734 104578 4786 104590
rect 4734 104514 4786 104526
rect 5630 104578 5682 104590
rect 5630 104514 5682 104526
rect 6078 104578 6130 104590
rect 17614 104578 17666 104590
rect 15474 104526 15486 104578
rect 15538 104526 15550 104578
rect 18498 104526 18510 104578
rect 18562 104526 18574 104578
rect 22194 104526 22206 104578
rect 22258 104526 22270 104578
rect 6078 104514 6130 104526
rect 17614 104514 17666 104526
rect 2930 104414 2942 104466
rect 2994 104463 3006 104466
rect 3378 104463 3390 104466
rect 2994 104417 3390 104463
rect 2994 104414 3006 104417
rect 3378 104414 3390 104417
rect 3442 104414 3454 104466
rect 1344 104298 28560 104332
rect 1344 104246 4616 104298
rect 4668 104246 4720 104298
rect 4772 104246 4824 104298
rect 4876 104246 11420 104298
rect 11472 104246 11524 104298
rect 11576 104246 11628 104298
rect 11680 104246 18224 104298
rect 18276 104246 18328 104298
rect 18380 104246 18432 104298
rect 18484 104246 25028 104298
rect 25080 104246 25132 104298
rect 25184 104246 25236 104298
rect 25288 104246 28560 104298
rect 1344 104212 28560 104246
rect 14702 104130 14754 104142
rect 14702 104066 14754 104078
rect 27582 104130 27634 104142
rect 27582 104066 27634 104078
rect 11230 104018 11282 104030
rect 23662 104018 23714 104030
rect 26014 104018 26066 104030
rect 1698 103966 1710 104018
rect 1762 103966 1774 104018
rect 5842 103966 5854 104018
rect 5906 103966 5918 104018
rect 12338 103966 12350 104018
rect 12402 103966 12414 104018
rect 13570 103966 13582 104018
rect 13634 103966 13646 104018
rect 24658 103966 24670 104018
rect 24722 103966 24734 104018
rect 11230 103954 11282 103966
rect 23662 103954 23714 103966
rect 26014 103954 26066 103966
rect 9886 103906 9938 103918
rect 12126 103906 12178 103918
rect 24446 103906 24498 103918
rect 27694 103906 27746 103918
rect 4498 103854 4510 103906
rect 4562 103854 4574 103906
rect 8642 103854 8654 103906
rect 8706 103854 8718 103906
rect 10658 103854 10670 103906
rect 10722 103854 10734 103906
rect 10882 103854 10894 103906
rect 10946 103854 10958 103906
rect 12226 103854 12238 103906
rect 12290 103854 12302 103906
rect 13906 103854 13918 103906
rect 13970 103854 13982 103906
rect 15026 103854 15038 103906
rect 15090 103854 15102 103906
rect 15474 103854 15486 103906
rect 15538 103854 15550 103906
rect 21410 103854 21422 103906
rect 21474 103854 21486 103906
rect 22306 103854 22318 103906
rect 22370 103854 22382 103906
rect 24882 103854 24894 103906
rect 24946 103854 24958 103906
rect 9886 103842 9938 103854
rect 12126 103842 12178 103854
rect 24446 103842 24498 103854
rect 27694 103842 27746 103854
rect 9326 103794 9378 103806
rect 3826 103742 3838 103794
rect 3890 103742 3902 103794
rect 7970 103742 7982 103794
rect 8034 103742 8046 103794
rect 9326 103730 9378 103742
rect 9662 103794 9714 103806
rect 9662 103730 9714 103742
rect 11118 103794 11170 103806
rect 26910 103794 26962 103806
rect 13794 103742 13806 103794
rect 13858 103742 13870 103794
rect 17490 103742 17502 103794
rect 17554 103742 17566 103794
rect 11118 103730 11170 103742
rect 26910 103730 26962 103742
rect 5070 103682 5122 103694
rect 5070 103618 5122 103630
rect 9214 103682 9266 103694
rect 11342 103682 11394 103694
rect 10210 103630 10222 103682
rect 10274 103630 10286 103682
rect 9214 103618 9266 103630
rect 11342 103618 11394 103630
rect 13022 103682 13074 103694
rect 13022 103618 13074 103630
rect 14142 103682 14194 103694
rect 14142 103618 14194 103630
rect 14366 103682 14418 103694
rect 14366 103618 14418 103630
rect 14814 103682 14866 103694
rect 14814 103618 14866 103630
rect 24110 103682 24162 103694
rect 24110 103618 24162 103630
rect 1344 103514 28720 103548
rect 1344 103462 8018 103514
rect 8070 103462 8122 103514
rect 8174 103462 8226 103514
rect 8278 103462 14822 103514
rect 14874 103462 14926 103514
rect 14978 103462 15030 103514
rect 15082 103462 21626 103514
rect 21678 103462 21730 103514
rect 21782 103462 21834 103514
rect 21886 103462 28430 103514
rect 28482 103462 28534 103514
rect 28586 103462 28638 103514
rect 28690 103462 28720 103514
rect 1344 103428 28720 103462
rect 4286 103346 4338 103358
rect 4286 103282 4338 103294
rect 5294 103346 5346 103358
rect 5294 103282 5346 103294
rect 6974 103346 7026 103358
rect 6974 103282 7026 103294
rect 7086 103346 7138 103358
rect 7086 103282 7138 103294
rect 7870 103346 7922 103358
rect 7870 103282 7922 103294
rect 8990 103346 9042 103358
rect 8990 103282 9042 103294
rect 9550 103346 9602 103358
rect 9550 103282 9602 103294
rect 17502 103346 17554 103358
rect 17502 103282 17554 103294
rect 18398 103346 18450 103358
rect 18398 103282 18450 103294
rect 22878 103346 22930 103358
rect 22878 103282 22930 103294
rect 23326 103346 23378 103358
rect 23650 103294 23662 103346
rect 23714 103294 23726 103346
rect 23986 103294 23998 103346
rect 24050 103294 24062 103346
rect 23326 103282 23378 103294
rect 3502 103234 3554 103246
rect 3502 103170 3554 103182
rect 3726 103234 3778 103246
rect 3726 103170 3778 103182
rect 4062 103234 4114 103246
rect 4062 103170 4114 103182
rect 7198 103234 7250 103246
rect 7198 103170 7250 103182
rect 7758 103234 7810 103246
rect 7758 103170 7810 103182
rect 18286 103234 18338 103246
rect 18286 103170 18338 103182
rect 2606 103122 2658 103134
rect 2606 103058 2658 103070
rect 3278 103122 3330 103134
rect 3278 103058 3330 103070
rect 3950 103122 4002 103134
rect 3950 103058 4002 103070
rect 4398 103122 4450 103134
rect 4398 103058 4450 103070
rect 7646 103122 7698 103134
rect 7646 103058 7698 103070
rect 8094 103122 8146 103134
rect 8094 103058 8146 103070
rect 8318 103122 8370 103134
rect 8318 103058 8370 103070
rect 8766 103122 8818 103134
rect 10222 103122 10274 103134
rect 9762 103070 9774 103122
rect 9826 103070 9838 103122
rect 9986 103070 9998 103122
rect 10050 103070 10062 103122
rect 8766 103058 8818 103070
rect 10222 103058 10274 103070
rect 10670 103122 10722 103134
rect 10670 103058 10722 103070
rect 10894 103122 10946 103134
rect 12574 103122 12626 103134
rect 17278 103122 17330 103134
rect 11778 103070 11790 103122
rect 11842 103070 11854 103122
rect 12114 103070 12126 103122
rect 12178 103070 12190 103122
rect 13122 103070 13134 103122
rect 13186 103070 13198 103122
rect 14018 103070 14030 103122
rect 14082 103070 14094 103122
rect 14914 103070 14926 103122
rect 14978 103070 14990 103122
rect 16146 103070 16158 103122
rect 16210 103070 16222 103122
rect 10894 103058 10946 103070
rect 12574 103058 12626 103070
rect 17278 103058 17330 103070
rect 17726 103122 17778 103134
rect 17726 103058 17778 103070
rect 17950 103122 18002 103134
rect 22206 103122 22258 103134
rect 18834 103070 18846 103122
rect 18898 103070 18910 103122
rect 24210 103070 24222 103122
rect 24274 103070 24286 103122
rect 17950 103058 18002 103070
rect 22206 103058 22258 103070
rect 2158 103010 2210 103022
rect 2158 102946 2210 102958
rect 2942 103010 2994 103022
rect 2942 102946 2994 102958
rect 5630 103010 5682 103022
rect 5630 102946 5682 102958
rect 6078 103010 6130 103022
rect 6078 102946 6130 102958
rect 6526 103010 6578 103022
rect 6526 102946 6578 102958
rect 8878 103010 8930 103022
rect 8878 102946 8930 102958
rect 10782 103010 10834 103022
rect 21982 103010 22034 103022
rect 12226 102958 12238 103010
rect 12290 102958 12302 103010
rect 14242 102958 14254 103010
rect 14306 102958 14318 103010
rect 19506 102958 19518 103010
rect 19570 102958 19582 103010
rect 21634 102958 21646 103010
rect 21698 102958 21710 103010
rect 10782 102946 10834 102958
rect 21982 102946 22034 102958
rect 22542 103010 22594 103022
rect 22542 102946 22594 102958
rect 22990 103010 23042 103022
rect 22990 102946 23042 102958
rect 25342 103010 25394 103022
rect 25342 102946 25394 102958
rect 9438 102898 9490 102910
rect 5058 102846 5070 102898
rect 5122 102895 5134 102898
rect 6066 102895 6078 102898
rect 5122 102849 6078 102895
rect 5122 102846 5134 102849
rect 6066 102846 6078 102849
rect 6130 102846 6142 102898
rect 12674 102846 12686 102898
rect 12738 102846 12750 102898
rect 9438 102834 9490 102846
rect 1344 102730 28560 102764
rect 1344 102678 4616 102730
rect 4668 102678 4720 102730
rect 4772 102678 4824 102730
rect 4876 102678 11420 102730
rect 11472 102678 11524 102730
rect 11576 102678 11628 102730
rect 11680 102678 18224 102730
rect 18276 102678 18328 102730
rect 18380 102678 18432 102730
rect 18484 102678 25028 102730
rect 25080 102678 25132 102730
rect 25184 102678 25236 102730
rect 25288 102678 28560 102730
rect 1344 102644 28560 102678
rect 12238 102562 12290 102574
rect 4162 102510 4174 102562
rect 4226 102559 4238 102562
rect 5058 102559 5070 102562
rect 4226 102513 5070 102559
rect 4226 102510 4238 102513
rect 5058 102510 5070 102513
rect 5122 102510 5134 102562
rect 8306 102510 8318 102562
rect 8370 102510 8382 102562
rect 12238 102498 12290 102510
rect 22542 102562 22594 102574
rect 22542 102498 22594 102510
rect 5966 102450 6018 102462
rect 5966 102386 6018 102398
rect 8654 102450 8706 102462
rect 20190 102450 20242 102462
rect 11106 102398 11118 102450
rect 11170 102398 11182 102450
rect 16818 102398 16830 102450
rect 16882 102398 16894 102450
rect 8654 102386 8706 102398
rect 20190 102386 20242 102398
rect 20638 102450 20690 102462
rect 20638 102386 20690 102398
rect 20750 102450 20802 102462
rect 20750 102386 20802 102398
rect 22766 102450 22818 102462
rect 22766 102386 22818 102398
rect 23662 102450 23714 102462
rect 23662 102386 23714 102398
rect 24222 102450 24274 102462
rect 24222 102386 24274 102398
rect 24782 102450 24834 102462
rect 24782 102386 24834 102398
rect 3390 102338 3442 102350
rect 8878 102338 8930 102350
rect 9550 102338 9602 102350
rect 12350 102338 12402 102350
rect 7634 102286 7646 102338
rect 7698 102286 7710 102338
rect 9202 102286 9214 102338
rect 9266 102286 9278 102338
rect 10098 102286 10110 102338
rect 10162 102286 10174 102338
rect 3390 102274 3442 102286
rect 8878 102274 8930 102286
rect 9550 102274 9602 102286
rect 12350 102274 12402 102286
rect 12574 102338 12626 102350
rect 12574 102274 12626 102286
rect 12798 102338 12850 102350
rect 12798 102274 12850 102286
rect 13806 102338 13858 102350
rect 20414 102338 20466 102350
rect 14242 102286 14254 102338
rect 14306 102286 14318 102338
rect 13806 102274 13858 102286
rect 20414 102274 20466 102286
rect 21534 102338 21586 102350
rect 23214 102338 23266 102350
rect 21858 102286 21870 102338
rect 21922 102286 21934 102338
rect 23986 102286 23998 102338
rect 24050 102286 24062 102338
rect 21534 102274 21586 102286
rect 23214 102274 23266 102286
rect 9662 102226 9714 102238
rect 9662 102162 9714 102174
rect 13470 102226 13522 102238
rect 13470 102162 13522 102174
rect 13582 102226 13634 102238
rect 13582 102162 13634 102174
rect 19742 102226 19794 102238
rect 19742 102162 19794 102174
rect 19966 102226 20018 102238
rect 19966 102162 20018 102174
rect 24334 102226 24386 102238
rect 24334 102162 24386 102174
rect 2606 102114 2658 102126
rect 2606 102050 2658 102062
rect 3054 102114 3106 102126
rect 3054 102050 3106 102062
rect 3502 102114 3554 102126
rect 3502 102050 3554 102062
rect 3726 102114 3778 102126
rect 3726 102050 3778 102062
rect 4286 102114 4338 102126
rect 4286 102050 4338 102062
rect 4734 102114 4786 102126
rect 4734 102050 4786 102062
rect 5070 102114 5122 102126
rect 5070 102050 5122 102062
rect 6526 102114 6578 102126
rect 6526 102050 6578 102062
rect 6862 102114 6914 102126
rect 6862 102050 6914 102062
rect 7310 102114 7362 102126
rect 7310 102050 7362 102062
rect 7758 102114 7810 102126
rect 7758 102050 7810 102062
rect 9774 102114 9826 102126
rect 9774 102050 9826 102062
rect 12238 102114 12290 102126
rect 12238 102050 12290 102062
rect 21310 102114 21362 102126
rect 21310 102050 21362 102062
rect 21422 102114 21474 102126
rect 22194 102062 22206 102114
rect 22258 102062 22270 102114
rect 21422 102050 21474 102062
rect 1344 101946 28720 101980
rect 1344 101894 8018 101946
rect 8070 101894 8122 101946
rect 8174 101894 8226 101946
rect 8278 101894 14822 101946
rect 14874 101894 14926 101946
rect 14978 101894 15030 101946
rect 15082 101894 21626 101946
rect 21678 101894 21730 101946
rect 21782 101894 21834 101946
rect 21886 101894 28430 101946
rect 28482 101894 28534 101946
rect 28586 101894 28638 101946
rect 28690 101894 28720 101946
rect 1344 101860 28720 101894
rect 17502 101778 17554 101790
rect 17502 101714 17554 101726
rect 24558 101666 24610 101678
rect 9874 101614 9886 101666
rect 9938 101614 9950 101666
rect 19394 101614 19406 101666
rect 19458 101614 19470 101666
rect 24558 101602 24610 101614
rect 23326 101554 23378 101566
rect 4498 101502 4510 101554
rect 4562 101502 4574 101554
rect 5842 101502 5854 101554
rect 5906 101502 5918 101554
rect 10210 101502 10222 101554
rect 10274 101502 10286 101554
rect 11106 101502 11118 101554
rect 11170 101502 11182 101554
rect 12226 101502 12238 101554
rect 12290 101502 12302 101554
rect 22194 101502 22206 101554
rect 22258 101502 22270 101554
rect 23326 101490 23378 101502
rect 23662 101554 23714 101566
rect 23662 101490 23714 101502
rect 23886 101554 23938 101566
rect 23886 101490 23938 101502
rect 5182 101442 5234 101454
rect 1698 101390 1710 101442
rect 1762 101390 1774 101442
rect 3826 101390 3838 101442
rect 3890 101390 3902 101442
rect 5182 101378 5234 101390
rect 5630 101442 5682 101454
rect 8766 101442 8818 101454
rect 23550 101442 23602 101454
rect 6626 101390 6638 101442
rect 6690 101390 6702 101442
rect 10658 101390 10670 101442
rect 10722 101390 10734 101442
rect 14242 101390 14254 101442
rect 14306 101390 14318 101442
rect 5630 101378 5682 101390
rect 8766 101378 8818 101390
rect 23550 101378 23602 101390
rect 25342 101442 25394 101454
rect 25342 101378 25394 101390
rect 24334 101330 24386 101342
rect 24334 101266 24386 101278
rect 24670 101330 24722 101342
rect 24670 101266 24722 101278
rect 1344 101162 28560 101196
rect 1344 101110 4616 101162
rect 4668 101110 4720 101162
rect 4772 101110 4824 101162
rect 4876 101110 11420 101162
rect 11472 101110 11524 101162
rect 11576 101110 11628 101162
rect 11680 101110 18224 101162
rect 18276 101110 18328 101162
rect 18380 101110 18432 101162
rect 18484 101110 25028 101162
rect 25080 101110 25132 101162
rect 25184 101110 25236 101162
rect 25288 101110 28560 101162
rect 1344 101076 28560 101110
rect 3726 100882 3778 100894
rect 3726 100818 3778 100830
rect 6302 100882 6354 100894
rect 7410 100830 7422 100882
rect 7474 100830 7486 100882
rect 10658 100830 10670 100882
rect 10722 100830 10734 100882
rect 12562 100830 12574 100882
rect 12626 100830 12638 100882
rect 21298 100830 21310 100882
rect 21362 100830 21374 100882
rect 24546 100830 24558 100882
rect 24610 100830 24622 100882
rect 6302 100818 6354 100830
rect 3278 100770 3330 100782
rect 3278 100706 3330 100718
rect 3502 100770 3554 100782
rect 3502 100706 3554 100718
rect 3950 100770 4002 100782
rect 3950 100706 4002 100718
rect 5742 100770 5794 100782
rect 20078 100770 20130 100782
rect 7298 100718 7310 100770
rect 7362 100718 7374 100770
rect 9314 100718 9326 100770
rect 9378 100718 9390 100770
rect 10434 100718 10446 100770
rect 10498 100718 10510 100770
rect 12898 100718 12910 100770
rect 12962 100718 12974 100770
rect 13458 100718 13470 100770
rect 13522 100718 13534 100770
rect 19730 100718 19742 100770
rect 19794 100718 19806 100770
rect 24210 100718 24222 100770
rect 24274 100718 24286 100770
rect 27346 100718 27358 100770
rect 27410 100718 27422 100770
rect 5742 100706 5794 100718
rect 20078 100706 20130 100718
rect 2606 100658 2658 100670
rect 2606 100594 2658 100606
rect 4846 100658 4898 100670
rect 4846 100594 4898 100606
rect 6414 100658 6466 100670
rect 6414 100594 6466 100606
rect 7758 100658 7810 100670
rect 20302 100658 20354 100670
rect 9538 100606 9550 100658
rect 9602 100606 9614 100658
rect 15474 100606 15486 100658
rect 15538 100606 15550 100658
rect 23426 100606 23438 100658
rect 23490 100606 23502 100658
rect 26674 100606 26686 100658
rect 26738 100606 26750 100658
rect 7758 100594 7810 100606
rect 20302 100594 20354 100606
rect 2158 100546 2210 100558
rect 2158 100482 2210 100494
rect 3054 100546 3106 100558
rect 3054 100482 3106 100494
rect 4510 100546 4562 100558
rect 4510 100482 4562 100494
rect 4958 100546 5010 100558
rect 4958 100482 5010 100494
rect 5182 100546 5234 100558
rect 5182 100482 5234 100494
rect 6190 100546 6242 100558
rect 6190 100482 6242 100494
rect 7422 100546 7474 100558
rect 7422 100482 7474 100494
rect 20750 100546 20802 100558
rect 20750 100482 20802 100494
rect 1344 100378 28720 100412
rect 1344 100326 8018 100378
rect 8070 100326 8122 100378
rect 8174 100326 8226 100378
rect 8278 100326 14822 100378
rect 14874 100326 14926 100378
rect 14978 100326 15030 100378
rect 15082 100326 21626 100378
rect 21678 100326 21730 100378
rect 21782 100326 21834 100378
rect 21886 100326 28430 100378
rect 28482 100326 28534 100378
rect 28586 100326 28638 100378
rect 28690 100326 28720 100378
rect 1344 100292 28720 100326
rect 4286 100210 4338 100222
rect 4286 100146 4338 100158
rect 8766 100210 8818 100222
rect 8766 100146 8818 100158
rect 8990 100210 9042 100222
rect 8990 100146 9042 100158
rect 23438 100210 23490 100222
rect 23438 100146 23490 100158
rect 23550 100210 23602 100222
rect 23550 100146 23602 100158
rect 25230 100210 25282 100222
rect 25230 100146 25282 100158
rect 25342 100210 25394 100222
rect 25342 100146 25394 100158
rect 3502 100098 3554 100110
rect 8542 100098 8594 100110
rect 25678 100098 25730 100110
rect 5282 100046 5294 100098
rect 5346 100046 5358 100098
rect 11106 100046 11118 100098
rect 11170 100046 11182 100098
rect 21186 100046 21198 100098
rect 21250 100046 21262 100098
rect 3502 100034 3554 100046
rect 8542 100034 8594 100046
rect 25678 100034 25730 100046
rect 2942 99986 2994 99998
rect 2942 99922 2994 99934
rect 3166 99986 3218 99998
rect 22878 99986 22930 99998
rect 4610 99934 4622 99986
rect 4674 99934 4686 99986
rect 10098 99934 10110 99986
rect 10162 99934 10174 99986
rect 11778 99934 11790 99986
rect 11842 99934 11854 99986
rect 18274 99934 18286 99986
rect 18338 99934 18350 99986
rect 3166 99922 3218 99934
rect 22878 99922 22930 99934
rect 23326 99986 23378 99998
rect 23326 99922 23378 99934
rect 24110 99986 24162 99998
rect 24110 99922 24162 99934
rect 25454 99986 25506 99998
rect 25454 99922 25506 99934
rect 2158 99874 2210 99886
rect 2158 99810 2210 99822
rect 2606 99874 2658 99886
rect 3390 99874 3442 99886
rect 2818 99822 2830 99874
rect 2882 99822 2894 99874
rect 2606 99810 2658 99822
rect 2146 99710 2158 99762
rect 2210 99759 2222 99762
rect 2833 99759 2879 99822
rect 3390 99810 3442 99822
rect 7422 99874 7474 99886
rect 7422 99810 7474 99822
rect 8206 99874 8258 99886
rect 8206 99810 8258 99822
rect 8878 99874 8930 99886
rect 23886 99874 23938 99886
rect 10770 99822 10782 99874
rect 10834 99822 10846 99874
rect 13570 99822 13582 99874
rect 13634 99822 13646 99874
rect 8878 99810 8930 99822
rect 23886 99810 23938 99822
rect 26238 99874 26290 99886
rect 26238 99810 26290 99822
rect 26686 99874 26738 99886
rect 26686 99810 26738 99822
rect 2210 99713 2879 99759
rect 2210 99710 2222 99713
rect 24434 99710 24446 99762
rect 24498 99710 24510 99762
rect 1344 99594 28560 99628
rect 1344 99542 4616 99594
rect 4668 99542 4720 99594
rect 4772 99542 4824 99594
rect 4876 99542 11420 99594
rect 11472 99542 11524 99594
rect 11576 99542 11628 99594
rect 11680 99542 18224 99594
rect 18276 99542 18328 99594
rect 18380 99542 18432 99594
rect 18484 99542 25028 99594
rect 25080 99542 25132 99594
rect 25184 99542 25236 99594
rect 25288 99542 28560 99594
rect 1344 99508 28560 99542
rect 22306 99374 22318 99426
rect 22370 99374 22382 99426
rect 5182 99314 5234 99326
rect 20638 99314 20690 99326
rect 1698 99262 1710 99314
rect 1762 99262 1774 99314
rect 3826 99262 3838 99314
rect 3890 99262 3902 99314
rect 11778 99262 11790 99314
rect 11842 99262 11854 99314
rect 15474 99262 15486 99314
rect 15538 99262 15550 99314
rect 24882 99262 24894 99314
rect 24946 99262 24958 99314
rect 5182 99250 5234 99262
rect 20638 99250 20690 99262
rect 5854 99202 5906 99214
rect 6638 99202 6690 99214
rect 4610 99150 4622 99202
rect 4674 99150 4686 99202
rect 6066 99150 6078 99202
rect 6130 99150 6142 99202
rect 6290 99150 6302 99202
rect 6354 99150 6366 99202
rect 5854 99138 5906 99150
rect 6638 99138 6690 99150
rect 6750 99202 6802 99214
rect 6750 99138 6802 99150
rect 7422 99202 7474 99214
rect 19182 99202 19234 99214
rect 7634 99150 7646 99202
rect 7698 99150 7710 99202
rect 14242 99150 14254 99202
rect 14306 99150 14318 99202
rect 7422 99138 7474 99150
rect 19182 99138 19234 99150
rect 19854 99202 19906 99214
rect 19854 99138 19906 99150
rect 20190 99202 20242 99214
rect 21758 99202 21810 99214
rect 21522 99150 21534 99202
rect 21586 99150 21598 99202
rect 20190 99138 20242 99150
rect 21758 99138 21810 99150
rect 21870 99202 21922 99214
rect 22866 99150 22878 99202
rect 22930 99150 22942 99202
rect 21870 99138 21922 99150
rect 6526 99090 6578 99102
rect 6526 99026 6578 99038
rect 7086 99090 7138 99102
rect 7086 99026 7138 99038
rect 6862 98978 6914 98990
rect 6862 98914 6914 98926
rect 19070 98978 19122 98990
rect 19070 98914 19122 98926
rect 19294 98978 19346 98990
rect 19294 98914 19346 98926
rect 19518 98978 19570 98990
rect 19518 98914 19570 98926
rect 20078 98978 20130 98990
rect 20078 98914 20130 98926
rect 1344 98810 28720 98844
rect 1344 98758 8018 98810
rect 8070 98758 8122 98810
rect 8174 98758 8226 98810
rect 8278 98758 14822 98810
rect 14874 98758 14926 98810
rect 14978 98758 15030 98810
rect 15082 98758 21626 98810
rect 21678 98758 21730 98810
rect 21782 98758 21834 98810
rect 21886 98758 28430 98810
rect 28482 98758 28534 98810
rect 28586 98758 28638 98810
rect 28690 98758 28720 98810
rect 1344 98724 28720 98758
rect 2830 98642 2882 98654
rect 2830 98578 2882 98590
rect 3054 98642 3106 98654
rect 3054 98578 3106 98590
rect 3278 98642 3330 98654
rect 3278 98578 3330 98590
rect 4398 98642 4450 98654
rect 4398 98578 4450 98590
rect 10894 98642 10946 98654
rect 10894 98578 10946 98590
rect 18062 98642 18114 98654
rect 18062 98578 18114 98590
rect 18174 98642 18226 98654
rect 18174 98578 18226 98590
rect 18734 98642 18786 98654
rect 18734 98578 18786 98590
rect 18846 98642 18898 98654
rect 18846 98578 18898 98590
rect 21870 98642 21922 98654
rect 21870 98578 21922 98590
rect 22766 98642 22818 98654
rect 22766 98578 22818 98590
rect 23886 98642 23938 98654
rect 23886 98578 23938 98590
rect 4062 98530 4114 98542
rect 9886 98530 9938 98542
rect 17950 98530 18002 98542
rect 24446 98530 24498 98542
rect 6626 98478 6638 98530
rect 6690 98478 6702 98530
rect 11778 98478 11790 98530
rect 11842 98478 11854 98530
rect 17826 98478 17838 98530
rect 17890 98478 17902 98530
rect 20850 98478 20862 98530
rect 20914 98478 20926 98530
rect 21186 98478 21198 98530
rect 21250 98478 21262 98530
rect 4062 98466 4114 98478
rect 9886 98466 9938 98478
rect 17950 98466 18002 98478
rect 24446 98466 24498 98478
rect 3390 98418 3442 98430
rect 9550 98418 9602 98430
rect 5170 98366 5182 98418
rect 5234 98366 5246 98418
rect 5954 98366 5966 98418
rect 6018 98366 6030 98418
rect 3390 98354 3442 98366
rect 9550 98354 9602 98366
rect 9774 98418 9826 98430
rect 9774 98354 9826 98366
rect 10110 98418 10162 98430
rect 10110 98354 10162 98366
rect 10334 98418 10386 98430
rect 10334 98354 10386 98366
rect 10782 98418 10834 98430
rect 18286 98418 18338 98430
rect 15586 98366 15598 98418
rect 15650 98366 15662 98418
rect 10782 98354 10834 98366
rect 18286 98354 18338 98366
rect 18622 98418 18674 98430
rect 20190 98418 20242 98430
rect 19170 98366 19182 98418
rect 19234 98366 19246 98418
rect 18622 98354 18674 98366
rect 20190 98354 20242 98366
rect 23998 98418 24050 98430
rect 23998 98354 24050 98366
rect 24558 98418 24610 98430
rect 28018 98366 28030 98418
rect 28082 98366 28094 98418
rect 24558 98354 24610 98366
rect 2382 98306 2434 98318
rect 2382 98242 2434 98254
rect 4846 98306 4898 98318
rect 4846 98242 4898 98254
rect 5406 98306 5458 98318
rect 19742 98306 19794 98318
rect 8754 98254 8766 98306
rect 8818 98254 8830 98306
rect 5406 98242 5458 98254
rect 19742 98242 19794 98254
rect 22318 98306 22370 98318
rect 22318 98242 22370 98254
rect 23550 98306 23602 98318
rect 25218 98254 25230 98306
rect 25282 98254 25294 98306
rect 27346 98254 27358 98306
rect 27410 98254 27422 98306
rect 23550 98242 23602 98254
rect 5518 98194 5570 98206
rect 5518 98130 5570 98142
rect 20526 98194 20578 98206
rect 23886 98194 23938 98206
rect 21858 98142 21870 98194
rect 21922 98191 21934 98194
rect 22306 98191 22318 98194
rect 21922 98145 22318 98191
rect 21922 98142 21934 98145
rect 22306 98142 22318 98145
rect 22370 98142 22382 98194
rect 20526 98130 20578 98142
rect 23886 98130 23938 98142
rect 24446 98194 24498 98206
rect 24446 98130 24498 98142
rect 1344 98026 28560 98060
rect 1344 97974 4616 98026
rect 4668 97974 4720 98026
rect 4772 97974 4824 98026
rect 4876 97974 11420 98026
rect 11472 97974 11524 98026
rect 11576 97974 11628 98026
rect 11680 97974 18224 98026
rect 18276 97974 18328 98026
rect 18380 97974 18432 98026
rect 18484 97974 25028 98026
rect 25080 97974 25132 98026
rect 25184 97974 25236 98026
rect 25288 97974 28560 98026
rect 1344 97940 28560 97974
rect 23438 97858 23490 97870
rect 15138 97806 15150 97858
rect 15202 97806 15214 97858
rect 25330 97806 25342 97858
rect 25394 97806 25406 97858
rect 23438 97794 23490 97806
rect 3278 97746 3330 97758
rect 3278 97682 3330 97694
rect 4622 97746 4674 97758
rect 21870 97746 21922 97758
rect 17714 97694 17726 97746
rect 17778 97694 17790 97746
rect 4622 97682 4674 97694
rect 21870 97682 21922 97694
rect 22542 97746 22594 97758
rect 24434 97694 24446 97746
rect 24498 97694 24510 97746
rect 25442 97694 25454 97746
rect 25506 97694 25518 97746
rect 22542 97682 22594 97694
rect 3838 97634 3890 97646
rect 3838 97570 3890 97582
rect 5742 97634 5794 97646
rect 5742 97570 5794 97582
rect 5854 97634 5906 97646
rect 5854 97570 5906 97582
rect 6078 97634 6130 97646
rect 6078 97570 6130 97582
rect 6190 97634 6242 97646
rect 6190 97570 6242 97582
rect 6750 97634 6802 97646
rect 6750 97570 6802 97582
rect 6862 97634 6914 97646
rect 14702 97634 14754 97646
rect 19294 97634 19346 97646
rect 23102 97634 23154 97646
rect 7858 97582 7870 97634
rect 7922 97582 7934 97634
rect 15026 97582 15038 97634
rect 15090 97582 15102 97634
rect 15922 97582 15934 97634
rect 15986 97582 15998 97634
rect 16594 97582 16606 97634
rect 16658 97582 16670 97634
rect 17490 97582 17502 97634
rect 17554 97582 17566 97634
rect 20066 97582 20078 97634
rect 20130 97582 20142 97634
rect 6862 97570 6914 97582
rect 14702 97570 14754 97582
rect 19294 97570 19346 97582
rect 23102 97570 23154 97582
rect 23550 97634 23602 97646
rect 27358 97634 27410 97646
rect 24210 97582 24222 97634
rect 24274 97582 24286 97634
rect 25666 97582 25678 97634
rect 25730 97582 25742 97634
rect 23550 97570 23602 97582
rect 27358 97570 27410 97582
rect 5070 97522 5122 97534
rect 5070 97458 5122 97470
rect 7198 97522 7250 97534
rect 14142 97522 14194 97534
rect 18958 97522 19010 97534
rect 21422 97522 21474 97534
rect 10434 97470 10446 97522
rect 10498 97470 10510 97522
rect 16706 97470 16718 97522
rect 16770 97470 16782 97522
rect 17378 97470 17390 97522
rect 17442 97470 17454 97522
rect 19954 97470 19966 97522
rect 20018 97470 20030 97522
rect 7198 97458 7250 97470
rect 14142 97458 14194 97470
rect 18958 97458 19010 97470
rect 21422 97458 21474 97470
rect 22878 97522 22930 97534
rect 22878 97458 22930 97470
rect 24894 97522 24946 97534
rect 24894 97458 24946 97470
rect 26686 97522 26738 97534
rect 26686 97458 26738 97470
rect 26798 97522 26850 97534
rect 26798 97458 26850 97470
rect 2830 97410 2882 97422
rect 2830 97346 2882 97358
rect 4174 97410 4226 97422
rect 4174 97346 4226 97358
rect 6974 97410 7026 97422
rect 6974 97346 7026 97358
rect 13806 97410 13858 97422
rect 13806 97346 13858 97358
rect 14030 97410 14082 97422
rect 14030 97346 14082 97358
rect 14254 97410 14306 97422
rect 14254 97346 14306 97358
rect 17726 97410 17778 97422
rect 17726 97346 17778 97358
rect 17950 97410 18002 97422
rect 17950 97346 18002 97358
rect 18398 97410 18450 97422
rect 18398 97346 18450 97358
rect 20638 97410 20690 97422
rect 20638 97346 20690 97358
rect 23326 97410 23378 97422
rect 23326 97346 23378 97358
rect 27022 97410 27074 97422
rect 27022 97346 27074 97358
rect 1344 97242 28720 97276
rect 1344 97190 8018 97242
rect 8070 97190 8122 97242
rect 8174 97190 8226 97242
rect 8278 97190 14822 97242
rect 14874 97190 14926 97242
rect 14978 97190 15030 97242
rect 15082 97190 21626 97242
rect 21678 97190 21730 97242
rect 21782 97190 21834 97242
rect 21886 97190 28430 97242
rect 28482 97190 28534 97242
rect 28586 97190 28638 97242
rect 28690 97190 28720 97242
rect 1344 97156 28720 97190
rect 8878 97074 8930 97086
rect 7522 97022 7534 97074
rect 7586 97022 7598 97074
rect 8878 97010 8930 97022
rect 13806 97074 13858 97086
rect 13806 97010 13858 97022
rect 18174 97074 18226 97086
rect 23550 97074 23602 97086
rect 18498 97022 18510 97074
rect 18562 97022 18574 97074
rect 18174 97010 18226 97022
rect 23550 97010 23602 97022
rect 2270 96962 2322 96974
rect 2270 96898 2322 96910
rect 2718 96962 2770 96974
rect 13470 96962 13522 96974
rect 6290 96910 6302 96962
rect 6354 96910 6366 96962
rect 11890 96910 11902 96962
rect 11954 96910 11966 96962
rect 2718 96898 2770 96910
rect 13470 96898 13522 96910
rect 13694 96962 13746 96974
rect 13694 96898 13746 96910
rect 14030 96962 14082 96974
rect 17950 96962 18002 96974
rect 15698 96910 15710 96962
rect 15762 96910 15774 96962
rect 14030 96898 14082 96910
rect 17950 96898 18002 96910
rect 20190 96962 20242 96974
rect 22654 96962 22706 96974
rect 20850 96910 20862 96962
rect 20914 96910 20926 96962
rect 21298 96910 21310 96962
rect 21362 96910 21374 96962
rect 27346 96910 27358 96962
rect 27410 96910 27422 96962
rect 20190 96898 20242 96910
rect 22654 96898 22706 96910
rect 1934 96850 1986 96862
rect 1934 96786 1986 96798
rect 2158 96850 2210 96862
rect 2158 96786 2210 96798
rect 2494 96850 2546 96862
rect 2494 96786 2546 96798
rect 2942 96850 2994 96862
rect 2942 96786 2994 96798
rect 3278 96850 3330 96862
rect 8542 96850 8594 96862
rect 6962 96798 6974 96850
rect 7026 96798 7038 96850
rect 3278 96786 3330 96798
rect 8542 96786 8594 96798
rect 8766 96850 8818 96862
rect 8766 96786 8818 96798
rect 9102 96850 9154 96862
rect 16494 96850 16546 96862
rect 18846 96850 18898 96862
rect 10882 96798 10894 96850
rect 10946 96798 10958 96850
rect 11778 96798 11790 96850
rect 11842 96798 11854 96850
rect 12338 96798 12350 96850
rect 12402 96798 12414 96850
rect 14354 96798 14366 96850
rect 14418 96798 14430 96850
rect 15138 96798 15150 96850
rect 15202 96798 15214 96850
rect 17378 96798 17390 96850
rect 17442 96798 17454 96850
rect 17714 96798 17726 96850
rect 17778 96798 17790 96850
rect 22082 96798 22094 96850
rect 22146 96798 22158 96850
rect 28018 96798 28030 96850
rect 28082 96798 28094 96850
rect 9102 96786 9154 96798
rect 16494 96786 16546 96798
rect 18846 96786 18898 96798
rect 3166 96738 3218 96750
rect 3166 96674 3218 96686
rect 4174 96738 4226 96750
rect 4174 96674 4226 96686
rect 8094 96738 8146 96750
rect 13134 96738 13186 96750
rect 16270 96738 16322 96750
rect 10210 96686 10222 96738
rect 10274 96686 10286 96738
rect 12002 96686 12014 96738
rect 12066 96686 12078 96738
rect 15026 96686 15038 96738
rect 15090 96686 15102 96738
rect 8094 96674 8146 96686
rect 13134 96674 13186 96686
rect 16270 96674 16322 96686
rect 16830 96738 16882 96750
rect 19070 96738 19122 96750
rect 17826 96686 17838 96738
rect 17890 96686 17902 96738
rect 16830 96674 16882 96686
rect 19070 96674 19122 96686
rect 19630 96738 19682 96750
rect 19630 96674 19682 96686
rect 23886 96738 23938 96750
rect 25218 96686 25230 96738
rect 25282 96686 25294 96738
rect 23886 96674 23938 96686
rect 7870 96626 7922 96638
rect 7870 96562 7922 96574
rect 20526 96626 20578 96638
rect 20526 96562 20578 96574
rect 1344 96458 28560 96492
rect 1344 96406 4616 96458
rect 4668 96406 4720 96458
rect 4772 96406 4824 96458
rect 4876 96406 11420 96458
rect 11472 96406 11524 96458
rect 11576 96406 11628 96458
rect 11680 96406 18224 96458
rect 18276 96406 18328 96458
rect 18380 96406 18432 96458
rect 18484 96406 25028 96458
rect 25080 96406 25132 96458
rect 25184 96406 25236 96458
rect 25288 96406 28560 96458
rect 1344 96372 28560 96406
rect 18286 96290 18338 96302
rect 18286 96226 18338 96238
rect 18622 96290 18674 96302
rect 18622 96226 18674 96238
rect 19518 96290 19570 96302
rect 19518 96226 19570 96238
rect 21870 96290 21922 96302
rect 21870 96226 21922 96238
rect 22094 96290 22146 96302
rect 22094 96226 22146 96238
rect 22766 96290 22818 96302
rect 22766 96226 22818 96238
rect 16718 96178 16770 96190
rect 1698 96126 1710 96178
rect 1762 96126 1774 96178
rect 3826 96126 3838 96178
rect 3890 96126 3902 96178
rect 6626 96126 6638 96178
rect 6690 96126 6702 96178
rect 12114 96126 12126 96178
rect 12178 96126 12190 96178
rect 14690 96126 14702 96178
rect 14754 96126 14766 96178
rect 24322 96126 24334 96178
rect 24386 96126 24398 96178
rect 16718 96114 16770 96126
rect 15934 96066 15986 96078
rect 4610 96014 4622 96066
rect 4674 96014 4686 96066
rect 11218 96014 11230 96066
rect 11282 96014 11294 96066
rect 12002 96014 12014 96066
rect 12066 96014 12078 96066
rect 14018 96014 14030 96066
rect 14082 96014 14094 96066
rect 14802 96014 14814 96066
rect 14866 96014 14878 96066
rect 15934 96002 15986 96014
rect 16382 96066 16434 96078
rect 16382 96002 16434 96014
rect 17502 96066 17554 96078
rect 17502 96002 17554 96014
rect 18062 96066 18114 96078
rect 18062 96002 18114 96014
rect 19854 96066 19906 96078
rect 19854 96002 19906 96014
rect 22318 96066 22370 96078
rect 25230 96066 25282 96078
rect 23650 96014 23662 96066
rect 23714 96014 23726 96066
rect 22318 96002 22370 96014
rect 25230 96002 25282 96014
rect 25902 96066 25954 96078
rect 25902 96002 25954 96014
rect 6078 95954 6130 95966
rect 17614 95954 17666 95966
rect 12114 95902 12126 95954
rect 12178 95902 12190 95954
rect 15362 95902 15374 95954
rect 15426 95902 15438 95954
rect 6078 95890 6130 95902
rect 17614 95890 17666 95902
rect 18846 95954 18898 95966
rect 21646 95954 21698 95966
rect 20066 95902 20078 95954
rect 20130 95902 20142 95954
rect 20626 95902 20638 95954
rect 20690 95902 20702 95954
rect 18846 95890 18898 95902
rect 21646 95890 21698 95902
rect 23214 95954 23266 95966
rect 23214 95890 23266 95902
rect 25342 95954 25394 95966
rect 25342 95890 25394 95902
rect 5070 95842 5122 95854
rect 5070 95778 5122 95790
rect 13694 95842 13746 95854
rect 13694 95778 13746 95790
rect 15710 95842 15762 95854
rect 15710 95778 15762 95790
rect 15822 95842 15874 95854
rect 15822 95778 15874 95790
rect 17726 95842 17778 95854
rect 17726 95778 17778 95790
rect 23326 95842 23378 95854
rect 23326 95778 23378 95790
rect 25454 95842 25506 95854
rect 25454 95778 25506 95790
rect 26238 95842 26290 95854
rect 26238 95778 26290 95790
rect 1344 95674 28720 95708
rect 1344 95622 8018 95674
rect 8070 95622 8122 95674
rect 8174 95622 8226 95674
rect 8278 95622 14822 95674
rect 14874 95622 14926 95674
rect 14978 95622 15030 95674
rect 15082 95622 21626 95674
rect 21678 95622 21730 95674
rect 21782 95622 21834 95674
rect 21886 95622 28430 95674
rect 28482 95622 28534 95674
rect 28586 95622 28638 95674
rect 28690 95622 28720 95674
rect 1344 95588 28720 95622
rect 2382 95506 2434 95518
rect 2382 95442 2434 95454
rect 3278 95506 3330 95518
rect 13246 95506 13298 95518
rect 6514 95454 6526 95506
rect 6578 95454 6590 95506
rect 3278 95442 3330 95454
rect 13246 95442 13298 95454
rect 15598 95506 15650 95518
rect 15598 95442 15650 95454
rect 16830 95506 16882 95518
rect 16830 95442 16882 95454
rect 18622 95506 18674 95518
rect 18622 95442 18674 95454
rect 20526 95506 20578 95518
rect 20526 95442 20578 95454
rect 24110 95506 24162 95518
rect 24110 95442 24162 95454
rect 24446 95506 24498 95518
rect 24446 95442 24498 95454
rect 2830 95394 2882 95406
rect 2830 95330 2882 95342
rect 5966 95394 6018 95406
rect 5966 95330 6018 95342
rect 6862 95394 6914 95406
rect 6862 95330 6914 95342
rect 9662 95394 9714 95406
rect 9662 95330 9714 95342
rect 10222 95394 10274 95406
rect 10222 95330 10274 95342
rect 13918 95394 13970 95406
rect 13918 95330 13970 95342
rect 15038 95394 15090 95406
rect 15038 95330 15090 95342
rect 15934 95394 15986 95406
rect 15934 95330 15986 95342
rect 16270 95394 16322 95406
rect 16270 95330 16322 95342
rect 18174 95394 18226 95406
rect 18174 95330 18226 95342
rect 18846 95394 18898 95406
rect 18846 95330 18898 95342
rect 20078 95394 20130 95406
rect 20078 95330 20130 95342
rect 24558 95394 24610 95406
rect 24558 95330 24610 95342
rect 25454 95394 25506 95406
rect 25454 95330 25506 95342
rect 5854 95282 5906 95294
rect 5854 95218 5906 95230
rect 6078 95282 6130 95294
rect 9550 95282 9602 95294
rect 7186 95230 7198 95282
rect 7250 95230 7262 95282
rect 8530 95230 8542 95282
rect 8594 95230 8606 95282
rect 6078 95218 6130 95230
rect 9550 95218 9602 95230
rect 10334 95282 10386 95294
rect 10334 95218 10386 95230
rect 10558 95282 10610 95294
rect 13582 95282 13634 95294
rect 10770 95230 10782 95282
rect 10834 95230 10846 95282
rect 10994 95230 11006 95282
rect 11058 95230 11070 95282
rect 12002 95230 12014 95282
rect 12066 95230 12078 95282
rect 12338 95230 12350 95282
rect 12402 95230 12414 95282
rect 10558 95218 10610 95230
rect 13582 95218 13634 95230
rect 14030 95282 14082 95294
rect 14030 95218 14082 95230
rect 14478 95282 14530 95294
rect 14478 95218 14530 95230
rect 14702 95282 14754 95294
rect 14702 95218 14754 95230
rect 15374 95282 15426 95294
rect 15374 95218 15426 95230
rect 15598 95282 15650 95294
rect 15598 95218 15650 95230
rect 16382 95282 16434 95294
rect 18398 95282 18450 95294
rect 17602 95230 17614 95282
rect 17666 95230 17678 95282
rect 16382 95218 16434 95230
rect 18398 95218 18450 95230
rect 19070 95282 19122 95294
rect 19070 95218 19122 95230
rect 24222 95282 24274 95294
rect 24222 95218 24274 95230
rect 25342 95282 25394 95294
rect 25342 95218 25394 95230
rect 25678 95282 25730 95294
rect 25678 95218 25730 95230
rect 26014 95282 26066 95294
rect 26014 95218 26066 95230
rect 3726 95170 3778 95182
rect 3726 95106 3778 95118
rect 4062 95170 4114 95182
rect 4062 95106 4114 95118
rect 4510 95170 4562 95182
rect 4510 95106 4562 95118
rect 4958 95170 5010 95182
rect 4958 95106 5010 95118
rect 5406 95170 5458 95182
rect 5406 95106 5458 95118
rect 6974 95170 7026 95182
rect 6974 95106 7026 95118
rect 7646 95170 7698 95182
rect 8990 95170 9042 95182
rect 8082 95118 8094 95170
rect 8146 95118 8158 95170
rect 7646 95106 7698 95118
rect 8990 95106 9042 95118
rect 13694 95170 13746 95182
rect 13694 95106 13746 95118
rect 14590 95170 14642 95182
rect 17490 95118 17502 95170
rect 17554 95118 17566 95170
rect 14590 95106 14642 95118
rect 9662 95058 9714 95070
rect 19518 95058 19570 95070
rect 4386 95006 4398 95058
rect 4450 95055 4462 95058
rect 4946 95055 4958 95058
rect 4450 95009 4958 95055
rect 4450 95006 4462 95009
rect 4946 95006 4958 95009
rect 5010 95055 5022 95058
rect 5394 95055 5406 95058
rect 5010 95009 5406 95055
rect 5010 95006 5022 95009
rect 5394 95006 5406 95009
rect 5458 95006 5470 95058
rect 11778 95006 11790 95058
rect 11842 95006 11854 95058
rect 9662 94994 9714 95006
rect 19518 94994 19570 95006
rect 19854 95058 19906 95070
rect 19854 94994 19906 95006
rect 1344 94890 28560 94924
rect 1344 94838 4616 94890
rect 4668 94838 4720 94890
rect 4772 94838 4824 94890
rect 4876 94838 11420 94890
rect 11472 94838 11524 94890
rect 11576 94838 11628 94890
rect 11680 94838 18224 94890
rect 18276 94838 18328 94890
rect 18380 94838 18432 94890
rect 18484 94838 25028 94890
rect 25080 94838 25132 94890
rect 25184 94838 25236 94890
rect 25288 94838 28560 94890
rect 1344 94804 28560 94838
rect 6414 94722 6466 94734
rect 6414 94658 6466 94670
rect 14142 94722 14194 94734
rect 14142 94658 14194 94670
rect 3054 94610 3106 94622
rect 4622 94610 4674 94622
rect 3378 94558 3390 94610
rect 3442 94558 3454 94610
rect 3054 94546 3106 94558
rect 4622 94546 4674 94558
rect 5070 94610 5122 94622
rect 5070 94546 5122 94558
rect 5742 94610 5794 94622
rect 5742 94546 5794 94558
rect 6638 94610 6690 94622
rect 11230 94610 11282 94622
rect 14366 94610 14418 94622
rect 9762 94558 9774 94610
rect 9826 94558 9838 94610
rect 12450 94558 12462 94610
rect 12514 94558 12526 94610
rect 6638 94546 6690 94558
rect 11230 94546 11282 94558
rect 14366 94546 14418 94558
rect 16606 94610 16658 94622
rect 16606 94546 16658 94558
rect 19630 94610 19682 94622
rect 25778 94558 25790 94610
rect 25842 94558 25854 94610
rect 19630 94546 19682 94558
rect 3726 94498 3778 94510
rect 11118 94498 11170 94510
rect 3938 94446 3950 94498
rect 4002 94446 4014 94498
rect 10434 94446 10446 94498
rect 10498 94446 10510 94498
rect 3726 94434 3778 94446
rect 11118 94434 11170 94446
rect 11342 94498 11394 94510
rect 16158 94498 16210 94510
rect 11666 94446 11678 94498
rect 11730 94446 11742 94498
rect 12786 94446 12798 94498
rect 12850 94446 12862 94498
rect 13682 94446 13694 94498
rect 13746 94446 13758 94498
rect 15586 94446 15598 94498
rect 15650 94446 15662 94498
rect 11342 94434 11394 94446
rect 16158 94434 16210 94446
rect 16382 94498 16434 94510
rect 16382 94434 16434 94446
rect 16942 94498 16994 94510
rect 19070 94498 19122 94510
rect 18722 94446 18734 94498
rect 18786 94446 18798 94498
rect 16942 94434 16994 94446
rect 19070 94434 19122 94446
rect 21198 94498 21250 94510
rect 21198 94434 21250 94446
rect 21646 94498 21698 94510
rect 24994 94446 25006 94498
rect 25058 94446 25070 94498
rect 21646 94434 21698 94446
rect 14590 94386 14642 94398
rect 13906 94334 13918 94386
rect 13970 94334 13982 94386
rect 14590 94322 14642 94334
rect 14926 94386 14978 94398
rect 14926 94322 14978 94334
rect 15038 94386 15090 94398
rect 15038 94322 15090 94334
rect 16718 94386 16770 94398
rect 16718 94322 16770 94334
rect 17390 94386 17442 94398
rect 17390 94322 17442 94334
rect 17614 94386 17666 94398
rect 17614 94322 17666 94334
rect 18062 94386 18114 94398
rect 18062 94322 18114 94334
rect 18174 94386 18226 94398
rect 18174 94322 18226 94334
rect 18286 94386 18338 94398
rect 18286 94322 18338 94334
rect 19182 94386 19234 94398
rect 19182 94322 19234 94334
rect 21870 94386 21922 94398
rect 21870 94322 21922 94334
rect 2494 94274 2546 94286
rect 2494 94210 2546 94222
rect 3390 94274 3442 94286
rect 3390 94210 3442 94222
rect 3502 94274 3554 94286
rect 7086 94274 7138 94286
rect 15262 94274 15314 94286
rect 6066 94222 6078 94274
rect 6130 94222 6142 94274
rect 7522 94222 7534 94274
rect 7586 94222 7598 94274
rect 14018 94222 14030 94274
rect 14082 94222 14094 94274
rect 3502 94210 3554 94222
rect 7086 94210 7138 94222
rect 15262 94210 15314 94222
rect 15710 94274 15762 94286
rect 15710 94210 15762 94222
rect 17166 94274 17218 94286
rect 17166 94210 17218 94222
rect 17950 94274 18002 94286
rect 17950 94210 18002 94222
rect 21422 94274 21474 94286
rect 21422 94210 21474 94222
rect 22430 94274 22482 94286
rect 28018 94222 28030 94274
rect 28082 94222 28094 94274
rect 22430 94210 22482 94222
rect 1344 94106 28720 94140
rect 1344 94054 8018 94106
rect 8070 94054 8122 94106
rect 8174 94054 8226 94106
rect 8278 94054 14822 94106
rect 14874 94054 14926 94106
rect 14978 94054 15030 94106
rect 15082 94054 21626 94106
rect 21678 94054 21730 94106
rect 21782 94054 21834 94106
rect 21886 94054 28430 94106
rect 28482 94054 28534 94106
rect 28586 94054 28638 94106
rect 28690 94054 28720 94106
rect 1344 94020 28720 94054
rect 4062 93938 4114 93950
rect 4062 93874 4114 93886
rect 8654 93938 8706 93950
rect 8654 93874 8706 93886
rect 11118 93938 11170 93950
rect 11118 93874 11170 93886
rect 12350 93938 12402 93950
rect 13918 93938 13970 93950
rect 12786 93886 12798 93938
rect 12850 93886 12862 93938
rect 12350 93874 12402 93886
rect 13918 93874 13970 93886
rect 14366 93938 14418 93950
rect 14366 93874 14418 93886
rect 15262 93938 15314 93950
rect 15262 93874 15314 93886
rect 16270 93938 16322 93950
rect 16270 93874 16322 93886
rect 16382 93938 16434 93950
rect 22318 93938 22370 93950
rect 20962 93886 20974 93938
rect 21026 93886 21038 93938
rect 16382 93874 16434 93886
rect 22318 93874 22370 93886
rect 26910 93938 26962 93950
rect 26910 93874 26962 93886
rect 2494 93826 2546 93838
rect 2494 93762 2546 93774
rect 2942 93826 2994 93838
rect 2942 93762 2994 93774
rect 3166 93826 3218 93838
rect 10782 93826 10834 93838
rect 9874 93774 9886 93826
rect 9938 93774 9950 93826
rect 10322 93774 10334 93826
rect 10386 93774 10398 93826
rect 3166 93762 3218 93774
rect 10782 93762 10834 93774
rect 15150 93826 15202 93838
rect 15150 93762 15202 93774
rect 15486 93826 15538 93838
rect 19058 93774 19070 93826
rect 19122 93774 19134 93826
rect 15486 93762 15538 93774
rect 8430 93714 8482 93726
rect 4834 93662 4846 93714
rect 4898 93662 4910 93714
rect 8430 93650 8482 93662
rect 8654 93714 8706 93726
rect 8654 93650 8706 93662
rect 8990 93714 9042 93726
rect 12462 93714 12514 93726
rect 9538 93662 9550 93714
rect 9602 93662 9614 93714
rect 12114 93662 12126 93714
rect 12178 93662 12190 93714
rect 8990 93650 9042 93662
rect 12462 93650 12514 93662
rect 13134 93714 13186 93726
rect 13134 93650 13186 93662
rect 14254 93714 14306 93726
rect 14254 93650 14306 93662
rect 14590 93714 14642 93726
rect 14590 93650 14642 93662
rect 14814 93714 14866 93726
rect 14814 93650 14866 93662
rect 15710 93714 15762 93726
rect 16158 93714 16210 93726
rect 16034 93662 16046 93714
rect 16098 93662 16110 93714
rect 15710 93650 15762 93662
rect 16158 93650 16210 93662
rect 17614 93714 17666 93726
rect 20302 93714 20354 93726
rect 18498 93662 18510 93714
rect 18562 93662 18574 93714
rect 20514 93662 20526 93714
rect 20578 93662 20590 93714
rect 22530 93662 22542 93714
rect 22594 93662 22606 93714
rect 27122 93662 27134 93714
rect 27186 93662 27198 93714
rect 17614 93650 17666 93662
rect 20302 93650 20354 93662
rect 3054 93602 3106 93614
rect 3054 93538 3106 93550
rect 4510 93602 4562 93614
rect 7646 93602 7698 93614
rect 5506 93550 5518 93602
rect 5570 93550 5582 93602
rect 4510 93538 4562 93550
rect 7646 93538 7698 93550
rect 13358 93602 13410 93614
rect 23102 93602 23154 93614
rect 19170 93550 19182 93602
rect 19234 93550 19246 93602
rect 13358 93538 13410 93550
rect 23102 93538 23154 93550
rect 27806 93602 27858 93614
rect 27806 93538 27858 93550
rect 1344 93322 28560 93356
rect 1344 93270 4616 93322
rect 4668 93270 4720 93322
rect 4772 93270 4824 93322
rect 4876 93270 11420 93322
rect 11472 93270 11524 93322
rect 11576 93270 11628 93322
rect 11680 93270 18224 93322
rect 18276 93270 18328 93322
rect 18380 93270 18432 93322
rect 18484 93270 25028 93322
rect 25080 93270 25132 93322
rect 25184 93270 25236 93322
rect 25288 93270 28560 93322
rect 1344 93236 28560 93270
rect 11566 93154 11618 93166
rect 11566 93090 11618 93102
rect 14926 93154 14978 93166
rect 22306 93102 22318 93154
rect 22370 93102 22382 93154
rect 14926 93090 14978 93102
rect 5182 93042 5234 93054
rect 1698 92990 1710 93042
rect 1762 92990 1774 93042
rect 3826 92990 3838 93042
rect 3890 92990 3902 93042
rect 5182 92978 5234 92990
rect 6190 93042 6242 93054
rect 15598 93042 15650 93054
rect 21646 93042 21698 93054
rect 9202 92990 9214 93042
rect 9266 92990 9278 93042
rect 11330 92990 11342 93042
rect 11394 92990 11406 93042
rect 17490 92990 17502 93042
rect 17554 92990 17566 93042
rect 19954 92990 19966 93042
rect 20018 92990 20030 93042
rect 6190 92978 6242 92990
rect 15598 92978 15650 92990
rect 21646 92978 21698 92990
rect 22878 93042 22930 93054
rect 25778 92990 25790 93042
rect 25842 92990 25854 93042
rect 22878 92978 22930 92990
rect 6078 92930 6130 92942
rect 4610 92878 4622 92930
rect 4674 92878 4686 92930
rect 6078 92866 6130 92878
rect 6302 92930 6354 92942
rect 6302 92866 6354 92878
rect 6974 92930 7026 92942
rect 6974 92866 7026 92878
rect 7758 92930 7810 92942
rect 12238 92930 12290 92942
rect 8418 92878 8430 92930
rect 8482 92878 8494 92930
rect 7758 92866 7810 92878
rect 12238 92866 12290 92878
rect 13694 92930 13746 92942
rect 13694 92866 13746 92878
rect 14590 92930 14642 92942
rect 21422 92930 21474 92942
rect 16482 92878 16494 92930
rect 16546 92878 16558 92930
rect 17602 92878 17614 92930
rect 17666 92878 17678 92930
rect 19730 92878 19742 92930
rect 19794 92878 19806 92930
rect 14590 92866 14642 92878
rect 21422 92866 21474 92878
rect 21758 92930 21810 92942
rect 22654 92930 22706 92942
rect 21970 92878 21982 92930
rect 22034 92878 22046 92930
rect 21758 92866 21810 92878
rect 22654 92866 22706 92878
rect 23662 92930 23714 92942
rect 23662 92866 23714 92878
rect 26238 92930 26290 92942
rect 26238 92866 26290 92878
rect 26350 92930 26402 92942
rect 26350 92866 26402 92878
rect 26574 92930 26626 92942
rect 26574 92866 26626 92878
rect 11678 92818 11730 92830
rect 11678 92754 11730 92766
rect 13918 92818 13970 92830
rect 13918 92754 13970 92766
rect 14030 92818 14082 92830
rect 14030 92754 14082 92766
rect 14366 92818 14418 92830
rect 19966 92818 20018 92830
rect 15922 92766 15934 92818
rect 15986 92766 15998 92818
rect 16594 92766 16606 92818
rect 16658 92766 16670 92818
rect 16930 92766 16942 92818
rect 16994 92766 17006 92818
rect 14366 92754 14418 92766
rect 19966 92754 20018 92766
rect 20414 92818 20466 92830
rect 20414 92754 20466 92766
rect 23326 92818 23378 92830
rect 23326 92754 23378 92766
rect 23998 92818 24050 92830
rect 23998 92754 24050 92766
rect 24110 92818 24162 92830
rect 24110 92754 24162 92766
rect 25454 92818 25506 92830
rect 25454 92754 25506 92766
rect 27134 92818 27186 92830
rect 27134 92754 27186 92766
rect 5854 92706 5906 92718
rect 5854 92642 5906 92654
rect 7534 92706 7586 92718
rect 11902 92706 11954 92718
rect 8082 92654 8094 92706
rect 8146 92654 8158 92706
rect 7534 92642 7586 92654
rect 11902 92642 11954 92654
rect 12686 92706 12738 92718
rect 12686 92642 12738 92654
rect 19406 92706 19458 92718
rect 19406 92642 19458 92654
rect 20190 92706 20242 92718
rect 20190 92642 20242 92654
rect 21534 92706 21586 92718
rect 21534 92642 21586 92654
rect 23438 92706 23490 92718
rect 23438 92642 23490 92654
rect 23774 92706 23826 92718
rect 23774 92642 23826 92654
rect 25678 92706 25730 92718
rect 25678 92642 25730 92654
rect 26238 92706 26290 92718
rect 26238 92642 26290 92654
rect 27022 92706 27074 92718
rect 27022 92642 27074 92654
rect 1344 92538 28720 92572
rect 1344 92486 8018 92538
rect 8070 92486 8122 92538
rect 8174 92486 8226 92538
rect 8278 92486 14822 92538
rect 14874 92486 14926 92538
rect 14978 92486 15030 92538
rect 15082 92486 21626 92538
rect 21678 92486 21730 92538
rect 21782 92486 21834 92538
rect 21886 92486 28430 92538
rect 28482 92486 28534 92538
rect 28586 92486 28638 92538
rect 28690 92486 28720 92538
rect 1344 92452 28720 92486
rect 10222 92370 10274 92382
rect 10222 92306 10274 92318
rect 10334 92370 10386 92382
rect 10334 92306 10386 92318
rect 10558 92370 10610 92382
rect 10558 92306 10610 92318
rect 16830 92370 16882 92382
rect 16830 92306 16882 92318
rect 17726 92370 17778 92382
rect 17726 92306 17778 92318
rect 18510 92370 18562 92382
rect 18510 92306 18562 92318
rect 20414 92370 20466 92382
rect 20414 92306 20466 92318
rect 21310 92370 21362 92382
rect 21310 92306 21362 92318
rect 22430 92370 22482 92382
rect 22430 92306 22482 92318
rect 23998 92370 24050 92382
rect 23998 92306 24050 92318
rect 2494 92258 2546 92270
rect 2494 92194 2546 92206
rect 3278 92258 3330 92270
rect 9774 92258 9826 92270
rect 6738 92206 6750 92258
rect 6802 92206 6814 92258
rect 3278 92194 3330 92206
rect 9774 92194 9826 92206
rect 20302 92258 20354 92270
rect 20302 92194 20354 92206
rect 20638 92258 20690 92270
rect 20638 92194 20690 92206
rect 22318 92258 22370 92270
rect 22318 92194 22370 92206
rect 23102 92258 23154 92270
rect 23102 92194 23154 92206
rect 23550 92258 23602 92270
rect 23550 92194 23602 92206
rect 24110 92258 24162 92270
rect 24110 92194 24162 92206
rect 25230 92258 25282 92270
rect 25230 92194 25282 92206
rect 25454 92258 25506 92270
rect 25454 92194 25506 92206
rect 26798 92258 26850 92270
rect 26798 92194 26850 92206
rect 3054 92146 3106 92158
rect 3054 92082 3106 92094
rect 3390 92146 3442 92158
rect 10110 92146 10162 92158
rect 17502 92146 17554 92158
rect 5058 92094 5070 92146
rect 5122 92094 5134 92146
rect 10994 92094 11006 92146
rect 11058 92094 11070 92146
rect 3390 92082 3442 92094
rect 10110 92082 10162 92094
rect 17502 92082 17554 92094
rect 17838 92146 17890 92158
rect 17838 92082 17890 92094
rect 17950 92146 18002 92158
rect 17950 92082 18002 92094
rect 20750 92146 20802 92158
rect 22542 92146 22594 92158
rect 21970 92094 21982 92146
rect 22034 92094 22046 92146
rect 20750 92082 20802 92094
rect 22542 92082 22594 92094
rect 22878 92146 22930 92158
rect 22878 92082 22930 92094
rect 23326 92146 23378 92158
rect 23326 92082 23378 92094
rect 23886 92146 23938 92158
rect 25790 92146 25842 92158
rect 24322 92094 24334 92146
rect 24386 92094 24398 92146
rect 24658 92094 24670 92146
rect 24722 92094 24734 92146
rect 23886 92082 23938 92094
rect 25790 92082 25842 92094
rect 26238 92146 26290 92158
rect 26238 92082 26290 92094
rect 26462 92146 26514 92158
rect 26462 92082 26514 92094
rect 27358 92146 27410 92158
rect 27358 92082 27410 92094
rect 27582 92146 27634 92158
rect 27582 92082 27634 92094
rect 28030 92146 28082 92158
rect 28030 92082 28082 92094
rect 2830 92034 2882 92046
rect 18958 92034 19010 92046
rect 13458 91982 13470 92034
rect 13522 91982 13534 92034
rect 2830 91970 2882 91982
rect 18958 91970 19010 91982
rect 25678 92034 25730 92046
rect 27470 92034 27522 92046
rect 26674 91982 26686 92034
rect 26738 91982 26750 92034
rect 25678 91970 25730 91982
rect 27470 91970 27522 91982
rect 23438 91922 23490 91934
rect 23438 91858 23490 91870
rect 27022 91922 27074 91934
rect 27022 91858 27074 91870
rect 1344 91754 28560 91788
rect 1344 91702 4616 91754
rect 4668 91702 4720 91754
rect 4772 91702 4824 91754
rect 4876 91702 11420 91754
rect 11472 91702 11524 91754
rect 11576 91702 11628 91754
rect 11680 91702 18224 91754
rect 18276 91702 18328 91754
rect 18380 91702 18432 91754
rect 18484 91702 25028 91754
rect 25080 91702 25132 91754
rect 25184 91702 25236 91754
rect 25288 91702 28560 91754
rect 1344 91668 28560 91702
rect 22878 91586 22930 91598
rect 5730 91534 5742 91586
rect 5794 91534 5806 91586
rect 22878 91522 22930 91534
rect 26126 91586 26178 91598
rect 26126 91522 26178 91534
rect 26350 91586 26402 91598
rect 26350 91522 26402 91534
rect 26462 91586 26514 91598
rect 26462 91522 26514 91534
rect 27246 91586 27298 91598
rect 27246 91522 27298 91534
rect 17278 91474 17330 91486
rect 18958 91474 19010 91486
rect 2482 91422 2494 91474
rect 2546 91422 2558 91474
rect 4610 91422 4622 91474
rect 4674 91422 4686 91474
rect 6066 91422 6078 91474
rect 6130 91422 6142 91474
rect 10770 91422 10782 91474
rect 10834 91422 10846 91474
rect 12674 91422 12686 91474
rect 12738 91422 12750 91474
rect 14578 91422 14590 91474
rect 14642 91422 14654 91474
rect 18050 91422 18062 91474
rect 18114 91422 18126 91474
rect 17278 91410 17330 91422
rect 18958 91410 19010 91422
rect 22990 91474 23042 91486
rect 22990 91410 23042 91422
rect 28142 91474 28194 91486
rect 28142 91410 28194 91422
rect 7310 91362 7362 91374
rect 18846 91362 18898 91374
rect 1810 91310 1822 91362
rect 1874 91310 1886 91362
rect 6514 91310 6526 91362
rect 6578 91310 6590 91362
rect 7970 91310 7982 91362
rect 8034 91310 8046 91362
rect 12786 91310 12798 91362
rect 12850 91310 12862 91362
rect 15474 91310 15486 91362
rect 15538 91310 15550 91362
rect 16034 91310 16046 91362
rect 16098 91310 16110 91362
rect 18498 91310 18510 91362
rect 18562 91310 18574 91362
rect 7310 91298 7362 91310
rect 18846 91298 18898 91310
rect 19182 91362 19234 91374
rect 19182 91298 19234 91310
rect 19406 91362 19458 91374
rect 19406 91298 19458 91310
rect 22206 91362 22258 91374
rect 25566 91362 25618 91374
rect 22306 91310 22318 91362
rect 22370 91310 22382 91362
rect 23538 91310 23550 91362
rect 23602 91310 23614 91362
rect 22206 91298 22258 91310
rect 25566 91298 25618 91310
rect 26910 91362 26962 91374
rect 26910 91298 26962 91310
rect 13582 91250 13634 91262
rect 8642 91198 8654 91250
rect 8706 91198 8718 91250
rect 12898 91198 12910 91250
rect 12962 91198 12974 91250
rect 13582 91186 13634 91198
rect 13694 91250 13746 91262
rect 18062 91250 18114 91262
rect 14242 91198 14254 91250
rect 14306 91198 14318 91250
rect 16370 91198 16382 91250
rect 16434 91198 16446 91250
rect 16818 91198 16830 91250
rect 16882 91198 16894 91250
rect 13694 91186 13746 91198
rect 18062 91186 18114 91198
rect 22094 91250 22146 91262
rect 22094 91186 22146 91198
rect 22542 91250 22594 91262
rect 22542 91186 22594 91198
rect 23774 91250 23826 91262
rect 23774 91186 23826 91198
rect 23998 91250 24050 91262
rect 23998 91186 24050 91198
rect 24222 91250 24274 91262
rect 24222 91186 24274 91198
rect 24334 91250 24386 91262
rect 24334 91186 24386 91198
rect 25118 91250 25170 91262
rect 25118 91186 25170 91198
rect 25678 91250 25730 91262
rect 25678 91186 25730 91198
rect 26014 91250 26066 91262
rect 26014 91186 26066 91198
rect 5070 91138 5122 91150
rect 5070 91074 5122 91086
rect 6974 91138 7026 91150
rect 6974 91074 7026 91086
rect 7198 91138 7250 91150
rect 7198 91074 7250 91086
rect 11454 91138 11506 91150
rect 11454 91074 11506 91086
rect 12014 91138 12066 91150
rect 12014 91074 12066 91086
rect 13358 91138 13410 91150
rect 13358 91074 13410 91086
rect 17950 91138 18002 91150
rect 17950 91074 18002 91086
rect 18286 91138 18338 91150
rect 18286 91074 18338 91086
rect 23214 91138 23266 91150
rect 23214 91074 23266 91086
rect 23326 91138 23378 91150
rect 23326 91074 23378 91086
rect 25230 91138 25282 91150
rect 25230 91074 25282 91086
rect 27134 91138 27186 91150
rect 27134 91074 27186 91086
rect 1344 90970 28720 91004
rect 1344 90918 8018 90970
rect 8070 90918 8122 90970
rect 8174 90918 8226 90970
rect 8278 90918 14822 90970
rect 14874 90918 14926 90970
rect 14978 90918 15030 90970
rect 15082 90918 21626 90970
rect 21678 90918 21730 90970
rect 21782 90918 21834 90970
rect 21886 90918 28430 90970
rect 28482 90918 28534 90970
rect 28586 90918 28638 90970
rect 28690 90918 28720 90970
rect 1344 90884 28720 90918
rect 4734 90802 4786 90814
rect 4734 90738 4786 90750
rect 8654 90802 8706 90814
rect 8654 90738 8706 90750
rect 11454 90802 11506 90814
rect 11454 90738 11506 90750
rect 15710 90802 15762 90814
rect 15710 90738 15762 90750
rect 19406 90802 19458 90814
rect 19406 90738 19458 90750
rect 19966 90802 20018 90814
rect 19966 90738 20018 90750
rect 22766 90802 22818 90814
rect 22766 90738 22818 90750
rect 4510 90690 4562 90702
rect 4510 90626 4562 90638
rect 5294 90690 5346 90702
rect 5294 90626 5346 90638
rect 5742 90690 5794 90702
rect 5742 90626 5794 90638
rect 7534 90690 7586 90702
rect 7534 90626 7586 90638
rect 8430 90690 8482 90702
rect 8430 90626 8482 90638
rect 8766 90690 8818 90702
rect 8766 90626 8818 90638
rect 9662 90690 9714 90702
rect 9662 90626 9714 90638
rect 10558 90690 10610 90702
rect 10558 90626 10610 90638
rect 10894 90690 10946 90702
rect 10894 90626 10946 90638
rect 11902 90690 11954 90702
rect 11902 90626 11954 90638
rect 14030 90690 14082 90702
rect 14030 90626 14082 90638
rect 14702 90690 14754 90702
rect 14702 90626 14754 90638
rect 14926 90690 14978 90702
rect 14926 90626 14978 90638
rect 20078 90690 20130 90702
rect 20078 90626 20130 90638
rect 21870 90690 21922 90702
rect 21870 90626 21922 90638
rect 22878 90690 22930 90702
rect 22878 90626 22930 90638
rect 23438 90690 23490 90702
rect 23438 90626 23490 90638
rect 23550 90690 23602 90702
rect 23550 90626 23602 90638
rect 6974 90578 7026 90590
rect 6402 90526 6414 90578
rect 6466 90526 6478 90578
rect 6974 90514 7026 90526
rect 7086 90578 7138 90590
rect 7086 90514 7138 90526
rect 7422 90578 7474 90590
rect 7422 90514 7474 90526
rect 7758 90578 7810 90590
rect 7758 90514 7810 90526
rect 8990 90578 9042 90590
rect 8990 90514 9042 90526
rect 9774 90578 9826 90590
rect 9774 90514 9826 90526
rect 9886 90578 9938 90590
rect 9886 90514 9938 90526
rect 10334 90578 10386 90590
rect 10334 90514 10386 90526
rect 11118 90578 11170 90590
rect 11118 90514 11170 90526
rect 11678 90578 11730 90590
rect 11678 90514 11730 90526
rect 12686 90578 12738 90590
rect 15150 90578 15202 90590
rect 13458 90526 13470 90578
rect 13522 90526 13534 90578
rect 12686 90514 12738 90526
rect 15150 90514 15202 90526
rect 15374 90578 15426 90590
rect 15374 90514 15426 90526
rect 15598 90578 15650 90590
rect 20190 90578 20242 90590
rect 20638 90578 20690 90590
rect 19730 90526 19742 90578
rect 19794 90526 19806 90578
rect 20402 90526 20414 90578
rect 20466 90526 20478 90578
rect 15598 90514 15650 90526
rect 20190 90514 20242 90526
rect 20638 90514 20690 90526
rect 21086 90578 21138 90590
rect 21086 90514 21138 90526
rect 21310 90578 21362 90590
rect 21310 90514 21362 90526
rect 21646 90578 21698 90590
rect 21646 90514 21698 90526
rect 21982 90578 22034 90590
rect 21982 90514 22034 90526
rect 22542 90578 22594 90590
rect 27582 90578 27634 90590
rect 27010 90526 27022 90578
rect 27074 90526 27086 90578
rect 22542 90514 22594 90526
rect 27582 90514 27634 90526
rect 8094 90466 8146 90478
rect 8094 90402 8146 90414
rect 10670 90466 10722 90478
rect 10670 90402 10722 90414
rect 11566 90466 11618 90478
rect 11566 90402 11618 90414
rect 12350 90466 12402 90478
rect 12350 90402 12402 90414
rect 12910 90466 12962 90478
rect 16270 90466 16322 90478
rect 13346 90414 13358 90466
rect 13410 90414 13422 90466
rect 12910 90402 12962 90414
rect 16270 90402 16322 90414
rect 16606 90466 16658 90478
rect 16606 90402 16658 90414
rect 17614 90466 17666 90478
rect 17614 90402 17666 90414
rect 17950 90466 18002 90478
rect 17950 90402 18002 90414
rect 18398 90466 18450 90478
rect 18398 90402 18450 90414
rect 20862 90466 20914 90478
rect 28018 90414 28030 90466
rect 28082 90414 28094 90466
rect 20862 90402 20914 90414
rect 23438 90354 23490 90366
rect 17938 90302 17950 90354
rect 18002 90351 18014 90354
rect 18386 90351 18398 90354
rect 18002 90305 18398 90351
rect 18002 90302 18014 90305
rect 18386 90302 18398 90305
rect 18450 90302 18462 90354
rect 23438 90290 23490 90302
rect 27134 90354 27186 90366
rect 27134 90290 27186 90302
rect 1344 90186 28560 90220
rect 1344 90134 4616 90186
rect 4668 90134 4720 90186
rect 4772 90134 4824 90186
rect 4876 90134 11420 90186
rect 11472 90134 11524 90186
rect 11576 90134 11628 90186
rect 11680 90134 18224 90186
rect 18276 90134 18328 90186
rect 18380 90134 18432 90186
rect 18484 90134 25028 90186
rect 25080 90134 25132 90186
rect 25184 90134 25236 90186
rect 25288 90134 28560 90186
rect 1344 90100 28560 90134
rect 18846 90018 18898 90030
rect 18846 89954 18898 89966
rect 23214 90018 23266 90030
rect 23214 89954 23266 89966
rect 4846 89906 4898 89918
rect 4846 89842 4898 89854
rect 5854 89906 5906 89918
rect 9550 89906 9602 89918
rect 7970 89854 7982 89906
rect 8034 89854 8046 89906
rect 5854 89842 5906 89854
rect 9550 89842 9602 89854
rect 9998 89906 10050 89918
rect 13918 89906 13970 89918
rect 12450 89854 12462 89906
rect 12514 89854 12526 89906
rect 9998 89842 10050 89854
rect 13918 89842 13970 89854
rect 15038 89906 15090 89918
rect 15474 89854 15486 89906
rect 15538 89854 15550 89906
rect 15038 89842 15090 89854
rect 13582 89794 13634 89806
rect 8642 89742 8654 89794
rect 8706 89742 8718 89794
rect 10770 89742 10782 89794
rect 10834 89742 10846 89794
rect 13582 89730 13634 89742
rect 13806 89794 13858 89806
rect 13806 89730 13858 89742
rect 14590 89794 14642 89806
rect 14590 89730 14642 89742
rect 15262 89794 15314 89806
rect 19630 89794 19682 89806
rect 15698 89742 15710 89794
rect 15762 89742 15774 89794
rect 16594 89742 16606 89794
rect 16658 89742 16670 89794
rect 17714 89742 17726 89794
rect 17778 89742 17790 89794
rect 15262 89730 15314 89742
rect 19630 89730 19682 89742
rect 20190 89794 20242 89806
rect 20190 89730 20242 89742
rect 21758 89794 21810 89806
rect 21758 89730 21810 89742
rect 22542 89794 22594 89806
rect 22542 89730 22594 89742
rect 22878 89794 22930 89806
rect 22878 89730 22930 89742
rect 24222 89794 24274 89806
rect 24222 89730 24274 89742
rect 24558 89794 24610 89806
rect 26114 89742 26126 89794
rect 26178 89742 26190 89794
rect 27010 89742 27022 89794
rect 27074 89742 27086 89794
rect 24558 89730 24610 89742
rect 14030 89682 14082 89694
rect 14030 89618 14082 89630
rect 14814 89682 14866 89694
rect 19966 89682 20018 89694
rect 15810 89630 15822 89682
rect 15874 89630 15886 89682
rect 16258 89630 16270 89682
rect 16322 89630 16334 89682
rect 14814 89618 14866 89630
rect 19966 89618 20018 89630
rect 21870 89682 21922 89694
rect 21870 89618 21922 89630
rect 22766 89682 22818 89694
rect 22766 89618 22818 89630
rect 23326 89682 23378 89694
rect 23326 89618 23378 89630
rect 23998 89682 24050 89694
rect 24882 89630 24894 89682
rect 24946 89630 24958 89682
rect 27234 89630 27246 89682
rect 27298 89630 27310 89682
rect 23998 89618 24050 89630
rect 18062 89570 18114 89582
rect 18062 89506 18114 89518
rect 19294 89570 19346 89582
rect 19294 89506 19346 89518
rect 19742 89570 19794 89582
rect 19742 89506 19794 89518
rect 21982 89570 22034 89582
rect 21982 89506 22034 89518
rect 22206 89570 22258 89582
rect 22206 89506 22258 89518
rect 24110 89570 24162 89582
rect 26002 89518 26014 89570
rect 26066 89518 26078 89570
rect 24110 89506 24162 89518
rect 1344 89402 28720 89436
rect 1344 89350 8018 89402
rect 8070 89350 8122 89402
rect 8174 89350 8226 89402
rect 8278 89350 14822 89402
rect 14874 89350 14926 89402
rect 14978 89350 15030 89402
rect 15082 89350 21626 89402
rect 21678 89350 21730 89402
rect 21782 89350 21834 89402
rect 21886 89350 28430 89402
rect 28482 89350 28534 89402
rect 28586 89350 28638 89402
rect 28690 89350 28720 89402
rect 1344 89316 28720 89350
rect 18622 89234 18674 89246
rect 18622 89170 18674 89182
rect 18846 89234 18898 89246
rect 18846 89170 18898 89182
rect 21646 89234 21698 89246
rect 21646 89170 21698 89182
rect 22430 89234 22482 89246
rect 22430 89170 22482 89182
rect 15710 89122 15762 89134
rect 15710 89058 15762 89070
rect 15822 89122 15874 89134
rect 25566 89122 25618 89134
rect 15822 89058 15874 89070
rect 15934 89066 15986 89078
rect 23314 89070 23326 89122
rect 23378 89070 23390 89122
rect 27122 89070 27134 89122
rect 27186 89070 27198 89122
rect 5070 89010 5122 89022
rect 4610 88958 4622 89010
rect 4674 88958 4686 89010
rect 5070 88946 5122 88958
rect 6862 89010 6914 89022
rect 6862 88946 6914 88958
rect 7198 89010 7250 89022
rect 7198 88946 7250 88958
rect 7758 89010 7810 89022
rect 7758 88946 7810 88958
rect 8654 89010 8706 89022
rect 25566 89058 25618 89070
rect 10098 88958 10110 89010
rect 10162 88958 10174 89010
rect 15934 89002 15986 89014
rect 16830 89010 16882 89022
rect 16370 88958 16382 89010
rect 16434 88958 16446 89010
rect 8654 88946 8706 88958
rect 16830 88946 16882 88958
rect 17502 89010 17554 89022
rect 17502 88946 17554 88958
rect 17950 89010 18002 89022
rect 17950 88946 18002 88958
rect 18174 89010 18226 89022
rect 18174 88946 18226 88958
rect 18734 89010 18786 89022
rect 18734 88946 18786 88958
rect 18958 89010 19010 89022
rect 21422 89010 21474 89022
rect 19170 88958 19182 89010
rect 19234 88958 19246 89010
rect 18958 88946 19010 88958
rect 21422 88946 21474 88958
rect 22094 89010 22146 89022
rect 25118 89010 25170 89022
rect 23538 88958 23550 89010
rect 23602 88958 23614 89010
rect 22094 88946 22146 88958
rect 25118 88946 25170 88958
rect 25342 89010 25394 89022
rect 25342 88946 25394 88958
rect 25790 89010 25842 89022
rect 25790 88946 25842 88958
rect 26350 89010 26402 89022
rect 28130 88958 28142 89010
rect 28194 88958 28206 89010
rect 26350 88946 26402 88958
rect 8094 88898 8146 88910
rect 1698 88846 1710 88898
rect 1762 88846 1774 88898
rect 3826 88846 3838 88898
rect 3890 88846 3902 88898
rect 8094 88834 8146 88846
rect 9102 88898 9154 88910
rect 17726 88898 17778 88910
rect 13346 88846 13358 88898
rect 13410 88846 13422 88898
rect 9102 88834 9154 88846
rect 17726 88834 17778 88846
rect 19630 88898 19682 88910
rect 19630 88834 19682 88846
rect 21534 88898 21586 88910
rect 21534 88834 21586 88846
rect 24558 88898 24610 88910
rect 24558 88834 24610 88846
rect 26238 88898 26290 88910
rect 27122 88846 27134 88898
rect 27186 88846 27198 88898
rect 26238 88834 26290 88846
rect 22766 88786 22818 88798
rect 7074 88734 7086 88786
rect 7138 88783 7150 88786
rect 8194 88783 8206 88786
rect 7138 88737 8206 88783
rect 7138 88734 7150 88737
rect 8194 88734 8206 88737
rect 8258 88734 8270 88786
rect 19394 88734 19406 88786
rect 19458 88783 19470 88786
rect 19730 88783 19742 88786
rect 19458 88737 19742 88783
rect 19458 88734 19470 88737
rect 19730 88734 19742 88737
rect 19794 88734 19806 88786
rect 22766 88722 22818 88734
rect 23998 88786 24050 88798
rect 23998 88722 24050 88734
rect 24334 88786 24386 88798
rect 24334 88722 24386 88734
rect 1344 88618 28560 88652
rect 1344 88566 4616 88618
rect 4668 88566 4720 88618
rect 4772 88566 4824 88618
rect 4876 88566 11420 88618
rect 11472 88566 11524 88618
rect 11576 88566 11628 88618
rect 11680 88566 18224 88618
rect 18276 88566 18328 88618
rect 18380 88566 18432 88618
rect 18484 88566 25028 88618
rect 25080 88566 25132 88618
rect 25184 88566 25236 88618
rect 25288 88566 28560 88618
rect 1344 88532 28560 88566
rect 22990 88450 23042 88462
rect 5618 88398 5630 88450
rect 5682 88447 5694 88450
rect 6626 88447 6638 88450
rect 5682 88401 6638 88447
rect 5682 88398 5694 88401
rect 6626 88398 6638 88401
rect 6690 88398 6702 88450
rect 6850 88398 6862 88450
rect 6914 88447 6926 88450
rect 7746 88447 7758 88450
rect 6914 88401 7758 88447
rect 6914 88398 6926 88401
rect 7746 88398 7758 88401
rect 7810 88398 7822 88450
rect 22642 88398 22654 88450
rect 22706 88398 22718 88450
rect 24770 88398 24782 88450
rect 24834 88398 24846 88450
rect 22990 88386 23042 88398
rect 5742 88338 5794 88350
rect 5742 88274 5794 88286
rect 6190 88338 6242 88350
rect 6190 88274 6242 88286
rect 6638 88338 6690 88350
rect 6638 88274 6690 88286
rect 7198 88338 7250 88350
rect 7198 88274 7250 88286
rect 8094 88338 8146 88350
rect 20078 88338 20130 88350
rect 10770 88286 10782 88338
rect 10834 88286 10846 88338
rect 12898 88286 12910 88338
rect 12962 88286 12974 88338
rect 16818 88286 16830 88338
rect 16882 88286 16894 88338
rect 19730 88286 19742 88338
rect 19794 88286 19806 88338
rect 8094 88274 8146 88286
rect 20078 88274 20130 88286
rect 20526 88338 20578 88350
rect 20526 88274 20578 88286
rect 23214 88338 23266 88350
rect 23214 88274 23266 88286
rect 8206 88226 8258 88238
rect 8206 88162 8258 88174
rect 8542 88226 8594 88238
rect 8542 88162 8594 88174
rect 9102 88226 9154 88238
rect 18286 88226 18338 88238
rect 9538 88174 9550 88226
rect 9602 88174 9614 88226
rect 10098 88174 10110 88226
rect 10162 88174 10174 88226
rect 13458 88174 13470 88226
rect 13522 88174 13534 88226
rect 9102 88162 9154 88174
rect 18286 88162 18338 88174
rect 19294 88226 19346 88238
rect 24558 88226 24610 88238
rect 26462 88226 26514 88238
rect 20738 88174 20750 88226
rect 20802 88174 20814 88226
rect 24994 88174 25006 88226
rect 25058 88174 25070 88226
rect 26786 88174 26798 88226
rect 26850 88174 26862 88226
rect 19294 88162 19346 88174
rect 24558 88162 24610 88174
rect 26462 88162 26514 88174
rect 1710 88114 1762 88126
rect 1710 88050 1762 88062
rect 2494 88114 2546 88126
rect 2494 88050 2546 88062
rect 2830 88114 2882 88126
rect 2830 88050 2882 88062
rect 7758 88114 7810 88126
rect 7758 88050 7810 88062
rect 7982 88114 8034 88126
rect 7982 88050 8034 88062
rect 9214 88114 9266 88126
rect 9214 88050 9266 88062
rect 17726 88114 17778 88126
rect 17726 88050 17778 88062
rect 18062 88114 18114 88126
rect 18062 88050 18114 88062
rect 18510 88114 18562 88126
rect 18510 88050 18562 88062
rect 18622 88114 18674 88126
rect 18622 88050 18674 88062
rect 19182 88114 19234 88126
rect 19182 88050 19234 88062
rect 19854 88114 19906 88126
rect 19854 88050 19906 88062
rect 20414 88114 20466 88126
rect 20414 88050 20466 88062
rect 3390 88002 3442 88014
rect 2034 87950 2046 88002
rect 2098 87950 2110 88002
rect 3390 87938 3442 87950
rect 8990 88002 9042 88014
rect 8990 87938 9042 87950
rect 1344 87834 28720 87868
rect 1344 87782 8018 87834
rect 8070 87782 8122 87834
rect 8174 87782 8226 87834
rect 8278 87782 14822 87834
rect 14874 87782 14926 87834
rect 14978 87782 15030 87834
rect 15082 87782 21626 87834
rect 21678 87782 21730 87834
rect 21782 87782 21834 87834
rect 21886 87782 28430 87834
rect 28482 87782 28534 87834
rect 28586 87782 28638 87834
rect 28690 87782 28720 87834
rect 1344 87748 28720 87782
rect 1822 87666 1874 87678
rect 1822 87602 1874 87614
rect 15150 87666 15202 87678
rect 15150 87602 15202 87614
rect 16606 87666 16658 87678
rect 16606 87602 16658 87614
rect 17502 87666 17554 87678
rect 17502 87602 17554 87614
rect 18846 87666 18898 87678
rect 18846 87602 18898 87614
rect 19966 87666 20018 87678
rect 27582 87666 27634 87678
rect 26114 87614 26126 87666
rect 26178 87614 26190 87666
rect 19966 87602 20018 87614
rect 27582 87602 27634 87614
rect 4734 87554 4786 87566
rect 13806 87554 13858 87566
rect 6850 87502 6862 87554
rect 6914 87502 6926 87554
rect 4734 87490 4786 87502
rect 13806 87490 13858 87502
rect 15262 87554 15314 87566
rect 15262 87490 15314 87502
rect 15822 87554 15874 87566
rect 15822 87490 15874 87502
rect 24670 87554 24722 87566
rect 24670 87490 24722 87502
rect 5630 87442 5682 87454
rect 14030 87442 14082 87454
rect 5394 87390 5406 87442
rect 5458 87390 5470 87442
rect 6066 87390 6078 87442
rect 6130 87390 6142 87442
rect 9538 87390 9550 87442
rect 9602 87390 9614 87442
rect 5630 87378 5682 87390
rect 14030 87378 14082 87390
rect 14478 87442 14530 87454
rect 14478 87378 14530 87390
rect 14702 87442 14754 87454
rect 14702 87378 14754 87390
rect 14926 87442 14978 87454
rect 25790 87442 25842 87454
rect 18386 87390 18398 87442
rect 18450 87390 18462 87442
rect 24098 87390 24110 87442
rect 24162 87390 24174 87442
rect 14926 87378 14978 87390
rect 25790 87378 25842 87390
rect 27134 87442 27186 87454
rect 27134 87378 27186 87390
rect 27358 87442 27410 87454
rect 27358 87378 27410 87390
rect 4510 87330 4562 87342
rect 13918 87330 13970 87342
rect 8978 87278 8990 87330
rect 9042 87278 9054 87330
rect 13234 87278 13246 87330
rect 13298 87278 13310 87330
rect 4510 87266 4562 87278
rect 13918 87266 13970 87278
rect 15934 87330 15986 87342
rect 15934 87266 15986 87278
rect 16046 87330 16098 87342
rect 17838 87330 17890 87342
rect 16706 87278 16718 87330
rect 16770 87278 16782 87330
rect 16046 87266 16098 87278
rect 17838 87266 17890 87278
rect 19518 87330 19570 87342
rect 19518 87266 19570 87278
rect 20302 87330 20354 87342
rect 20302 87266 20354 87278
rect 20862 87330 20914 87342
rect 20862 87266 20914 87278
rect 21310 87330 21362 87342
rect 21310 87266 21362 87278
rect 21758 87330 21810 87342
rect 25566 87330 25618 87342
rect 28142 87330 28194 87342
rect 24322 87278 24334 87330
rect 24386 87278 24398 87330
rect 27458 87278 27470 87330
rect 27522 87278 27534 87330
rect 21758 87266 21810 87278
rect 25566 87266 25618 87278
rect 28142 87266 28194 87278
rect 16382 87218 16434 87230
rect 16382 87154 16434 87166
rect 18062 87218 18114 87230
rect 26686 87218 26738 87230
rect 20850 87166 20862 87218
rect 20914 87215 20926 87218
rect 21746 87215 21758 87218
rect 20914 87169 21758 87215
rect 20914 87166 20926 87169
rect 21746 87166 21758 87169
rect 21810 87166 21822 87218
rect 18062 87154 18114 87166
rect 26686 87154 26738 87166
rect 26910 87218 26962 87230
rect 26910 87154 26962 87166
rect 1344 87050 28560 87084
rect 1344 86998 4616 87050
rect 4668 86998 4720 87050
rect 4772 86998 4824 87050
rect 4876 86998 11420 87050
rect 11472 86998 11524 87050
rect 11576 86998 11628 87050
rect 11680 86998 18224 87050
rect 18276 86998 18328 87050
rect 18380 86998 18432 87050
rect 18484 86998 25028 87050
rect 25080 86998 25132 87050
rect 25184 86998 25236 87050
rect 25288 86998 28560 87050
rect 1344 86964 28560 86998
rect 4510 86882 4562 86894
rect 18958 86882 19010 86894
rect 7074 86830 7086 86882
rect 7138 86879 7150 86882
rect 7858 86879 7870 86882
rect 7138 86833 7870 86879
rect 7138 86830 7150 86833
rect 7858 86830 7870 86833
rect 7922 86830 7934 86882
rect 4510 86818 4562 86830
rect 18958 86818 19010 86830
rect 19742 86882 19794 86894
rect 23986 86830 23998 86882
rect 24050 86830 24062 86882
rect 19742 86818 19794 86830
rect 4734 86770 4786 86782
rect 4734 86706 4786 86718
rect 6078 86770 6130 86782
rect 6078 86706 6130 86718
rect 6526 86770 6578 86782
rect 6526 86706 6578 86718
rect 7086 86770 7138 86782
rect 7086 86706 7138 86718
rect 7870 86770 7922 86782
rect 7870 86706 7922 86718
rect 8430 86770 8482 86782
rect 16482 86718 16494 86770
rect 16546 86718 16558 86770
rect 24098 86718 24110 86770
rect 24162 86718 24174 86770
rect 8430 86706 8482 86718
rect 7534 86658 7586 86670
rect 7534 86594 7586 86606
rect 8990 86658 9042 86670
rect 12238 86658 12290 86670
rect 19182 86658 19234 86670
rect 10098 86606 10110 86658
rect 10162 86606 10174 86658
rect 12562 86606 12574 86658
rect 12626 86606 12638 86658
rect 15026 86606 15038 86658
rect 15090 86606 15102 86658
rect 15698 86606 15710 86658
rect 15762 86606 15774 86658
rect 17266 86606 17278 86658
rect 17330 86606 17342 86658
rect 21298 86606 21310 86658
rect 21362 86606 21374 86658
rect 21858 86606 21870 86658
rect 21922 86606 21934 86658
rect 24994 86606 25006 86658
rect 25058 86606 25070 86658
rect 26002 86606 26014 86658
rect 26066 86606 26078 86658
rect 27234 86606 27246 86658
rect 27298 86606 27310 86658
rect 27906 86606 27918 86658
rect 27970 86606 27982 86658
rect 8990 86594 9042 86606
rect 12238 86594 12290 86606
rect 19182 86594 19234 86606
rect 3838 86546 3890 86558
rect 3838 86482 3890 86494
rect 8654 86546 8706 86558
rect 8654 86482 8706 86494
rect 9214 86546 9266 86558
rect 9214 86482 9266 86494
rect 10894 86546 10946 86558
rect 10894 86482 10946 86494
rect 11230 86546 11282 86558
rect 19518 86546 19570 86558
rect 16370 86494 16382 86546
rect 16434 86494 16446 86546
rect 11230 86482 11282 86494
rect 19518 86482 19570 86494
rect 20078 86546 20130 86558
rect 22878 86546 22930 86558
rect 21970 86494 21982 86546
rect 22034 86494 22046 86546
rect 20078 86482 20130 86494
rect 22878 86482 22930 86494
rect 3502 86434 3554 86446
rect 8766 86434 8818 86446
rect 4162 86382 4174 86434
rect 4226 86382 4238 86434
rect 3502 86370 3554 86382
rect 8766 86370 8818 86382
rect 9550 86434 9602 86446
rect 9550 86370 9602 86382
rect 9662 86434 9714 86446
rect 9662 86370 9714 86382
rect 9774 86434 9826 86446
rect 9774 86370 9826 86382
rect 10782 86434 10834 86446
rect 10782 86370 10834 86382
rect 11006 86434 11058 86446
rect 11006 86370 11058 86382
rect 12014 86434 12066 86446
rect 12014 86370 12066 86382
rect 12126 86434 12178 86446
rect 18846 86434 18898 86446
rect 15026 86382 15038 86434
rect 15090 86382 15102 86434
rect 12126 86370 12178 86382
rect 18846 86370 18898 86382
rect 20190 86434 20242 86446
rect 20190 86370 20242 86382
rect 20414 86434 20466 86446
rect 20414 86370 20466 86382
rect 20750 86434 20802 86446
rect 21522 86382 21534 86434
rect 21586 86382 21598 86434
rect 20750 86370 20802 86382
rect 1344 86266 28720 86300
rect 1344 86214 8018 86266
rect 8070 86214 8122 86266
rect 8174 86214 8226 86266
rect 8278 86214 14822 86266
rect 14874 86214 14926 86266
rect 14978 86214 15030 86266
rect 15082 86214 21626 86266
rect 21678 86214 21730 86266
rect 21782 86214 21834 86266
rect 21886 86214 28430 86266
rect 28482 86214 28534 86266
rect 28586 86214 28638 86266
rect 28690 86214 28720 86266
rect 1344 86180 28720 86214
rect 7310 86098 7362 86110
rect 7310 86034 7362 86046
rect 15262 86098 15314 86110
rect 15262 86034 15314 86046
rect 24446 86098 24498 86110
rect 24446 86034 24498 86046
rect 25678 86098 25730 86110
rect 25778 86046 25790 86098
rect 25842 86046 25854 86098
rect 25678 86034 25730 86046
rect 8094 85986 8146 85998
rect 2034 85934 2046 85986
rect 2098 85934 2110 85986
rect 3714 85934 3726 85986
rect 3778 85934 3790 85986
rect 8094 85922 8146 85934
rect 8654 85986 8706 85998
rect 15934 85986 15986 85998
rect 10770 85934 10782 85986
rect 10834 85934 10846 85986
rect 8654 85922 8706 85934
rect 15934 85922 15986 85934
rect 16158 85986 16210 85998
rect 16158 85922 16210 85934
rect 16382 85986 16434 85998
rect 23886 85986 23938 85998
rect 27806 85986 27858 85998
rect 22978 85934 22990 85986
rect 23042 85934 23054 85986
rect 26450 85934 26462 85986
rect 26514 85934 26526 85986
rect 16382 85922 16434 85934
rect 23886 85922 23938 85934
rect 27806 85922 27858 85934
rect 1710 85874 1762 85886
rect 7758 85874 7810 85886
rect 3042 85822 3054 85874
rect 3106 85822 3118 85874
rect 1710 85810 1762 85822
rect 7758 85810 7810 85822
rect 8318 85874 8370 85886
rect 13458 85822 13470 85874
rect 13522 85822 13534 85874
rect 19394 85822 19406 85874
rect 19458 85822 19470 85874
rect 25442 85822 25454 85874
rect 25506 85822 25518 85874
rect 26338 85822 26350 85874
rect 26402 85822 26414 85874
rect 27234 85822 27246 85874
rect 27298 85822 27310 85874
rect 8318 85810 8370 85822
rect 2494 85762 2546 85774
rect 2494 85698 2546 85710
rect 5854 85762 5906 85774
rect 5854 85698 5906 85710
rect 6974 85762 7026 85774
rect 6974 85698 7026 85710
rect 8206 85762 8258 85774
rect 8206 85698 8258 85710
rect 17838 85762 17890 85774
rect 17838 85698 17890 85710
rect 24558 85762 24610 85774
rect 24558 85698 24610 85710
rect 24670 85762 24722 85774
rect 24670 85698 24722 85710
rect 23998 85650 24050 85662
rect 7186 85598 7198 85650
rect 7250 85647 7262 85650
rect 7858 85647 7870 85650
rect 7250 85601 7870 85647
rect 7250 85598 7262 85601
rect 7858 85598 7870 85601
rect 7922 85598 7934 85650
rect 16706 85598 16718 85650
rect 16770 85598 16782 85650
rect 23998 85586 24050 85598
rect 27470 85650 27522 85662
rect 27470 85586 27522 85598
rect 27694 85650 27746 85662
rect 27694 85586 27746 85598
rect 1344 85482 28560 85516
rect 1344 85430 4616 85482
rect 4668 85430 4720 85482
rect 4772 85430 4824 85482
rect 4876 85430 11420 85482
rect 11472 85430 11524 85482
rect 11576 85430 11628 85482
rect 11680 85430 18224 85482
rect 18276 85430 18328 85482
rect 18380 85430 18432 85482
rect 18484 85430 25028 85482
rect 25080 85430 25132 85482
rect 25184 85430 25236 85482
rect 25288 85430 28560 85482
rect 1344 85396 28560 85430
rect 17390 85314 17442 85326
rect 17390 85250 17442 85262
rect 18174 85314 18226 85326
rect 18174 85250 18226 85262
rect 19182 85314 19234 85326
rect 19182 85250 19234 85262
rect 20638 85314 20690 85326
rect 24670 85314 24722 85326
rect 25454 85314 25506 85326
rect 22978 85262 22990 85314
rect 23042 85311 23054 85314
rect 23314 85311 23326 85314
rect 23042 85265 23326 85311
rect 23042 85262 23054 85265
rect 23314 85262 23326 85265
rect 23378 85262 23390 85314
rect 25106 85262 25118 85314
rect 25170 85262 25182 85314
rect 20638 85250 20690 85262
rect 24670 85250 24722 85262
rect 25454 85250 25506 85262
rect 23326 85202 23378 85214
rect 3938 85150 3950 85202
rect 4002 85150 4014 85202
rect 7186 85150 7198 85202
rect 7250 85150 7262 85202
rect 9314 85150 9326 85202
rect 9378 85150 9390 85202
rect 14466 85150 14478 85202
rect 14530 85150 14542 85202
rect 16594 85150 16606 85202
rect 16658 85150 16670 85202
rect 17602 85150 17614 85202
rect 17666 85150 17678 85202
rect 21970 85150 21982 85202
rect 22034 85150 22046 85202
rect 23326 85138 23378 85150
rect 24222 85202 24274 85214
rect 26562 85150 26574 85202
rect 26626 85150 26638 85202
rect 24222 85138 24274 85150
rect 12574 85090 12626 85102
rect 17950 85090 18002 85102
rect 25678 85090 25730 85102
rect 3042 85038 3054 85090
rect 3106 85038 3118 85090
rect 6514 85038 6526 85090
rect 6578 85038 6590 85090
rect 9650 85038 9662 85090
rect 9714 85038 9726 85090
rect 13794 85038 13806 85090
rect 13858 85038 13870 85090
rect 18610 85038 18622 85090
rect 18674 85038 18686 85090
rect 22306 85038 22318 85090
rect 22370 85038 22382 85090
rect 26226 85038 26238 85090
rect 26290 85038 26302 85090
rect 27010 85038 27022 85090
rect 27074 85038 27086 85090
rect 12574 85026 12626 85038
rect 17950 85026 18002 85038
rect 25678 85026 25730 85038
rect 12798 84978 12850 84990
rect 11442 84926 11454 84978
rect 11506 84926 11518 84978
rect 12798 84914 12850 84926
rect 12910 84978 12962 84990
rect 12910 84914 12962 84926
rect 17166 84978 17218 84990
rect 17166 84914 17218 84926
rect 17614 84978 17666 84990
rect 17614 84914 17666 84926
rect 20750 84978 20802 84990
rect 20750 84914 20802 84926
rect 21310 84978 21362 84990
rect 21310 84914 21362 84926
rect 22766 84978 22818 84990
rect 22766 84914 22818 84926
rect 24782 84978 24834 84990
rect 27358 84978 27410 84990
rect 27122 84926 27134 84978
rect 27186 84926 27198 84978
rect 24782 84914 24834 84926
rect 27358 84914 27410 84926
rect 27470 84978 27522 84990
rect 27470 84914 27522 84926
rect 27918 84978 27970 84990
rect 27918 84914 27970 84926
rect 6078 84866 6130 84878
rect 6078 84802 6130 84814
rect 20638 84866 20690 84878
rect 20638 84802 20690 84814
rect 21422 84866 21474 84878
rect 21422 84802 21474 84814
rect 23662 84866 23714 84878
rect 23662 84802 23714 84814
rect 24670 84866 24722 84878
rect 24670 84802 24722 84814
rect 27694 84866 27746 84878
rect 27694 84802 27746 84814
rect 1344 84698 28720 84732
rect 1344 84646 8018 84698
rect 8070 84646 8122 84698
rect 8174 84646 8226 84698
rect 8278 84646 14822 84698
rect 14874 84646 14926 84698
rect 14978 84646 15030 84698
rect 15082 84646 21626 84698
rect 21678 84646 21730 84698
rect 21782 84646 21834 84698
rect 21886 84646 28430 84698
rect 28482 84646 28534 84698
rect 28586 84646 28638 84698
rect 28690 84646 28720 84698
rect 1344 84612 28720 84646
rect 5742 84530 5794 84542
rect 5742 84466 5794 84478
rect 8990 84530 9042 84542
rect 19854 84530 19906 84542
rect 14018 84478 14030 84530
rect 14082 84478 14094 84530
rect 8990 84466 9042 84478
rect 19854 84466 19906 84478
rect 19966 84530 20018 84542
rect 19966 84466 20018 84478
rect 10222 84418 10274 84430
rect 20078 84418 20130 84430
rect 26238 84418 26290 84430
rect 11778 84366 11790 84418
rect 11842 84366 11854 84418
rect 15362 84366 15374 84418
rect 15426 84366 15438 84418
rect 20178 84366 20190 84418
rect 20242 84366 20254 84418
rect 22866 84366 22878 84418
rect 22930 84366 22942 84418
rect 10222 84354 10274 84366
rect 20078 84354 20130 84366
rect 26238 84354 26290 84366
rect 26574 84418 26626 84430
rect 26574 84354 26626 84366
rect 10670 84306 10722 84318
rect 19742 84306 19794 84318
rect 11106 84254 11118 84306
rect 11170 84254 11182 84306
rect 14466 84254 14478 84306
rect 14530 84254 14542 84306
rect 17602 84254 17614 84306
rect 17666 84254 17678 84306
rect 10670 84242 10722 84254
rect 19742 84242 19794 84254
rect 20862 84306 20914 84318
rect 20862 84242 20914 84254
rect 21086 84306 21138 84318
rect 24446 84306 24498 84318
rect 26126 84306 26178 84318
rect 27470 84306 27522 84318
rect 21746 84254 21758 84306
rect 21810 84254 21822 84306
rect 22530 84254 22542 84306
rect 22594 84254 22606 84306
rect 23762 84254 23774 84306
rect 23826 84254 23838 84306
rect 25554 84254 25566 84306
rect 25618 84254 25630 84306
rect 27122 84254 27134 84306
rect 27186 84254 27198 84306
rect 21086 84242 21138 84254
rect 24446 84242 24498 84254
rect 26126 84242 26178 84254
rect 27470 84242 27522 84254
rect 27582 84306 27634 84318
rect 27582 84242 27634 84254
rect 2494 84194 2546 84206
rect 2494 84130 2546 84142
rect 5406 84194 5458 84206
rect 5406 84130 5458 84142
rect 9774 84194 9826 84206
rect 9774 84130 9826 84142
rect 16830 84194 16882 84206
rect 21422 84194 21474 84206
rect 26686 84194 26738 84206
rect 18610 84142 18622 84194
rect 18674 84142 18686 84194
rect 22642 84142 22654 84194
rect 22706 84142 22718 84194
rect 23538 84142 23550 84194
rect 23602 84142 23614 84194
rect 16830 84130 16882 84142
rect 21422 84130 21474 84142
rect 26686 84130 26738 84142
rect 28030 84194 28082 84206
rect 28030 84130 28082 84142
rect 26910 84082 26962 84094
rect 28018 84030 28030 84082
rect 28082 84079 28094 84082
rect 28242 84079 28254 84082
rect 28082 84033 28254 84079
rect 28082 84030 28094 84033
rect 28242 84030 28254 84033
rect 28306 84030 28318 84082
rect 26910 84018 26962 84030
rect 1344 83914 28560 83948
rect 1344 83862 4616 83914
rect 4668 83862 4720 83914
rect 4772 83862 4824 83914
rect 4876 83862 11420 83914
rect 11472 83862 11524 83914
rect 11576 83862 11628 83914
rect 11680 83862 18224 83914
rect 18276 83862 18328 83914
rect 18380 83862 18432 83914
rect 18484 83862 25028 83914
rect 25080 83862 25132 83914
rect 25184 83862 25236 83914
rect 25288 83862 28560 83914
rect 1344 83828 28560 83862
rect 26350 83746 26402 83758
rect 7410 83694 7422 83746
rect 7474 83743 7486 83746
rect 7746 83743 7758 83746
rect 7474 83697 7758 83743
rect 7474 83694 7486 83697
rect 7746 83694 7758 83697
rect 7810 83694 7822 83746
rect 26350 83682 26402 83694
rect 27470 83746 27522 83758
rect 27470 83682 27522 83694
rect 15598 83634 15650 83646
rect 12338 83582 12350 83634
rect 12402 83582 12414 83634
rect 15598 83570 15650 83582
rect 18398 83634 18450 83646
rect 18398 83570 18450 83582
rect 18958 83634 19010 83646
rect 19506 83582 19518 83634
rect 19570 83582 19582 83634
rect 20290 83582 20302 83634
rect 20354 83582 20366 83634
rect 21522 83582 21534 83634
rect 21586 83582 21598 83634
rect 22642 83582 22654 83634
rect 22706 83582 22718 83634
rect 24322 83582 24334 83634
rect 24386 83582 24398 83634
rect 18958 83570 19010 83582
rect 5966 83522 6018 83534
rect 14478 83522 14530 83534
rect 5730 83470 5742 83522
rect 5794 83470 5806 83522
rect 9538 83470 9550 83522
rect 9602 83470 9614 83522
rect 5966 83458 6018 83470
rect 14478 83458 14530 83470
rect 14590 83522 14642 83534
rect 14590 83458 14642 83470
rect 14926 83522 14978 83534
rect 14926 83458 14978 83470
rect 18062 83522 18114 83534
rect 20750 83522 20802 83534
rect 26014 83522 26066 83534
rect 19282 83470 19294 83522
rect 19346 83470 19358 83522
rect 21970 83470 21982 83522
rect 22034 83470 22046 83522
rect 22754 83470 22766 83522
rect 22818 83470 22830 83522
rect 23650 83470 23662 83522
rect 23714 83470 23726 83522
rect 24434 83470 24446 83522
rect 24498 83470 24510 83522
rect 18062 83458 18114 83470
rect 20750 83458 20802 83470
rect 26014 83458 26066 83470
rect 1710 83410 1762 83422
rect 1710 83346 1762 83358
rect 3278 83410 3330 83422
rect 6414 83410 6466 83422
rect 6178 83358 6190 83410
rect 6242 83358 6254 83410
rect 3278 83346 3330 83358
rect 6414 83346 6466 83358
rect 6862 83410 6914 83422
rect 12910 83410 12962 83422
rect 10210 83358 10222 83410
rect 10274 83358 10286 83410
rect 6862 83346 6914 83358
rect 12910 83346 12962 83358
rect 14814 83410 14866 83422
rect 14814 83346 14866 83358
rect 17838 83410 17890 83422
rect 17838 83346 17890 83358
rect 18846 83410 18898 83422
rect 18846 83346 18898 83358
rect 21310 83410 21362 83422
rect 25790 83410 25842 83422
rect 23426 83358 23438 83410
rect 23490 83358 23502 83410
rect 24546 83358 24558 83410
rect 24610 83358 24622 83410
rect 21310 83346 21362 83358
rect 25790 83346 25842 83358
rect 27134 83410 27186 83422
rect 27134 83346 27186 83358
rect 2046 83298 2098 83310
rect 2046 83234 2098 83246
rect 2830 83298 2882 83310
rect 2830 83234 2882 83246
rect 3838 83298 3890 83310
rect 3838 83234 3890 83246
rect 4174 83298 4226 83310
rect 4174 83234 4226 83246
rect 4622 83298 4674 83310
rect 4622 83234 4674 83246
rect 5070 83298 5122 83310
rect 5070 83234 5122 83246
rect 5630 83298 5682 83310
rect 5630 83234 5682 83246
rect 6750 83298 6802 83310
rect 6750 83234 6802 83246
rect 7310 83298 7362 83310
rect 7310 83234 7362 83246
rect 7758 83298 7810 83310
rect 7758 83234 7810 83246
rect 12574 83298 12626 83310
rect 12574 83234 12626 83246
rect 12798 83298 12850 83310
rect 12798 83234 12850 83246
rect 13918 83298 13970 83310
rect 13918 83234 13970 83246
rect 15934 83298 15986 83310
rect 15934 83234 15986 83246
rect 16382 83298 16434 83310
rect 16382 83234 16434 83246
rect 17166 83298 17218 83310
rect 17166 83234 17218 83246
rect 17614 83298 17666 83310
rect 17614 83234 17666 83246
rect 21534 83298 21586 83310
rect 21534 83234 21586 83246
rect 26798 83298 26850 83310
rect 26798 83234 26850 83246
rect 27358 83298 27410 83310
rect 27358 83234 27410 83246
rect 28030 83298 28082 83310
rect 28030 83234 28082 83246
rect 1344 83130 28720 83164
rect 1344 83078 8018 83130
rect 8070 83078 8122 83130
rect 8174 83078 8226 83130
rect 8278 83078 14822 83130
rect 14874 83078 14926 83130
rect 14978 83078 15030 83130
rect 15082 83078 21626 83130
rect 21678 83078 21730 83130
rect 21782 83078 21834 83130
rect 21886 83078 28430 83130
rect 28482 83078 28534 83130
rect 28586 83078 28638 83130
rect 28690 83078 28720 83130
rect 1344 83044 28720 83078
rect 7422 82962 7474 82974
rect 7422 82898 7474 82910
rect 9886 82962 9938 82974
rect 9886 82898 9938 82910
rect 10334 82962 10386 82974
rect 10334 82898 10386 82910
rect 10782 82962 10834 82974
rect 10782 82898 10834 82910
rect 11118 82962 11170 82974
rect 11118 82898 11170 82910
rect 11230 82962 11282 82974
rect 11230 82898 11282 82910
rect 11566 82962 11618 82974
rect 11566 82898 11618 82910
rect 16606 82962 16658 82974
rect 16606 82898 16658 82910
rect 17502 82962 17554 82974
rect 17502 82898 17554 82910
rect 19966 82962 20018 82974
rect 25454 82962 25506 82974
rect 23538 82910 23550 82962
rect 23602 82910 23614 82962
rect 19966 82898 20018 82910
rect 25454 82898 25506 82910
rect 16382 82850 16434 82862
rect 4834 82798 4846 82850
rect 4898 82798 4910 82850
rect 16382 82786 16434 82798
rect 21086 82850 21138 82862
rect 27470 82850 27522 82862
rect 22082 82798 22094 82850
rect 22146 82798 22158 82850
rect 24210 82798 24222 82850
rect 24274 82798 24286 82850
rect 26226 82798 26238 82850
rect 26290 82798 26302 82850
rect 21086 82786 21138 82798
rect 27470 82786 27522 82798
rect 2270 82738 2322 82750
rect 2270 82674 2322 82686
rect 2606 82738 2658 82750
rect 11342 82738 11394 82750
rect 15598 82738 15650 82750
rect 3042 82686 3054 82738
rect 3106 82686 3118 82738
rect 3378 82686 3390 82738
rect 3442 82686 3454 82738
rect 4050 82686 4062 82738
rect 4114 82686 4126 82738
rect 12338 82686 12350 82738
rect 12402 82686 12414 82738
rect 2606 82674 2658 82686
rect 11342 82674 11394 82686
rect 15598 82674 15650 82686
rect 15822 82738 15874 82750
rect 15822 82674 15874 82686
rect 16270 82738 16322 82750
rect 16270 82674 16322 82686
rect 16718 82738 16770 82750
rect 16718 82674 16770 82686
rect 20302 82738 20354 82750
rect 27022 82738 27074 82750
rect 20514 82686 20526 82738
rect 20578 82686 20590 82738
rect 22530 82686 22542 82738
rect 22594 82686 22606 82738
rect 23426 82686 23438 82738
rect 23490 82686 23502 82738
rect 25442 82686 25454 82738
rect 25506 82686 25518 82738
rect 26114 82686 26126 82738
rect 26178 82686 26190 82738
rect 20302 82674 20354 82686
rect 27022 82674 27074 82686
rect 27246 82738 27298 82750
rect 27246 82674 27298 82686
rect 2382 82626 2434 82638
rect 8094 82626 8146 82638
rect 15710 82626 15762 82638
rect 6962 82574 6974 82626
rect 7026 82574 7038 82626
rect 7410 82574 7422 82626
rect 7474 82574 7486 82626
rect 13458 82574 13470 82626
rect 13522 82574 13534 82626
rect 2382 82562 2434 82574
rect 8094 82562 8146 82574
rect 15710 82562 15762 82574
rect 18062 82626 18114 82638
rect 18062 82562 18114 82574
rect 18510 82626 18562 82638
rect 18510 82562 18562 82574
rect 18958 82626 19010 82638
rect 18958 82562 19010 82574
rect 19406 82626 19458 82638
rect 19406 82562 19458 82574
rect 19854 82626 19906 82638
rect 27134 82626 27186 82638
rect 26338 82574 26350 82626
rect 26402 82574 26414 82626
rect 19854 82562 19906 82574
rect 27134 82562 27186 82574
rect 28030 82626 28082 82638
rect 28030 82562 28082 82574
rect 3390 82514 3442 82526
rect 2818 82462 2830 82514
rect 2882 82462 2894 82514
rect 3390 82450 3442 82462
rect 3726 82514 3778 82526
rect 3726 82450 3778 82462
rect 7646 82514 7698 82526
rect 18050 82462 18062 82514
rect 18114 82511 18126 82514
rect 18946 82511 18958 82514
rect 18114 82465 18958 82511
rect 18114 82462 18126 82465
rect 18946 82462 18958 82465
rect 19010 82462 19022 82514
rect 7646 82450 7698 82462
rect 1344 82346 28560 82380
rect 1344 82294 4616 82346
rect 4668 82294 4720 82346
rect 4772 82294 4824 82346
rect 4876 82294 11420 82346
rect 11472 82294 11524 82346
rect 11576 82294 11628 82346
rect 11680 82294 18224 82346
rect 18276 82294 18328 82346
rect 18380 82294 18432 82346
rect 18484 82294 25028 82346
rect 25080 82294 25132 82346
rect 25184 82294 25236 82346
rect 25288 82294 28560 82346
rect 1344 82260 28560 82294
rect 5966 82178 6018 82190
rect 26014 82178 26066 82190
rect 10210 82126 10222 82178
rect 10274 82175 10286 82178
rect 11218 82175 11230 82178
rect 10274 82129 11230 82175
rect 10274 82126 10286 82129
rect 11218 82126 11230 82129
rect 11282 82126 11294 82178
rect 21970 82126 21982 82178
rect 22034 82126 22046 82178
rect 25218 82126 25230 82178
rect 25282 82126 25294 82178
rect 5966 82114 6018 82126
rect 26014 82114 26066 82126
rect 27694 82178 27746 82190
rect 27694 82114 27746 82126
rect 4958 82066 5010 82078
rect 9662 82066 9714 82078
rect 2482 82014 2494 82066
rect 2546 82014 2558 82066
rect 4610 82014 4622 82066
rect 4674 82014 4686 82066
rect 9314 82014 9326 82066
rect 9378 82014 9390 82066
rect 4958 82002 5010 82014
rect 9662 82002 9714 82014
rect 10222 82066 10274 82078
rect 17726 82066 17778 82078
rect 15586 82014 15598 82066
rect 15650 82014 15662 82066
rect 10222 82002 10274 82014
rect 17726 82002 17778 82014
rect 18398 82066 18450 82078
rect 27246 82066 27298 82078
rect 18398 82002 18450 82014
rect 24782 82010 24834 82022
rect 26562 82014 26574 82066
rect 26626 82014 26638 82066
rect 21310 81954 21362 81966
rect 27246 82002 27298 82014
rect 1810 81902 1822 81954
rect 1874 81902 1886 81954
rect 5954 81902 5966 81954
rect 6018 81902 6030 81954
rect 6514 81902 6526 81954
rect 6578 81902 6590 81954
rect 14802 81902 14814 81954
rect 14866 81902 14878 81954
rect 20178 81902 20190 81954
rect 20242 81902 20254 81954
rect 21522 81902 21534 81954
rect 21586 81902 21598 81954
rect 23202 81902 23214 81954
rect 23266 81902 23278 81954
rect 24434 81902 24446 81954
rect 24498 81902 24510 81954
rect 24782 81946 24834 81958
rect 27470 81954 27522 81966
rect 25442 81902 25454 81954
rect 25506 81902 25518 81954
rect 26226 81902 26238 81954
rect 26290 81902 26302 81954
rect 21310 81890 21362 81902
rect 27470 81890 27522 81902
rect 5630 81842 5682 81854
rect 20526 81842 20578 81854
rect 7186 81790 7198 81842
rect 7250 81790 7262 81842
rect 5630 81778 5682 81790
rect 20526 81778 20578 81790
rect 24670 81842 24722 81854
rect 24670 81778 24722 81790
rect 5070 81730 5122 81742
rect 5070 81666 5122 81678
rect 9774 81730 9826 81742
rect 9774 81666 9826 81678
rect 10670 81730 10722 81742
rect 10670 81666 10722 81678
rect 11118 81730 11170 81742
rect 11118 81666 11170 81678
rect 11566 81730 11618 81742
rect 11566 81666 11618 81678
rect 12014 81730 12066 81742
rect 12014 81666 12066 81678
rect 12462 81730 12514 81742
rect 12462 81666 12514 81678
rect 13022 81730 13074 81742
rect 13022 81666 13074 81678
rect 13582 81730 13634 81742
rect 13582 81666 13634 81678
rect 14030 81730 14082 81742
rect 14030 81666 14082 81678
rect 14478 81730 14530 81742
rect 14478 81666 14530 81678
rect 18846 81730 18898 81742
rect 18846 81666 18898 81678
rect 19294 81730 19346 81742
rect 19294 81666 19346 81678
rect 19742 81730 19794 81742
rect 19742 81666 19794 81678
rect 20638 81730 20690 81742
rect 20638 81666 20690 81678
rect 20750 81730 20802 81742
rect 20750 81666 20802 81678
rect 28142 81730 28194 81742
rect 28142 81666 28194 81678
rect 1344 81562 28720 81596
rect 1344 81510 8018 81562
rect 8070 81510 8122 81562
rect 8174 81510 8226 81562
rect 8278 81510 14822 81562
rect 14874 81510 14926 81562
rect 14978 81510 15030 81562
rect 15082 81510 21626 81562
rect 21678 81510 21730 81562
rect 21782 81510 21834 81562
rect 21886 81510 28430 81562
rect 28482 81510 28534 81562
rect 28586 81510 28638 81562
rect 28690 81510 28720 81562
rect 1344 81476 28720 81510
rect 10222 81394 10274 81406
rect 7186 81342 7198 81394
rect 7250 81342 7262 81394
rect 10222 81330 10274 81342
rect 11902 81394 11954 81406
rect 11902 81330 11954 81342
rect 17502 81394 17554 81406
rect 17502 81330 17554 81342
rect 17838 81394 17890 81406
rect 17838 81330 17890 81342
rect 19294 81394 19346 81406
rect 19294 81330 19346 81342
rect 22878 81394 22930 81406
rect 22878 81330 22930 81342
rect 23438 81394 23490 81406
rect 23438 81330 23490 81342
rect 23662 81394 23714 81406
rect 23662 81330 23714 81342
rect 23774 81394 23826 81406
rect 23774 81330 23826 81342
rect 24558 81394 24610 81406
rect 24558 81330 24610 81342
rect 26126 81394 26178 81406
rect 26126 81330 26178 81342
rect 16606 81282 16658 81294
rect 16606 81218 16658 81230
rect 16830 81282 16882 81294
rect 16830 81218 16882 81230
rect 18398 81282 18450 81294
rect 18398 81218 18450 81230
rect 18510 81282 18562 81294
rect 22654 81282 22706 81294
rect 19954 81230 19966 81282
rect 20018 81230 20030 81282
rect 18510 81218 18562 81230
rect 22654 81218 22706 81230
rect 23886 81282 23938 81294
rect 23886 81218 23938 81230
rect 24446 81282 24498 81294
rect 24446 81218 24498 81230
rect 26350 81282 26402 81294
rect 26350 81218 26402 81230
rect 6974 81170 7026 81182
rect 3042 81118 3054 81170
rect 3106 81118 3118 81170
rect 6974 81106 7026 81118
rect 7310 81170 7362 81182
rect 7310 81106 7362 81118
rect 7422 81170 7474 81182
rect 10782 81170 10834 81182
rect 17726 81170 17778 81182
rect 7746 81118 7758 81170
rect 7810 81118 7822 81170
rect 10546 81118 10558 81170
rect 10610 81118 10622 81170
rect 12226 81118 12238 81170
rect 12290 81118 12302 81170
rect 7422 81106 7474 81118
rect 10782 81106 10834 81118
rect 17726 81106 17778 81118
rect 17950 81170 18002 81182
rect 17950 81106 18002 81118
rect 18174 81170 18226 81182
rect 18174 81106 18226 81118
rect 19406 81170 19458 81182
rect 22542 81170 22594 81182
rect 20738 81118 20750 81170
rect 20802 81118 20814 81170
rect 21634 81118 21646 81170
rect 21698 81118 21710 81170
rect 19406 81106 19458 81118
rect 22542 81106 22594 81118
rect 22990 81170 23042 81182
rect 26898 81118 26910 81170
rect 26962 81118 26974 81170
rect 27122 81118 27134 81170
rect 27186 81118 27198 81170
rect 28130 81118 28142 81170
rect 28194 81118 28206 81170
rect 22990 81106 23042 81118
rect 5742 81058 5794 81070
rect 4834 81006 4846 81058
rect 4898 81006 4910 81058
rect 5742 80994 5794 81006
rect 6190 81058 6242 81070
rect 6190 80994 6242 81006
rect 6638 81058 6690 81070
rect 25230 81058 25282 81070
rect 14018 81006 14030 81058
rect 14082 81006 14094 81058
rect 20514 81006 20526 81058
rect 20578 81006 20590 81058
rect 28018 81006 28030 81058
rect 28082 81006 28094 81058
rect 6638 80994 6690 81006
rect 25230 80994 25282 81006
rect 11006 80946 11058 80958
rect 11006 80882 11058 80894
rect 11118 80946 11170 80958
rect 11118 80882 11170 80894
rect 16494 80946 16546 80958
rect 16494 80882 16546 80894
rect 19294 80946 19346 80958
rect 19294 80882 19346 80894
rect 24558 80946 24610 80958
rect 24558 80882 24610 80894
rect 25454 80946 25506 80958
rect 25454 80882 25506 80894
rect 25678 80946 25730 80958
rect 25678 80882 25730 80894
rect 26462 80946 26514 80958
rect 26462 80882 26514 80894
rect 1344 80778 28560 80812
rect 1344 80726 4616 80778
rect 4668 80726 4720 80778
rect 4772 80726 4824 80778
rect 4876 80726 11420 80778
rect 11472 80726 11524 80778
rect 11576 80726 11628 80778
rect 11680 80726 18224 80778
rect 18276 80726 18328 80778
rect 18380 80726 18432 80778
rect 18484 80726 25028 80778
rect 25080 80726 25132 80778
rect 25184 80726 25236 80778
rect 25288 80726 28560 80778
rect 1344 80692 28560 80726
rect 21646 80610 21698 80622
rect 20178 80558 20190 80610
rect 20242 80558 20254 80610
rect 21646 80546 21698 80558
rect 24110 80610 24162 80622
rect 24110 80546 24162 80558
rect 24558 80610 24610 80622
rect 24558 80546 24610 80558
rect 26238 80610 26290 80622
rect 26238 80546 26290 80558
rect 26574 80610 26626 80622
rect 26574 80546 26626 80558
rect 27246 80610 27298 80622
rect 27570 80558 27582 80610
rect 27634 80558 27646 80610
rect 27246 80546 27298 80558
rect 2830 80498 2882 80510
rect 2830 80434 2882 80446
rect 4062 80498 4114 80510
rect 4062 80434 4114 80446
rect 7086 80498 7138 80510
rect 27022 80498 27074 80510
rect 10098 80446 10110 80498
rect 10162 80446 10174 80498
rect 12226 80446 12238 80498
rect 12290 80446 12302 80498
rect 16482 80446 16494 80498
rect 16546 80446 16558 80498
rect 17490 80446 17502 80498
rect 17554 80446 17566 80498
rect 18274 80446 18286 80498
rect 18338 80446 18350 80498
rect 23426 80446 23438 80498
rect 23490 80446 23502 80498
rect 7086 80434 7138 80446
rect 27022 80434 27074 80446
rect 28030 80498 28082 80510
rect 28030 80434 28082 80446
rect 17838 80386 17890 80398
rect 18846 80386 18898 80398
rect 21310 80386 21362 80398
rect 24446 80386 24498 80398
rect 3042 80334 3054 80386
rect 3106 80334 3118 80386
rect 6066 80334 6078 80386
rect 6130 80334 6142 80386
rect 9426 80334 9438 80386
rect 9490 80334 9502 80386
rect 13570 80334 13582 80386
rect 13634 80334 13646 80386
rect 17378 80334 17390 80386
rect 17442 80334 17454 80386
rect 18050 80334 18062 80386
rect 18114 80334 18126 80386
rect 19282 80334 19294 80386
rect 19346 80334 19358 80386
rect 19954 80334 19966 80386
rect 20018 80334 20030 80386
rect 22082 80334 22094 80386
rect 22146 80334 22158 80386
rect 17838 80322 17890 80334
rect 18846 80322 18898 80334
rect 21310 80322 21362 80334
rect 24446 80322 24498 80334
rect 25230 80386 25282 80398
rect 25230 80322 25282 80334
rect 25566 80386 25618 80398
rect 25566 80322 25618 80334
rect 25902 80386 25954 80398
rect 25902 80322 25954 80334
rect 5742 80274 5794 80286
rect 20526 80274 20578 80286
rect 14354 80222 14366 80274
rect 14418 80222 14430 80274
rect 5742 80210 5794 80222
rect 20526 80210 20578 80222
rect 22430 80274 22482 80286
rect 22430 80210 22482 80222
rect 23102 80274 23154 80286
rect 23102 80210 23154 80222
rect 23998 80274 24050 80286
rect 23998 80210 24050 80222
rect 26462 80274 26514 80286
rect 26462 80210 26514 80222
rect 1710 80162 1762 80174
rect 5070 80162 5122 80174
rect 2034 80110 2046 80162
rect 2098 80110 2110 80162
rect 1710 80098 1762 80110
rect 5070 80098 5122 80110
rect 5854 80162 5906 80174
rect 5854 80098 5906 80110
rect 6526 80162 6578 80174
rect 6526 80098 6578 80110
rect 13022 80162 13074 80174
rect 13022 80098 13074 80110
rect 21534 80162 21586 80174
rect 21534 80098 21586 80110
rect 23326 80162 23378 80174
rect 23326 80098 23378 80110
rect 25006 80162 25058 80174
rect 25006 80098 25058 80110
rect 25566 80162 25618 80174
rect 25566 80098 25618 80110
rect 1344 79994 28720 80028
rect 1344 79942 8018 79994
rect 8070 79942 8122 79994
rect 8174 79942 8226 79994
rect 8278 79942 14822 79994
rect 14874 79942 14926 79994
rect 14978 79942 15030 79994
rect 15082 79942 21626 79994
rect 21678 79942 21730 79994
rect 21782 79942 21834 79994
rect 21886 79942 28430 79994
rect 28482 79942 28534 79994
rect 28586 79942 28638 79994
rect 28690 79942 28720 79994
rect 1344 79908 28720 79942
rect 2494 79826 2546 79838
rect 2494 79762 2546 79774
rect 17726 79826 17778 79838
rect 17726 79762 17778 79774
rect 24670 79826 24722 79838
rect 24670 79762 24722 79774
rect 26238 79826 26290 79838
rect 26238 79762 26290 79774
rect 26686 79826 26738 79838
rect 26686 79762 26738 79774
rect 27134 79826 27186 79838
rect 27134 79762 27186 79774
rect 28030 79826 28082 79838
rect 28030 79762 28082 79774
rect 17614 79714 17666 79726
rect 12674 79662 12686 79714
rect 12738 79662 12750 79714
rect 14802 79662 14814 79714
rect 14866 79662 14878 79714
rect 15810 79662 15822 79714
rect 15874 79662 15886 79714
rect 17614 79650 17666 79662
rect 19518 79714 19570 79726
rect 19518 79650 19570 79662
rect 7758 79602 7810 79614
rect 3266 79550 3278 79602
rect 3330 79550 3342 79602
rect 4498 79550 4510 79602
rect 4562 79550 4574 79602
rect 7758 79538 7810 79550
rect 10110 79602 10162 79614
rect 17950 79602 18002 79614
rect 10322 79550 10334 79602
rect 10386 79550 10398 79602
rect 11666 79550 11678 79602
rect 11730 79550 11742 79602
rect 14914 79550 14926 79602
rect 14978 79550 14990 79602
rect 16370 79550 16382 79602
rect 16434 79550 16446 79602
rect 10110 79538 10162 79550
rect 17950 79538 18002 79550
rect 18174 79602 18226 79614
rect 23774 79602 23826 79614
rect 19058 79550 19070 79602
rect 19122 79550 19134 79602
rect 19730 79550 19742 79602
rect 19794 79550 19806 79602
rect 21074 79550 21086 79602
rect 21138 79550 21150 79602
rect 21522 79550 21534 79602
rect 21586 79550 21598 79602
rect 21858 79550 21870 79602
rect 21922 79550 21934 79602
rect 18174 79538 18226 79550
rect 23774 79538 23826 79550
rect 24222 79602 24274 79614
rect 24222 79538 24274 79550
rect 25790 79602 25842 79614
rect 25790 79538 25842 79550
rect 4062 79490 4114 79502
rect 8318 79490 8370 79502
rect 5282 79438 5294 79490
rect 5346 79438 5358 79490
rect 7410 79438 7422 79490
rect 7474 79438 7486 79490
rect 4062 79426 4114 79438
rect 8318 79426 8370 79438
rect 9102 79490 9154 79502
rect 23326 79490 23378 79502
rect 10546 79438 10558 79490
rect 10610 79438 10622 79490
rect 13122 79438 13134 79490
rect 13186 79438 13198 79490
rect 19170 79438 19182 79490
rect 19234 79438 19246 79490
rect 19954 79438 19966 79490
rect 20018 79438 20030 79490
rect 22642 79438 22654 79490
rect 22706 79438 22718 79490
rect 9102 79426 9154 79438
rect 23326 79426 23378 79438
rect 25454 79490 25506 79502
rect 25454 79426 25506 79438
rect 27582 79490 27634 79502
rect 27582 79426 27634 79438
rect 7870 79378 7922 79390
rect 3602 79326 3614 79378
rect 3666 79326 3678 79378
rect 10658 79326 10670 79378
rect 10722 79326 10734 79378
rect 27346 79326 27358 79378
rect 27410 79375 27422 79378
rect 28018 79375 28030 79378
rect 27410 79329 28030 79375
rect 27410 79326 27422 79329
rect 28018 79326 28030 79329
rect 28082 79326 28094 79378
rect 7870 79314 7922 79326
rect 1344 79210 28560 79244
rect 1344 79158 4616 79210
rect 4668 79158 4720 79210
rect 4772 79158 4824 79210
rect 4876 79158 11420 79210
rect 11472 79158 11524 79210
rect 11576 79158 11628 79210
rect 11680 79158 18224 79210
rect 18276 79158 18328 79210
rect 18380 79158 18432 79210
rect 18484 79158 25028 79210
rect 25080 79158 25132 79210
rect 25184 79158 25236 79210
rect 25288 79158 28560 79210
rect 1344 79124 28560 79158
rect 18958 79042 19010 79054
rect 5842 78990 5854 79042
rect 5906 78990 5918 79042
rect 14242 78990 14254 79042
rect 14306 78990 14318 79042
rect 18958 78978 19010 78990
rect 19742 79042 19794 79054
rect 25330 78990 25342 79042
rect 25394 79039 25406 79042
rect 25554 79039 25566 79042
rect 25394 78993 25566 79039
rect 25394 78990 25406 78993
rect 25554 78990 25566 78993
rect 25618 78990 25630 79042
rect 19742 78978 19794 78990
rect 19070 78930 19122 78942
rect 4610 78878 4622 78930
rect 4674 78878 4686 78930
rect 11218 78878 11230 78930
rect 11282 78878 11294 78930
rect 12002 78878 12014 78930
rect 12066 78878 12078 78930
rect 17714 78878 17726 78930
rect 17778 78878 17790 78930
rect 19070 78866 19122 78878
rect 21422 78930 21474 78942
rect 21422 78866 21474 78878
rect 24222 78930 24274 78942
rect 24222 78866 24274 78878
rect 26462 78930 26514 78942
rect 26462 78866 26514 78878
rect 26910 78930 26962 78942
rect 26910 78866 26962 78878
rect 27358 78930 27410 78942
rect 27358 78866 27410 78878
rect 28142 78930 28194 78942
rect 28142 78866 28194 78878
rect 12126 78818 12178 78830
rect 13694 78818 13746 78830
rect 23774 78818 23826 78830
rect 1810 78766 1822 78818
rect 1874 78766 1886 78818
rect 5842 78766 5854 78818
rect 5906 78766 5918 78818
rect 6178 78766 6190 78818
rect 6242 78766 6254 78818
rect 8418 78766 8430 78818
rect 8482 78766 8494 78818
rect 12226 78766 12238 78818
rect 12290 78766 12302 78818
rect 13906 78766 13918 78818
rect 13970 78766 13982 78818
rect 14242 78766 14254 78818
rect 14306 78766 14318 78818
rect 14802 78766 14814 78818
rect 14866 78766 14878 78818
rect 18050 78766 18062 78818
rect 18114 78766 18126 78818
rect 19282 78766 19294 78818
rect 19346 78766 19358 78818
rect 20178 78766 20190 78818
rect 20242 78766 20254 78818
rect 12126 78754 12178 78766
rect 13694 78754 13746 78766
rect 23774 78754 23826 78766
rect 6414 78706 6466 78718
rect 19630 78706 19682 78718
rect 2482 78654 2494 78706
rect 2546 78654 2558 78706
rect 9090 78654 9102 78706
rect 9154 78654 9166 78706
rect 15586 78654 15598 78706
rect 15650 78654 15662 78706
rect 6414 78642 6466 78654
rect 19630 78642 19682 78654
rect 19742 78706 19794 78718
rect 19742 78642 19794 78654
rect 20526 78706 20578 78718
rect 20526 78642 20578 78654
rect 21310 78706 21362 78718
rect 21310 78642 21362 78654
rect 22542 78706 22594 78718
rect 22542 78642 22594 78654
rect 23326 78706 23378 78718
rect 23326 78642 23378 78654
rect 5070 78594 5122 78606
rect 5070 78530 5122 78542
rect 5630 78594 5682 78606
rect 5630 78530 5682 78542
rect 6862 78594 6914 78606
rect 6862 78530 6914 78542
rect 7870 78594 7922 78606
rect 7870 78530 7922 78542
rect 13022 78594 13074 78606
rect 13022 78530 13074 78542
rect 14478 78594 14530 78606
rect 21534 78594 21586 78606
rect 18610 78542 18622 78594
rect 18674 78542 18686 78594
rect 14478 78530 14530 78542
rect 21534 78530 21586 78542
rect 22094 78594 22146 78606
rect 22094 78530 22146 78542
rect 22654 78594 22706 78606
rect 22654 78530 22706 78542
rect 22766 78594 22818 78606
rect 22766 78530 22818 78542
rect 24670 78594 24722 78606
rect 24670 78530 24722 78542
rect 25118 78594 25170 78606
rect 25118 78530 25170 78542
rect 25678 78594 25730 78606
rect 25678 78530 25730 78542
rect 26126 78594 26178 78606
rect 26126 78530 26178 78542
rect 1344 78426 28720 78460
rect 1344 78374 8018 78426
rect 8070 78374 8122 78426
rect 8174 78374 8226 78426
rect 8278 78374 14822 78426
rect 14874 78374 14926 78426
rect 14978 78374 15030 78426
rect 15082 78374 21626 78426
rect 21678 78374 21730 78426
rect 21782 78374 21834 78426
rect 21886 78374 28430 78426
rect 28482 78374 28534 78426
rect 28586 78374 28638 78426
rect 28690 78374 28720 78426
rect 1344 78340 28720 78374
rect 2382 78258 2434 78270
rect 2382 78194 2434 78206
rect 4846 78258 4898 78270
rect 4846 78194 4898 78206
rect 5294 78258 5346 78270
rect 5294 78194 5346 78206
rect 6414 78258 6466 78270
rect 6414 78194 6466 78206
rect 8990 78258 9042 78270
rect 17502 78258 17554 78270
rect 10994 78206 11006 78258
rect 11058 78206 11070 78258
rect 8990 78194 9042 78206
rect 17502 78194 17554 78206
rect 2046 78146 2098 78158
rect 2046 78082 2098 78094
rect 3166 78146 3218 78158
rect 3166 78082 3218 78094
rect 18846 78146 18898 78158
rect 18846 78082 18898 78094
rect 20190 78146 20242 78158
rect 20190 78082 20242 78094
rect 1710 78034 1762 78046
rect 3502 78034 3554 78046
rect 7870 78034 7922 78046
rect 2594 77982 2606 78034
rect 2658 77982 2670 78034
rect 2930 77982 2942 78034
rect 2994 77982 3006 78034
rect 3714 77982 3726 78034
rect 3778 78031 3790 78034
rect 3778 77985 3999 78031
rect 3778 77982 3790 77985
rect 1710 77970 1762 77982
rect 3502 77970 3554 77982
rect 3614 77922 3666 77934
rect 3614 77858 3666 77870
rect 2718 77810 2770 77822
rect 3953 77807 3999 77985
rect 7870 77970 7922 77982
rect 8206 78034 8258 78046
rect 8206 77970 8258 77982
rect 8542 78034 8594 78046
rect 17390 78034 17442 78046
rect 19742 78034 19794 78046
rect 8754 77982 8766 78034
rect 8818 77982 8830 78034
rect 9874 77982 9886 78034
rect 9938 77982 9950 78034
rect 13010 77982 13022 78034
rect 13074 77982 13086 78034
rect 17602 77982 17614 78034
rect 17666 77982 17678 78034
rect 17938 77982 17950 78034
rect 18002 77982 18014 78034
rect 18498 77982 18510 78034
rect 18562 77982 18574 78034
rect 21858 77982 21870 78034
rect 21922 77982 21934 78034
rect 25330 77982 25342 78034
rect 25394 77982 25406 78034
rect 8542 77970 8594 77982
rect 17390 77970 17442 77982
rect 19742 77970 19794 77982
rect 4062 77922 4114 77934
rect 4062 77858 4114 77870
rect 6078 77922 6130 77934
rect 6078 77858 6130 77870
rect 6974 77922 7026 77934
rect 6974 77858 7026 77870
rect 7422 77922 7474 77934
rect 19294 77922 19346 77934
rect 13570 77870 13582 77922
rect 13634 77870 13646 77922
rect 7422 77858 7474 77870
rect 19294 77858 19346 77870
rect 20638 77922 20690 77934
rect 20638 77858 20690 77870
rect 21086 77922 21138 77934
rect 22530 77870 22542 77922
rect 22594 77870 22606 77922
rect 24658 77870 24670 77922
rect 24722 77870 24734 77922
rect 26002 77870 26014 77922
rect 26066 77870 26078 77922
rect 28130 77870 28142 77922
rect 28194 77870 28206 77922
rect 21086 77858 21138 77870
rect 17838 77810 17890 77822
rect 4050 77807 4062 77810
rect 3953 77761 4062 77807
rect 4050 77758 4062 77761
rect 4114 77758 4126 77810
rect 7410 77758 7422 77810
rect 7474 77807 7486 77810
rect 7970 77807 7982 77810
rect 7474 77761 7982 77807
rect 7474 77758 7486 77761
rect 7970 77758 7982 77761
rect 8034 77758 8046 77810
rect 8754 77758 8766 77810
rect 8818 77758 8830 77810
rect 2718 77746 2770 77758
rect 17838 77746 17890 77758
rect 18510 77810 18562 77822
rect 20626 77758 20638 77810
rect 20690 77807 20702 77810
rect 21410 77807 21422 77810
rect 20690 77761 21422 77807
rect 20690 77758 20702 77761
rect 21410 77758 21422 77761
rect 21474 77758 21486 77810
rect 18510 77746 18562 77758
rect 1344 77642 28560 77676
rect 1344 77590 4616 77642
rect 4668 77590 4720 77642
rect 4772 77590 4824 77642
rect 4876 77590 11420 77642
rect 11472 77590 11524 77642
rect 11576 77590 11628 77642
rect 11680 77590 18224 77642
rect 18276 77590 18328 77642
rect 18380 77590 18432 77642
rect 18484 77590 25028 77642
rect 25080 77590 25132 77642
rect 25184 77590 25236 77642
rect 25288 77590 28560 77642
rect 1344 77556 28560 77590
rect 20414 77474 20466 77486
rect 22530 77422 22542 77474
rect 22594 77422 22606 77474
rect 20414 77410 20466 77422
rect 21422 77362 21474 77374
rect 2706 77310 2718 77362
rect 2770 77310 2782 77362
rect 8530 77310 8542 77362
rect 8594 77310 8606 77362
rect 12898 77310 12910 77362
rect 12962 77310 12974 77362
rect 21422 77298 21474 77310
rect 23214 77362 23266 77374
rect 25218 77310 25230 77362
rect 25282 77310 25294 77362
rect 23214 77298 23266 77310
rect 9662 77250 9714 77262
rect 21982 77250 22034 77262
rect 24446 77250 24498 77262
rect 3490 77198 3502 77250
rect 3554 77198 3566 77250
rect 5618 77198 5630 77250
rect 5682 77198 5694 77250
rect 10098 77198 10110 77250
rect 10162 77198 10174 77250
rect 15026 77198 15038 77250
rect 15090 77198 15102 77250
rect 22530 77198 22542 77250
rect 22594 77198 22606 77250
rect 28018 77198 28030 77250
rect 28082 77198 28094 77250
rect 9662 77186 9714 77198
rect 21982 77186 22034 77198
rect 24446 77186 24498 77198
rect 2494 77138 2546 77150
rect 2494 77074 2546 77086
rect 2718 77138 2770 77150
rect 13582 77138 13634 77150
rect 23662 77138 23714 77150
rect 6402 77086 6414 77138
rect 6466 77086 6478 77138
rect 10770 77086 10782 77138
rect 10834 77086 10846 77138
rect 18386 77086 18398 77138
rect 18450 77086 18462 77138
rect 22194 77086 22206 77138
rect 22258 77086 22270 77138
rect 2718 77074 2770 77086
rect 13582 77074 13634 77086
rect 23662 77074 23714 77086
rect 24334 77138 24386 77150
rect 24334 77074 24386 77086
rect 24670 77138 24722 77150
rect 24670 77074 24722 77086
rect 24894 77138 24946 77150
rect 27346 77086 27358 77138
rect 27410 77086 27422 77138
rect 24894 77074 24946 77086
rect 2158 77026 2210 77038
rect 4734 77026 4786 77038
rect 4050 76974 4062 77026
rect 4114 76974 4126 77026
rect 2158 76962 2210 76974
rect 4734 76962 4786 76974
rect 5070 77026 5122 77038
rect 5070 76962 5122 76974
rect 9326 77026 9378 77038
rect 9326 76962 9378 76974
rect 13694 77026 13746 77038
rect 13694 76962 13746 76974
rect 19966 77026 20018 77038
rect 19966 76962 20018 76974
rect 20526 77026 20578 77038
rect 20526 76962 20578 76974
rect 20638 77026 20690 77038
rect 23102 77026 23154 77038
rect 22418 76974 22430 77026
rect 22482 76974 22494 77026
rect 20638 76962 20690 76974
rect 23102 76962 23154 76974
rect 1344 76858 28720 76892
rect 1344 76806 8018 76858
rect 8070 76806 8122 76858
rect 8174 76806 8226 76858
rect 8278 76806 14822 76858
rect 14874 76806 14926 76858
rect 14978 76806 15030 76858
rect 15082 76806 21626 76858
rect 21678 76806 21730 76858
rect 21782 76806 21834 76858
rect 21886 76806 28430 76858
rect 28482 76806 28534 76858
rect 28586 76806 28638 76858
rect 28690 76806 28720 76858
rect 1344 76772 28720 76806
rect 6638 76690 6690 76702
rect 6638 76626 6690 76638
rect 11118 76690 11170 76702
rect 11118 76626 11170 76638
rect 11230 76690 11282 76702
rect 11230 76626 11282 76638
rect 11902 76690 11954 76702
rect 11902 76626 11954 76638
rect 13134 76690 13186 76702
rect 13134 76626 13186 76638
rect 17502 76690 17554 76702
rect 17502 76626 17554 76638
rect 22206 76690 22258 76702
rect 22206 76626 22258 76638
rect 22654 76690 22706 76702
rect 22654 76626 22706 76638
rect 24446 76690 24498 76702
rect 24446 76626 24498 76638
rect 25342 76690 25394 76702
rect 25342 76626 25394 76638
rect 26238 76690 26290 76702
rect 26238 76626 26290 76638
rect 26910 76690 26962 76702
rect 26910 76626 26962 76638
rect 27022 76690 27074 76702
rect 27022 76626 27074 76638
rect 28142 76690 28194 76702
rect 28142 76626 28194 76638
rect 2830 76578 2882 76590
rect 2830 76514 2882 76526
rect 10446 76578 10498 76590
rect 18174 76578 18226 76590
rect 15250 76526 15262 76578
rect 15314 76526 15326 76578
rect 10446 76514 10498 76526
rect 18174 76514 18226 76526
rect 27358 76578 27410 76590
rect 27358 76514 27410 76526
rect 5294 76466 5346 76478
rect 3714 76414 3726 76466
rect 3778 76414 3790 76466
rect 5294 76402 5346 76414
rect 6526 76466 6578 76478
rect 6526 76402 6578 76414
rect 6862 76466 6914 76478
rect 9774 76466 9826 76478
rect 7074 76414 7086 76466
rect 7138 76414 7150 76466
rect 7970 76414 7982 76466
rect 8034 76414 8046 76466
rect 6862 76402 6914 76414
rect 9774 76402 9826 76414
rect 10110 76466 10162 76478
rect 10110 76402 10162 76414
rect 10670 76466 10722 76478
rect 10670 76402 10722 76414
rect 11790 76466 11842 76478
rect 11790 76402 11842 76414
rect 12126 76466 12178 76478
rect 12126 76402 12178 76414
rect 12350 76466 12402 76478
rect 16494 76466 16546 76478
rect 25902 76466 25954 76478
rect 14018 76414 14030 76466
rect 14082 76414 14094 76466
rect 18946 76414 18958 76466
rect 19010 76414 19022 76466
rect 12350 76402 12402 76414
rect 16494 76402 16546 76414
rect 25902 76402 25954 76414
rect 26350 76466 26402 76478
rect 26350 76402 26402 76414
rect 26462 76466 26514 76478
rect 26462 76402 26514 76414
rect 27134 76466 27186 76478
rect 27134 76402 27186 76414
rect 1822 76354 1874 76366
rect 1822 76290 1874 76302
rect 2270 76354 2322 76366
rect 2270 76290 2322 76302
rect 2718 76354 2770 76366
rect 2718 76290 2770 76302
rect 4622 76354 4674 76366
rect 4622 76290 4674 76302
rect 5742 76354 5794 76366
rect 5742 76290 5794 76302
rect 6302 76354 6354 76366
rect 6302 76290 6354 76302
rect 7758 76354 7810 76366
rect 7758 76290 7810 76302
rect 8542 76354 8594 76366
rect 8542 76290 8594 76302
rect 8990 76354 9042 76366
rect 8990 76290 9042 76302
rect 10222 76354 10274 76366
rect 23214 76354 23266 76366
rect 19618 76302 19630 76354
rect 19682 76302 19694 76354
rect 21746 76302 21758 76354
rect 21810 76302 21822 76354
rect 10222 76290 10274 76302
rect 23214 76290 23266 76302
rect 23550 76354 23602 76366
rect 23550 76290 23602 76302
rect 24110 76354 24162 76366
rect 24110 76290 24162 76302
rect 2606 76242 2658 76254
rect 7646 76242 7698 76254
rect 7074 76190 7086 76242
rect 7138 76190 7150 76242
rect 2606 76178 2658 76190
rect 7646 76178 7698 76190
rect 11006 76242 11058 76254
rect 11006 76178 11058 76190
rect 18062 76242 18114 76254
rect 21970 76190 21982 76242
rect 22034 76239 22046 76242
rect 22866 76239 22878 76242
rect 22034 76193 22878 76239
rect 22034 76190 22046 76193
rect 22866 76190 22878 76193
rect 22930 76239 22942 76242
rect 24434 76239 24446 76242
rect 22930 76193 24446 76239
rect 22930 76190 22942 76193
rect 24434 76190 24446 76193
rect 24498 76190 24510 76242
rect 18062 76178 18114 76190
rect 1344 76074 28560 76108
rect 1344 76022 4616 76074
rect 4668 76022 4720 76074
rect 4772 76022 4824 76074
rect 4876 76022 11420 76074
rect 11472 76022 11524 76074
rect 11576 76022 11628 76074
rect 11680 76022 18224 76074
rect 18276 76022 18328 76074
rect 18380 76022 18432 76074
rect 18484 76022 25028 76074
rect 25080 76022 25132 76074
rect 25184 76022 25236 76074
rect 25288 76022 28560 76074
rect 1344 75988 28560 76022
rect 18274 75854 18286 75906
rect 18338 75854 18350 75906
rect 20178 75854 20190 75906
rect 20242 75854 20254 75906
rect 21858 75854 21870 75906
rect 21922 75903 21934 75906
rect 22082 75903 22094 75906
rect 21922 75857 22094 75903
rect 21922 75854 21934 75857
rect 22082 75854 22094 75857
rect 22146 75854 22158 75906
rect 12462 75794 12514 75806
rect 16830 75794 16882 75806
rect 4610 75742 4622 75794
rect 4674 75742 4686 75794
rect 8530 75742 8542 75794
rect 8594 75742 8606 75794
rect 9762 75742 9774 75794
rect 9826 75742 9838 75794
rect 11890 75742 11902 75794
rect 11954 75742 11966 75794
rect 16370 75742 16382 75794
rect 16434 75742 16446 75794
rect 12462 75730 12514 75742
rect 16830 75730 16882 75742
rect 19182 75794 19234 75806
rect 19182 75730 19234 75742
rect 19742 75794 19794 75806
rect 19742 75730 19794 75742
rect 21422 75794 21474 75806
rect 21422 75730 21474 75742
rect 21870 75794 21922 75806
rect 21870 75730 21922 75742
rect 22318 75794 22370 75806
rect 26462 75794 26514 75806
rect 25666 75742 25678 75794
rect 25730 75742 25742 75794
rect 22318 75730 22370 75742
rect 26462 75730 26514 75742
rect 27358 75794 27410 75806
rect 27358 75730 27410 75742
rect 4958 75682 5010 75694
rect 1698 75630 1710 75682
rect 1762 75630 1774 75682
rect 4958 75618 5010 75630
rect 5070 75682 5122 75694
rect 12574 75682 12626 75694
rect 19966 75682 20018 75694
rect 27022 75682 27074 75694
rect 5618 75630 5630 75682
rect 5682 75630 5694 75682
rect 9090 75630 9102 75682
rect 9154 75630 9166 75682
rect 12898 75630 12910 75682
rect 12962 75630 12974 75682
rect 13570 75630 13582 75682
rect 13634 75630 13646 75682
rect 18274 75630 18286 75682
rect 18338 75630 18350 75682
rect 20178 75630 20190 75682
rect 20242 75630 20254 75682
rect 22866 75630 22878 75682
rect 22930 75630 22942 75682
rect 5070 75618 5122 75630
rect 12574 75618 12626 75630
rect 19966 75618 20018 75630
rect 27022 75618 27074 75630
rect 17726 75570 17778 75582
rect 19630 75570 19682 75582
rect 2482 75518 2494 75570
rect 2546 75518 2558 75570
rect 6402 75518 6414 75570
rect 6466 75518 6478 75570
rect 14242 75518 14254 75570
rect 14306 75518 14318 75570
rect 17938 75518 17950 75570
rect 18002 75518 18014 75570
rect 23538 75518 23550 75570
rect 23602 75518 23614 75570
rect 17726 75506 17778 75518
rect 19630 75506 19682 75518
rect 12350 75458 12402 75470
rect 12350 75394 12402 75406
rect 17278 75458 17330 75470
rect 21310 75458 21362 75470
rect 18162 75406 18174 75458
rect 18226 75406 18238 75458
rect 17278 75394 17330 75406
rect 21310 75394 21362 75406
rect 26350 75458 26402 75470
rect 26350 75394 26402 75406
rect 26574 75458 26626 75470
rect 26574 75394 26626 75406
rect 27806 75458 27858 75470
rect 27806 75394 27858 75406
rect 1344 75290 28720 75324
rect 1344 75238 8018 75290
rect 8070 75238 8122 75290
rect 8174 75238 8226 75290
rect 8278 75238 14822 75290
rect 14874 75238 14926 75290
rect 14978 75238 15030 75290
rect 15082 75238 21626 75290
rect 21678 75238 21730 75290
rect 21782 75238 21834 75290
rect 21886 75238 28430 75290
rect 28482 75238 28534 75290
rect 28586 75238 28638 75290
rect 28690 75238 28720 75290
rect 1344 75204 28720 75238
rect 2382 75122 2434 75134
rect 2382 75058 2434 75070
rect 4846 75122 4898 75134
rect 4846 75058 4898 75070
rect 6414 75122 6466 75134
rect 6414 75058 6466 75070
rect 6974 75122 7026 75134
rect 6974 75058 7026 75070
rect 7534 75122 7586 75134
rect 7534 75058 7586 75070
rect 7982 75122 8034 75134
rect 7982 75058 8034 75070
rect 8542 75122 8594 75134
rect 8542 75058 8594 75070
rect 8766 75122 8818 75134
rect 8766 75058 8818 75070
rect 9774 75122 9826 75134
rect 9774 75058 9826 75070
rect 9998 75122 10050 75134
rect 9998 75058 10050 75070
rect 11006 75122 11058 75134
rect 11006 75058 11058 75070
rect 11230 75122 11282 75134
rect 11230 75058 11282 75070
rect 11342 75122 11394 75134
rect 11342 75058 11394 75070
rect 12350 75122 12402 75134
rect 12350 75058 12402 75070
rect 14254 75122 14306 75134
rect 14254 75058 14306 75070
rect 15150 75122 15202 75134
rect 15150 75058 15202 75070
rect 15934 75122 15986 75134
rect 15934 75058 15986 75070
rect 20750 75122 20802 75134
rect 20750 75058 20802 75070
rect 23774 75122 23826 75134
rect 23774 75058 23826 75070
rect 24670 75122 24722 75134
rect 24670 75058 24722 75070
rect 26686 75122 26738 75134
rect 26686 75058 26738 75070
rect 28142 75122 28194 75134
rect 28142 75058 28194 75070
rect 2046 75010 2098 75022
rect 3166 75010 3218 75022
rect 2930 74958 2942 75010
rect 2994 74958 3006 75010
rect 2046 74946 2098 74958
rect 3166 74946 3218 74958
rect 5630 75010 5682 75022
rect 5630 74946 5682 74958
rect 10222 75010 10274 75022
rect 10222 74946 10274 74958
rect 13582 75010 13634 75022
rect 18162 74958 18174 75010
rect 18226 74958 18238 75010
rect 13582 74946 13634 74958
rect 1710 74898 1762 74910
rect 2718 74898 2770 74910
rect 5966 74898 6018 74910
rect 2482 74846 2494 74898
rect 2546 74846 2558 74898
rect 3602 74846 3614 74898
rect 3666 74846 3678 74898
rect 1710 74834 1762 74846
rect 2718 74834 2770 74846
rect 5966 74834 6018 74846
rect 6078 74898 6130 74910
rect 6862 74898 6914 74910
rect 6178 74846 6190 74898
rect 6242 74846 6254 74898
rect 6078 74834 6130 74846
rect 6862 74834 6914 74846
rect 8430 74898 8482 74910
rect 8430 74834 8482 74846
rect 8990 74898 9042 74910
rect 8990 74834 9042 74846
rect 9550 74898 9602 74910
rect 9550 74834 9602 74846
rect 11454 74898 11506 74910
rect 13246 74898 13298 74910
rect 11778 74846 11790 74898
rect 11842 74846 11854 74898
rect 11454 74834 11506 74846
rect 13246 74834 13298 74846
rect 14030 74898 14082 74910
rect 14030 74834 14082 74846
rect 14254 74898 14306 74910
rect 14254 74834 14306 74846
rect 14590 74898 14642 74910
rect 14590 74834 14642 74846
rect 14926 74898 14978 74910
rect 14926 74834 14978 74846
rect 15038 74898 15090 74910
rect 15038 74834 15090 74846
rect 15598 74898 15650 74910
rect 15598 74834 15650 74846
rect 16382 74898 16434 74910
rect 16382 74834 16434 74846
rect 16830 74898 16882 74910
rect 21982 74898 22034 74910
rect 17490 74846 17502 74898
rect 17554 74846 17566 74898
rect 16830 74834 16882 74846
rect 21982 74834 22034 74846
rect 5294 74786 5346 74798
rect 4162 74734 4174 74786
rect 4226 74734 4238 74786
rect 5294 74722 5346 74734
rect 10334 74786 10386 74798
rect 10334 74722 10386 74734
rect 12798 74786 12850 74798
rect 21310 74786 21362 74798
rect 20290 74734 20302 74786
rect 20354 74734 20366 74786
rect 12798 74722 12850 74734
rect 21310 74722 21362 74734
rect 22542 74786 22594 74798
rect 22542 74722 22594 74734
rect 22990 74786 23042 74798
rect 22990 74722 23042 74734
rect 23326 74786 23378 74798
rect 23326 74722 23378 74734
rect 24222 74786 24274 74798
rect 24222 74722 24274 74734
rect 25790 74786 25842 74798
rect 25790 74722 25842 74734
rect 26126 74786 26178 74798
rect 26126 74722 26178 74734
rect 27134 74786 27186 74798
rect 27134 74722 27186 74734
rect 27582 74786 27634 74798
rect 27582 74722 27634 74734
rect 6750 74674 6802 74686
rect 6750 74610 6802 74622
rect 8878 74674 8930 74686
rect 13694 74674 13746 74686
rect 12562 74622 12574 74674
rect 12626 74671 12638 74674
rect 13346 74671 13358 74674
rect 12626 74625 13358 74671
rect 12626 74622 12638 74625
rect 13346 74622 13358 74625
rect 13410 74622 13422 74674
rect 15698 74622 15710 74674
rect 15762 74671 15774 74674
rect 16258 74671 16270 74674
rect 15762 74625 16270 74671
rect 15762 74622 15774 74625
rect 16258 74622 16270 74625
rect 16322 74622 16334 74674
rect 22194 74622 22206 74674
rect 22258 74671 22270 74674
rect 23314 74671 23326 74674
rect 22258 74625 23326 74671
rect 22258 74622 22270 74625
rect 23314 74622 23326 74625
rect 23378 74622 23390 74674
rect 25890 74622 25902 74674
rect 25954 74671 25966 74674
rect 26674 74671 26686 74674
rect 25954 74625 26686 74671
rect 25954 74622 25966 74625
rect 26674 74622 26686 74625
rect 26738 74671 26750 74674
rect 27122 74671 27134 74674
rect 26738 74625 27134 74671
rect 26738 74622 26750 74625
rect 27122 74622 27134 74625
rect 27186 74671 27198 74674
rect 27570 74671 27582 74674
rect 27186 74625 27582 74671
rect 27186 74622 27198 74625
rect 27570 74622 27582 74625
rect 27634 74622 27646 74674
rect 8878 74610 8930 74622
rect 13694 74610 13746 74622
rect 1344 74506 28560 74540
rect 1344 74454 4616 74506
rect 4668 74454 4720 74506
rect 4772 74454 4824 74506
rect 4876 74454 11420 74506
rect 11472 74454 11524 74506
rect 11576 74454 11628 74506
rect 11680 74454 18224 74506
rect 18276 74454 18328 74506
rect 18380 74454 18432 74506
rect 18484 74454 25028 74506
rect 25080 74454 25132 74506
rect 25184 74454 25236 74506
rect 25288 74454 28560 74506
rect 1344 74420 28560 74454
rect 12574 74338 12626 74350
rect 9090 74286 9102 74338
rect 9154 74335 9166 74338
rect 10098 74335 10110 74338
rect 9154 74289 10110 74335
rect 9154 74286 9166 74289
rect 10098 74286 10110 74289
rect 10162 74286 10174 74338
rect 12574 74274 12626 74286
rect 18622 74338 18674 74350
rect 19282 74286 19294 74338
rect 19346 74335 19358 74338
rect 20290 74335 20302 74338
rect 19346 74289 20302 74335
rect 19346 74286 19358 74289
rect 20290 74286 20302 74289
rect 20354 74286 20366 74338
rect 18622 74274 18674 74286
rect 2270 74226 2322 74238
rect 2270 74162 2322 74174
rect 5742 74226 5794 74238
rect 5742 74162 5794 74174
rect 8654 74226 8706 74238
rect 8654 74162 8706 74174
rect 9102 74226 9154 74238
rect 9102 74162 9154 74174
rect 9998 74226 10050 74238
rect 9998 74162 10050 74174
rect 10446 74226 10498 74238
rect 10446 74162 10498 74174
rect 12126 74226 12178 74238
rect 12126 74162 12178 74174
rect 12462 74226 12514 74238
rect 12462 74162 12514 74174
rect 14030 74226 14082 74238
rect 14030 74162 14082 74174
rect 17278 74226 17330 74238
rect 17278 74162 17330 74174
rect 18734 74226 18786 74238
rect 24210 74174 24222 74226
rect 24274 74174 24286 74226
rect 18734 74162 18786 74174
rect 3614 74114 3666 74126
rect 3614 74050 3666 74062
rect 15598 74114 15650 74126
rect 19854 74114 19906 74126
rect 18946 74062 18958 74114
rect 19010 74062 19022 74114
rect 15598 74050 15650 74062
rect 19854 74050 19906 74062
rect 20302 74114 20354 74126
rect 24782 74114 24834 74126
rect 21410 74062 21422 74114
rect 21474 74062 21486 74114
rect 20302 74050 20354 74062
rect 24782 74050 24834 74062
rect 25902 74114 25954 74126
rect 25902 74050 25954 74062
rect 26238 74114 26290 74126
rect 26238 74050 26290 74062
rect 26574 74114 26626 74126
rect 26574 74050 26626 74062
rect 27022 74114 27074 74126
rect 27022 74050 27074 74062
rect 27918 74114 27970 74126
rect 27918 74050 27970 74062
rect 7198 74002 7250 74014
rect 7198 73938 7250 73950
rect 10894 74002 10946 74014
rect 10894 73938 10946 73950
rect 11678 74002 11730 74014
rect 11678 73938 11730 73950
rect 14926 74002 14978 74014
rect 14926 73938 14978 73950
rect 16046 74002 16098 74014
rect 16046 73938 16098 73950
rect 19518 74002 19570 74014
rect 19518 73938 19570 73950
rect 20750 74002 20802 74014
rect 25006 74002 25058 74014
rect 22082 73950 22094 74002
rect 22146 73950 22158 74002
rect 20750 73938 20802 73950
rect 25006 73938 25058 73950
rect 25678 74002 25730 74014
rect 25678 73938 25730 73950
rect 27134 74002 27186 74014
rect 27134 73938 27186 73950
rect 27358 74002 27410 74014
rect 27358 73938 27410 73950
rect 1822 73890 1874 73902
rect 1822 73826 1874 73838
rect 2942 73890 2994 73902
rect 2942 73826 2994 73838
rect 4062 73890 4114 73902
rect 4062 73826 4114 73838
rect 4846 73890 4898 73902
rect 4846 73826 4898 73838
rect 6750 73890 6802 73902
rect 6750 73826 6802 73838
rect 9550 73890 9602 73902
rect 9550 73826 9602 73838
rect 13582 73890 13634 73902
rect 13582 73826 13634 73838
rect 14590 73890 14642 73902
rect 14590 73826 14642 73838
rect 14814 73890 14866 73902
rect 14814 73826 14866 73838
rect 15598 73890 15650 73902
rect 15598 73826 15650 73838
rect 24558 73890 24610 73902
rect 24558 73826 24610 73838
rect 24670 73890 24722 73902
rect 24670 73826 24722 73838
rect 25566 73890 25618 73902
rect 25566 73826 25618 73838
rect 26126 73890 26178 73902
rect 26126 73826 26178 73838
rect 26910 73890 26962 73902
rect 26910 73826 26962 73838
rect 1344 73722 28720 73756
rect 1344 73670 8018 73722
rect 8070 73670 8122 73722
rect 8174 73670 8226 73722
rect 8278 73670 14822 73722
rect 14874 73670 14926 73722
rect 14978 73670 15030 73722
rect 15082 73670 21626 73722
rect 21678 73670 21730 73722
rect 21782 73670 21834 73722
rect 21886 73670 28430 73722
rect 28482 73670 28534 73722
rect 28586 73670 28638 73722
rect 28690 73670 28720 73722
rect 1344 73636 28720 73670
rect 8990 73554 9042 73566
rect 8990 73490 9042 73502
rect 9662 73554 9714 73566
rect 9662 73490 9714 73502
rect 10110 73554 10162 73566
rect 10110 73490 10162 73502
rect 20302 73554 20354 73566
rect 20302 73490 20354 73502
rect 21870 73554 21922 73566
rect 21870 73490 21922 73502
rect 23550 73554 23602 73566
rect 23550 73490 23602 73502
rect 2046 73442 2098 73454
rect 2046 73378 2098 73390
rect 14030 73442 14082 73454
rect 14030 73378 14082 73390
rect 18062 73442 18114 73454
rect 18062 73378 18114 73390
rect 19294 73442 19346 73454
rect 19294 73378 19346 73390
rect 20750 73442 20802 73454
rect 20750 73378 20802 73390
rect 23998 73442 24050 73454
rect 26002 73390 26014 73442
rect 26066 73390 26078 73442
rect 23998 73378 24050 73390
rect 1710 73330 1762 73342
rect 13134 73330 13186 73342
rect 2706 73278 2718 73330
rect 2770 73278 2782 73330
rect 3154 73278 3166 73330
rect 3218 73278 3230 73330
rect 4946 73278 4958 73330
rect 5010 73278 5022 73330
rect 1710 73266 1762 73278
rect 13134 73266 13186 73278
rect 13358 73330 13410 73342
rect 13806 73330 13858 73342
rect 13682 73278 13694 73330
rect 13746 73278 13758 73330
rect 13358 73266 13410 73278
rect 13806 73266 13858 73278
rect 15934 73330 15986 73342
rect 15934 73266 15986 73278
rect 17502 73330 17554 73342
rect 17502 73266 17554 73278
rect 17950 73330 18002 73342
rect 17950 73266 18002 73278
rect 18286 73330 18338 73342
rect 18286 73266 18338 73278
rect 21086 73330 21138 73342
rect 23438 73330 23490 73342
rect 21298 73278 21310 73330
rect 21362 73278 21374 73330
rect 21858 73278 21870 73330
rect 21922 73278 21934 73330
rect 22530 73278 22542 73330
rect 22594 73278 22606 73330
rect 21086 73266 21138 73278
rect 23438 73266 23490 73278
rect 23774 73330 23826 73342
rect 25330 73278 25342 73330
rect 25394 73278 25406 73330
rect 23774 73266 23826 73278
rect 4174 73218 4226 73230
rect 3490 73166 3502 73218
rect 3554 73166 3566 73218
rect 4174 73154 4226 73166
rect 4622 73218 4674 73230
rect 8318 73218 8370 73230
rect 14590 73218 14642 73230
rect 5730 73166 5742 73218
rect 5794 73166 5806 73218
rect 7858 73166 7870 73218
rect 7922 73166 7934 73218
rect 13906 73166 13918 73218
rect 13970 73166 13982 73218
rect 4622 73154 4674 73166
rect 8318 73154 8370 73166
rect 14590 73154 14642 73166
rect 15150 73218 15202 73230
rect 15150 73154 15202 73166
rect 16382 73218 16434 73230
rect 16382 73154 16434 73166
rect 16718 73218 16770 73230
rect 16718 73154 16770 73166
rect 18734 73218 18786 73230
rect 18734 73154 18786 73166
rect 19854 73218 19906 73230
rect 19854 73154 19906 73166
rect 22318 73218 22370 73230
rect 22318 73154 22370 73166
rect 22990 73218 23042 73230
rect 22990 73154 23042 73166
rect 24446 73218 24498 73230
rect 28130 73166 28142 73218
rect 28194 73166 28206 73218
rect 24446 73154 24498 73166
rect 2382 73106 2434 73118
rect 2382 73042 2434 73054
rect 2718 73106 2770 73118
rect 2718 73042 2770 73054
rect 17278 73106 17330 73118
rect 17278 73042 17330 73054
rect 19406 73106 19458 73118
rect 22206 73106 22258 73118
rect 21634 73054 21646 73106
rect 21698 73054 21710 73106
rect 19406 73042 19458 73054
rect 22206 73042 22258 73054
rect 24334 73106 24386 73118
rect 24334 73042 24386 73054
rect 1344 72938 28560 72972
rect 1344 72886 4616 72938
rect 4668 72886 4720 72938
rect 4772 72886 4824 72938
rect 4876 72886 11420 72938
rect 11472 72886 11524 72938
rect 11576 72886 11628 72938
rect 11680 72886 18224 72938
rect 18276 72886 18328 72938
rect 18380 72886 18432 72938
rect 18484 72886 25028 72938
rect 25080 72886 25132 72938
rect 25184 72886 25236 72938
rect 25288 72886 28560 72938
rect 1344 72852 28560 72886
rect 8430 72770 8482 72782
rect 8430 72706 8482 72718
rect 13694 72770 13746 72782
rect 13694 72706 13746 72718
rect 14254 72770 14306 72782
rect 14254 72706 14306 72718
rect 5854 72658 5906 72670
rect 4610 72606 4622 72658
rect 4674 72606 4686 72658
rect 5854 72594 5906 72606
rect 6190 72658 6242 72670
rect 6190 72594 6242 72606
rect 6974 72658 7026 72670
rect 6974 72594 7026 72606
rect 7982 72658 8034 72670
rect 12910 72658 12962 72670
rect 12226 72606 12238 72658
rect 12290 72606 12302 72658
rect 7982 72594 8034 72606
rect 12910 72594 12962 72606
rect 13918 72658 13970 72670
rect 21422 72658 21474 72670
rect 17826 72606 17838 72658
rect 17890 72606 17902 72658
rect 18946 72606 18958 72658
rect 19010 72606 19022 72658
rect 27682 72606 27694 72658
rect 27746 72606 27758 72658
rect 13918 72594 13970 72606
rect 21422 72594 21474 72606
rect 6078 72546 6130 72558
rect 8318 72546 8370 72558
rect 1810 72494 1822 72546
rect 1874 72494 1886 72546
rect 6290 72494 6302 72546
rect 6354 72494 6366 72546
rect 7186 72494 7198 72546
rect 7250 72494 7262 72546
rect 6078 72482 6130 72494
rect 8318 72482 8370 72494
rect 8542 72546 8594 72558
rect 8542 72482 8594 72494
rect 8766 72546 8818 72558
rect 8766 72482 8818 72494
rect 8990 72546 9042 72558
rect 13582 72546 13634 72558
rect 9314 72494 9326 72546
rect 9378 72494 9390 72546
rect 8990 72482 9042 72494
rect 13582 72482 13634 72494
rect 14142 72546 14194 72558
rect 22318 72546 22370 72558
rect 23214 72546 23266 72558
rect 15586 72494 15598 72546
rect 15650 72494 15662 72546
rect 16370 72494 16382 72546
rect 16434 72494 16446 72546
rect 18610 72494 18622 72546
rect 18674 72494 18686 72546
rect 19170 72494 19182 72546
rect 19234 72494 19246 72546
rect 22418 72494 22430 72546
rect 22482 72494 22494 72546
rect 22978 72494 22990 72546
rect 23042 72494 23054 72546
rect 14142 72482 14194 72494
rect 22318 72482 22370 72494
rect 23214 72482 23266 72494
rect 23438 72546 23490 72558
rect 25666 72494 25678 72546
rect 25730 72494 25742 72546
rect 23438 72482 23490 72494
rect 5070 72434 5122 72446
rect 2482 72382 2494 72434
rect 2546 72382 2558 72434
rect 5070 72370 5122 72382
rect 5742 72434 5794 72446
rect 5742 72370 5794 72382
rect 6862 72434 6914 72446
rect 21870 72434 21922 72446
rect 10098 72382 10110 72434
rect 10162 72382 10174 72434
rect 15250 72382 15262 72434
rect 15314 72382 15326 72434
rect 16258 72382 16270 72434
rect 16322 72382 16334 72434
rect 18498 72382 18510 72434
rect 18562 72382 18574 72434
rect 22082 72382 22094 72434
rect 22146 72382 22158 72434
rect 6862 72370 6914 72382
rect 21870 72370 21922 72382
rect 19518 72322 19570 72334
rect 19518 72258 19570 72270
rect 20190 72322 20242 72334
rect 20190 72258 20242 72270
rect 20638 72322 20690 72334
rect 23326 72322 23378 72334
rect 22194 72270 22206 72322
rect 22258 72270 22270 72322
rect 20638 72258 20690 72270
rect 23326 72258 23378 72270
rect 23550 72322 23602 72334
rect 23550 72258 23602 72270
rect 24110 72322 24162 72334
rect 24110 72258 24162 72270
rect 24558 72322 24610 72334
rect 24558 72258 24610 72270
rect 25006 72322 25058 72334
rect 25006 72258 25058 72270
rect 1344 72154 28720 72188
rect 1344 72102 8018 72154
rect 8070 72102 8122 72154
rect 8174 72102 8226 72154
rect 8278 72102 14822 72154
rect 14874 72102 14926 72154
rect 14978 72102 15030 72154
rect 15082 72102 21626 72154
rect 21678 72102 21730 72154
rect 21782 72102 21834 72154
rect 21886 72102 28430 72154
rect 28482 72102 28534 72154
rect 28586 72102 28638 72154
rect 28690 72102 28720 72154
rect 1344 72068 28720 72102
rect 7646 71986 7698 71998
rect 2482 71934 2494 71986
rect 2546 71934 2558 71986
rect 7646 71922 7698 71934
rect 8542 71986 8594 71998
rect 8542 71922 8594 71934
rect 8878 71986 8930 71998
rect 8878 71922 8930 71934
rect 10558 71986 10610 71998
rect 10558 71922 10610 71934
rect 11678 71986 11730 71998
rect 11678 71922 11730 71934
rect 12462 71986 12514 71998
rect 12462 71922 12514 71934
rect 12910 71986 12962 71998
rect 12910 71922 12962 71934
rect 14366 71986 14418 71998
rect 14366 71922 14418 71934
rect 15150 71986 15202 71998
rect 23550 71986 23602 71998
rect 18834 71934 18846 71986
rect 18898 71934 18910 71986
rect 15150 71922 15202 71934
rect 23550 71922 23602 71934
rect 24558 71986 24610 71998
rect 24558 71922 24610 71934
rect 26462 71986 26514 71998
rect 26462 71922 26514 71934
rect 27470 71986 27522 71998
rect 27470 71922 27522 71934
rect 28142 71986 28194 71998
rect 28142 71922 28194 71934
rect 2270 71874 2322 71886
rect 2270 71810 2322 71822
rect 10446 71874 10498 71886
rect 10446 71810 10498 71822
rect 11006 71874 11058 71886
rect 11006 71810 11058 71822
rect 11566 71874 11618 71886
rect 11566 71810 11618 71822
rect 14254 71874 14306 71886
rect 14254 71810 14306 71822
rect 16382 71874 16434 71886
rect 19394 71822 19406 71874
rect 19458 71822 19470 71874
rect 21970 71822 21982 71874
rect 22034 71822 22046 71874
rect 16382 71810 16434 71822
rect 2606 71762 2658 71774
rect 2606 71698 2658 71710
rect 2718 71762 2770 71774
rect 3390 71762 3442 71774
rect 8766 71762 8818 71774
rect 3042 71710 3054 71762
rect 3106 71710 3118 71762
rect 4386 71710 4398 71762
rect 4450 71710 4462 71762
rect 5058 71710 5070 71762
rect 5122 71710 5134 71762
rect 2718 71698 2770 71710
rect 3390 71698 3442 71710
rect 8766 71698 8818 71710
rect 8990 71762 9042 71774
rect 8990 71698 9042 71710
rect 9550 71762 9602 71774
rect 9550 71698 9602 71710
rect 9774 71762 9826 71774
rect 9774 71698 9826 71710
rect 10222 71762 10274 71774
rect 10222 71698 10274 71710
rect 10782 71762 10834 71774
rect 10782 71698 10834 71710
rect 11454 71762 11506 71774
rect 11454 71698 11506 71710
rect 12126 71762 12178 71774
rect 12126 71698 12178 71710
rect 15710 71762 15762 71774
rect 15710 71698 15762 71710
rect 15934 71762 15986 71774
rect 15934 71698 15986 71710
rect 16158 71762 16210 71774
rect 16158 71698 16210 71710
rect 17502 71762 17554 71774
rect 17502 71698 17554 71710
rect 17950 71762 18002 71774
rect 17950 71698 18002 71710
rect 18062 71762 18114 71774
rect 23438 71762 23490 71774
rect 19058 71710 19070 71762
rect 19122 71710 19134 71762
rect 20402 71710 20414 71762
rect 20466 71710 20478 71762
rect 22642 71710 22654 71762
rect 22706 71710 22718 71762
rect 18062 71698 18114 71710
rect 23438 71698 23490 71710
rect 23774 71762 23826 71774
rect 26686 71762 26738 71774
rect 23986 71710 23998 71762
rect 24050 71710 24062 71762
rect 24322 71710 24334 71762
rect 24386 71710 24398 71762
rect 23774 71698 23826 71710
rect 26686 71698 26738 71710
rect 27134 71762 27186 71774
rect 27134 71698 27186 71710
rect 3502 71650 3554 71662
rect 3502 71586 3554 71598
rect 3950 71650 4002 71662
rect 8094 71650 8146 71662
rect 7186 71598 7198 71650
rect 7250 71598 7262 71650
rect 3950 71586 4002 71598
rect 8094 71586 8146 71598
rect 9662 71650 9714 71662
rect 18286 71650 18338 71662
rect 16258 71598 16270 71650
rect 16322 71598 16334 71650
rect 9662 71586 9714 71598
rect 18286 71586 18338 71598
rect 23662 71650 23714 71662
rect 23662 71586 23714 71598
rect 25342 71650 25394 71662
rect 25342 71586 25394 71598
rect 26014 71650 26066 71662
rect 26014 71586 26066 71598
rect 26574 71650 26626 71662
rect 26574 71586 26626 71598
rect 13470 71538 13522 71550
rect 7522 71486 7534 71538
rect 7586 71535 7598 71538
rect 8082 71535 8094 71538
rect 7586 71489 8094 71535
rect 7586 71486 7598 71489
rect 8082 71486 8094 71489
rect 8146 71486 8158 71538
rect 13470 71474 13522 71486
rect 13582 71538 13634 71550
rect 13582 71474 13634 71486
rect 13806 71538 13858 71550
rect 13806 71474 13858 71486
rect 13918 71538 13970 71550
rect 13918 71474 13970 71486
rect 15486 71538 15538 71550
rect 15486 71474 15538 71486
rect 17278 71538 17330 71550
rect 17278 71474 17330 71486
rect 24670 71538 24722 71550
rect 24670 71474 24722 71486
rect 1344 71370 28560 71404
rect 1344 71318 4616 71370
rect 4668 71318 4720 71370
rect 4772 71318 4824 71370
rect 4876 71318 11420 71370
rect 11472 71318 11524 71370
rect 11576 71318 11628 71370
rect 11680 71318 18224 71370
rect 18276 71318 18328 71370
rect 18380 71318 18432 71370
rect 18484 71318 25028 71370
rect 25080 71318 25132 71370
rect 25184 71318 25236 71370
rect 25288 71318 28560 71370
rect 1344 71284 28560 71318
rect 8430 71202 8482 71214
rect 3490 71150 3502 71202
rect 3554 71199 3566 71202
rect 3938 71199 3950 71202
rect 3554 71153 3950 71199
rect 3554 71150 3566 71153
rect 3938 71150 3950 71153
rect 4002 71150 4014 71202
rect 7298 71150 7310 71202
rect 7362 71199 7374 71202
rect 8082 71199 8094 71202
rect 7362 71153 8094 71199
rect 7362 71150 7374 71153
rect 8082 71150 8094 71153
rect 8146 71150 8158 71202
rect 8430 71138 8482 71150
rect 14926 71202 14978 71214
rect 14926 71138 14978 71150
rect 15150 71202 15202 71214
rect 15150 71138 15202 71150
rect 5742 71090 5794 71102
rect 5742 71026 5794 71038
rect 8318 71090 8370 71102
rect 8318 71026 8370 71038
rect 8878 71090 8930 71102
rect 8878 71026 8930 71038
rect 9550 71090 9602 71102
rect 9550 71026 9602 71038
rect 13582 71090 13634 71102
rect 15374 71090 15426 71102
rect 14242 71038 14254 71090
rect 14306 71038 14318 71090
rect 13582 71026 13634 71038
rect 15374 71026 15426 71038
rect 18846 71090 18898 71102
rect 22194 71038 22206 71090
rect 22258 71038 22270 71090
rect 24322 71038 24334 71090
rect 24386 71038 24398 71090
rect 28130 71038 28142 71090
rect 28194 71038 28206 71090
rect 18846 71026 18898 71038
rect 3502 70978 3554 70990
rect 1810 70926 1822 70978
rect 1874 70926 1886 70978
rect 3502 70914 3554 70926
rect 6078 70978 6130 70990
rect 6862 70978 6914 70990
rect 11230 70978 11282 70990
rect 6178 70926 6190 70978
rect 6242 70926 6254 70978
rect 7074 70926 7086 70978
rect 7138 70926 7150 70978
rect 9986 70926 9998 70978
rect 10050 70926 10062 70978
rect 6078 70914 6130 70926
rect 6862 70914 6914 70926
rect 11230 70914 11282 70926
rect 13806 70978 13858 70990
rect 13806 70914 13858 70926
rect 14030 70978 14082 70990
rect 14030 70914 14082 70926
rect 14478 70978 14530 70990
rect 16818 70926 16830 70978
rect 16882 70926 16894 70978
rect 17266 70926 17278 70978
rect 17330 70926 17342 70978
rect 19282 70926 19294 70978
rect 19346 70926 19358 70978
rect 20178 70926 20190 70978
rect 20242 70926 20254 70978
rect 21522 70926 21534 70978
rect 21586 70926 21598 70978
rect 25330 70926 25342 70978
rect 25394 70926 25406 70978
rect 14478 70914 14530 70926
rect 4622 70866 4674 70878
rect 4622 70802 4674 70814
rect 5630 70866 5682 70878
rect 6750 70866 6802 70878
rect 5842 70814 5854 70866
rect 5906 70814 5918 70866
rect 5630 70802 5682 70814
rect 6750 70802 6802 70814
rect 14254 70866 14306 70878
rect 18398 70866 18450 70878
rect 16258 70814 16270 70866
rect 16322 70814 16334 70866
rect 17938 70814 17950 70866
rect 18002 70814 18014 70866
rect 20738 70814 20750 70866
rect 20802 70814 20814 70866
rect 26002 70814 26014 70866
rect 26066 70814 26078 70866
rect 14254 70802 14306 70814
rect 18398 70802 18450 70814
rect 2046 70754 2098 70766
rect 2046 70690 2098 70702
rect 2606 70754 2658 70766
rect 2606 70690 2658 70702
rect 3054 70754 3106 70766
rect 3054 70690 3106 70702
rect 3950 70754 4002 70766
rect 3950 70690 4002 70702
rect 5182 70754 5234 70766
rect 5182 70690 5234 70702
rect 7534 70754 7586 70766
rect 7534 70690 7586 70702
rect 7982 70754 8034 70766
rect 7982 70690 8034 70702
rect 9438 70754 9490 70766
rect 9438 70690 9490 70702
rect 9662 70754 9714 70766
rect 9662 70690 9714 70702
rect 10446 70754 10498 70766
rect 10446 70690 10498 70702
rect 12462 70754 12514 70766
rect 12462 70690 12514 70702
rect 12910 70754 12962 70766
rect 12910 70690 12962 70702
rect 15598 70754 15650 70766
rect 15598 70690 15650 70702
rect 15710 70754 15762 70766
rect 15710 70690 15762 70702
rect 15822 70754 15874 70766
rect 18286 70754 18338 70766
rect 17826 70702 17838 70754
rect 17890 70702 17902 70754
rect 15822 70690 15874 70702
rect 18286 70690 18338 70702
rect 19518 70754 19570 70766
rect 24782 70754 24834 70766
rect 19618 70702 19630 70754
rect 19682 70702 19694 70754
rect 19518 70690 19570 70702
rect 24782 70690 24834 70702
rect 1344 70586 28720 70620
rect 1344 70534 8018 70586
rect 8070 70534 8122 70586
rect 8174 70534 8226 70586
rect 8278 70534 14822 70586
rect 14874 70534 14926 70586
rect 14978 70534 15030 70586
rect 15082 70534 21626 70586
rect 21678 70534 21730 70586
rect 21782 70534 21834 70586
rect 21886 70534 28430 70586
rect 28482 70534 28534 70586
rect 28586 70534 28638 70586
rect 28690 70534 28720 70586
rect 1344 70500 28720 70534
rect 2270 70418 2322 70430
rect 2270 70354 2322 70366
rect 9774 70418 9826 70430
rect 10894 70418 10946 70430
rect 10210 70366 10222 70418
rect 10274 70366 10286 70418
rect 9774 70354 9826 70366
rect 10894 70354 10946 70366
rect 11342 70418 11394 70430
rect 11342 70354 11394 70366
rect 13022 70418 13074 70430
rect 13022 70354 13074 70366
rect 21310 70418 21362 70430
rect 21310 70354 21362 70366
rect 25678 70418 25730 70430
rect 25678 70354 25730 70366
rect 26126 70418 26178 70430
rect 26126 70354 26178 70366
rect 27918 70418 27970 70430
rect 27918 70354 27970 70366
rect 9550 70306 9602 70318
rect 26350 70306 26402 70318
rect 15026 70254 15038 70306
rect 15090 70254 15102 70306
rect 15922 70254 15934 70306
rect 15986 70254 15998 70306
rect 9550 70242 9602 70254
rect 26350 70242 26402 70254
rect 26574 70306 26626 70318
rect 26574 70242 26626 70254
rect 27022 70306 27074 70318
rect 27022 70242 27074 70254
rect 9998 70194 10050 70206
rect 2706 70142 2718 70194
rect 2770 70142 2782 70194
rect 7858 70142 7870 70194
rect 7922 70142 7934 70194
rect 9998 70130 10050 70142
rect 10222 70194 10274 70206
rect 10222 70130 10274 70142
rect 12238 70194 12290 70206
rect 12238 70130 12290 70142
rect 12462 70194 12514 70206
rect 12462 70130 12514 70142
rect 12910 70194 12962 70206
rect 12910 70130 12962 70142
rect 13134 70194 13186 70206
rect 25902 70194 25954 70206
rect 15250 70142 15262 70194
rect 15314 70142 15326 70194
rect 15586 70142 15598 70194
rect 15650 70142 15662 70194
rect 17378 70142 17390 70194
rect 17442 70142 17454 70194
rect 22082 70142 22094 70194
rect 22146 70142 22158 70194
rect 13134 70130 13186 70142
rect 25902 70130 25954 70142
rect 11902 70082 11954 70094
rect 3042 70030 3054 70082
rect 3106 70030 3118 70082
rect 5058 70030 5070 70082
rect 5122 70030 5134 70082
rect 11902 70018 11954 70030
rect 12686 70082 12738 70094
rect 20750 70082 20802 70094
rect 14242 70030 14254 70082
rect 14306 70030 14318 70082
rect 18162 70030 18174 70082
rect 18226 70030 18238 70082
rect 20290 70030 20302 70082
rect 20354 70030 20366 70082
rect 12686 70018 12738 70030
rect 20750 70018 20802 70030
rect 21758 70082 21810 70094
rect 27470 70082 27522 70094
rect 23874 70030 23886 70082
rect 23938 70030 23950 70082
rect 21758 70018 21810 70030
rect 27470 70018 27522 70030
rect 2046 69970 2098 69982
rect 2046 69906 2098 69918
rect 2382 69970 2434 69982
rect 2382 69906 2434 69918
rect 26910 69970 26962 69982
rect 26910 69906 26962 69918
rect 1344 69802 28560 69836
rect 1344 69750 4616 69802
rect 4668 69750 4720 69802
rect 4772 69750 4824 69802
rect 4876 69750 11420 69802
rect 11472 69750 11524 69802
rect 11576 69750 11628 69802
rect 11680 69750 18224 69802
rect 18276 69750 18328 69802
rect 18380 69750 18432 69802
rect 18484 69750 25028 69802
rect 25080 69750 25132 69802
rect 25184 69750 25236 69802
rect 25288 69750 28560 69802
rect 1344 69716 28560 69750
rect 8318 69634 8370 69646
rect 12686 69634 12738 69646
rect 11778 69582 11790 69634
rect 11842 69631 11854 69634
rect 12338 69631 12350 69634
rect 11842 69585 12350 69631
rect 11842 69582 11854 69585
rect 12338 69582 12350 69585
rect 12402 69582 12414 69634
rect 8318 69570 8370 69582
rect 12686 69570 12738 69582
rect 13358 69522 13410 69534
rect 19406 69522 19458 69534
rect 4610 69470 4622 69522
rect 4674 69470 4686 69522
rect 16482 69470 16494 69522
rect 16546 69470 16558 69522
rect 13358 69458 13410 69470
rect 19406 69458 19458 69470
rect 21646 69522 21698 69534
rect 25342 69522 25394 69534
rect 21970 69470 21982 69522
rect 22034 69470 22046 69522
rect 23538 69470 23550 69522
rect 23602 69470 23614 69522
rect 21646 69458 21698 69470
rect 25342 69458 25394 69470
rect 25790 69522 25842 69534
rect 25790 69458 25842 69470
rect 8206 69410 8258 69422
rect 1698 69358 1710 69410
rect 1762 69358 1774 69410
rect 8206 69346 8258 69358
rect 8766 69410 8818 69422
rect 8766 69346 8818 69358
rect 13470 69410 13522 69422
rect 13470 69346 13522 69358
rect 14030 69410 14082 69422
rect 14030 69346 14082 69358
rect 14814 69410 14866 69422
rect 18286 69410 18338 69422
rect 15810 69358 15822 69410
rect 15874 69358 15886 69410
rect 16258 69358 16270 69410
rect 16322 69358 16334 69410
rect 14814 69346 14866 69358
rect 18286 69346 18338 69358
rect 18958 69410 19010 69422
rect 18958 69346 19010 69358
rect 19518 69410 19570 69422
rect 26686 69410 26738 69422
rect 19842 69358 19854 69410
rect 19906 69358 19918 69410
rect 22306 69358 22318 69410
rect 22370 69358 22382 69410
rect 19518 69346 19570 69358
rect 26686 69346 26738 69358
rect 27582 69410 27634 69422
rect 27582 69346 27634 69358
rect 9326 69298 9378 69310
rect 2482 69246 2494 69298
rect 2546 69246 2558 69298
rect 9326 69234 9378 69246
rect 12574 69298 12626 69310
rect 18734 69298 18786 69310
rect 15250 69246 15262 69298
rect 15314 69246 15326 69298
rect 16818 69246 16830 69298
rect 16882 69246 16894 69298
rect 12574 69234 12626 69246
rect 18734 69234 18786 69246
rect 26350 69298 26402 69310
rect 26350 69234 26402 69246
rect 26910 69298 26962 69310
rect 26910 69234 26962 69246
rect 27246 69298 27298 69310
rect 27246 69234 27298 69246
rect 27806 69298 27858 69310
rect 27806 69234 27858 69246
rect 5070 69186 5122 69198
rect 5070 69122 5122 69134
rect 7870 69186 7922 69198
rect 7870 69122 7922 69134
rect 9214 69186 9266 69198
rect 9214 69122 9266 69134
rect 9438 69186 9490 69198
rect 9438 69122 9490 69134
rect 10446 69186 10498 69198
rect 10446 69122 10498 69134
rect 11790 69186 11842 69198
rect 11790 69122 11842 69134
rect 12238 69186 12290 69198
rect 12238 69122 12290 69134
rect 13694 69186 13746 69198
rect 13694 69122 13746 69134
rect 13918 69186 13970 69198
rect 13918 69122 13970 69134
rect 17390 69186 17442 69198
rect 17390 69122 17442 69134
rect 17838 69186 17890 69198
rect 17838 69122 17890 69134
rect 18622 69186 18674 69198
rect 18622 69122 18674 69134
rect 19294 69186 19346 69198
rect 19294 69122 19346 69134
rect 20414 69186 20466 69198
rect 20414 69122 20466 69134
rect 20750 69186 20802 69198
rect 20750 69122 20802 69134
rect 26574 69186 26626 69198
rect 26574 69122 26626 69134
rect 27582 69186 27634 69198
rect 27582 69122 27634 69134
rect 1344 69018 28720 69052
rect 1344 68966 8018 69018
rect 8070 68966 8122 69018
rect 8174 68966 8226 69018
rect 8278 68966 14822 69018
rect 14874 68966 14926 69018
rect 14978 68966 15030 69018
rect 15082 68966 21626 69018
rect 21678 68966 21730 69018
rect 21782 68966 21834 69018
rect 21886 68966 28430 69018
rect 28482 68966 28534 69018
rect 28586 68966 28638 69018
rect 28690 68966 28720 69018
rect 1344 68932 28720 68966
rect 8430 68850 8482 68862
rect 2594 68798 2606 68850
rect 2658 68798 2670 68850
rect 8430 68786 8482 68798
rect 8990 68850 9042 68862
rect 8990 68786 9042 68798
rect 14926 68850 14978 68862
rect 14926 68786 14978 68798
rect 15374 68850 15426 68862
rect 15374 68786 15426 68798
rect 16830 68850 16882 68862
rect 16830 68786 16882 68798
rect 19406 68850 19458 68862
rect 19406 68786 19458 68798
rect 20302 68850 20354 68862
rect 20302 68786 20354 68798
rect 20750 68850 20802 68862
rect 20750 68786 20802 68798
rect 3054 68738 3106 68750
rect 17838 68738 17890 68750
rect 12786 68686 12798 68738
rect 12850 68686 12862 68738
rect 27346 68686 27358 68738
rect 27410 68686 27422 68738
rect 3054 68674 3106 68686
rect 17838 68674 17890 68686
rect 3390 68626 3442 68638
rect 17390 68626 17442 68638
rect 2482 68574 2494 68626
rect 2546 68574 2558 68626
rect 2818 68574 2830 68626
rect 2882 68574 2894 68626
rect 4834 68574 4846 68626
rect 4898 68574 4910 68626
rect 9538 68574 9550 68626
rect 9602 68574 9614 68626
rect 14018 68574 14030 68626
rect 14082 68574 14094 68626
rect 3390 68562 3442 68574
rect 17390 68562 17442 68574
rect 17614 68626 17666 68638
rect 22306 68574 22318 68626
rect 22370 68574 22382 68626
rect 28130 68574 28142 68626
rect 28194 68574 28206 68626
rect 17614 68562 17666 68574
rect 3502 68514 3554 68526
rect 3502 68450 3554 68462
rect 3950 68514 4002 68526
rect 3950 68450 4002 68462
rect 4398 68514 4450 68526
rect 8318 68514 8370 68526
rect 17502 68514 17554 68526
rect 5506 68462 5518 68514
rect 5570 68462 5582 68514
rect 7634 68462 7646 68514
rect 7698 68462 7710 68514
rect 10322 68462 10334 68514
rect 10386 68462 10398 68514
rect 12450 68462 12462 68514
rect 12514 68462 12526 68514
rect 14242 68462 14254 68514
rect 14306 68462 14318 68514
rect 4398 68450 4450 68462
rect 8318 68450 8370 68462
rect 17502 68450 17554 68462
rect 18510 68514 18562 68526
rect 18510 68450 18562 68462
rect 18958 68514 19010 68526
rect 18958 68450 19010 68462
rect 19854 68514 19906 68526
rect 19854 68450 19906 68462
rect 21198 68514 21250 68526
rect 21198 68450 21250 68462
rect 21758 68514 21810 68526
rect 24210 68462 24222 68514
rect 24274 68462 24286 68514
rect 25218 68462 25230 68514
rect 25282 68462 25294 68514
rect 21758 68450 21810 68462
rect 2482 68350 2494 68402
rect 2546 68350 2558 68402
rect 3938 68350 3950 68402
rect 4002 68399 4014 68402
rect 4498 68399 4510 68402
rect 4002 68353 4510 68399
rect 4002 68350 4014 68353
rect 4498 68350 4510 68353
rect 4562 68350 4574 68402
rect 19282 68350 19294 68402
rect 19346 68399 19358 68402
rect 19954 68399 19966 68402
rect 19346 68353 19966 68399
rect 19346 68350 19358 68353
rect 19954 68350 19966 68353
rect 20018 68399 20030 68402
rect 21186 68399 21198 68402
rect 20018 68353 21198 68399
rect 20018 68350 20030 68353
rect 21186 68350 21198 68353
rect 21250 68350 21262 68402
rect 1344 68234 28560 68268
rect 1344 68182 4616 68234
rect 4668 68182 4720 68234
rect 4772 68182 4824 68234
rect 4876 68182 11420 68234
rect 11472 68182 11524 68234
rect 11576 68182 11628 68234
rect 11680 68182 18224 68234
rect 18276 68182 18328 68234
rect 18380 68182 18432 68234
rect 18484 68182 25028 68234
rect 25080 68182 25132 68234
rect 25184 68182 25236 68234
rect 25288 68182 28560 68234
rect 1344 68148 28560 68182
rect 3278 67954 3330 67966
rect 3278 67890 3330 67902
rect 6078 67954 6130 67966
rect 6078 67890 6130 67902
rect 7758 67954 7810 67966
rect 7758 67890 7810 67902
rect 10446 67954 10498 67966
rect 10446 67890 10498 67902
rect 12910 67954 12962 67966
rect 12910 67890 12962 67902
rect 13470 67954 13522 67966
rect 21646 67954 21698 67966
rect 27022 67954 27074 67966
rect 16034 67902 16046 67954
rect 16098 67902 16110 67954
rect 24210 67902 24222 67954
rect 24274 67902 24286 67954
rect 13470 67890 13522 67902
rect 21646 67890 21698 67902
rect 27022 67890 27074 67902
rect 28142 67954 28194 67966
rect 28142 67890 28194 67902
rect 10222 67842 10274 67854
rect 10222 67778 10274 67790
rect 10894 67842 10946 67854
rect 10894 67778 10946 67790
rect 11566 67842 11618 67854
rect 11566 67778 11618 67790
rect 11678 67842 11730 67854
rect 13694 67842 13746 67854
rect 22878 67842 22930 67854
rect 12002 67790 12014 67842
rect 12066 67790 12078 67842
rect 18946 67790 18958 67842
rect 19010 67790 19022 67842
rect 19282 67790 19294 67842
rect 19346 67790 19358 67842
rect 20178 67790 20190 67842
rect 20242 67790 20254 67842
rect 21858 67790 21870 67842
rect 21922 67790 21934 67842
rect 26002 67790 26014 67842
rect 26066 67790 26078 67842
rect 11678 67778 11730 67790
rect 13694 67778 13746 67790
rect 22878 67778 22930 67790
rect 5182 67730 5234 67742
rect 5182 67666 5234 67678
rect 5966 67730 6018 67742
rect 5966 67666 6018 67678
rect 6302 67730 6354 67742
rect 6302 67666 6354 67678
rect 6526 67730 6578 67742
rect 6526 67666 6578 67678
rect 10670 67730 10722 67742
rect 21534 67730 21586 67742
rect 14018 67678 14030 67730
rect 14082 67678 14094 67730
rect 18162 67678 18174 67730
rect 18226 67678 18238 67730
rect 20514 67678 20526 67730
rect 20578 67678 20590 67730
rect 10670 67666 10722 67678
rect 21534 67666 21586 67678
rect 23214 67730 23266 67742
rect 23214 67666 23266 67678
rect 27358 67730 27410 67742
rect 27358 67666 27410 67678
rect 1822 67618 1874 67630
rect 1822 67554 1874 67566
rect 7086 67618 7138 67630
rect 7086 67554 7138 67566
rect 9662 67618 9714 67630
rect 9662 67554 9714 67566
rect 9998 67618 10050 67630
rect 9998 67554 10050 67566
rect 11454 67618 11506 67630
rect 11454 67554 11506 67566
rect 12462 67618 12514 67630
rect 12462 67554 12514 67566
rect 14478 67618 14530 67630
rect 22318 67618 22370 67630
rect 19394 67566 19406 67618
rect 19458 67566 19470 67618
rect 19618 67566 19630 67618
rect 19682 67566 19694 67618
rect 14478 67554 14530 67566
rect 22318 67554 22370 67566
rect 22990 67618 23042 67630
rect 22990 67554 23042 67566
rect 23102 67618 23154 67630
rect 23102 67554 23154 67566
rect 23326 67618 23378 67630
rect 23326 67554 23378 67566
rect 26910 67618 26962 67630
rect 26910 67554 26962 67566
rect 27134 67618 27186 67630
rect 27134 67554 27186 67566
rect 1344 67450 28720 67484
rect 1344 67398 8018 67450
rect 8070 67398 8122 67450
rect 8174 67398 8226 67450
rect 8278 67398 14822 67450
rect 14874 67398 14926 67450
rect 14978 67398 15030 67450
rect 15082 67398 21626 67450
rect 21678 67398 21730 67450
rect 21782 67398 21834 67450
rect 21886 67398 28430 67450
rect 28482 67398 28534 67450
rect 28586 67398 28638 67450
rect 28690 67398 28720 67450
rect 1344 67364 28720 67398
rect 8094 67282 8146 67294
rect 8094 67218 8146 67230
rect 11342 67282 11394 67294
rect 14030 67282 14082 67294
rect 13122 67230 13134 67282
rect 13186 67230 13198 67282
rect 11342 67218 11394 67230
rect 14030 67218 14082 67230
rect 17838 67282 17890 67294
rect 17838 67218 17890 67230
rect 18734 67282 18786 67294
rect 18734 67218 18786 67230
rect 2046 67170 2098 67182
rect 17950 67170 18002 67182
rect 15810 67118 15822 67170
rect 15874 67118 15886 67170
rect 16706 67118 16718 67170
rect 16770 67118 16782 67170
rect 2046 67106 2098 67118
rect 17950 67106 18002 67118
rect 19406 67170 19458 67182
rect 19406 67106 19458 67118
rect 24446 67170 24498 67182
rect 24446 67106 24498 67118
rect 24558 67170 24610 67182
rect 24558 67106 24610 67118
rect 24670 67170 24722 67182
rect 27346 67118 27358 67170
rect 27410 67118 27422 67170
rect 24670 67106 24722 67118
rect 1710 67058 1762 67070
rect 7870 67058 7922 67070
rect 8878 67058 8930 67070
rect 2706 67006 2718 67058
rect 2770 67006 2782 67058
rect 3042 67006 3054 67058
rect 3106 67006 3118 67058
rect 4722 67006 4734 67058
rect 4786 67006 4798 67058
rect 8418 67006 8430 67058
rect 8482 67006 8494 67058
rect 1710 66994 1762 67006
rect 7870 66994 7922 67006
rect 8878 66994 8930 67006
rect 11566 67058 11618 67070
rect 11566 66994 11618 67006
rect 12014 67058 12066 67070
rect 12014 66994 12066 67006
rect 12574 67058 12626 67070
rect 12574 66994 12626 67006
rect 16158 67058 16210 67070
rect 16158 66994 16210 67006
rect 17502 67058 17554 67070
rect 17502 66994 17554 67006
rect 17614 67058 17666 67070
rect 17614 66994 17666 67006
rect 18398 67058 18450 67070
rect 19518 67058 19570 67070
rect 19058 67006 19070 67058
rect 19122 67006 19134 67058
rect 18398 66994 18450 67006
rect 19518 66994 19570 67006
rect 19630 67058 19682 67070
rect 23998 67058 24050 67070
rect 20178 67006 20190 67058
rect 20242 67006 20254 67058
rect 28130 67006 28142 67058
rect 28194 67006 28206 67058
rect 19630 66994 19682 67006
rect 23998 66994 24050 67006
rect 3838 66946 3890 66958
rect 7982 66946 8034 66958
rect 9662 66946 9714 66958
rect 5394 66894 5406 66946
rect 5458 66894 5470 66946
rect 7522 66894 7534 66946
rect 7586 66894 7598 66946
rect 8418 66894 8430 66946
rect 8482 66943 8494 66946
rect 8754 66943 8766 66946
rect 8482 66897 8766 66943
rect 8482 66894 8494 66897
rect 8754 66894 8766 66897
rect 8818 66894 8830 66946
rect 3838 66882 3890 66894
rect 7982 66882 8034 66894
rect 9662 66882 9714 66894
rect 11006 66946 11058 66958
rect 11006 66882 11058 66894
rect 11454 66946 11506 66958
rect 11454 66882 11506 66894
rect 13582 66946 13634 66958
rect 13582 66882 13634 66894
rect 15262 66946 15314 66958
rect 23438 66946 23490 66958
rect 20850 66894 20862 66946
rect 20914 66894 20926 66946
rect 22978 66894 22990 66946
rect 23042 66894 23054 66946
rect 25218 66894 25230 66946
rect 25282 66894 25294 66946
rect 15262 66882 15314 66894
rect 23438 66882 23490 66894
rect 2382 66834 2434 66846
rect 2382 66770 2434 66782
rect 2718 66834 2770 66846
rect 2718 66770 2770 66782
rect 3166 66834 3218 66846
rect 12798 66834 12850 66846
rect 10770 66782 10782 66834
rect 10834 66831 10846 66834
rect 11106 66831 11118 66834
rect 10834 66785 11118 66831
rect 10834 66782 10846 66785
rect 11106 66782 11118 66785
rect 11170 66782 11182 66834
rect 3166 66770 3218 66782
rect 12798 66770 12850 66782
rect 15486 66834 15538 66846
rect 15486 66770 15538 66782
rect 16382 66834 16434 66846
rect 16382 66770 16434 66782
rect 1344 66666 28560 66700
rect 1344 66614 4616 66666
rect 4668 66614 4720 66666
rect 4772 66614 4824 66666
rect 4876 66614 11420 66666
rect 11472 66614 11524 66666
rect 11576 66614 11628 66666
rect 11680 66614 18224 66666
rect 18276 66614 18328 66666
rect 18380 66614 18432 66666
rect 18484 66614 25028 66666
rect 25080 66614 25132 66666
rect 25184 66614 25236 66666
rect 25288 66614 28560 66666
rect 1344 66580 28560 66614
rect 21522 66446 21534 66498
rect 21586 66446 21598 66498
rect 5966 66386 6018 66398
rect 12910 66386 12962 66398
rect 4610 66334 4622 66386
rect 4674 66334 4686 66386
rect 9538 66334 9550 66386
rect 9602 66334 9614 66386
rect 16370 66334 16382 66386
rect 16434 66334 16446 66386
rect 17826 66334 17838 66386
rect 17890 66334 17902 66386
rect 27906 66334 27918 66386
rect 27970 66334 27982 66386
rect 5966 66322 6018 66334
rect 12910 66322 12962 66334
rect 6078 66274 6130 66286
rect 1698 66222 1710 66274
rect 1762 66222 1774 66274
rect 6078 66210 6130 66222
rect 6414 66274 6466 66286
rect 8306 66222 8318 66274
rect 8370 66222 8382 66274
rect 13458 66222 13470 66274
rect 13522 66222 13534 66274
rect 14242 66222 14254 66274
rect 14306 66222 14318 66274
rect 17490 66222 17502 66274
rect 17554 66222 17566 66274
rect 18498 66222 18510 66274
rect 18562 66222 18574 66274
rect 21522 66222 21534 66274
rect 21586 66222 21598 66274
rect 22866 66222 22878 66274
rect 22930 66222 22942 66274
rect 6414 66210 6466 66222
rect 5182 66162 5234 66174
rect 2482 66110 2494 66162
rect 2546 66110 2558 66162
rect 5182 66098 5234 66110
rect 5854 66162 5906 66174
rect 5854 66098 5906 66110
rect 16830 66162 16882 66174
rect 22094 66162 22146 66174
rect 17602 66110 17614 66162
rect 17666 66110 17678 66162
rect 21858 66110 21870 66162
rect 21922 66110 21934 66162
rect 16830 66098 16882 66110
rect 22094 66098 22146 66110
rect 22542 66162 22594 66174
rect 22542 66098 22594 66110
rect 6862 66050 6914 66062
rect 19406 66050 19458 66062
rect 18834 65998 18846 66050
rect 18898 65998 18910 66050
rect 6862 65986 6914 65998
rect 19406 65986 19458 65998
rect 19966 66050 20018 66062
rect 19966 65986 20018 65998
rect 20750 66050 20802 66062
rect 20750 65986 20802 65998
rect 21310 66050 21362 66062
rect 21310 65986 21362 65998
rect 1344 65882 28720 65916
rect 1344 65830 8018 65882
rect 8070 65830 8122 65882
rect 8174 65830 8226 65882
rect 8278 65830 14822 65882
rect 14874 65830 14926 65882
rect 14978 65830 15030 65882
rect 15082 65830 21626 65882
rect 21678 65830 21730 65882
rect 21782 65830 21834 65882
rect 21886 65830 28430 65882
rect 28482 65830 28534 65882
rect 28586 65830 28638 65882
rect 28690 65830 28720 65882
rect 1344 65796 28720 65830
rect 3390 65714 3442 65726
rect 2594 65662 2606 65714
rect 2658 65662 2670 65714
rect 3390 65650 3442 65662
rect 7534 65714 7586 65726
rect 7534 65650 7586 65662
rect 13582 65714 13634 65726
rect 13582 65650 13634 65662
rect 14702 65714 14754 65726
rect 14702 65650 14754 65662
rect 15934 65714 15986 65726
rect 15934 65650 15986 65662
rect 23326 65714 23378 65726
rect 23326 65650 23378 65662
rect 3054 65602 3106 65614
rect 2818 65550 2830 65602
rect 2882 65550 2894 65602
rect 3054 65538 3106 65550
rect 4398 65602 4450 65614
rect 4398 65538 4450 65550
rect 13470 65602 13522 65614
rect 13470 65538 13522 65550
rect 14478 65602 14530 65614
rect 14478 65538 14530 65550
rect 17950 65602 18002 65614
rect 17950 65538 18002 65550
rect 18062 65602 18114 65614
rect 18062 65538 18114 65550
rect 18734 65602 18786 65614
rect 18734 65538 18786 65550
rect 23102 65602 23154 65614
rect 23102 65538 23154 65550
rect 2606 65490 2658 65502
rect 2482 65438 2494 65490
rect 2546 65438 2558 65490
rect 2606 65426 2658 65438
rect 7310 65490 7362 65502
rect 7310 65426 7362 65438
rect 7422 65490 7474 65502
rect 7422 65426 7474 65438
rect 7982 65490 8034 65502
rect 13806 65490 13858 65502
rect 9650 65438 9662 65490
rect 9714 65438 9726 65490
rect 7982 65426 8034 65438
rect 13806 65426 13858 65438
rect 14030 65490 14082 65502
rect 14030 65426 14082 65438
rect 14590 65490 14642 65502
rect 14590 65426 14642 65438
rect 15150 65490 15202 65502
rect 15150 65426 15202 65438
rect 17278 65490 17330 65502
rect 17278 65426 17330 65438
rect 17502 65490 17554 65502
rect 17502 65426 17554 65438
rect 21422 65490 21474 65502
rect 23998 65490 24050 65502
rect 22866 65438 22878 65490
rect 22930 65438 22942 65490
rect 23538 65438 23550 65490
rect 23602 65438 23614 65490
rect 21422 65426 21474 65438
rect 23998 65426 24050 65438
rect 24446 65490 24498 65502
rect 24446 65426 24498 65438
rect 25342 65490 25394 65502
rect 25342 65426 25394 65438
rect 25790 65490 25842 65502
rect 25790 65426 25842 65438
rect 26126 65490 26178 65502
rect 26126 65426 26178 65438
rect 26350 65490 26402 65502
rect 26350 65426 26402 65438
rect 26910 65490 26962 65502
rect 26910 65426 26962 65438
rect 27806 65490 27858 65502
rect 27806 65426 27858 65438
rect 3502 65378 3554 65390
rect 3502 65314 3554 65326
rect 3950 65378 4002 65390
rect 3950 65314 4002 65326
rect 4846 65378 4898 65390
rect 4846 65314 4898 65326
rect 8318 65378 8370 65390
rect 8318 65314 8370 65326
rect 8766 65378 8818 65390
rect 13134 65378 13186 65390
rect 10322 65326 10334 65378
rect 10386 65326 10398 65378
rect 12450 65326 12462 65378
rect 12514 65326 12526 65378
rect 8766 65314 8818 65326
rect 13134 65314 13186 65326
rect 15486 65378 15538 65390
rect 15486 65314 15538 65326
rect 16382 65378 16434 65390
rect 16382 65314 16434 65326
rect 16942 65378 16994 65390
rect 16942 65314 16994 65326
rect 18286 65378 18338 65390
rect 18286 65314 18338 65326
rect 19406 65378 19458 65390
rect 19406 65314 19458 65326
rect 19966 65378 20018 65390
rect 19966 65314 20018 65326
rect 20974 65378 21026 65390
rect 20974 65314 21026 65326
rect 21870 65378 21922 65390
rect 21870 65314 21922 65326
rect 22318 65378 22370 65390
rect 22318 65314 22370 65326
rect 23214 65378 23266 65390
rect 23214 65314 23266 65326
rect 25902 65378 25954 65390
rect 25902 65314 25954 65326
rect 27358 65378 27410 65390
rect 27358 65314 27410 65326
rect 15474 65214 15486 65266
rect 15538 65263 15550 65266
rect 16146 65263 16158 65266
rect 15538 65217 16158 65263
rect 15538 65214 15550 65217
rect 16146 65214 16158 65217
rect 16210 65263 16222 65266
rect 16818 65263 16830 65266
rect 16210 65217 16830 65263
rect 16210 65214 16222 65217
rect 16818 65214 16830 65217
rect 16882 65214 16894 65266
rect 20962 65214 20974 65266
rect 21026 65263 21038 65266
rect 22082 65263 22094 65266
rect 21026 65217 22094 65263
rect 21026 65214 21038 65217
rect 22082 65214 22094 65217
rect 22146 65214 22158 65266
rect 1344 65098 28560 65132
rect 1344 65046 4616 65098
rect 4668 65046 4720 65098
rect 4772 65046 4824 65098
rect 4876 65046 11420 65098
rect 11472 65046 11524 65098
rect 11576 65046 11628 65098
rect 11680 65046 18224 65098
rect 18276 65046 18328 65098
rect 18380 65046 18432 65098
rect 18484 65046 25028 65098
rect 25080 65046 25132 65098
rect 25184 65046 25236 65098
rect 25288 65046 28560 65098
rect 1344 65012 28560 65046
rect 3714 64878 3726 64930
rect 3778 64927 3790 64930
rect 3938 64927 3950 64930
rect 3778 64881 3950 64927
rect 3778 64878 3790 64881
rect 3938 64878 3950 64881
rect 4002 64878 4014 64930
rect 12338 64878 12350 64930
rect 12402 64927 12414 64930
rect 13010 64927 13022 64930
rect 12402 64881 13022 64927
rect 12402 64878 12414 64881
rect 13010 64878 13022 64881
rect 13074 64878 13086 64930
rect 16930 64878 16942 64930
rect 16994 64927 17006 64930
rect 17154 64927 17166 64930
rect 16994 64881 17166 64927
rect 16994 64878 17006 64881
rect 17154 64878 17166 64881
rect 17218 64927 17230 64930
rect 17490 64927 17502 64930
rect 17218 64881 17502 64927
rect 17218 64878 17230 64881
rect 17490 64878 17502 64881
rect 17554 64878 17566 64930
rect 8990 64818 9042 64830
rect 8530 64766 8542 64818
rect 8594 64766 8606 64818
rect 8990 64754 9042 64766
rect 10334 64818 10386 64830
rect 24670 64818 24722 64830
rect 18834 64766 18846 64818
rect 18898 64766 18910 64818
rect 24210 64766 24222 64818
rect 24274 64766 24286 64818
rect 26002 64766 26014 64818
rect 26066 64766 26078 64818
rect 28130 64766 28142 64818
rect 28194 64766 28206 64818
rect 10334 64754 10386 64766
rect 24670 64754 24722 64766
rect 4174 64706 4226 64718
rect 10446 64706 10498 64718
rect 5730 64654 5742 64706
rect 5794 64654 5806 64706
rect 4174 64642 4226 64654
rect 10446 64642 10498 64654
rect 10782 64706 10834 64718
rect 10782 64642 10834 64654
rect 16942 64706 16994 64718
rect 16942 64642 16994 64654
rect 20414 64706 20466 64718
rect 20514 64654 20526 64706
rect 20578 64654 20590 64706
rect 21298 64654 21310 64706
rect 21362 64654 21374 64706
rect 25330 64654 25342 64706
rect 25394 64654 25406 64706
rect 20414 64642 20466 64654
rect 1710 64594 1762 64606
rect 1710 64530 1762 64542
rect 3054 64594 3106 64606
rect 3054 64530 3106 64542
rect 4622 64594 4674 64606
rect 10222 64594 10274 64606
rect 6402 64542 6414 64594
rect 6466 64542 6478 64594
rect 4622 64530 4674 64542
rect 10222 64530 10274 64542
rect 11230 64594 11282 64606
rect 11230 64530 11282 64542
rect 19182 64594 19234 64606
rect 19182 64530 19234 64542
rect 19966 64594 20018 64606
rect 20178 64542 20190 64594
rect 20242 64542 20254 64594
rect 22082 64542 22094 64594
rect 22146 64542 22158 64594
rect 19966 64530 20018 64542
rect 2046 64482 2098 64494
rect 2046 64418 2098 64430
rect 2830 64482 2882 64494
rect 2830 64418 2882 64430
rect 2942 64482 2994 64494
rect 2942 64418 2994 64430
rect 3726 64482 3778 64494
rect 3726 64418 3778 64430
rect 9886 64482 9938 64494
rect 9886 64418 9938 64430
rect 12686 64482 12738 64494
rect 12686 64418 12738 64430
rect 13582 64482 13634 64494
rect 13582 64418 13634 64430
rect 14254 64482 14306 64494
rect 14254 64418 14306 64430
rect 17390 64482 17442 64494
rect 17390 64418 17442 64430
rect 18958 64482 19010 64494
rect 18958 64418 19010 64430
rect 19630 64482 19682 64494
rect 19630 64418 19682 64430
rect 20750 64482 20802 64494
rect 20750 64418 20802 64430
rect 1344 64314 28720 64348
rect 1344 64262 8018 64314
rect 8070 64262 8122 64314
rect 8174 64262 8226 64314
rect 8278 64262 14822 64314
rect 14874 64262 14926 64314
rect 14978 64262 15030 64314
rect 15082 64262 21626 64314
rect 21678 64262 21730 64314
rect 21782 64262 21834 64314
rect 21886 64262 28430 64314
rect 28482 64262 28534 64314
rect 28586 64262 28638 64314
rect 28690 64262 28720 64314
rect 1344 64228 28720 64262
rect 2494 64146 2546 64158
rect 2494 64082 2546 64094
rect 6302 64146 6354 64158
rect 6302 64082 6354 64094
rect 7646 64146 7698 64158
rect 7646 64082 7698 64094
rect 13582 64146 13634 64158
rect 13582 64082 13634 64094
rect 20974 64146 21026 64158
rect 20974 64082 21026 64094
rect 21870 64146 21922 64158
rect 21870 64082 21922 64094
rect 24670 64146 24722 64158
rect 24670 64082 24722 64094
rect 25566 64146 25618 64158
rect 25566 64082 25618 64094
rect 25678 64146 25730 64158
rect 25678 64082 25730 64094
rect 27022 64146 27074 64158
rect 27022 64082 27074 64094
rect 3278 64034 3330 64046
rect 3278 63970 3330 63982
rect 22430 64034 22482 64046
rect 22430 63970 22482 63982
rect 26126 64034 26178 64046
rect 26126 63970 26178 63982
rect 26350 64034 26402 64046
rect 26350 63970 26402 63982
rect 27470 64034 27522 64046
rect 27470 63970 27522 63982
rect 28030 64034 28082 64046
rect 28030 63970 28082 63982
rect 1822 63922 1874 63934
rect 2830 63922 2882 63934
rect 4510 63922 4562 63934
rect 2706 63870 2718 63922
rect 2770 63870 2782 63922
rect 3042 63870 3054 63922
rect 3106 63870 3118 63922
rect 3938 63870 3950 63922
rect 4002 63870 4014 63922
rect 1822 63858 1874 63870
rect 2830 63858 2882 63870
rect 4510 63858 4562 63870
rect 5742 63922 5794 63934
rect 5742 63858 5794 63870
rect 6078 63922 6130 63934
rect 6078 63858 6130 63870
rect 6302 63922 6354 63934
rect 6302 63858 6354 63870
rect 6638 63922 6690 63934
rect 6638 63858 6690 63870
rect 7422 63922 7474 63934
rect 7422 63858 7474 63870
rect 8094 63922 8146 63934
rect 8094 63858 8146 63870
rect 8430 63922 8482 63934
rect 21758 63922 21810 63934
rect 10098 63870 10110 63922
rect 10162 63870 10174 63922
rect 13906 63870 13918 63922
rect 13970 63870 13982 63922
rect 20402 63870 20414 63922
rect 20466 63870 20478 63922
rect 8430 63858 8482 63870
rect 21758 63858 21810 63870
rect 23102 63922 23154 63934
rect 23102 63858 23154 63870
rect 23550 63922 23602 63934
rect 23550 63858 23602 63870
rect 23774 63922 23826 63934
rect 23774 63858 23826 63870
rect 24222 63922 24274 63934
rect 24222 63858 24274 63870
rect 25118 63922 25170 63934
rect 25118 63858 25170 63870
rect 25790 63922 25842 63934
rect 25790 63858 25842 63870
rect 26798 63922 26850 63934
rect 26798 63858 26850 63870
rect 27246 63922 27298 63934
rect 27246 63858 27298 63870
rect 7086 63810 7138 63822
rect 7086 63746 7138 63758
rect 7534 63810 7586 63822
rect 7534 63746 7586 63758
rect 8878 63810 8930 63822
rect 8878 63746 8930 63758
rect 9550 63810 9602 63822
rect 22878 63810 22930 63822
rect 10882 63758 10894 63810
rect 10946 63758 10958 63810
rect 13010 63758 13022 63810
rect 13074 63758 13086 63810
rect 14690 63758 14702 63810
rect 14754 63758 14766 63810
rect 16818 63758 16830 63810
rect 16882 63758 16894 63810
rect 17602 63758 17614 63810
rect 17666 63758 17678 63810
rect 19730 63758 19742 63810
rect 19794 63758 19806 63810
rect 9550 63746 9602 63758
rect 22878 63746 22930 63758
rect 23662 63810 23714 63822
rect 23662 63746 23714 63758
rect 26574 63810 26626 63822
rect 26574 63746 26626 63758
rect 27134 63810 27186 63822
rect 27134 63746 27186 63758
rect 9662 63698 9714 63710
rect 21646 63698 21698 63710
rect 21074 63646 21086 63698
rect 21138 63695 21150 63698
rect 21410 63695 21422 63698
rect 21138 63649 21422 63695
rect 21138 63646 21150 63649
rect 21410 63646 21422 63649
rect 21474 63646 21486 63698
rect 23986 63646 23998 63698
rect 24050 63695 24062 63698
rect 24658 63695 24670 63698
rect 24050 63649 24670 63695
rect 24050 63646 24062 63649
rect 24658 63646 24670 63649
rect 24722 63646 24734 63698
rect 9662 63634 9714 63646
rect 21646 63634 21698 63646
rect 1344 63530 28560 63564
rect 1344 63478 4616 63530
rect 4668 63478 4720 63530
rect 4772 63478 4824 63530
rect 4876 63478 11420 63530
rect 11472 63478 11524 63530
rect 11576 63478 11628 63530
rect 11680 63478 18224 63530
rect 18276 63478 18328 63530
rect 18380 63478 18432 63530
rect 18484 63478 25028 63530
rect 25080 63478 25132 63530
rect 25184 63478 25236 63530
rect 25288 63478 28560 63530
rect 1344 63444 28560 63478
rect 18846 63362 18898 63374
rect 17602 63310 17614 63362
rect 17666 63359 17678 63362
rect 18162 63359 18174 63362
rect 17666 63313 18174 63359
rect 17666 63310 17678 63313
rect 18162 63310 18174 63313
rect 18226 63310 18238 63362
rect 19282 63310 19294 63362
rect 19346 63359 19358 63362
rect 19730 63359 19742 63362
rect 19346 63313 19742 63359
rect 19346 63310 19358 63313
rect 19730 63310 19742 63313
rect 19794 63310 19806 63362
rect 18846 63298 18898 63310
rect 5070 63250 5122 63262
rect 11342 63250 11394 63262
rect 2482 63198 2494 63250
rect 2546 63198 2558 63250
rect 4610 63198 4622 63250
rect 4674 63198 4686 63250
rect 9650 63198 9662 63250
rect 9714 63198 9726 63250
rect 5070 63186 5122 63198
rect 11342 63186 11394 63198
rect 14478 63250 14530 63262
rect 14478 63186 14530 63198
rect 14926 63250 14978 63262
rect 14926 63186 14978 63198
rect 15374 63250 15426 63262
rect 15374 63186 15426 63198
rect 16270 63250 16322 63262
rect 16270 63186 16322 63198
rect 17726 63250 17778 63262
rect 27022 63250 27074 63262
rect 23986 63198 23998 63250
rect 24050 63198 24062 63250
rect 17726 63186 17778 63198
rect 27022 63186 27074 63198
rect 27470 63250 27522 63262
rect 27470 63186 27522 63198
rect 28142 63250 28194 63262
rect 28142 63186 28194 63198
rect 10222 63138 10274 63150
rect 11566 63138 11618 63150
rect 1698 63086 1710 63138
rect 1762 63086 1774 63138
rect 6738 63086 6750 63138
rect 6802 63086 6814 63138
rect 10546 63086 10558 63138
rect 10610 63086 10622 63138
rect 10222 63074 10274 63086
rect 11566 63074 11618 63086
rect 11790 63138 11842 63150
rect 11790 63074 11842 63086
rect 12462 63138 12514 63150
rect 12462 63074 12514 63086
rect 13470 63138 13522 63150
rect 13470 63074 13522 63086
rect 15262 63138 15314 63150
rect 15262 63074 15314 63086
rect 15486 63138 15538 63150
rect 15486 63074 15538 63086
rect 15822 63138 15874 63150
rect 15822 63074 15874 63086
rect 16158 63138 16210 63150
rect 16158 63074 16210 63086
rect 16382 63138 16434 63150
rect 16382 63074 16434 63086
rect 17166 63138 17218 63150
rect 19630 63138 19682 63150
rect 19170 63086 19182 63138
rect 19234 63086 19246 63138
rect 17166 63074 17218 63086
rect 19630 63074 19682 63086
rect 20078 63138 20130 63150
rect 21410 63086 21422 63138
rect 21474 63086 21486 63138
rect 20078 63074 20130 63086
rect 11230 63026 11282 63038
rect 7522 62974 7534 63026
rect 7586 62974 7598 63026
rect 11230 62962 11282 62974
rect 12350 63026 12402 63038
rect 12350 62962 12402 62974
rect 16606 63026 16658 63038
rect 16606 62962 16658 62974
rect 18398 63026 18450 63038
rect 18610 62974 18622 63026
rect 18674 62974 18686 63026
rect 18398 62962 18450 62974
rect 9998 62914 10050 62926
rect 9998 62850 10050 62862
rect 10110 62914 10162 62926
rect 10110 62850 10162 62862
rect 12238 62914 12290 62926
rect 12238 62850 12290 62862
rect 12686 62914 12738 62926
rect 12686 62850 12738 62862
rect 13582 62914 13634 62926
rect 13582 62850 13634 62862
rect 14030 62914 14082 62926
rect 14030 62850 14082 62862
rect 19182 62914 19234 62926
rect 19182 62850 19234 62862
rect 20526 62914 20578 62926
rect 20526 62850 20578 62862
rect 1344 62746 28720 62780
rect 1344 62694 8018 62746
rect 8070 62694 8122 62746
rect 8174 62694 8226 62746
rect 8278 62694 14822 62746
rect 14874 62694 14926 62746
rect 14978 62694 15030 62746
rect 15082 62694 21626 62746
rect 21678 62694 21730 62746
rect 21782 62694 21834 62746
rect 21886 62694 28430 62746
rect 28482 62694 28534 62746
rect 28586 62694 28638 62746
rect 28690 62694 28720 62746
rect 1344 62660 28720 62694
rect 3502 62578 3554 62590
rect 3502 62514 3554 62526
rect 7870 62578 7922 62590
rect 7870 62514 7922 62526
rect 8766 62578 8818 62590
rect 8766 62514 8818 62526
rect 9886 62578 9938 62590
rect 9886 62514 9938 62526
rect 10558 62578 10610 62590
rect 10558 62514 10610 62526
rect 11006 62578 11058 62590
rect 11006 62514 11058 62526
rect 11454 62578 11506 62590
rect 11454 62514 11506 62526
rect 12014 62578 12066 62590
rect 12014 62514 12066 62526
rect 12462 62578 12514 62590
rect 12462 62514 12514 62526
rect 13022 62578 13074 62590
rect 13022 62514 13074 62526
rect 13582 62578 13634 62590
rect 13582 62514 13634 62526
rect 19294 62578 19346 62590
rect 19294 62514 19346 62526
rect 19742 62578 19794 62590
rect 19742 62514 19794 62526
rect 20190 62578 20242 62590
rect 20190 62514 20242 62526
rect 20638 62578 20690 62590
rect 20638 62514 20690 62526
rect 24670 62578 24722 62590
rect 24670 62514 24722 62526
rect 3614 62466 3666 62478
rect 3614 62402 3666 62414
rect 8318 62466 8370 62478
rect 8318 62402 8370 62414
rect 14478 62466 14530 62478
rect 14478 62402 14530 62414
rect 16270 62466 16322 62478
rect 18622 62466 18674 62478
rect 17490 62414 17502 62466
rect 17554 62414 17566 62466
rect 27346 62414 27358 62466
rect 27410 62414 27422 62466
rect 16270 62402 16322 62414
rect 18622 62402 18674 62414
rect 7758 62354 7810 62366
rect 7758 62290 7810 62302
rect 8094 62354 8146 62366
rect 8094 62290 8146 62302
rect 14366 62354 14418 62366
rect 14366 62290 14418 62302
rect 14702 62354 14754 62366
rect 14702 62290 14754 62302
rect 15374 62354 15426 62366
rect 15374 62290 15426 62302
rect 16830 62354 16882 62366
rect 17602 62302 17614 62354
rect 17666 62302 17678 62354
rect 18274 62302 18286 62354
rect 18338 62302 18350 62354
rect 21298 62302 21310 62354
rect 21362 62302 21374 62354
rect 28018 62302 28030 62354
rect 28082 62302 28094 62354
rect 16830 62290 16882 62302
rect 2494 62242 2546 62254
rect 2494 62178 2546 62190
rect 6638 62242 6690 62254
rect 6638 62178 6690 62190
rect 7422 62242 7474 62254
rect 7422 62178 7474 62190
rect 15822 62242 15874 62254
rect 17490 62190 17502 62242
rect 17554 62190 17566 62242
rect 22082 62190 22094 62242
rect 22146 62190 22158 62242
rect 24210 62190 24222 62242
rect 24274 62190 24286 62242
rect 25218 62190 25230 62242
rect 25282 62190 25294 62242
rect 15822 62178 15874 62190
rect 15362 62078 15374 62130
rect 15426 62127 15438 62130
rect 16034 62127 16046 62130
rect 15426 62081 16046 62127
rect 15426 62078 15438 62081
rect 16034 62078 16046 62081
rect 16098 62078 16110 62130
rect 1344 61962 28560 61996
rect 1344 61910 4616 61962
rect 4668 61910 4720 61962
rect 4772 61910 4824 61962
rect 4876 61910 11420 61962
rect 11472 61910 11524 61962
rect 11576 61910 11628 61962
rect 11680 61910 18224 61962
rect 18276 61910 18328 61962
rect 18380 61910 18432 61962
rect 18484 61910 25028 61962
rect 25080 61910 25132 61962
rect 25184 61910 25236 61962
rect 25288 61910 28560 61962
rect 1344 61876 28560 61910
rect 14466 61742 14478 61794
rect 14530 61742 14542 61794
rect 2830 61682 2882 61694
rect 4622 61682 4674 61694
rect 3490 61630 3502 61682
rect 3554 61630 3566 61682
rect 2830 61618 2882 61630
rect 4622 61618 4674 61630
rect 5070 61682 5122 61694
rect 5070 61618 5122 61630
rect 7982 61682 8034 61694
rect 13582 61682 13634 61694
rect 21422 61682 21474 61694
rect 11778 61630 11790 61682
rect 11842 61630 11854 61682
rect 12674 61630 12686 61682
rect 12738 61630 12750 61682
rect 17826 61630 17838 61682
rect 17890 61630 17902 61682
rect 7982 61618 8034 61630
rect 13582 61618 13634 61630
rect 21422 61618 21474 61630
rect 22430 61682 22482 61694
rect 26898 61630 26910 61682
rect 26962 61630 26974 61682
rect 22430 61618 22482 61630
rect 5966 61570 6018 61582
rect 3266 61518 3278 61570
rect 3330 61518 3342 61570
rect 5966 61506 6018 61518
rect 6078 61570 6130 61582
rect 6862 61570 6914 61582
rect 12350 61570 12402 61582
rect 14926 61570 14978 61582
rect 22654 61570 22706 61582
rect 6178 61518 6190 61570
rect 6242 61518 6254 61570
rect 7074 61518 7086 61570
rect 7138 61518 7150 61570
rect 8978 61518 8990 61570
rect 9042 61518 9054 61570
rect 14130 61518 14142 61570
rect 14194 61518 14206 61570
rect 15250 61518 15262 61570
rect 15314 61518 15326 61570
rect 16034 61518 16046 61570
rect 16098 61518 16110 61570
rect 16818 61518 16830 61570
rect 16882 61518 16894 61570
rect 17266 61518 17278 61570
rect 17330 61518 17342 61570
rect 20738 61518 20750 61570
rect 20802 61518 20814 61570
rect 6078 61506 6130 61518
rect 6862 61506 6914 61518
rect 12350 61506 12402 61518
rect 14926 61506 14978 61518
rect 22654 61506 22706 61518
rect 22878 61570 22930 61582
rect 22878 61506 22930 61518
rect 23326 61570 23378 61582
rect 24222 61570 24274 61582
rect 23986 61518 23998 61570
rect 24050 61518 24062 61570
rect 24658 61518 24670 61570
rect 24722 61518 24734 61570
rect 25666 61518 25678 61570
rect 25730 61518 25742 61570
rect 23326 61506 23378 61518
rect 24222 61506 24274 61518
rect 1710 61458 1762 61470
rect 1710 61394 1762 61406
rect 2046 61458 2098 61470
rect 2046 61394 2098 61406
rect 5630 61458 5682 61470
rect 5630 61394 5682 61406
rect 6750 61458 6802 61470
rect 12126 61458 12178 61470
rect 9650 61406 9662 61458
rect 9714 61406 9726 61458
rect 6750 61394 6802 61406
rect 12126 61394 12178 61406
rect 13918 61458 13970 61470
rect 22318 61458 22370 61470
rect 16146 61406 16158 61458
rect 16210 61406 16222 61458
rect 19954 61406 19966 61458
rect 20018 61406 20030 61458
rect 13918 61394 13970 61406
rect 22318 61394 22370 61406
rect 4174 61346 4226 61358
rect 4174 61282 4226 61294
rect 5742 61346 5794 61358
rect 5742 61282 5794 61294
rect 7534 61346 7586 61358
rect 7534 61282 7586 61294
rect 12574 61346 12626 61358
rect 12574 61282 12626 61294
rect 12686 61346 12738 61358
rect 12686 61282 12738 61294
rect 17390 61346 17442 61358
rect 17390 61282 17442 61294
rect 21982 61346 22034 61358
rect 21982 61282 22034 61294
rect 24334 61346 24386 61358
rect 24334 61282 24386 61294
rect 24446 61346 24498 61358
rect 24446 61282 24498 61294
rect 25118 61346 25170 61358
rect 25118 61282 25170 61294
rect 1344 61178 28720 61212
rect 1344 61126 8018 61178
rect 8070 61126 8122 61178
rect 8174 61126 8226 61178
rect 8278 61126 14822 61178
rect 14874 61126 14926 61178
rect 14978 61126 15030 61178
rect 15082 61126 21626 61178
rect 21678 61126 21730 61178
rect 21782 61126 21834 61178
rect 21886 61126 28430 61178
rect 28482 61126 28534 61178
rect 28586 61126 28638 61178
rect 28690 61126 28720 61178
rect 1344 61092 28720 61126
rect 2046 61010 2098 61022
rect 10334 61010 10386 61022
rect 2594 60958 2606 61010
rect 2658 60958 2670 61010
rect 2046 60946 2098 60958
rect 10334 60946 10386 60958
rect 19966 61010 20018 61022
rect 19966 60946 20018 60958
rect 20414 61010 20466 61022
rect 20414 60946 20466 60958
rect 25454 61010 25506 61022
rect 25454 60946 25506 60958
rect 27582 61010 27634 61022
rect 27582 60946 27634 60958
rect 3054 60898 3106 60910
rect 19182 60898 19234 60910
rect 5058 60846 5070 60898
rect 5122 60846 5134 60898
rect 11442 60846 11454 60898
rect 11506 60846 11518 60898
rect 13794 60846 13806 60898
rect 13858 60846 13870 60898
rect 14914 60846 14926 60898
rect 14978 60846 14990 60898
rect 17602 60846 17614 60898
rect 17666 60846 17678 60898
rect 19394 60846 19406 60898
rect 19458 60846 19470 60898
rect 3054 60834 3106 60846
rect 19182 60834 19234 60846
rect 8318 60786 8370 60798
rect 2370 60734 2382 60786
rect 2434 60734 2446 60786
rect 2818 60734 2830 60786
rect 2882 60734 2894 60786
rect 3378 60734 3390 60786
rect 3442 60734 3454 60786
rect 4386 60734 4398 60786
rect 4450 60734 4462 60786
rect 7858 60734 7870 60786
rect 7922 60734 7934 60786
rect 8318 60722 8370 60734
rect 10110 60786 10162 60798
rect 10110 60722 10162 60734
rect 10334 60786 10386 60798
rect 10334 60722 10386 60734
rect 10670 60786 10722 60798
rect 16382 60786 16434 60798
rect 12450 60734 12462 60786
rect 12514 60734 12526 60786
rect 14130 60734 14142 60786
rect 14194 60734 14206 60786
rect 10670 60722 10722 60734
rect 16382 60722 16434 60734
rect 17390 60786 17442 60798
rect 26574 60786 26626 60798
rect 17938 60734 17950 60786
rect 18002 60734 18014 60786
rect 18610 60734 18622 60786
rect 18674 60734 18686 60786
rect 19730 60734 19742 60786
rect 19794 60734 19806 60786
rect 21858 60734 21870 60786
rect 21922 60734 21934 60786
rect 17390 60722 17442 60734
rect 26574 60722 26626 60734
rect 26798 60786 26850 60798
rect 26798 60722 26850 60734
rect 27246 60786 27298 60798
rect 27246 60722 27298 60734
rect 3726 60674 3778 60686
rect 7646 60674 7698 60686
rect 7186 60622 7198 60674
rect 7250 60622 7262 60674
rect 3726 60610 3778 60622
rect 7646 60610 7698 60622
rect 8990 60674 9042 60686
rect 8990 60610 9042 60622
rect 9774 60674 9826 60686
rect 24334 60674 24386 60686
rect 10882 60622 10894 60674
rect 10946 60671 10958 60674
rect 11106 60671 11118 60674
rect 10946 60625 11118 60671
rect 10946 60622 10958 60625
rect 11106 60622 11118 60625
rect 11170 60622 11182 60674
rect 12338 60622 12350 60674
rect 12402 60622 12414 60674
rect 13906 60622 13918 60674
rect 13970 60622 13982 60674
rect 22418 60622 22430 60674
rect 22482 60622 22494 60674
rect 9774 60610 9826 60622
rect 24334 60610 24386 60622
rect 26238 60674 26290 60686
rect 26238 60610 26290 60622
rect 26686 60674 26738 60686
rect 26686 60610 26738 60622
rect 2606 60562 2658 60574
rect 2606 60498 2658 60510
rect 3390 60562 3442 60574
rect 3390 60498 3442 60510
rect 7534 60562 7586 60574
rect 7534 60498 7586 60510
rect 17278 60562 17330 60574
rect 17278 60498 17330 60510
rect 19630 60562 19682 60574
rect 19630 60498 19682 60510
rect 20302 60562 20354 60574
rect 20302 60498 20354 60510
rect 20638 60562 20690 60574
rect 20638 60498 20690 60510
rect 1344 60394 28560 60428
rect 1344 60342 4616 60394
rect 4668 60342 4720 60394
rect 4772 60342 4824 60394
rect 4876 60342 11420 60394
rect 11472 60342 11524 60394
rect 11576 60342 11628 60394
rect 11680 60342 18224 60394
rect 18276 60342 18328 60394
rect 18380 60342 18432 60394
rect 18484 60342 25028 60394
rect 25080 60342 25132 60394
rect 25184 60342 25236 60394
rect 25288 60342 28560 60394
rect 1344 60308 28560 60342
rect 14366 60226 14418 60238
rect 20078 60226 20130 60238
rect 19506 60174 19518 60226
rect 19570 60174 19582 60226
rect 14366 60162 14418 60174
rect 20078 60162 20130 60174
rect 20414 60226 20466 60238
rect 20414 60162 20466 60174
rect 8990 60114 9042 60126
rect 2482 60062 2494 60114
rect 2546 60062 2558 60114
rect 4610 60062 4622 60114
rect 4674 60062 4686 60114
rect 8530 60062 8542 60114
rect 8594 60062 8606 60114
rect 8990 60050 9042 60062
rect 11342 60114 11394 60126
rect 11342 60050 11394 60062
rect 12910 60114 12962 60126
rect 21634 60062 21646 60114
rect 21698 60062 21710 60114
rect 28130 60062 28142 60114
rect 28194 60062 28206 60114
rect 12910 60050 12962 60062
rect 11454 60002 11506 60014
rect 1810 59950 1822 60002
rect 1874 59950 1886 60002
rect 5730 59950 5742 60002
rect 5794 59950 5806 60002
rect 11454 59938 11506 59950
rect 11902 60002 11954 60014
rect 11902 59938 11954 59950
rect 13470 60002 13522 60014
rect 13470 59938 13522 59950
rect 13806 60002 13858 60014
rect 14590 60002 14642 60014
rect 16942 60002 16994 60014
rect 14242 59950 14254 60002
rect 14306 59950 14318 60002
rect 16370 59950 16382 60002
rect 16434 59950 16446 60002
rect 13806 59938 13858 59950
rect 14590 59938 14642 59950
rect 16942 59938 16994 59950
rect 18958 60002 19010 60014
rect 19506 59950 19518 60002
rect 19570 59950 19582 60002
rect 20066 59950 20078 60002
rect 20130 59950 20142 60002
rect 24546 59950 24558 60002
rect 24610 59950 24622 60002
rect 25330 59950 25342 60002
rect 25394 59950 25406 60002
rect 18958 59938 19010 59950
rect 17390 59890 17442 59902
rect 6402 59838 6414 59890
rect 6466 59838 6478 59890
rect 14802 59838 14814 59890
rect 14866 59838 14878 59890
rect 19170 59838 19182 59890
rect 19234 59838 19246 59890
rect 23762 59838 23774 59890
rect 23826 59838 23838 59890
rect 26002 59838 26014 59890
rect 26066 59838 26078 59890
rect 17390 59826 17442 59838
rect 5070 59778 5122 59790
rect 5070 59714 5122 59726
rect 10446 59778 10498 59790
rect 10446 59714 10498 59726
rect 10894 59778 10946 59790
rect 10894 59714 10946 59726
rect 11230 59778 11282 59790
rect 11230 59714 11282 59726
rect 12462 59778 12514 59790
rect 12462 59714 12514 59726
rect 13582 59778 13634 59790
rect 13582 59714 13634 59726
rect 14030 59778 14082 59790
rect 19070 59778 19122 59790
rect 18498 59726 18510 59778
rect 18562 59726 18574 59778
rect 14030 59714 14082 59726
rect 19070 59714 19122 59726
rect 1344 59610 28720 59644
rect 1344 59558 8018 59610
rect 8070 59558 8122 59610
rect 8174 59558 8226 59610
rect 8278 59558 14822 59610
rect 14874 59558 14926 59610
rect 14978 59558 15030 59610
rect 15082 59558 21626 59610
rect 21678 59558 21730 59610
rect 21782 59558 21834 59610
rect 21886 59558 28430 59610
rect 28482 59558 28534 59610
rect 28586 59558 28638 59610
rect 28690 59558 28720 59610
rect 1344 59524 28720 59558
rect 3166 59442 3218 59454
rect 3166 59378 3218 59390
rect 5742 59442 5794 59454
rect 5742 59378 5794 59390
rect 6638 59442 6690 59454
rect 6638 59378 6690 59390
rect 9886 59442 9938 59454
rect 9886 59378 9938 59390
rect 13806 59442 13858 59454
rect 13806 59378 13858 59390
rect 22766 59442 22818 59454
rect 22766 59378 22818 59390
rect 23662 59442 23714 59454
rect 23662 59378 23714 59390
rect 26014 59442 26066 59454
rect 26014 59378 26066 59390
rect 28142 59442 28194 59454
rect 28142 59378 28194 59390
rect 2046 59330 2098 59342
rect 2046 59266 2098 59278
rect 3278 59330 3330 59342
rect 15822 59330 15874 59342
rect 22878 59330 22930 59342
rect 14466 59278 14478 59330
rect 14530 59278 14542 59330
rect 14802 59278 14814 59330
rect 14866 59278 14878 59330
rect 20290 59278 20302 59330
rect 20354 59278 20366 59330
rect 3278 59266 3330 59278
rect 15822 59266 15874 59278
rect 22878 59266 22930 59278
rect 25902 59330 25954 59342
rect 25902 59266 25954 59278
rect 26462 59330 26514 59342
rect 26462 59266 26514 59278
rect 26910 59330 26962 59342
rect 26910 59266 26962 59278
rect 27358 59330 27410 59342
rect 27358 59266 27410 59278
rect 1710 59218 1762 59230
rect 1710 59154 1762 59166
rect 6526 59218 6578 59230
rect 7758 59218 7810 59230
rect 6738 59166 6750 59218
rect 6802 59166 6814 59218
rect 7298 59166 7310 59218
rect 7362 59166 7374 59218
rect 6526 59154 6578 59166
rect 7758 59154 7810 59166
rect 9774 59218 9826 59230
rect 16830 59218 16882 59230
rect 22542 59218 22594 59230
rect 10434 59166 10446 59218
rect 10498 59166 10510 59218
rect 14130 59166 14142 59218
rect 14194 59166 14206 59218
rect 15474 59166 15486 59218
rect 15538 59166 15550 59218
rect 16594 59166 16606 59218
rect 16658 59166 16670 59218
rect 21074 59166 21086 59218
rect 21138 59166 21150 59218
rect 9774 59154 9826 59166
rect 16830 59154 16882 59166
rect 22542 59154 22594 59166
rect 22990 59218 23042 59230
rect 22990 59154 23042 59166
rect 23438 59218 23490 59230
rect 23438 59154 23490 59166
rect 23550 59218 23602 59230
rect 26238 59218 26290 59230
rect 23986 59166 23998 59218
rect 24050 59166 24062 59218
rect 23550 59154 23602 59166
rect 26238 59154 26290 59166
rect 2494 59106 2546 59118
rect 2494 59042 2546 59054
rect 3726 59106 3778 59118
rect 3726 59042 3778 59054
rect 6190 59106 6242 59118
rect 17502 59106 17554 59118
rect 21534 59106 21586 59118
rect 11218 59054 11230 59106
rect 11282 59054 11294 59106
rect 13346 59054 13358 59106
rect 13410 59054 13422 59106
rect 18162 59054 18174 59106
rect 18226 59054 18238 59106
rect 6190 59042 6242 59054
rect 17502 59042 17554 59054
rect 21534 59042 21586 59054
rect 21982 59106 22034 59118
rect 21982 59042 22034 59054
rect 24446 59106 24498 59118
rect 24446 59042 24498 59054
rect 25342 59106 25394 59118
rect 25342 59042 25394 59054
rect 9886 58994 9938 59006
rect 7074 58942 7086 58994
rect 7138 58942 7150 58994
rect 7410 58942 7422 58994
rect 7474 58991 7486 58994
rect 7634 58991 7646 58994
rect 7474 58945 7646 58991
rect 7474 58942 7486 58945
rect 7634 58942 7646 58945
rect 7698 58942 7710 58994
rect 15698 58942 15710 58994
rect 15762 58942 15774 58994
rect 17490 58942 17502 58994
rect 17554 58991 17566 58994
rect 17826 58991 17838 58994
rect 17554 58945 17838 58991
rect 17554 58942 17566 58945
rect 17826 58942 17838 58945
rect 17890 58942 17902 58994
rect 9886 58930 9938 58942
rect 1344 58826 28560 58860
rect 1344 58774 4616 58826
rect 4668 58774 4720 58826
rect 4772 58774 4824 58826
rect 4876 58774 11420 58826
rect 11472 58774 11524 58826
rect 11576 58774 11628 58826
rect 11680 58774 18224 58826
rect 18276 58774 18328 58826
rect 18380 58774 18432 58826
rect 18484 58774 25028 58826
rect 25080 58774 25132 58826
rect 25184 58774 25236 58826
rect 25288 58774 28560 58826
rect 1344 58740 28560 58774
rect 2942 58658 2994 58670
rect 2942 58594 2994 58606
rect 3726 58658 3778 58670
rect 11790 58658 11842 58670
rect 10098 58606 10110 58658
rect 10162 58655 10174 58658
rect 10322 58655 10334 58658
rect 10162 58609 10334 58655
rect 10162 58606 10174 58609
rect 10322 58606 10334 58609
rect 10386 58606 10398 58658
rect 14578 58606 14590 58658
rect 14642 58655 14654 58658
rect 14914 58655 14926 58658
rect 14642 58609 14926 58655
rect 14642 58606 14654 58609
rect 14914 58606 14926 58609
rect 14978 58606 14990 58658
rect 22530 58655 22542 58658
rect 22209 58609 22542 58655
rect 3726 58594 3778 58606
rect 11790 58594 11842 58606
rect 4622 58546 4674 58558
rect 10558 58546 10610 58558
rect 6066 58494 6078 58546
rect 6130 58494 6142 58546
rect 4622 58482 4674 58494
rect 10558 58482 10610 58494
rect 11454 58546 11506 58558
rect 11454 58482 11506 58494
rect 12686 58546 12738 58558
rect 12686 58482 12738 58494
rect 14926 58546 14978 58558
rect 14926 58482 14978 58494
rect 15598 58546 15650 58558
rect 15598 58482 15650 58494
rect 16158 58546 16210 58558
rect 20638 58546 20690 58558
rect 22209 58546 22255 58609
rect 22530 58606 22542 58609
rect 22594 58655 22606 58658
rect 23314 58655 23326 58658
rect 22594 58609 23326 58655
rect 22594 58606 22606 58609
rect 23314 58606 23326 58609
rect 23378 58606 23390 58658
rect 23326 58546 23378 58558
rect 19394 58494 19406 58546
rect 19458 58494 19470 58546
rect 22194 58494 22206 58546
rect 22258 58494 22270 58546
rect 16158 58482 16210 58494
rect 20638 58482 20690 58494
rect 23326 58482 23378 58494
rect 23774 58546 23826 58558
rect 28130 58494 28142 58546
rect 28194 58494 28206 58546
rect 23774 58482 23826 58494
rect 2818 58382 2830 58434
rect 2882 58382 2894 58434
rect 5618 58382 5630 58434
rect 5682 58382 5694 58434
rect 12002 58382 12014 58434
rect 12066 58382 12078 58434
rect 12898 58382 12910 58434
rect 12962 58382 12974 58434
rect 16370 58382 16382 58434
rect 16434 58382 16446 58434
rect 18386 58382 18398 58434
rect 18450 58382 18462 58434
rect 25330 58382 25342 58434
rect 25394 58382 25406 58434
rect 3390 58322 3442 58334
rect 3154 58270 3166 58322
rect 3218 58270 3230 58322
rect 3390 58258 3442 58270
rect 4062 58322 4114 58334
rect 4062 58258 4114 58270
rect 9214 58322 9266 58334
rect 9214 58258 9266 58270
rect 11342 58322 11394 58334
rect 12574 58322 12626 58334
rect 11554 58270 11566 58322
rect 11618 58270 11630 58322
rect 11342 58258 11394 58270
rect 12574 58258 12626 58270
rect 14030 58322 14082 58334
rect 19518 58322 19570 58334
rect 16482 58270 16494 58322
rect 16546 58270 16558 58322
rect 26002 58270 26014 58322
rect 26066 58270 26078 58322
rect 14030 58258 14082 58270
rect 19518 58258 19570 58270
rect 2270 58210 2322 58222
rect 2270 58146 2322 58158
rect 2606 58210 2658 58222
rect 2606 58146 2658 58158
rect 3838 58210 3890 58222
rect 3838 58146 3890 58158
rect 9662 58210 9714 58222
rect 9662 58146 9714 58158
rect 10110 58210 10162 58222
rect 10110 58146 10162 58158
rect 11006 58210 11058 58222
rect 11006 58146 11058 58158
rect 13582 58210 13634 58222
rect 13582 58146 13634 58158
rect 14478 58210 14530 58222
rect 14478 58146 14530 58158
rect 21422 58210 21474 58222
rect 21422 58146 21474 58158
rect 21870 58210 21922 58222
rect 21870 58146 21922 58158
rect 22318 58210 22370 58222
rect 22318 58146 22370 58158
rect 22766 58210 22818 58222
rect 22766 58146 22818 58158
rect 24446 58210 24498 58222
rect 24446 58146 24498 58158
rect 24894 58210 24946 58222
rect 24894 58146 24946 58158
rect 1344 58042 28720 58076
rect 1344 57990 8018 58042
rect 8070 57990 8122 58042
rect 8174 57990 8226 58042
rect 8278 57990 14822 58042
rect 14874 57990 14926 58042
rect 14978 57990 15030 58042
rect 15082 57990 21626 58042
rect 21678 57990 21730 58042
rect 21782 57990 21834 58042
rect 21886 57990 28430 58042
rect 28482 57990 28534 58042
rect 28586 57990 28638 58042
rect 28690 57990 28720 58042
rect 1344 57956 28720 57990
rect 5070 57874 5122 57886
rect 5070 57810 5122 57822
rect 5966 57874 6018 57886
rect 5966 57810 6018 57822
rect 7086 57874 7138 57886
rect 7086 57810 7138 57822
rect 7534 57874 7586 57886
rect 7534 57810 7586 57822
rect 8094 57874 8146 57886
rect 8094 57810 8146 57822
rect 8542 57874 8594 57886
rect 8542 57810 8594 57822
rect 8990 57874 9042 57886
rect 8990 57810 9042 57822
rect 9550 57874 9602 57886
rect 9550 57810 9602 57822
rect 13022 57874 13074 57886
rect 13022 57810 13074 57822
rect 13470 57874 13522 57886
rect 24222 57874 24274 57886
rect 17490 57822 17502 57874
rect 17554 57822 17566 57874
rect 13470 57810 13522 57822
rect 24222 57810 24274 57822
rect 26014 57874 26066 57886
rect 26014 57810 26066 57822
rect 27246 57874 27298 57886
rect 27246 57810 27298 57822
rect 27806 57874 27858 57886
rect 27806 57810 27858 57822
rect 6302 57762 6354 57774
rect 17950 57762 18002 57774
rect 2482 57710 2494 57762
rect 2546 57710 2558 57762
rect 15474 57710 15486 57762
rect 15538 57710 15550 57762
rect 6302 57698 6354 57710
rect 17950 57698 18002 57710
rect 19966 57762 20018 57774
rect 19966 57698 20018 57710
rect 21646 57762 21698 57774
rect 21646 57698 21698 57710
rect 22878 57762 22930 57774
rect 22878 57698 22930 57710
rect 23886 57762 23938 57774
rect 23886 57698 23938 57710
rect 25902 57762 25954 57774
rect 25902 57698 25954 57710
rect 26238 57762 26290 57774
rect 26238 57698 26290 57710
rect 9774 57650 9826 57662
rect 10670 57650 10722 57662
rect 1810 57598 1822 57650
rect 1874 57598 1886 57650
rect 6626 57598 6638 57650
rect 6690 57598 6702 57650
rect 10098 57598 10110 57650
rect 10162 57598 10174 57650
rect 9774 57586 9826 57598
rect 10670 57586 10722 57598
rect 11902 57650 11954 57662
rect 11902 57586 11954 57598
rect 12238 57650 12290 57662
rect 12238 57586 12290 57598
rect 12462 57650 12514 57662
rect 12462 57586 12514 57598
rect 15150 57650 15202 57662
rect 23214 57650 23266 57662
rect 15586 57598 15598 57650
rect 15650 57598 15662 57650
rect 17378 57598 17390 57650
rect 17442 57598 17454 57650
rect 21186 57598 21198 57650
rect 21250 57598 21262 57650
rect 15150 57586 15202 57598
rect 23214 57586 23266 57598
rect 23438 57650 23490 57662
rect 23438 57586 23490 57598
rect 23774 57650 23826 57662
rect 23774 57586 23826 57598
rect 23998 57650 24050 57662
rect 23998 57586 24050 57598
rect 26462 57650 26514 57662
rect 26462 57586 26514 57598
rect 26798 57650 26850 57662
rect 26798 57586 26850 57598
rect 26910 57650 26962 57662
rect 26910 57586 26962 57598
rect 27022 57650 27074 57662
rect 27022 57586 27074 57598
rect 6414 57538 6466 57550
rect 4610 57486 4622 57538
rect 4674 57486 4686 57538
rect 6414 57474 6466 57486
rect 9662 57538 9714 57550
rect 9662 57474 9714 57486
rect 11118 57538 11170 57550
rect 11118 57474 11170 57486
rect 11566 57538 11618 57550
rect 11566 57474 11618 57486
rect 12014 57538 12066 57550
rect 12014 57474 12066 57486
rect 13918 57538 13970 57550
rect 13918 57474 13970 57486
rect 14590 57538 14642 57550
rect 22542 57538 22594 57550
rect 16818 57486 16830 57538
rect 16882 57486 16894 57538
rect 14590 57474 14642 57486
rect 22542 57474 22594 57486
rect 22990 57538 23042 57550
rect 22990 57474 23042 57486
rect 25342 57538 25394 57550
rect 25342 57474 25394 57486
rect 6850 57374 6862 57426
rect 6914 57423 6926 57426
rect 7186 57423 7198 57426
rect 6914 57377 7198 57423
rect 6914 57374 6926 57377
rect 7186 57374 7198 57377
rect 7250 57423 7262 57426
rect 8082 57423 8094 57426
rect 7250 57377 8094 57423
rect 7250 57374 7262 57377
rect 8082 57374 8094 57377
rect 8146 57374 8158 57426
rect 10994 57374 11006 57426
rect 11058 57423 11070 57426
rect 11554 57423 11566 57426
rect 11058 57377 11566 57423
rect 11058 57374 11070 57377
rect 11554 57374 11566 57377
rect 11618 57374 11630 57426
rect 1344 57258 28560 57292
rect 1344 57206 4616 57258
rect 4668 57206 4720 57258
rect 4772 57206 4824 57258
rect 4876 57206 11420 57258
rect 11472 57206 11524 57258
rect 11576 57206 11628 57258
rect 11680 57206 18224 57258
rect 18276 57206 18328 57258
rect 18380 57206 18432 57258
rect 18484 57206 25028 57258
rect 25080 57206 25132 57258
rect 25184 57206 25236 57258
rect 25288 57206 28560 57258
rect 1344 57172 28560 57206
rect 3502 57090 3554 57102
rect 20190 57090 20242 57102
rect 6178 57038 6190 57090
rect 6242 57038 6254 57090
rect 3502 57026 3554 57038
rect 20190 57026 20242 57038
rect 5070 56978 5122 56990
rect 13582 56978 13634 56990
rect 9650 56926 9662 56978
rect 9714 56926 9726 56978
rect 10770 56926 10782 56978
rect 10834 56926 10846 56978
rect 12898 56926 12910 56978
rect 12962 56926 12974 56978
rect 5070 56914 5122 56926
rect 13582 56914 13634 56926
rect 14590 56978 14642 56990
rect 25566 56978 25618 56990
rect 22642 56926 22654 56978
rect 22706 56926 22718 56978
rect 24770 56926 24782 56978
rect 24834 56926 24846 56978
rect 14590 56914 14642 56926
rect 25566 56914 25618 56926
rect 27694 56978 27746 56990
rect 27694 56914 27746 56926
rect 28142 56978 28194 56990
rect 28142 56914 28194 56926
rect 5630 56866 5682 56878
rect 13470 56866 13522 56878
rect 6178 56814 6190 56866
rect 6242 56814 6254 56866
rect 6850 56814 6862 56866
rect 6914 56814 6926 56866
rect 10098 56814 10110 56866
rect 10162 56814 10174 56866
rect 5630 56802 5682 56814
rect 13470 56802 13522 56814
rect 14142 56866 14194 56878
rect 14142 56802 14194 56814
rect 16606 56866 16658 56878
rect 16606 56802 16658 56814
rect 17054 56866 17106 56878
rect 21970 56814 21982 56866
rect 22034 56814 22046 56866
rect 17054 56802 17106 56814
rect 3614 56754 3666 56766
rect 3614 56690 3666 56702
rect 4062 56754 4114 56766
rect 15598 56754 15650 56766
rect 5842 56702 5854 56754
rect 5906 56702 5918 56754
rect 7522 56702 7534 56754
rect 7586 56702 7598 56754
rect 4062 56690 4114 56702
rect 15598 56690 15650 56702
rect 18174 56754 18226 56766
rect 18174 56690 18226 56702
rect 19518 56754 19570 56766
rect 19518 56690 19570 56702
rect 21422 56754 21474 56766
rect 21422 56690 21474 56702
rect 26910 56754 26962 56766
rect 26910 56690 26962 56702
rect 5742 56642 5794 56654
rect 5742 56578 5794 56590
rect 13694 56642 13746 56654
rect 18958 56642 19010 56654
rect 15026 56590 15038 56642
rect 15090 56590 15102 56642
rect 13694 56578 13746 56590
rect 18958 56578 19010 56590
rect 19070 56642 19122 56654
rect 19070 56578 19122 56590
rect 19294 56642 19346 56654
rect 19294 56578 19346 56590
rect 19966 56642 20018 56654
rect 19966 56578 20018 56590
rect 20078 56642 20130 56654
rect 20078 56578 20130 56590
rect 20638 56642 20690 56654
rect 20638 56578 20690 56590
rect 26014 56642 26066 56654
rect 26014 56578 26066 56590
rect 26462 56642 26514 56654
rect 26462 56578 26514 56590
rect 1344 56474 28720 56508
rect 1344 56422 8018 56474
rect 8070 56422 8122 56474
rect 8174 56422 8226 56474
rect 8278 56422 14822 56474
rect 14874 56422 14926 56474
rect 14978 56422 15030 56474
rect 15082 56422 21626 56474
rect 21678 56422 21730 56474
rect 21782 56422 21834 56474
rect 21886 56422 28430 56474
rect 28482 56422 28534 56474
rect 28586 56422 28638 56474
rect 28690 56422 28720 56474
rect 1344 56388 28720 56422
rect 8430 56306 8482 56318
rect 8430 56242 8482 56254
rect 11790 56306 11842 56318
rect 11790 56242 11842 56254
rect 11902 56306 11954 56318
rect 11902 56242 11954 56254
rect 13134 56306 13186 56318
rect 23438 56306 23490 56318
rect 17826 56254 17838 56306
rect 17890 56254 17902 56306
rect 13134 56242 13186 56254
rect 23438 56242 23490 56254
rect 2046 56194 2098 56206
rect 2046 56130 2098 56142
rect 3614 56194 3666 56206
rect 3614 56130 3666 56142
rect 3838 56194 3890 56206
rect 8654 56194 8706 56206
rect 5282 56142 5294 56194
rect 5346 56142 5358 56194
rect 3838 56130 3890 56142
rect 8654 56130 8706 56142
rect 8878 56194 8930 56206
rect 8878 56130 8930 56142
rect 10222 56194 10274 56206
rect 10222 56130 10274 56142
rect 11230 56194 11282 56206
rect 11230 56130 11282 56142
rect 12238 56194 12290 56206
rect 15598 56194 15650 56206
rect 13570 56142 13582 56194
rect 13634 56142 13646 56194
rect 15026 56142 15038 56194
rect 15090 56142 15102 56194
rect 12238 56130 12290 56142
rect 15598 56130 15650 56142
rect 23886 56194 23938 56206
rect 23886 56130 23938 56142
rect 1710 56082 1762 56094
rect 8318 56082 8370 56094
rect 9998 56082 10050 56094
rect 11678 56082 11730 56094
rect 4162 56030 4174 56082
rect 4226 56030 4238 56082
rect 4610 56030 4622 56082
rect 4674 56030 4686 56082
rect 9762 56030 9774 56082
rect 9826 56030 9838 56082
rect 10434 56030 10446 56082
rect 10498 56030 10510 56082
rect 10882 56030 10894 56082
rect 10946 56030 10958 56082
rect 1710 56018 1762 56030
rect 8318 56018 8370 56030
rect 9998 56018 10050 56030
rect 11678 56018 11730 56030
rect 12014 56082 12066 56094
rect 12798 56082 12850 56094
rect 12562 56030 12574 56082
rect 12626 56030 12638 56082
rect 12014 56018 12066 56030
rect 12798 56018 12850 56030
rect 12910 56082 12962 56094
rect 12910 56018 12962 56030
rect 13022 56082 13074 56094
rect 23326 56082 23378 56094
rect 13682 56030 13694 56082
rect 13746 56030 13758 56082
rect 14466 56030 14478 56082
rect 14530 56030 14542 56082
rect 14802 56030 14814 56082
rect 14866 56030 14878 56082
rect 15474 56030 15486 56082
rect 15538 56030 15550 56082
rect 16146 56030 16158 56082
rect 16210 56030 16222 56082
rect 16594 56030 16606 56082
rect 16658 56030 16670 56082
rect 17938 56030 17950 56082
rect 18002 56030 18014 56082
rect 18274 56030 18286 56082
rect 18338 56030 18350 56082
rect 19506 56030 19518 56082
rect 19570 56030 19582 56082
rect 13022 56018 13074 56030
rect 23326 56018 23378 56030
rect 23662 56082 23714 56094
rect 25330 56030 25342 56082
rect 25394 56030 25406 56082
rect 23662 56018 23714 56030
rect 2494 55970 2546 55982
rect 2494 55906 2546 55918
rect 3950 55970 4002 55982
rect 8094 55970 8146 55982
rect 16942 55970 16994 55982
rect 19070 55970 19122 55982
rect 22766 55970 22818 55982
rect 24334 55970 24386 55982
rect 7410 55918 7422 55970
rect 7474 55918 7486 55970
rect 10322 55918 10334 55970
rect 10386 55918 10398 55970
rect 17602 55918 17614 55970
rect 17666 55918 17678 55970
rect 20178 55918 20190 55970
rect 20242 55918 20254 55970
rect 22306 55918 22318 55970
rect 22370 55918 22382 55970
rect 23426 55918 23438 55970
rect 23490 55918 23502 55970
rect 26002 55918 26014 55970
rect 26066 55918 26078 55970
rect 28130 55918 28142 55970
rect 28194 55918 28206 55970
rect 3950 55906 4002 55918
rect 8094 55906 8146 55918
rect 16942 55906 16994 55918
rect 19070 55906 19122 55918
rect 22766 55906 22818 55918
rect 24334 55906 24386 55918
rect 10894 55858 10946 55870
rect 10894 55794 10946 55806
rect 1344 55690 28560 55724
rect 1344 55638 4616 55690
rect 4668 55638 4720 55690
rect 4772 55638 4824 55690
rect 4876 55638 11420 55690
rect 11472 55638 11524 55690
rect 11576 55638 11628 55690
rect 11680 55638 18224 55690
rect 18276 55638 18328 55690
rect 18380 55638 18432 55690
rect 18484 55638 25028 55690
rect 25080 55638 25132 55690
rect 25184 55638 25236 55690
rect 25288 55638 28560 55690
rect 1344 55604 28560 55638
rect 20302 55522 20354 55534
rect 10210 55470 10222 55522
rect 10274 55519 10286 55522
rect 11666 55519 11678 55522
rect 10274 55473 11678 55519
rect 10274 55470 10286 55473
rect 11666 55470 11678 55473
rect 11730 55470 11742 55522
rect 12450 55470 12462 55522
rect 12514 55519 12526 55522
rect 13010 55519 13022 55522
rect 12514 55473 13022 55519
rect 12514 55470 12526 55473
rect 13010 55470 13022 55473
rect 13074 55470 13086 55522
rect 13570 55470 13582 55522
rect 13634 55519 13646 55522
rect 13634 55473 14191 55519
rect 13634 55470 13646 55473
rect 6638 55410 6690 55422
rect 4610 55358 4622 55410
rect 4674 55358 4686 55410
rect 6638 55346 6690 55358
rect 7198 55410 7250 55422
rect 7198 55346 7250 55358
rect 7982 55410 8034 55422
rect 7982 55346 8034 55358
rect 8878 55410 8930 55422
rect 8878 55346 8930 55358
rect 9438 55410 9490 55422
rect 9438 55346 9490 55358
rect 12574 55410 12626 55422
rect 14145 55407 14191 55473
rect 20302 55458 20354 55470
rect 21422 55410 21474 55422
rect 14242 55407 14254 55410
rect 14145 55361 14254 55407
rect 14242 55358 14254 55361
rect 14306 55358 14318 55410
rect 12574 55346 12626 55358
rect 21422 55346 21474 55358
rect 23214 55410 23266 55422
rect 23214 55346 23266 55358
rect 21310 55298 21362 55310
rect 1810 55246 1822 55298
rect 1874 55246 1886 55298
rect 14354 55246 14366 55298
rect 14418 55246 14430 55298
rect 20066 55246 20078 55298
rect 20130 55246 20142 55298
rect 21310 55234 21362 55246
rect 21870 55298 21922 55310
rect 21870 55234 21922 55246
rect 22318 55298 22370 55310
rect 22318 55234 22370 55246
rect 22878 55298 22930 55310
rect 22878 55234 22930 55246
rect 25118 55298 25170 55310
rect 25118 55234 25170 55246
rect 25566 55298 25618 55310
rect 25566 55234 25618 55246
rect 26350 55298 26402 55310
rect 27358 55298 27410 55310
rect 26786 55246 26798 55298
rect 26850 55246 26862 55298
rect 27682 55246 27694 55298
rect 27746 55246 27758 55298
rect 26350 55234 26402 55246
rect 27358 55234 27410 55246
rect 11230 55186 11282 55198
rect 2482 55134 2494 55186
rect 2546 55134 2558 55186
rect 11230 55122 11282 55134
rect 11566 55186 11618 55198
rect 11566 55122 11618 55134
rect 12014 55186 12066 55198
rect 20750 55186 20802 55198
rect 17154 55134 17166 55186
rect 17218 55134 17230 55186
rect 20514 55134 20526 55186
rect 20578 55134 20590 55186
rect 12014 55122 12066 55134
rect 20750 55122 20802 55134
rect 21646 55186 21698 55198
rect 21646 55122 21698 55134
rect 25790 55186 25842 55198
rect 25790 55122 25842 55134
rect 27246 55186 27298 55198
rect 27246 55122 27298 55134
rect 5070 55074 5122 55086
rect 5070 55010 5122 55022
rect 6078 55074 6130 55086
rect 6078 55010 6130 55022
rect 7646 55074 7698 55086
rect 7646 55010 7698 55022
rect 8430 55074 8482 55086
rect 8430 55010 8482 55022
rect 9886 55074 9938 55086
rect 9886 55010 9938 55022
rect 10222 55074 10274 55086
rect 10222 55010 10274 55022
rect 10670 55074 10722 55086
rect 10670 55010 10722 55022
rect 12910 55074 12962 55086
rect 12910 55010 12962 55022
rect 13582 55074 13634 55086
rect 13582 55010 13634 55022
rect 14030 55074 14082 55086
rect 14030 55010 14082 55022
rect 19966 55074 20018 55086
rect 19966 55010 20018 55022
rect 22206 55074 22258 55086
rect 22206 55010 22258 55022
rect 22430 55074 22482 55086
rect 22430 55010 22482 55022
rect 23662 55074 23714 55086
rect 23662 55010 23714 55022
rect 24110 55074 24162 55086
rect 24110 55010 24162 55022
rect 24558 55074 24610 55086
rect 24558 55010 24610 55022
rect 25454 55074 25506 55086
rect 25454 55010 25506 55022
rect 26238 55074 26290 55086
rect 26238 55010 26290 55022
rect 26462 55074 26514 55086
rect 26462 55010 26514 55022
rect 26574 55074 26626 55086
rect 26574 55010 26626 55022
rect 27134 55074 27186 55086
rect 27134 55010 27186 55022
rect 28142 55074 28194 55086
rect 28142 55010 28194 55022
rect 1344 54906 28720 54940
rect 1344 54854 8018 54906
rect 8070 54854 8122 54906
rect 8174 54854 8226 54906
rect 8278 54854 14822 54906
rect 14874 54854 14926 54906
rect 14978 54854 15030 54906
rect 15082 54854 21626 54906
rect 21678 54854 21730 54906
rect 21782 54854 21834 54906
rect 21886 54854 28430 54906
rect 28482 54854 28534 54906
rect 28586 54854 28638 54906
rect 28690 54854 28720 54906
rect 1344 54820 28720 54854
rect 2942 54738 2994 54750
rect 2942 54674 2994 54686
rect 5294 54738 5346 54750
rect 5294 54674 5346 54686
rect 5742 54738 5794 54750
rect 5742 54674 5794 54686
rect 15374 54738 15426 54750
rect 15374 54674 15426 54686
rect 22878 54738 22930 54750
rect 22878 54674 22930 54686
rect 24222 54738 24274 54750
rect 24222 54674 24274 54686
rect 24670 54738 24722 54750
rect 24670 54674 24722 54686
rect 25790 54738 25842 54750
rect 25790 54674 25842 54686
rect 2606 54626 2658 54638
rect 2606 54562 2658 54574
rect 2830 54626 2882 54638
rect 4398 54626 4450 54638
rect 3042 54574 3054 54626
rect 3106 54574 3118 54626
rect 2830 54562 2882 54574
rect 4398 54562 4450 54574
rect 12798 54626 12850 54638
rect 12798 54562 12850 54574
rect 15822 54626 15874 54638
rect 19506 54574 19518 54626
rect 19570 54574 19582 54626
rect 15822 54562 15874 54574
rect 2158 54514 2210 54526
rect 13134 54514 13186 54526
rect 20974 54514 21026 54526
rect 3378 54462 3390 54514
rect 3442 54462 3454 54514
rect 7298 54462 7310 54514
rect 7362 54462 7374 54514
rect 9650 54462 9662 54514
rect 9714 54462 9726 54514
rect 10322 54462 10334 54514
rect 10386 54462 10398 54514
rect 15250 54462 15262 54514
rect 15314 54462 15326 54514
rect 20178 54462 20190 54514
rect 20242 54462 20254 54514
rect 2158 54450 2210 54462
rect 13134 54450 13186 54462
rect 20974 54450 21026 54462
rect 21198 54514 21250 54526
rect 21198 54450 21250 54462
rect 4958 54402 5010 54414
rect 4958 54338 5010 54350
rect 6190 54402 6242 54414
rect 6190 54338 6242 54350
rect 6638 54402 6690 54414
rect 6638 54338 6690 54350
rect 6974 54402 7026 54414
rect 6974 54338 7026 54350
rect 7086 54402 7138 54414
rect 7086 54338 7138 54350
rect 8206 54402 8258 54414
rect 8206 54338 8258 54350
rect 8542 54402 8594 54414
rect 8542 54338 8594 54350
rect 9102 54402 9154 54414
rect 15038 54402 15090 54414
rect 21982 54402 22034 54414
rect 12450 54350 12462 54402
rect 12514 54350 12526 54402
rect 13234 54350 13246 54402
rect 13298 54350 13310 54402
rect 17378 54350 17390 54402
rect 17442 54350 17454 54402
rect 9102 54338 9154 54350
rect 15038 54338 15090 54350
rect 21982 54338 22034 54350
rect 22430 54402 22482 54414
rect 22430 54338 22482 54350
rect 23326 54402 23378 54414
rect 23326 54338 23378 54350
rect 23774 54402 23826 54414
rect 23774 54338 23826 54350
rect 25342 54402 25394 54414
rect 25342 54338 25394 54350
rect 26238 54402 26290 54414
rect 26238 54338 26290 54350
rect 26686 54402 26738 54414
rect 26686 54338 26738 54350
rect 27134 54402 27186 54414
rect 27134 54338 27186 54350
rect 27582 54402 27634 54414
rect 27582 54338 27634 54350
rect 28030 54402 28082 54414
rect 28030 54338 28082 54350
rect 3278 54290 3330 54302
rect 5058 54238 5070 54290
rect 5122 54287 5134 54290
rect 5618 54287 5630 54290
rect 5122 54241 5630 54287
rect 5122 54238 5134 54241
rect 5618 54238 5630 54241
rect 5682 54238 5694 54290
rect 21522 54238 21534 54290
rect 21586 54238 21598 54290
rect 22754 54238 22766 54290
rect 22818 54287 22830 54290
rect 24546 54287 24558 54290
rect 22818 54241 24558 54287
rect 22818 54238 22830 54241
rect 24546 54238 24558 54241
rect 24610 54238 24622 54290
rect 25106 54238 25118 54290
rect 25170 54287 25182 54290
rect 25442 54287 25454 54290
rect 25170 54241 25454 54287
rect 25170 54238 25182 54241
rect 25442 54238 25454 54241
rect 25506 54287 25518 54290
rect 25778 54287 25790 54290
rect 25506 54241 25790 54287
rect 25506 54238 25518 54241
rect 25778 54238 25790 54241
rect 25842 54287 25854 54290
rect 26674 54287 26686 54290
rect 25842 54241 26686 54287
rect 25842 54238 25854 54241
rect 26674 54238 26686 54241
rect 26738 54287 26750 54290
rect 28130 54287 28142 54290
rect 26738 54241 28142 54287
rect 26738 54238 26750 54241
rect 28130 54238 28142 54241
rect 28194 54238 28206 54290
rect 3278 54226 3330 54238
rect 1344 54122 28560 54156
rect 1344 54070 4616 54122
rect 4668 54070 4720 54122
rect 4772 54070 4824 54122
rect 4876 54070 11420 54122
rect 11472 54070 11524 54122
rect 11576 54070 11628 54122
rect 11680 54070 18224 54122
rect 18276 54070 18328 54122
rect 18380 54070 18432 54122
rect 18484 54070 25028 54122
rect 25080 54070 25132 54122
rect 25184 54070 25236 54122
rect 25288 54070 28560 54122
rect 1344 54036 28560 54070
rect 18722 53902 18734 53954
rect 18786 53951 18798 53954
rect 19058 53951 19070 53954
rect 18786 53905 19070 53951
rect 18786 53902 18798 53905
rect 19058 53902 19070 53905
rect 19122 53902 19134 53954
rect 3390 53842 3442 53854
rect 10222 53842 10274 53854
rect 4722 53790 4734 53842
rect 4786 53790 4798 53842
rect 8530 53790 8542 53842
rect 8594 53790 8606 53842
rect 3390 53778 3442 53790
rect 10222 53778 10274 53790
rect 10670 53842 10722 53854
rect 10670 53778 10722 53790
rect 11790 53842 11842 53854
rect 11790 53778 11842 53790
rect 12910 53842 12962 53854
rect 12910 53778 12962 53790
rect 13918 53842 13970 53854
rect 13918 53778 13970 53790
rect 16494 53842 16546 53854
rect 24110 53842 24162 53854
rect 21634 53790 21646 53842
rect 21698 53790 21710 53842
rect 16494 53778 16546 53790
rect 24110 53778 24162 53790
rect 2494 53730 2546 53742
rect 2494 53666 2546 53678
rect 3838 53730 3890 53742
rect 3838 53666 3890 53678
rect 4398 53730 4450 53742
rect 4398 53666 4450 53678
rect 4622 53730 4674 53742
rect 8766 53730 8818 53742
rect 5618 53678 5630 53730
rect 5682 53678 5694 53730
rect 4622 53666 4674 53678
rect 8766 53666 8818 53678
rect 9102 53730 9154 53742
rect 9102 53666 9154 53678
rect 10782 53730 10834 53742
rect 10782 53666 10834 53678
rect 11118 53730 11170 53742
rect 11118 53666 11170 53678
rect 11902 53730 11954 53742
rect 18398 53730 18450 53742
rect 12562 53678 12574 53730
rect 12626 53678 12638 53730
rect 16258 53678 16270 53730
rect 16322 53678 16334 53730
rect 11902 53666 11954 53678
rect 18398 53666 18450 53678
rect 19630 53730 19682 53742
rect 20302 53730 20354 53742
rect 20066 53678 20078 53730
rect 20130 53678 20142 53730
rect 19630 53666 19682 53678
rect 20302 53666 20354 53678
rect 20638 53730 20690 53742
rect 21758 53730 21810 53742
rect 21522 53678 21534 53730
rect 21586 53678 21598 53730
rect 20638 53666 20690 53678
rect 21758 53666 21810 53678
rect 23102 53730 23154 53742
rect 23102 53666 23154 53678
rect 23326 53730 23378 53742
rect 23326 53666 23378 53678
rect 25790 53730 25842 53742
rect 25790 53666 25842 53678
rect 26350 53730 26402 53742
rect 26350 53666 26402 53678
rect 26798 53730 26850 53742
rect 27234 53678 27246 53730
rect 27298 53678 27310 53730
rect 26798 53666 26850 53678
rect 1710 53618 1762 53630
rect 4174 53618 4226 53630
rect 9438 53618 9490 53630
rect 2818 53566 2830 53618
rect 2882 53566 2894 53618
rect 6402 53566 6414 53618
rect 6466 53566 6478 53618
rect 1710 53554 1762 53566
rect 4174 53554 4226 53566
rect 9438 53554 9490 53566
rect 10558 53618 10610 53630
rect 10558 53554 10610 53566
rect 15262 53618 15314 53630
rect 22206 53618 22258 53630
rect 18498 53566 18510 53618
rect 18562 53566 18574 53618
rect 20514 53566 20526 53618
rect 20578 53566 20590 53618
rect 15262 53554 15314 53566
rect 22206 53554 22258 53566
rect 22766 53618 22818 53630
rect 22766 53554 22818 53566
rect 23774 53618 23826 53630
rect 23774 53554 23826 53566
rect 23998 53618 24050 53630
rect 23998 53554 24050 53566
rect 26126 53618 26178 53630
rect 26126 53554 26178 53566
rect 26686 53618 26738 53630
rect 26686 53554 26738 53566
rect 27694 53618 27746 53630
rect 27694 53554 27746 53566
rect 2046 53506 2098 53518
rect 2046 53442 2098 53454
rect 4734 53506 4786 53518
rect 4734 53442 4786 53454
rect 8990 53506 9042 53518
rect 8990 53442 9042 53454
rect 11678 53506 11730 53518
rect 11678 53442 11730 53454
rect 12126 53506 12178 53518
rect 12126 53442 12178 53454
rect 12798 53506 12850 53518
rect 12798 53442 12850 53454
rect 14366 53506 14418 53518
rect 14366 53442 14418 53454
rect 18958 53506 19010 53518
rect 18958 53442 19010 53454
rect 19406 53506 19458 53518
rect 19406 53442 19458 53454
rect 21982 53506 22034 53518
rect 21982 53442 22034 53454
rect 22990 53506 23042 53518
rect 22990 53442 23042 53454
rect 24222 53506 24274 53518
rect 24222 53442 24274 53454
rect 24670 53506 24722 53518
rect 24670 53442 24722 53454
rect 25118 53506 25170 53518
rect 25118 53442 25170 53454
rect 26014 53506 26066 53518
rect 26014 53442 26066 53454
rect 26910 53506 26962 53518
rect 26910 53442 26962 53454
rect 28142 53506 28194 53518
rect 28142 53442 28194 53454
rect 1344 53338 28720 53372
rect 1344 53286 8018 53338
rect 8070 53286 8122 53338
rect 8174 53286 8226 53338
rect 8278 53286 14822 53338
rect 14874 53286 14926 53338
rect 14978 53286 15030 53338
rect 15082 53286 21626 53338
rect 21678 53286 21730 53338
rect 21782 53286 21834 53338
rect 21886 53286 28430 53338
rect 28482 53286 28534 53338
rect 28586 53286 28638 53338
rect 28690 53286 28720 53338
rect 1344 53252 28720 53286
rect 2494 53170 2546 53182
rect 2494 53106 2546 53118
rect 3278 53170 3330 53182
rect 3278 53106 3330 53118
rect 3838 53170 3890 53182
rect 3838 53106 3890 53118
rect 4286 53170 4338 53182
rect 4286 53106 4338 53118
rect 4510 53170 4562 53182
rect 4510 53106 4562 53118
rect 4622 53170 4674 53182
rect 4622 53106 4674 53118
rect 5294 53170 5346 53182
rect 5294 53106 5346 53118
rect 5518 53170 5570 53182
rect 5518 53106 5570 53118
rect 5630 53170 5682 53182
rect 8654 53170 8706 53182
rect 6402 53118 6414 53170
rect 6466 53118 6478 53170
rect 5630 53106 5682 53118
rect 8654 53106 8706 53118
rect 9102 53170 9154 53182
rect 9102 53106 9154 53118
rect 9774 53170 9826 53182
rect 9774 53106 9826 53118
rect 11230 53170 11282 53182
rect 11230 53106 11282 53118
rect 19742 53170 19794 53182
rect 19742 53106 19794 53118
rect 21310 53170 21362 53182
rect 21310 53106 21362 53118
rect 6078 53058 6130 53070
rect 9662 53058 9714 53070
rect 13694 53058 13746 53070
rect 6290 53006 6302 53058
rect 6354 53006 6366 53058
rect 11890 53006 11902 53058
rect 11954 53006 11966 53058
rect 12114 53006 12126 53058
rect 12178 53006 12190 53058
rect 6078 52994 6130 53006
rect 9662 52994 9714 53006
rect 13694 52994 13746 53006
rect 15710 53058 15762 53070
rect 15710 52994 15762 53006
rect 17950 53058 18002 53070
rect 17950 52994 18002 53006
rect 20526 53058 20578 53070
rect 20526 52994 20578 53006
rect 20638 53058 20690 53070
rect 23874 53006 23886 53058
rect 23938 53006 23950 53058
rect 26002 53006 26014 53058
rect 26066 53006 26078 53058
rect 20638 52994 20690 53006
rect 9886 52946 9938 52958
rect 12574 52946 12626 52958
rect 15150 52946 15202 52958
rect 20302 52946 20354 52958
rect 4050 52894 4062 52946
rect 4114 52894 4126 52946
rect 5058 52894 5070 52946
rect 5122 52894 5134 52946
rect 6626 52894 6638 52946
rect 6690 52894 6702 52946
rect 10210 52894 10222 52946
rect 10274 52894 10286 52946
rect 14802 52894 14814 52946
rect 14866 52894 14878 52946
rect 17378 52894 17390 52946
rect 17442 52894 17454 52946
rect 9886 52882 9938 52894
rect 12574 52882 12626 52894
rect 15150 52882 15202 52894
rect 20302 52882 20354 52894
rect 21086 52946 21138 52958
rect 24546 52894 24558 52946
rect 24610 52894 24622 52946
rect 25218 52894 25230 52946
rect 25282 52894 25294 52946
rect 21086 52882 21138 52894
rect 2158 52834 2210 52846
rect 2158 52770 2210 52782
rect 2606 52834 2658 52846
rect 7646 52834 7698 52846
rect 4610 52782 4622 52834
rect 4674 52782 4686 52834
rect 5618 52782 5630 52834
rect 5682 52782 5694 52834
rect 2606 52770 2658 52782
rect 7646 52770 7698 52782
rect 8094 52834 8146 52846
rect 8094 52770 8146 52782
rect 10894 52834 10946 52846
rect 10894 52770 10946 52782
rect 12798 52834 12850 52846
rect 19182 52834 19234 52846
rect 13570 52782 13582 52834
rect 13634 52782 13646 52834
rect 21746 52782 21758 52834
rect 21810 52782 21822 52834
rect 28130 52782 28142 52834
rect 28194 52782 28206 52834
rect 12798 52770 12850 52782
rect 19182 52770 19234 52782
rect 2718 52722 2770 52734
rect 6626 52670 6638 52722
rect 6690 52670 6702 52722
rect 8194 52670 8206 52722
rect 8258 52719 8270 52722
rect 8978 52719 8990 52722
rect 8258 52673 8990 52719
rect 8258 52670 8270 52673
rect 8978 52670 8990 52673
rect 9042 52670 9054 52722
rect 10434 52670 10446 52722
rect 10498 52719 10510 52722
rect 11330 52719 11342 52722
rect 10498 52673 11342 52719
rect 10498 52670 10510 52673
rect 11330 52670 11342 52673
rect 11394 52670 11406 52722
rect 2718 52658 2770 52670
rect 1344 52554 28560 52588
rect 1344 52502 4616 52554
rect 4668 52502 4720 52554
rect 4772 52502 4824 52554
rect 4876 52502 11420 52554
rect 11472 52502 11524 52554
rect 11576 52502 11628 52554
rect 11680 52502 18224 52554
rect 18276 52502 18328 52554
rect 18380 52502 18432 52554
rect 18484 52502 25028 52554
rect 25080 52502 25132 52554
rect 25184 52502 25236 52554
rect 25288 52502 28560 52554
rect 1344 52468 28560 52502
rect 11006 52386 11058 52398
rect 5954 52334 5966 52386
rect 6018 52383 6030 52386
rect 6514 52383 6526 52386
rect 6018 52337 6526 52383
rect 6018 52334 6030 52337
rect 6514 52334 6526 52337
rect 6578 52334 6590 52386
rect 10658 52334 10670 52386
rect 10722 52334 10734 52386
rect 11006 52322 11058 52334
rect 20750 52386 20802 52398
rect 21858 52334 21870 52386
rect 21922 52334 21934 52386
rect 20750 52322 20802 52334
rect 3390 52274 3442 52286
rect 2818 52222 2830 52274
rect 2882 52222 2894 52274
rect 3390 52210 3442 52222
rect 5854 52274 5906 52286
rect 5854 52210 5906 52222
rect 6750 52274 6802 52286
rect 6750 52210 6802 52222
rect 7086 52274 7138 52286
rect 11230 52274 11282 52286
rect 8194 52222 8206 52274
rect 8258 52222 8270 52274
rect 10322 52222 10334 52274
rect 10386 52222 10398 52274
rect 7086 52210 7138 52222
rect 11230 52210 11282 52222
rect 13022 52274 13074 52286
rect 19742 52274 19794 52286
rect 14130 52222 14142 52274
rect 14194 52222 14206 52274
rect 13022 52210 13074 52222
rect 19742 52210 19794 52222
rect 23886 52274 23938 52286
rect 23886 52210 23938 52222
rect 24334 52274 24386 52286
rect 24334 52210 24386 52222
rect 24782 52274 24834 52286
rect 27470 52274 27522 52286
rect 26226 52222 26238 52274
rect 26290 52222 26302 52274
rect 24782 52210 24834 52222
rect 27470 52210 27522 52222
rect 3726 52162 3778 52174
rect 2482 52110 2494 52162
rect 2546 52110 2558 52162
rect 3726 52098 3778 52110
rect 4174 52162 4226 52174
rect 4174 52098 4226 52110
rect 4286 52162 4338 52174
rect 12014 52162 12066 52174
rect 4722 52110 4734 52162
rect 4786 52110 4798 52162
rect 7522 52110 7534 52162
rect 7586 52110 7598 52162
rect 4286 52098 4338 52110
rect 12014 52098 12066 52110
rect 12126 52162 12178 52174
rect 19966 52162 20018 52174
rect 14018 52110 14030 52162
rect 14082 52110 14094 52162
rect 15586 52110 15598 52162
rect 15650 52110 15662 52162
rect 17602 52110 17614 52162
rect 17666 52110 17678 52162
rect 12126 52098 12178 52110
rect 19966 52098 20018 52110
rect 20078 52162 20130 52174
rect 20078 52098 20130 52110
rect 20526 52162 20578 52174
rect 22766 52162 22818 52174
rect 21522 52110 21534 52162
rect 21586 52110 21598 52162
rect 21858 52110 21870 52162
rect 21922 52110 21934 52162
rect 22418 52110 22430 52162
rect 22482 52110 22494 52162
rect 20526 52098 20578 52110
rect 22766 52098 22818 52110
rect 22990 52162 23042 52174
rect 22990 52098 23042 52110
rect 25230 52162 25282 52174
rect 25230 52098 25282 52110
rect 26350 52162 26402 52174
rect 26786 52110 26798 52162
rect 26850 52110 26862 52162
rect 27122 52110 27134 52162
rect 27186 52110 27198 52162
rect 26350 52098 26402 52110
rect 2270 52050 2322 52062
rect 2270 51986 2322 51998
rect 6190 52050 6242 52062
rect 6190 51986 6242 51998
rect 12350 52050 12402 52062
rect 16718 52050 16770 52062
rect 15026 51998 15038 52050
rect 15090 51998 15102 52050
rect 12350 51986 12402 51998
rect 16718 51986 16770 51998
rect 18174 52050 18226 52062
rect 18174 51986 18226 51998
rect 21310 52050 21362 52062
rect 21310 51986 21362 51998
rect 26238 52050 26290 52062
rect 26238 51986 26290 51998
rect 26574 52050 26626 52062
rect 26574 51986 26626 51998
rect 27582 52050 27634 52062
rect 27582 51986 27634 51998
rect 27806 52050 27858 52062
rect 27806 51986 27858 51998
rect 4398 51938 4450 51950
rect 4398 51874 4450 51886
rect 4510 51938 4562 51950
rect 23438 51938 23490 51950
rect 17714 51886 17726 51938
rect 17778 51886 17790 51938
rect 21634 51886 21646 51938
rect 21698 51886 21710 51938
rect 4510 51874 4562 51886
rect 23438 51874 23490 51886
rect 25678 51938 25730 51950
rect 25678 51874 25730 51886
rect 27358 51938 27410 51950
rect 27358 51874 27410 51886
rect 1344 51770 28720 51804
rect 1344 51718 8018 51770
rect 8070 51718 8122 51770
rect 8174 51718 8226 51770
rect 8278 51718 14822 51770
rect 14874 51718 14926 51770
rect 14978 51718 15030 51770
rect 15082 51718 21626 51770
rect 21678 51718 21730 51770
rect 21782 51718 21834 51770
rect 21886 51718 28430 51770
rect 28482 51718 28534 51770
rect 28586 51718 28638 51770
rect 28690 51718 28720 51770
rect 1344 51684 28720 51718
rect 2494 51602 2546 51614
rect 2494 51538 2546 51550
rect 4734 51602 4786 51614
rect 4734 51538 4786 51550
rect 5630 51602 5682 51614
rect 5630 51538 5682 51550
rect 7310 51602 7362 51614
rect 7310 51538 7362 51550
rect 7758 51602 7810 51614
rect 7758 51538 7810 51550
rect 8990 51602 9042 51614
rect 8990 51538 9042 51550
rect 16830 51602 16882 51614
rect 16830 51538 16882 51550
rect 17502 51602 17554 51614
rect 17502 51538 17554 51550
rect 19406 51602 19458 51614
rect 19406 51538 19458 51550
rect 19742 51602 19794 51614
rect 19742 51538 19794 51550
rect 23214 51602 23266 51614
rect 23214 51538 23266 51550
rect 24334 51602 24386 51614
rect 24334 51538 24386 51550
rect 27694 51602 27746 51614
rect 27694 51538 27746 51550
rect 4062 51490 4114 51502
rect 4062 51426 4114 51438
rect 5182 51490 5234 51502
rect 5182 51426 5234 51438
rect 5854 51490 5906 51502
rect 18622 51490 18674 51502
rect 10098 51438 10110 51490
rect 10162 51438 10174 51490
rect 5854 51426 5906 51438
rect 18622 51426 18674 51438
rect 18734 51490 18786 51502
rect 23326 51490 23378 51502
rect 20850 51438 20862 51490
rect 20914 51438 20926 51490
rect 18734 51426 18786 51438
rect 23326 51426 23378 51438
rect 25790 51490 25842 51502
rect 25790 51426 25842 51438
rect 26238 51490 26290 51502
rect 26238 51426 26290 51438
rect 3614 51378 3666 51390
rect 3614 51314 3666 51326
rect 6190 51378 6242 51390
rect 6190 51314 6242 51326
rect 6414 51378 6466 51390
rect 8766 51378 8818 51390
rect 16158 51378 16210 51390
rect 8418 51326 8430 51378
rect 8482 51326 8494 51378
rect 13458 51326 13470 51378
rect 13522 51326 13534 51378
rect 6414 51314 6466 51326
rect 8766 51314 8818 51326
rect 16158 51314 16210 51326
rect 16270 51378 16322 51390
rect 16270 51314 16322 51326
rect 18398 51378 18450 51390
rect 18398 51314 18450 51326
rect 19182 51378 19234 51390
rect 23886 51378 23938 51390
rect 26462 51378 26514 51390
rect 20178 51326 20190 51378
rect 20242 51326 20254 51378
rect 23538 51326 23550 51378
rect 23602 51326 23614 51378
rect 24098 51326 24110 51378
rect 24162 51326 24174 51378
rect 26786 51326 26798 51378
rect 26850 51326 26862 51378
rect 19182 51314 19234 51326
rect 23886 51314 23938 51326
rect 26462 51314 26514 51326
rect 2046 51266 2098 51278
rect 2046 51202 2098 51214
rect 3950 51266 4002 51278
rect 3950 51202 4002 51214
rect 5966 51266 6018 51278
rect 5966 51202 6018 51214
rect 8206 51266 8258 51278
rect 8206 51202 8258 51214
rect 8878 51266 8930 51278
rect 17950 51266 18002 51278
rect 25342 51266 25394 51278
rect 15362 51214 15374 51266
rect 15426 51214 15438 51266
rect 22978 51214 22990 51266
rect 23042 51214 23054 51266
rect 8878 51202 8930 51214
rect 17950 51202 18002 51214
rect 25342 51202 25394 51214
rect 26350 51266 26402 51278
rect 26350 51202 26402 51214
rect 27246 51266 27298 51278
rect 27246 51202 27298 51214
rect 28142 51266 28194 51278
rect 28142 51202 28194 51214
rect 2382 51154 2434 51166
rect 2382 51090 2434 51102
rect 2718 51154 2770 51166
rect 2718 51090 2770 51102
rect 3838 51154 3890 51166
rect 3838 51090 3890 51102
rect 15934 51154 15986 51166
rect 15934 51090 15986 51102
rect 24446 51154 24498 51166
rect 27346 51102 27358 51154
rect 27410 51151 27422 51154
rect 28018 51151 28030 51154
rect 27410 51105 28030 51151
rect 27410 51102 27422 51105
rect 28018 51102 28030 51105
rect 28082 51102 28094 51154
rect 24446 51090 24498 51102
rect 1344 50986 28560 51020
rect 1344 50934 4616 50986
rect 4668 50934 4720 50986
rect 4772 50934 4824 50986
rect 4876 50934 11420 50986
rect 11472 50934 11524 50986
rect 11576 50934 11628 50986
rect 11680 50934 18224 50986
rect 18276 50934 18328 50986
rect 18380 50934 18432 50986
rect 18484 50934 25028 50986
rect 25080 50934 25132 50986
rect 25184 50934 25236 50986
rect 25288 50934 28560 50986
rect 1344 50900 28560 50934
rect 22318 50818 22370 50830
rect 20178 50766 20190 50818
rect 20242 50815 20254 50818
rect 20738 50815 20750 50818
rect 20242 50769 20750 50815
rect 20242 50766 20254 50769
rect 20738 50766 20750 50769
rect 20802 50766 20814 50818
rect 22318 50754 22370 50766
rect 5182 50706 5234 50718
rect 4610 50654 4622 50706
rect 4674 50654 4686 50706
rect 5182 50642 5234 50654
rect 6526 50706 6578 50718
rect 10670 50706 10722 50718
rect 10210 50654 10222 50706
rect 10274 50654 10286 50706
rect 6526 50642 6578 50654
rect 10670 50642 10722 50654
rect 11118 50706 11170 50718
rect 11118 50642 11170 50654
rect 19630 50706 19682 50718
rect 19630 50642 19682 50654
rect 24334 50706 24386 50718
rect 27794 50654 27806 50706
rect 27858 50654 27870 50706
rect 24334 50642 24386 50654
rect 6190 50594 6242 50606
rect 1810 50542 1822 50594
rect 1874 50542 1886 50594
rect 6190 50530 6242 50542
rect 6414 50594 6466 50606
rect 6414 50530 6466 50542
rect 6638 50594 6690 50606
rect 7298 50542 7310 50594
rect 7362 50542 7374 50594
rect 11442 50542 11454 50594
rect 11506 50542 11518 50594
rect 6638 50530 6690 50542
rect 12462 50538 12514 50550
rect 12674 50542 12686 50594
rect 12738 50542 12750 50594
rect 13570 50542 13582 50594
rect 13634 50542 13646 50594
rect 15362 50542 15374 50594
rect 15426 50542 15438 50594
rect 17378 50542 17390 50594
rect 17442 50542 17454 50594
rect 21410 50542 21422 50594
rect 21474 50542 21486 50594
rect 24882 50542 24894 50594
rect 24946 50542 24958 50594
rect 6862 50482 6914 50494
rect 2482 50430 2494 50482
rect 2546 50430 2558 50482
rect 8082 50430 8094 50482
rect 8146 50430 8158 50482
rect 11554 50430 11566 50482
rect 11618 50430 11630 50482
rect 12462 50474 12514 50486
rect 13022 50482 13074 50494
rect 16494 50482 16546 50494
rect 14802 50430 14814 50482
rect 14866 50430 14878 50482
rect 15026 50430 15038 50482
rect 15090 50430 15102 50482
rect 19170 50430 19182 50482
rect 19234 50430 19246 50482
rect 25666 50430 25678 50482
rect 25730 50430 25742 50482
rect 6862 50418 6914 50430
rect 13022 50418 13074 50430
rect 16494 50418 16546 50430
rect 20078 50370 20130 50382
rect 15586 50318 15598 50370
rect 15650 50318 15662 50370
rect 20078 50306 20130 50318
rect 20526 50370 20578 50382
rect 20526 50306 20578 50318
rect 1344 50202 28720 50236
rect 1344 50150 8018 50202
rect 8070 50150 8122 50202
rect 8174 50150 8226 50202
rect 8278 50150 14822 50202
rect 14874 50150 14926 50202
rect 14978 50150 15030 50202
rect 15082 50150 21626 50202
rect 21678 50150 21730 50202
rect 21782 50150 21834 50202
rect 21886 50150 28430 50202
rect 28482 50150 28534 50202
rect 28586 50150 28638 50202
rect 28690 50150 28720 50202
rect 1344 50116 28720 50150
rect 8094 50034 8146 50046
rect 3154 49982 3166 50034
rect 3218 49982 3230 50034
rect 8094 49970 8146 49982
rect 8542 50034 8594 50046
rect 8542 49970 8594 49982
rect 9998 50034 10050 50046
rect 9998 49970 10050 49982
rect 11006 50034 11058 50046
rect 25678 50034 25730 50046
rect 16706 49982 16718 50034
rect 16770 49982 16782 50034
rect 11006 49970 11058 49982
rect 25678 49970 25730 49982
rect 2046 49922 2098 49934
rect 2046 49858 2098 49870
rect 2830 49922 2882 49934
rect 9550 49922 9602 49934
rect 5282 49870 5294 49922
rect 5346 49870 5358 49922
rect 2830 49858 2882 49870
rect 9550 49858 9602 49870
rect 10558 49922 10610 49934
rect 10558 49858 10610 49870
rect 12238 49922 12290 49934
rect 12238 49858 12290 49870
rect 13582 49922 13634 49934
rect 18510 49922 18562 49934
rect 16818 49870 16830 49922
rect 16882 49870 16894 49922
rect 13582 49858 13634 49870
rect 18510 49858 18562 49870
rect 19966 49922 20018 49934
rect 19966 49858 20018 49870
rect 26126 49922 26178 49934
rect 26126 49858 26178 49870
rect 1710 49810 1762 49822
rect 1710 49746 1762 49758
rect 3166 49810 3218 49822
rect 8430 49810 8482 49822
rect 3378 49758 3390 49810
rect 3442 49758 3454 49810
rect 4610 49758 4622 49810
rect 4674 49758 4686 49810
rect 3166 49746 3218 49758
rect 8430 49746 8482 49758
rect 8654 49810 8706 49822
rect 8654 49746 8706 49758
rect 8878 49810 8930 49822
rect 8878 49746 8930 49758
rect 9774 49810 9826 49822
rect 9774 49746 9826 49758
rect 10110 49810 10162 49822
rect 10110 49746 10162 49758
rect 10782 49810 10834 49822
rect 12462 49810 12514 49822
rect 11218 49758 11230 49810
rect 11282 49758 11294 49810
rect 10782 49746 10834 49758
rect 12462 49746 12514 49758
rect 12686 49810 12738 49822
rect 15150 49810 15202 49822
rect 19518 49810 19570 49822
rect 25566 49810 25618 49822
rect 13010 49758 13022 49810
rect 13074 49758 13086 49810
rect 18946 49758 18958 49810
rect 19010 49758 19022 49810
rect 21858 49758 21870 49810
rect 21922 49758 21934 49810
rect 12686 49746 12738 49758
rect 15150 49746 15202 49758
rect 19518 49746 19570 49758
rect 25566 49746 25618 49758
rect 25902 49810 25954 49822
rect 25902 49746 25954 49758
rect 2494 49698 2546 49710
rect 2494 49634 2546 49646
rect 4174 49698 4226 49710
rect 9886 49698 9938 49710
rect 26574 49698 26626 49710
rect 7410 49646 7422 49698
rect 7474 49646 7486 49698
rect 10994 49646 11006 49698
rect 11058 49646 11070 49698
rect 19730 49646 19742 49698
rect 19794 49646 19806 49698
rect 22530 49646 22542 49698
rect 22594 49646 22606 49698
rect 24658 49646 24670 49698
rect 24722 49646 24734 49698
rect 4174 49634 4226 49646
rect 9886 49634 9938 49646
rect 26574 49634 26626 49646
rect 27022 49698 27074 49710
rect 27022 49634 27074 49646
rect 27470 49698 27522 49710
rect 27470 49634 27522 49646
rect 27918 49698 27970 49710
rect 27918 49634 27970 49646
rect 3378 49534 3390 49586
rect 3442 49534 3454 49586
rect 11890 49534 11902 49586
rect 11954 49534 11966 49586
rect 26898 49534 26910 49586
rect 26962 49583 26974 49586
rect 27906 49583 27918 49586
rect 26962 49537 27918 49583
rect 26962 49534 26974 49537
rect 27906 49534 27918 49537
rect 27970 49534 27982 49586
rect 1344 49418 28560 49452
rect 1344 49366 4616 49418
rect 4668 49366 4720 49418
rect 4772 49366 4824 49418
rect 4876 49366 11420 49418
rect 11472 49366 11524 49418
rect 11576 49366 11628 49418
rect 11680 49366 18224 49418
rect 18276 49366 18328 49418
rect 18380 49366 18432 49418
rect 18484 49366 25028 49418
rect 25080 49366 25132 49418
rect 25184 49366 25236 49418
rect 25288 49366 28560 49418
rect 1344 49332 28560 49366
rect 25230 49250 25282 49262
rect 7410 49198 7422 49250
rect 7474 49247 7486 49250
rect 8194 49247 8206 49250
rect 7474 49201 8206 49247
rect 7474 49198 7486 49201
rect 8194 49198 8206 49201
rect 8258 49198 8270 49250
rect 13570 49198 13582 49250
rect 13634 49198 13646 49250
rect 23874 49198 23886 49250
rect 23938 49198 23950 49250
rect 25230 49186 25282 49198
rect 1822 49138 1874 49150
rect 1822 49074 1874 49086
rect 2606 49138 2658 49150
rect 2606 49074 2658 49086
rect 5630 49138 5682 49150
rect 5630 49074 5682 49086
rect 6526 49138 6578 49150
rect 6526 49074 6578 49086
rect 6862 49138 6914 49150
rect 6862 49074 6914 49086
rect 7422 49138 7474 49150
rect 7422 49074 7474 49086
rect 7870 49138 7922 49150
rect 7870 49074 7922 49086
rect 8206 49138 8258 49150
rect 8206 49074 8258 49086
rect 8654 49138 8706 49150
rect 8654 49074 8706 49086
rect 9102 49138 9154 49150
rect 9102 49074 9154 49086
rect 9550 49138 9602 49150
rect 9550 49074 9602 49086
rect 10894 49138 10946 49150
rect 10894 49074 10946 49086
rect 11342 49138 11394 49150
rect 23438 49138 23490 49150
rect 15362 49086 15374 49138
rect 15426 49086 15438 49138
rect 21410 49086 21422 49138
rect 21474 49086 21486 49138
rect 11342 49074 11394 49086
rect 23438 49074 23490 49086
rect 27134 49138 27186 49150
rect 27134 49074 27186 49086
rect 27582 49138 27634 49150
rect 27582 49074 27634 49086
rect 3614 49026 3666 49038
rect 3614 48962 3666 48974
rect 3950 49026 4002 49038
rect 12126 49026 12178 49038
rect 11778 48974 11790 49026
rect 11842 48974 11854 49026
rect 3950 48962 4002 48974
rect 12126 48962 12178 48974
rect 12350 49026 12402 49038
rect 14142 49026 14194 49038
rect 18622 49026 18674 49038
rect 21870 49026 21922 49038
rect 13906 48974 13918 49026
rect 13970 48974 13982 49026
rect 15922 48974 15934 49026
rect 15986 48974 15998 49026
rect 18946 48974 18958 49026
rect 19010 48974 19022 49026
rect 12350 48962 12402 48974
rect 14142 48962 14194 48974
rect 18622 48962 18674 48974
rect 21870 48962 21922 48974
rect 23662 49026 23714 49038
rect 26014 49026 26066 49038
rect 24098 48974 24110 49026
rect 24162 48974 24174 49026
rect 24658 48974 24670 49026
rect 24722 48974 24734 49026
rect 25218 48974 25230 49026
rect 25282 48974 25294 49026
rect 23662 48962 23714 48974
rect 26014 48962 26066 48974
rect 26350 49026 26402 49038
rect 26350 48962 26402 48974
rect 12574 48914 12626 48926
rect 12574 48850 12626 48862
rect 14366 48914 14418 48926
rect 14366 48850 14418 48862
rect 14590 48914 14642 48926
rect 23326 48914 23378 48926
rect 14914 48862 14926 48914
rect 14978 48862 14990 48914
rect 17042 48862 17054 48914
rect 17106 48862 17118 48914
rect 18834 48862 18846 48914
rect 18898 48862 18910 48914
rect 20626 48862 20638 48914
rect 20690 48862 20702 48914
rect 14590 48850 14642 48862
rect 23326 48850 23378 48862
rect 24446 48914 24498 48926
rect 24446 48850 24498 48862
rect 24894 48914 24946 48926
rect 24894 48850 24946 48862
rect 25566 48914 25618 48926
rect 25566 48850 25618 48862
rect 26686 48914 26738 48926
rect 26686 48850 26738 48862
rect 2942 48802 2994 48814
rect 2942 48738 2994 48750
rect 4062 48802 4114 48814
rect 4062 48738 4114 48750
rect 4174 48802 4226 48814
rect 4174 48738 4226 48750
rect 4958 48802 5010 48814
rect 4958 48738 5010 48750
rect 5742 48802 5794 48814
rect 5742 48738 5794 48750
rect 9998 48802 10050 48814
rect 9998 48738 10050 48750
rect 10558 48802 10610 48814
rect 10558 48738 10610 48750
rect 24334 48802 24386 48814
rect 24334 48738 24386 48750
rect 26238 48802 26290 48814
rect 26238 48738 26290 48750
rect 28030 48802 28082 48814
rect 28030 48738 28082 48750
rect 1344 48634 28720 48668
rect 1344 48582 8018 48634
rect 8070 48582 8122 48634
rect 8174 48582 8226 48634
rect 8278 48582 14822 48634
rect 14874 48582 14926 48634
rect 14978 48582 15030 48634
rect 15082 48582 21626 48634
rect 21678 48582 21730 48634
rect 21782 48582 21834 48634
rect 21886 48582 28430 48634
rect 28482 48582 28534 48634
rect 28586 48582 28638 48634
rect 28690 48582 28720 48634
rect 1344 48548 28720 48582
rect 6190 48466 6242 48478
rect 6190 48402 6242 48414
rect 7534 48466 7586 48478
rect 7534 48402 7586 48414
rect 9550 48466 9602 48478
rect 9550 48402 9602 48414
rect 9998 48466 10050 48478
rect 9998 48402 10050 48414
rect 11790 48466 11842 48478
rect 11790 48402 11842 48414
rect 12238 48466 12290 48478
rect 12238 48402 12290 48414
rect 12686 48466 12738 48478
rect 16594 48414 16606 48466
rect 16658 48414 16670 48466
rect 12686 48402 12738 48414
rect 5854 48354 5906 48366
rect 5854 48290 5906 48302
rect 11342 48354 11394 48366
rect 11342 48290 11394 48302
rect 14142 48354 14194 48366
rect 20526 48354 20578 48366
rect 16818 48302 16830 48354
rect 16882 48302 16894 48354
rect 17490 48302 17502 48354
rect 17554 48302 17566 48354
rect 14142 48290 14194 48302
rect 20526 48290 20578 48302
rect 22094 48354 22146 48366
rect 26002 48302 26014 48354
rect 26066 48302 26078 48354
rect 22094 48290 22146 48302
rect 8318 48242 8370 48254
rect 1810 48190 1822 48242
rect 1874 48190 1886 48242
rect 5282 48190 5294 48242
rect 5346 48190 5358 48242
rect 8318 48178 8370 48190
rect 8542 48242 8594 48254
rect 8542 48178 8594 48190
rect 8878 48242 8930 48254
rect 8878 48178 8930 48190
rect 9774 48242 9826 48254
rect 19518 48242 19570 48254
rect 14578 48190 14590 48242
rect 14642 48190 14654 48242
rect 15026 48190 15038 48242
rect 15090 48190 15102 48242
rect 17378 48190 17390 48242
rect 17442 48190 17454 48242
rect 9774 48178 9826 48190
rect 19518 48178 19570 48190
rect 21646 48242 21698 48254
rect 25330 48190 25342 48242
rect 25394 48190 25406 48242
rect 21646 48178 21698 48190
rect 6638 48130 6690 48142
rect 2482 48078 2494 48130
rect 2546 48078 2558 48130
rect 4610 48078 4622 48130
rect 4674 48078 4686 48130
rect 6638 48066 6690 48078
rect 7086 48130 7138 48142
rect 7086 48066 7138 48078
rect 8094 48130 8146 48142
rect 8094 48066 8146 48078
rect 8430 48130 8482 48142
rect 8430 48066 8482 48078
rect 9662 48130 9714 48142
rect 9662 48066 9714 48078
rect 10782 48130 10834 48142
rect 23326 48130 23378 48142
rect 19954 48078 19966 48130
rect 20018 48078 20030 48130
rect 10782 48066 10834 48078
rect 23326 48066 23378 48078
rect 23438 48130 23490 48142
rect 23438 48066 23490 48078
rect 24558 48130 24610 48142
rect 28130 48078 28142 48130
rect 28194 48078 28206 48130
rect 24558 48066 24610 48078
rect 4958 48018 5010 48030
rect 4958 47954 5010 47966
rect 5294 48018 5346 48030
rect 6066 47966 6078 48018
rect 6130 48015 6142 48018
rect 6626 48015 6638 48018
rect 6130 47969 6638 48015
rect 6130 47966 6142 47969
rect 6626 47966 6638 47969
rect 6690 47966 6702 48018
rect 11778 47966 11790 48018
rect 11842 48015 11854 48018
rect 12114 48015 12126 48018
rect 11842 47969 12126 48015
rect 11842 47966 11854 47969
rect 12114 47966 12126 47969
rect 12178 47966 12190 48018
rect 5294 47954 5346 47966
rect 1344 47850 28560 47884
rect 1344 47798 4616 47850
rect 4668 47798 4720 47850
rect 4772 47798 4824 47850
rect 4876 47798 11420 47850
rect 11472 47798 11524 47850
rect 11576 47798 11628 47850
rect 11680 47798 18224 47850
rect 18276 47798 18328 47850
rect 18380 47798 18432 47850
rect 18484 47798 25028 47850
rect 25080 47798 25132 47850
rect 25184 47798 25236 47850
rect 25288 47798 28560 47850
rect 1344 47764 28560 47798
rect 20862 47682 20914 47694
rect 3490 47630 3502 47682
rect 3554 47630 3566 47682
rect 10994 47630 11006 47682
rect 11058 47679 11070 47682
rect 11554 47679 11566 47682
rect 11058 47633 11566 47679
rect 11058 47630 11070 47633
rect 11554 47630 11566 47633
rect 11618 47630 11630 47682
rect 21298 47630 21310 47682
rect 21362 47630 21374 47682
rect 28018 47679 28030 47682
rect 27361 47633 28030 47679
rect 20862 47618 20914 47630
rect 2494 47570 2546 47582
rect 2494 47506 2546 47518
rect 3054 47570 3106 47582
rect 3054 47506 3106 47518
rect 4286 47570 4338 47582
rect 4286 47506 4338 47518
rect 4734 47570 4786 47582
rect 10334 47570 10386 47582
rect 7410 47518 7422 47570
rect 7474 47518 7486 47570
rect 9538 47518 9550 47570
rect 9602 47518 9614 47570
rect 4734 47506 4786 47518
rect 10334 47506 10386 47518
rect 11230 47570 11282 47582
rect 11230 47506 11282 47518
rect 11566 47570 11618 47582
rect 11566 47506 11618 47518
rect 12462 47570 12514 47582
rect 12462 47506 12514 47518
rect 19518 47570 19570 47582
rect 19518 47506 19570 47518
rect 20078 47570 20130 47582
rect 20078 47506 20130 47518
rect 21646 47570 21698 47582
rect 26798 47570 26850 47582
rect 26338 47518 26350 47570
rect 26402 47518 26414 47570
rect 27234 47518 27246 47570
rect 27298 47567 27310 47570
rect 27361 47567 27407 47633
rect 28018 47630 28030 47633
rect 28082 47630 28094 47682
rect 27298 47521 27407 47567
rect 27694 47570 27746 47582
rect 27298 47518 27310 47521
rect 21646 47506 21698 47518
rect 26798 47506 26850 47518
rect 27694 47506 27746 47518
rect 28142 47570 28194 47582
rect 28142 47506 28194 47518
rect 2942 47458 2994 47470
rect 10222 47458 10274 47470
rect 3154 47406 3166 47458
rect 3218 47406 3230 47458
rect 3490 47406 3502 47458
rect 3554 47406 3566 47458
rect 5730 47406 5742 47458
rect 5794 47406 5806 47458
rect 6738 47406 6750 47458
rect 6802 47406 6814 47458
rect 2942 47394 2994 47406
rect 10222 47394 10274 47406
rect 10558 47458 10610 47470
rect 14142 47458 14194 47470
rect 13906 47406 13918 47458
rect 13970 47406 13982 47458
rect 10558 47394 10610 47406
rect 14142 47394 14194 47406
rect 14702 47458 14754 47470
rect 18958 47458 19010 47470
rect 15250 47406 15262 47458
rect 15314 47406 15326 47458
rect 14702 47394 14754 47406
rect 18958 47394 19010 47406
rect 21870 47458 21922 47470
rect 26686 47458 26738 47470
rect 23538 47406 23550 47458
rect 23602 47406 23614 47458
rect 21870 47394 21922 47406
rect 26686 47394 26738 47406
rect 1710 47346 1762 47358
rect 1710 47282 1762 47294
rect 9998 47346 10050 47358
rect 9998 47282 10050 47294
rect 10446 47346 10498 47358
rect 10446 47282 10498 47294
rect 14366 47346 14418 47358
rect 14366 47282 14418 47294
rect 16382 47346 16434 47358
rect 16382 47282 16434 47294
rect 17054 47346 17106 47358
rect 17054 47282 17106 47294
rect 18398 47346 18450 47358
rect 18398 47282 18450 47294
rect 20302 47346 20354 47358
rect 20302 47282 20354 47294
rect 22318 47346 22370 47358
rect 22318 47282 22370 47294
rect 22766 47346 22818 47358
rect 26910 47346 26962 47358
rect 24210 47294 24222 47346
rect 24274 47294 24286 47346
rect 22766 47282 22818 47294
rect 26910 47282 26962 47294
rect 2046 47234 2098 47246
rect 2046 47170 2098 47182
rect 5854 47234 5906 47246
rect 5854 47170 5906 47182
rect 12014 47234 12066 47246
rect 12014 47170 12066 47182
rect 12910 47234 12962 47246
rect 20526 47234 20578 47246
rect 13570 47182 13582 47234
rect 13634 47182 13646 47234
rect 12910 47170 12962 47182
rect 20526 47170 20578 47182
rect 20750 47234 20802 47246
rect 20750 47170 20802 47182
rect 27134 47234 27186 47246
rect 27134 47170 27186 47182
rect 1344 47066 28720 47100
rect 1344 47014 8018 47066
rect 8070 47014 8122 47066
rect 8174 47014 8226 47066
rect 8278 47014 14822 47066
rect 14874 47014 14926 47066
rect 14978 47014 15030 47066
rect 15082 47014 21626 47066
rect 21678 47014 21730 47066
rect 21782 47014 21834 47066
rect 21886 47014 28430 47066
rect 28482 47014 28534 47066
rect 28586 47014 28638 47066
rect 28690 47014 28720 47066
rect 1344 46980 28720 47014
rect 4062 46898 4114 46910
rect 4062 46834 4114 46846
rect 5070 46898 5122 46910
rect 5070 46834 5122 46846
rect 9998 46898 10050 46910
rect 9998 46834 10050 46846
rect 13918 46898 13970 46910
rect 13918 46834 13970 46846
rect 15262 46898 15314 46910
rect 15262 46834 15314 46846
rect 18958 46898 19010 46910
rect 18958 46834 19010 46846
rect 21646 46898 21698 46910
rect 21646 46834 21698 46846
rect 22878 46898 22930 46910
rect 22878 46834 22930 46846
rect 24222 46898 24274 46910
rect 24222 46834 24274 46846
rect 25454 46898 25506 46910
rect 25454 46834 25506 46846
rect 26686 46898 26738 46910
rect 26686 46834 26738 46846
rect 27134 46898 27186 46910
rect 27134 46834 27186 46846
rect 28142 46898 28194 46910
rect 28142 46834 28194 46846
rect 2046 46786 2098 46798
rect 2046 46722 2098 46734
rect 4846 46786 4898 46798
rect 4846 46722 4898 46734
rect 16270 46786 16322 46798
rect 16270 46722 16322 46734
rect 17950 46786 18002 46798
rect 17950 46722 18002 46734
rect 22094 46786 22146 46798
rect 22094 46722 22146 46734
rect 1710 46674 1762 46686
rect 15038 46674 15090 46686
rect 20302 46674 20354 46686
rect 5506 46622 5518 46674
rect 5570 46622 5582 46674
rect 10322 46622 10334 46674
rect 10386 46622 10398 46674
rect 15250 46622 15262 46674
rect 15314 46622 15326 46674
rect 17378 46622 17390 46674
rect 17442 46622 17454 46674
rect 1710 46610 1762 46622
rect 15038 46610 15090 46622
rect 20302 46610 20354 46622
rect 20526 46674 20578 46686
rect 23102 46674 23154 46686
rect 20850 46622 20862 46674
rect 20914 46622 20926 46674
rect 21186 46622 21198 46674
rect 21250 46622 21262 46674
rect 21410 46622 21422 46674
rect 21474 46622 21486 46674
rect 20526 46610 20578 46622
rect 23102 46610 23154 46622
rect 23326 46674 23378 46686
rect 23326 46610 23378 46622
rect 23886 46674 23938 46686
rect 23886 46610 23938 46622
rect 24334 46674 24386 46686
rect 24334 46610 24386 46622
rect 24558 46674 24610 46686
rect 24558 46610 24610 46622
rect 25230 46674 25282 46686
rect 25230 46610 25282 46622
rect 25342 46674 25394 46686
rect 25778 46622 25790 46674
rect 25842 46622 25854 46674
rect 25342 46610 25394 46622
rect 2718 46562 2770 46574
rect 2718 46498 2770 46510
rect 3166 46562 3218 46574
rect 3166 46498 3218 46510
rect 3614 46562 3666 46574
rect 3614 46498 3666 46510
rect 4510 46562 4562 46574
rect 8990 46562 9042 46574
rect 19182 46562 19234 46574
rect 6290 46510 6302 46562
rect 6354 46510 6366 46562
rect 8418 46510 8430 46562
rect 8482 46510 8494 46562
rect 11106 46510 11118 46562
rect 11170 46510 11182 46562
rect 13234 46510 13246 46562
rect 13298 46510 13310 46562
rect 4510 46498 4562 46510
rect 8990 46498 9042 46510
rect 19182 46498 19234 46510
rect 20414 46562 20466 46574
rect 23214 46562 23266 46574
rect 21522 46510 21534 46562
rect 21586 46510 21598 46562
rect 20414 46498 20466 46510
rect 23214 46498 23266 46510
rect 26238 46562 26290 46574
rect 26238 46498 26290 46510
rect 27582 46562 27634 46574
rect 27582 46498 27634 46510
rect 5182 46450 5234 46462
rect 5182 46386 5234 46398
rect 1344 46282 28560 46316
rect 1344 46230 4616 46282
rect 4668 46230 4720 46282
rect 4772 46230 4824 46282
rect 4876 46230 11420 46282
rect 11472 46230 11524 46282
rect 11576 46230 11628 46282
rect 11680 46230 18224 46282
rect 18276 46230 18328 46282
rect 18380 46230 18432 46282
rect 18484 46230 25028 46282
rect 25080 46230 25132 46282
rect 25184 46230 25236 46282
rect 25288 46230 28560 46282
rect 1344 46196 28560 46230
rect 9426 46062 9438 46114
rect 9490 46111 9502 46114
rect 9986 46111 9998 46114
rect 9490 46065 9998 46111
rect 9490 46062 9502 46065
rect 9986 46062 9998 46065
rect 10050 46062 10062 46114
rect 10322 46062 10334 46114
rect 10386 46111 10398 46114
rect 10770 46111 10782 46114
rect 10386 46065 10782 46111
rect 10386 46062 10398 46065
rect 10770 46062 10782 46065
rect 10834 46062 10846 46114
rect 6862 46002 6914 46014
rect 4610 45950 4622 46002
rect 4674 45950 4686 46002
rect 6862 45938 6914 45950
rect 8990 46002 9042 46014
rect 8990 45938 9042 45950
rect 10334 46002 10386 46014
rect 10334 45938 10386 45950
rect 10782 46002 10834 46014
rect 25118 46002 25170 46014
rect 24210 45950 24222 46002
rect 24274 45950 24286 46002
rect 26562 45950 26574 46002
rect 26626 45950 26638 46002
rect 10782 45938 10834 45950
rect 25118 45938 25170 45950
rect 7310 45890 7362 45902
rect 1810 45838 1822 45890
rect 1874 45838 1886 45890
rect 7310 45826 7362 45838
rect 7870 45890 7922 45902
rect 7870 45826 7922 45838
rect 7982 45890 8034 45902
rect 9438 45890 9490 45902
rect 8306 45838 8318 45890
rect 8370 45838 8382 45890
rect 7982 45826 8034 45838
rect 9438 45826 9490 45838
rect 11230 45890 11282 45902
rect 15822 45890 15874 45902
rect 14354 45838 14366 45890
rect 14418 45838 14430 45890
rect 11230 45826 11282 45838
rect 15822 45826 15874 45838
rect 17838 45890 17890 45902
rect 17838 45826 17890 45838
rect 18286 45890 18338 45902
rect 21298 45838 21310 45890
rect 21362 45838 21374 45890
rect 27794 45838 27806 45890
rect 27858 45838 27870 45890
rect 18286 45826 18338 45838
rect 6414 45778 6466 45790
rect 2482 45726 2494 45778
rect 2546 45726 2558 45778
rect 6414 45714 6466 45726
rect 6750 45778 6802 45790
rect 6750 45714 6802 45726
rect 7086 45778 7138 45790
rect 7086 45714 7138 45726
rect 11118 45778 11170 45790
rect 11118 45714 11170 45726
rect 11454 45778 11506 45790
rect 11454 45714 11506 45726
rect 11678 45778 11730 45790
rect 11678 45714 11730 45726
rect 12238 45778 12290 45790
rect 19294 45778 19346 45790
rect 16258 45726 16270 45778
rect 16322 45726 16334 45778
rect 22082 45726 22094 45778
rect 22146 45726 22158 45778
rect 12238 45714 12290 45726
rect 19294 45714 19346 45726
rect 5182 45666 5234 45678
rect 5182 45602 5234 45614
rect 6078 45666 6130 45678
rect 6078 45602 6130 45614
rect 7758 45666 7810 45678
rect 7758 45602 7810 45614
rect 9886 45666 9938 45678
rect 9886 45602 9938 45614
rect 12126 45666 12178 45678
rect 12126 45602 12178 45614
rect 12350 45666 12402 45678
rect 12350 45602 12402 45614
rect 12574 45666 12626 45678
rect 12574 45602 12626 45614
rect 13806 45666 13858 45678
rect 20414 45666 20466 45678
rect 14690 45614 14702 45666
rect 14754 45614 14766 45666
rect 17154 45614 17166 45666
rect 17218 45614 17230 45666
rect 13806 45602 13858 45614
rect 20414 45602 20466 45614
rect 24670 45666 24722 45678
rect 24670 45602 24722 45614
rect 1344 45498 28720 45532
rect 1344 45446 8018 45498
rect 8070 45446 8122 45498
rect 8174 45446 8226 45498
rect 8278 45446 14822 45498
rect 14874 45446 14926 45498
rect 14978 45446 15030 45498
rect 15082 45446 21626 45498
rect 21678 45446 21730 45498
rect 21782 45446 21834 45498
rect 21886 45446 28430 45498
rect 28482 45446 28534 45498
rect 28586 45446 28638 45498
rect 28690 45446 28720 45498
rect 1344 45412 28720 45446
rect 4286 45330 4338 45342
rect 2594 45278 2606 45330
rect 2658 45278 2670 45330
rect 4286 45266 4338 45278
rect 5182 45330 5234 45342
rect 5182 45266 5234 45278
rect 5742 45330 5794 45342
rect 5742 45266 5794 45278
rect 11454 45330 11506 45342
rect 11454 45266 11506 45278
rect 11902 45330 11954 45342
rect 11902 45266 11954 45278
rect 12798 45330 12850 45342
rect 12798 45266 12850 45278
rect 15934 45330 15986 45342
rect 15934 45266 15986 45278
rect 17502 45330 17554 45342
rect 17502 45266 17554 45278
rect 22206 45330 22258 45342
rect 22206 45266 22258 45278
rect 23214 45330 23266 45342
rect 23214 45266 23266 45278
rect 23662 45330 23714 45342
rect 23662 45266 23714 45278
rect 23998 45330 24050 45342
rect 23998 45266 24050 45278
rect 7646 45218 7698 45230
rect 7646 45154 7698 45166
rect 9550 45218 9602 45230
rect 9550 45154 9602 45166
rect 13918 45218 13970 45230
rect 13918 45154 13970 45166
rect 14030 45218 14082 45230
rect 15486 45218 15538 45230
rect 14354 45166 14366 45218
rect 14418 45166 14430 45218
rect 14802 45166 14814 45218
rect 14866 45166 14878 45218
rect 14030 45154 14082 45166
rect 15486 45154 15538 45166
rect 16830 45218 16882 45230
rect 16830 45154 16882 45166
rect 22094 45218 22146 45230
rect 22094 45154 22146 45166
rect 22430 45218 22482 45230
rect 22430 45154 22482 45166
rect 22654 45218 22706 45230
rect 22654 45154 22706 45166
rect 3054 45106 3106 45118
rect 2258 45054 2270 45106
rect 2322 45054 2334 45106
rect 2818 45054 2830 45106
rect 2882 45054 2894 45106
rect 3054 45042 3106 45054
rect 3502 45106 3554 45118
rect 3502 45042 3554 45054
rect 9102 45106 9154 45118
rect 9102 45042 9154 45054
rect 9774 45106 9826 45118
rect 9774 45042 9826 45054
rect 9998 45106 10050 45118
rect 9998 45042 10050 45054
rect 10110 45106 10162 45118
rect 15262 45106 15314 45118
rect 16382 45106 16434 45118
rect 13458 45054 13470 45106
rect 13522 45054 13534 45106
rect 13682 45054 13694 45106
rect 13746 45054 13758 45106
rect 16146 45054 16158 45106
rect 16210 45054 16222 45106
rect 10110 45042 10162 45054
rect 15262 45042 15314 45054
rect 16382 45042 16434 45054
rect 16606 45106 16658 45118
rect 21186 45054 21198 45106
rect 21250 45054 21262 45106
rect 28130 45054 28142 45106
rect 28194 45054 28206 45106
rect 16606 45042 16658 45054
rect 2046 44994 2098 45006
rect 2046 44930 2098 44942
rect 3390 44994 3442 45006
rect 3390 44930 3442 44942
rect 4846 44994 4898 45006
rect 4846 44930 4898 44942
rect 6190 44994 6242 45006
rect 6190 44930 6242 44942
rect 6750 44994 6802 45006
rect 6750 44930 6802 44942
rect 7198 44994 7250 45006
rect 7198 44930 7250 44942
rect 7982 44994 8034 45006
rect 7982 44930 8034 44942
rect 8542 44994 8594 45006
rect 8542 44930 8594 44942
rect 9886 44994 9938 45006
rect 9886 44930 9938 44942
rect 11006 44994 11058 45006
rect 11006 44930 11058 44942
rect 12350 44994 12402 45006
rect 12350 44930 12402 44942
rect 13246 44994 13298 45006
rect 17950 44994 18002 45006
rect 21758 44994 21810 45006
rect 16258 44942 16270 44994
rect 16322 44942 16334 44994
rect 18386 44942 18398 44994
rect 18450 44942 18462 44994
rect 20514 44942 20526 44994
rect 20578 44942 20590 44994
rect 13246 44930 13298 44942
rect 17950 44930 18002 44942
rect 21758 44930 21810 44942
rect 24446 44994 24498 45006
rect 25218 44942 25230 44994
rect 25282 44942 25294 44994
rect 27346 44942 27358 44994
rect 27410 44942 27422 44994
rect 24446 44930 24498 44942
rect 2482 44830 2494 44882
rect 2546 44830 2558 44882
rect 6178 44830 6190 44882
rect 6242 44879 6254 44882
rect 7746 44879 7758 44882
rect 6242 44833 7758 44879
rect 6242 44830 6254 44833
rect 7746 44830 7758 44833
rect 7810 44830 7822 44882
rect 8530 44830 8542 44882
rect 8594 44879 8606 44882
rect 8866 44879 8878 44882
rect 8594 44833 8878 44879
rect 8594 44830 8606 44833
rect 8866 44830 8878 44833
rect 8930 44830 8942 44882
rect 11890 44830 11902 44882
rect 11954 44879 11966 44882
rect 12338 44879 12350 44882
rect 11954 44833 12350 44879
rect 11954 44830 11966 44833
rect 12338 44830 12350 44833
rect 12402 44879 12414 44882
rect 13234 44879 13246 44882
rect 12402 44833 13246 44879
rect 12402 44830 12414 44833
rect 13234 44830 13246 44833
rect 13298 44830 13310 44882
rect 1344 44714 28560 44748
rect 1344 44662 4616 44714
rect 4668 44662 4720 44714
rect 4772 44662 4824 44714
rect 4876 44662 11420 44714
rect 11472 44662 11524 44714
rect 11576 44662 11628 44714
rect 11680 44662 18224 44714
rect 18276 44662 18328 44714
rect 18380 44662 18432 44714
rect 18484 44662 25028 44714
rect 25080 44662 25132 44714
rect 25184 44662 25236 44714
rect 25288 44662 28560 44714
rect 1344 44628 28560 44662
rect 2258 44494 2270 44546
rect 2322 44543 2334 44546
rect 3154 44543 3166 44546
rect 2322 44497 3166 44543
rect 2322 44494 2334 44497
rect 3154 44494 3166 44497
rect 3218 44494 3230 44546
rect 6178 44494 6190 44546
rect 6242 44494 6254 44546
rect 9426 44494 9438 44546
rect 9490 44543 9502 44546
rect 9986 44543 9998 44546
rect 9490 44497 9998 44543
rect 9490 44494 9502 44497
rect 9986 44494 9998 44497
rect 10050 44494 10062 44546
rect 2494 44434 2546 44446
rect 2494 44370 2546 44382
rect 3726 44434 3778 44446
rect 9662 44434 9714 44446
rect 8418 44382 8430 44434
rect 8482 44382 8494 44434
rect 3726 44370 3778 44382
rect 9662 44370 9714 44382
rect 10110 44434 10162 44446
rect 15250 44382 15262 44434
rect 15314 44382 15326 44434
rect 26786 44382 26798 44434
rect 26850 44382 26862 44434
rect 10110 44370 10162 44382
rect 6750 44322 6802 44334
rect 6402 44270 6414 44322
rect 6466 44270 6478 44322
rect 6750 44258 6802 44270
rect 6862 44322 6914 44334
rect 10670 44322 10722 44334
rect 7746 44270 7758 44322
rect 7810 44270 7822 44322
rect 8642 44270 8654 44322
rect 8706 44270 8718 44322
rect 10434 44270 10446 44322
rect 10498 44270 10510 44322
rect 6862 44258 6914 44270
rect 10670 44258 10722 44270
rect 12238 44322 12290 44334
rect 12238 44258 12290 44270
rect 12574 44322 12626 44334
rect 12574 44258 12626 44270
rect 13470 44322 13522 44334
rect 13470 44258 13522 44270
rect 13582 44322 13634 44334
rect 14926 44322 14978 44334
rect 17502 44322 17554 44334
rect 20190 44322 20242 44334
rect 14690 44270 14702 44322
rect 14754 44270 14766 44322
rect 15362 44270 15374 44322
rect 15426 44270 15438 44322
rect 19618 44270 19630 44322
rect 19682 44270 19694 44322
rect 13582 44258 13634 44270
rect 14926 44258 14978 44270
rect 17502 44258 17554 44270
rect 20190 44258 20242 44270
rect 20414 44322 20466 44334
rect 20414 44258 20466 44270
rect 21422 44322 21474 44334
rect 23762 44270 23774 44322
rect 23826 44270 23838 44322
rect 21422 44258 21474 44270
rect 3390 44210 3442 44222
rect 3390 44146 3442 44158
rect 4510 44210 4562 44222
rect 4510 44146 4562 44158
rect 5630 44210 5682 44222
rect 8990 44210 9042 44222
rect 5842 44158 5854 44210
rect 5906 44158 5918 44210
rect 7858 44158 7870 44210
rect 7922 44158 7934 44210
rect 5630 44146 5682 44158
rect 8990 44146 9042 44158
rect 12014 44210 12066 44222
rect 19966 44210 20018 44222
rect 15810 44158 15822 44210
rect 15874 44158 15886 44210
rect 19506 44158 19518 44210
rect 19570 44158 19582 44210
rect 12014 44146 12066 44158
rect 19966 44146 20018 44158
rect 21198 44210 21250 44222
rect 21746 44158 21758 44210
rect 21810 44158 21822 44210
rect 22306 44158 22318 44210
rect 22370 44158 22382 44210
rect 21198 44146 21250 44158
rect 2158 44098 2210 44110
rect 2158 44034 2210 44046
rect 3054 44098 3106 44110
rect 3054 44034 3106 44046
rect 3838 44098 3890 44110
rect 3838 44034 3890 44046
rect 4398 44098 4450 44110
rect 4398 44034 4450 44046
rect 5182 44098 5234 44110
rect 5182 44034 5234 44046
rect 5742 44098 5794 44110
rect 5742 44034 5794 44046
rect 6974 44098 7026 44110
rect 6974 44034 7026 44046
rect 10782 44098 10834 44110
rect 10782 44034 10834 44046
rect 10894 44098 10946 44110
rect 10894 44034 10946 44046
rect 11006 44098 11058 44110
rect 11006 44034 11058 44046
rect 11790 44098 11842 44110
rect 11790 44034 11842 44046
rect 12126 44098 12178 44110
rect 12126 44034 12178 44046
rect 13694 44098 13746 44110
rect 13694 44034 13746 44046
rect 13918 44098 13970 44110
rect 13918 44034 13970 44046
rect 15150 44098 15202 44110
rect 20190 44098 20242 44110
rect 16034 44046 16046 44098
rect 16098 44046 16110 44098
rect 15150 44034 15202 44046
rect 20190 44034 20242 44046
rect 1344 43930 28720 43964
rect 1344 43878 8018 43930
rect 8070 43878 8122 43930
rect 8174 43878 8226 43930
rect 8278 43878 14822 43930
rect 14874 43878 14926 43930
rect 14978 43878 15030 43930
rect 15082 43878 21626 43930
rect 21678 43878 21730 43930
rect 21782 43878 21834 43930
rect 21886 43878 28430 43930
rect 28482 43878 28534 43930
rect 28586 43878 28638 43930
rect 28690 43878 28720 43930
rect 1344 43844 28720 43878
rect 2158 43762 2210 43774
rect 2158 43698 2210 43710
rect 19182 43762 19234 43774
rect 19182 43698 19234 43710
rect 20190 43762 20242 43774
rect 20190 43698 20242 43710
rect 22094 43762 22146 43774
rect 22094 43698 22146 43710
rect 23438 43762 23490 43774
rect 23438 43698 23490 43710
rect 25790 43762 25842 43774
rect 25790 43698 25842 43710
rect 26462 43762 26514 43774
rect 26462 43698 26514 43710
rect 2494 43650 2546 43662
rect 11006 43650 11058 43662
rect 17614 43650 17666 43662
rect 19406 43650 19458 43662
rect 5394 43598 5406 43650
rect 5458 43598 5470 43650
rect 10098 43598 10110 43650
rect 10162 43598 10174 43650
rect 10434 43598 10446 43650
rect 10498 43598 10510 43650
rect 12114 43598 12126 43650
rect 12178 43598 12190 43650
rect 18834 43598 18846 43650
rect 18898 43598 18910 43650
rect 2494 43586 2546 43598
rect 11006 43586 11058 43598
rect 17614 43586 17666 43598
rect 19406 43586 19458 43598
rect 21310 43650 21362 43662
rect 21310 43586 21362 43598
rect 23102 43650 23154 43662
rect 23102 43586 23154 43598
rect 27358 43650 27410 43662
rect 27358 43586 27410 43598
rect 28142 43650 28194 43662
rect 28142 43586 28194 43598
rect 10782 43538 10834 43550
rect 15038 43538 15090 43550
rect 2818 43486 2830 43538
rect 2882 43486 2894 43538
rect 4834 43486 4846 43538
rect 4898 43486 4910 43538
rect 11330 43486 11342 43538
rect 11394 43486 11406 43538
rect 10782 43474 10834 43486
rect 15038 43474 15090 43486
rect 15598 43538 15650 43550
rect 15598 43474 15650 43486
rect 15934 43538 15986 43550
rect 15934 43474 15986 43486
rect 16158 43538 16210 43550
rect 19294 43538 19346 43550
rect 23998 43538 24050 43550
rect 16818 43486 16830 43538
rect 16882 43486 16894 43538
rect 17826 43486 17838 43538
rect 17890 43486 17902 43538
rect 18498 43486 18510 43538
rect 18562 43486 18574 43538
rect 19730 43486 19742 43538
rect 19794 43486 19806 43538
rect 16158 43474 16210 43486
rect 19294 43474 19346 43486
rect 23998 43474 24050 43486
rect 24222 43538 24274 43550
rect 26238 43538 26290 43550
rect 24546 43486 24558 43538
rect 24610 43486 24622 43538
rect 24222 43474 24274 43486
rect 26238 43474 26290 43486
rect 26574 43538 26626 43550
rect 26574 43474 26626 43486
rect 26798 43538 26850 43550
rect 26798 43474 26850 43486
rect 27134 43538 27186 43550
rect 27134 43474 27186 43486
rect 27246 43538 27298 43550
rect 27246 43474 27298 43486
rect 27806 43538 27858 43550
rect 27806 43474 27858 43486
rect 2606 43426 2658 43438
rect 2606 43362 2658 43374
rect 9662 43426 9714 43438
rect 9662 43362 9714 43374
rect 9998 43426 10050 43438
rect 15710 43426 15762 43438
rect 14242 43374 14254 43426
rect 14306 43374 14318 43426
rect 9998 43362 10050 43374
rect 15710 43362 15762 43374
rect 16606 43426 16658 43438
rect 20638 43426 20690 43438
rect 18162 43374 18174 43426
rect 18226 43374 18238 43426
rect 16606 43362 16658 43374
rect 20638 43362 20690 43374
rect 21646 43426 21698 43438
rect 21646 43362 21698 43374
rect 22542 43426 22594 43438
rect 22542 43362 22594 43374
rect 24110 43426 24162 43438
rect 24110 43362 24162 43374
rect 16494 43314 16546 43326
rect 25566 43314 25618 43326
rect 19954 43262 19966 43314
rect 20018 43311 20030 43314
rect 20850 43311 20862 43314
rect 20018 43265 20862 43311
rect 20018 43262 20030 43265
rect 20850 43262 20862 43265
rect 20914 43262 20926 43314
rect 22306 43262 22318 43314
rect 22370 43311 22382 43314
rect 23426 43311 23438 43314
rect 22370 43265 23438 43311
rect 22370 43262 22382 43265
rect 23426 43262 23438 43265
rect 23490 43262 23502 43314
rect 16494 43250 16546 43262
rect 25566 43250 25618 43262
rect 25902 43314 25954 43326
rect 25902 43250 25954 43262
rect 1344 43146 28560 43180
rect 1344 43094 4616 43146
rect 4668 43094 4720 43146
rect 4772 43094 4824 43146
rect 4876 43094 11420 43146
rect 11472 43094 11524 43146
rect 11576 43094 11628 43146
rect 11680 43094 18224 43146
rect 18276 43094 18328 43146
rect 18380 43094 18432 43146
rect 18484 43094 25028 43146
rect 25080 43094 25132 43146
rect 25184 43094 25236 43146
rect 25288 43094 28560 43146
rect 1344 43060 28560 43094
rect 19294 42978 19346 42990
rect 19294 42914 19346 42926
rect 5070 42866 5122 42878
rect 4610 42814 4622 42866
rect 4674 42814 4686 42866
rect 5070 42802 5122 42814
rect 6078 42866 6130 42878
rect 10782 42866 10834 42878
rect 7186 42814 7198 42866
rect 7250 42814 7262 42866
rect 9314 42814 9326 42866
rect 9378 42814 9390 42866
rect 6078 42802 6130 42814
rect 10782 42802 10834 42814
rect 12014 42866 12066 42878
rect 12014 42802 12066 42814
rect 12910 42866 12962 42878
rect 12910 42802 12962 42814
rect 13918 42866 13970 42878
rect 18622 42866 18674 42878
rect 27918 42866 27970 42878
rect 15810 42814 15822 42866
rect 15874 42814 15886 42866
rect 17938 42814 17950 42866
rect 18002 42814 18014 42866
rect 21298 42814 21310 42866
rect 21362 42814 21374 42866
rect 24546 42814 24558 42866
rect 24610 42814 24622 42866
rect 13918 42802 13970 42814
rect 18622 42802 18674 42814
rect 27918 42802 27970 42814
rect 19518 42754 19570 42766
rect 1810 42702 1822 42754
rect 1874 42702 1886 42754
rect 6514 42702 6526 42754
rect 6578 42702 6590 42754
rect 9650 42702 9662 42754
rect 9714 42702 9726 42754
rect 15138 42702 15150 42754
rect 15202 42702 15214 42754
rect 19518 42690 19570 42702
rect 20078 42754 20130 42766
rect 20078 42690 20130 42702
rect 20302 42754 20354 42766
rect 20302 42690 20354 42702
rect 20750 42754 20802 42766
rect 24098 42702 24110 42754
rect 24162 42702 24174 42754
rect 27458 42702 27470 42754
rect 27522 42702 27534 42754
rect 20750 42690 20802 42702
rect 9998 42642 10050 42654
rect 2482 42590 2494 42642
rect 2546 42590 2558 42642
rect 9998 42578 10050 42590
rect 10446 42642 10498 42654
rect 10446 42578 10498 42590
rect 14590 42642 14642 42654
rect 14590 42578 14642 42590
rect 18286 42642 18338 42654
rect 18286 42578 18338 42590
rect 18846 42642 18898 42654
rect 18846 42578 18898 42590
rect 19966 42642 20018 42654
rect 23426 42590 23438 42642
rect 23490 42590 23502 42642
rect 26674 42590 26686 42642
rect 26738 42590 26750 42642
rect 19966 42578 20018 42590
rect 9886 42530 9938 42542
rect 9886 42466 9938 42478
rect 10670 42530 10722 42542
rect 10670 42466 10722 42478
rect 10894 42530 10946 42542
rect 10894 42466 10946 42478
rect 11006 42530 11058 42542
rect 11006 42466 11058 42478
rect 11566 42530 11618 42542
rect 11566 42466 11618 42478
rect 12462 42530 12514 42542
rect 12462 42466 12514 42478
rect 14142 42530 14194 42542
rect 14142 42466 14194 42478
rect 14254 42530 14306 42542
rect 14254 42466 14306 42478
rect 14366 42530 14418 42542
rect 14366 42466 14418 42478
rect 18510 42530 18562 42542
rect 18510 42466 18562 42478
rect 18734 42530 18786 42542
rect 18734 42466 18786 42478
rect 1344 42362 28720 42396
rect 1344 42310 8018 42362
rect 8070 42310 8122 42362
rect 8174 42310 8226 42362
rect 8278 42310 14822 42362
rect 14874 42310 14926 42362
rect 14978 42310 15030 42362
rect 15082 42310 21626 42362
rect 21678 42310 21730 42362
rect 21782 42310 21834 42362
rect 21886 42310 28430 42362
rect 28482 42310 28534 42362
rect 28586 42310 28638 42362
rect 28690 42310 28720 42362
rect 1344 42276 28720 42310
rect 2494 42194 2546 42206
rect 2494 42130 2546 42142
rect 8542 42194 8594 42206
rect 8542 42130 8594 42142
rect 11230 42194 11282 42206
rect 11230 42130 11282 42142
rect 19182 42194 19234 42206
rect 19182 42130 19234 42142
rect 21870 42194 21922 42206
rect 21870 42130 21922 42142
rect 23102 42194 23154 42206
rect 23102 42130 23154 42142
rect 23886 42194 23938 42206
rect 23886 42130 23938 42142
rect 2046 42082 2098 42094
rect 3278 42082 3330 42094
rect 3042 42030 3054 42082
rect 3106 42030 3118 42082
rect 2046 42018 2098 42030
rect 3278 42018 3330 42030
rect 10558 42082 10610 42094
rect 10558 42018 10610 42030
rect 11678 42082 11730 42094
rect 11678 42018 11730 42030
rect 15710 42082 15762 42094
rect 15710 42018 15762 42030
rect 19294 42082 19346 42094
rect 19294 42018 19346 42030
rect 19406 42082 19458 42094
rect 19406 42018 19458 42030
rect 22542 42082 22594 42094
rect 22542 42018 22594 42030
rect 24222 42082 24274 42094
rect 24222 42018 24274 42030
rect 1710 41970 1762 41982
rect 3726 41970 3778 41982
rect 7758 41970 7810 41982
rect 2706 41918 2718 41970
rect 2770 41918 2782 41970
rect 4162 41918 4174 41970
rect 4226 41918 4238 41970
rect 4834 41918 4846 41970
rect 4898 41918 4910 41970
rect 1710 41906 1762 41918
rect 3726 41906 3778 41918
rect 7758 41906 7810 41918
rect 8094 41970 8146 41982
rect 8094 41906 8146 41918
rect 8206 41970 8258 41982
rect 8990 41970 9042 41982
rect 8530 41918 8542 41970
rect 8594 41918 8606 41970
rect 8206 41906 8258 41918
rect 8990 41906 9042 41918
rect 10222 41970 10274 41982
rect 10222 41906 10274 41918
rect 10334 41970 10386 41982
rect 10334 41906 10386 41918
rect 10782 41970 10834 41982
rect 17502 41970 17554 41982
rect 12338 41918 12350 41970
rect 12402 41918 12414 41970
rect 15922 41918 15934 41970
rect 15986 41918 15998 41970
rect 16482 41918 16494 41970
rect 16546 41918 16558 41970
rect 10782 41906 10834 41918
rect 17502 41906 17554 41918
rect 17614 41970 17666 41982
rect 17614 41906 17666 41918
rect 17726 41970 17778 41982
rect 17726 41906 17778 41918
rect 18174 41970 18226 41982
rect 18174 41906 18226 41918
rect 18398 41970 18450 41982
rect 18398 41906 18450 41918
rect 19070 41970 19122 41982
rect 20078 41970 20130 41982
rect 19618 41918 19630 41970
rect 19682 41918 19694 41970
rect 19070 41906 19122 41918
rect 20078 41906 20130 41918
rect 20190 41970 20242 41982
rect 20190 41906 20242 41918
rect 20302 41970 20354 41982
rect 20302 41906 20354 41918
rect 20414 41970 20466 41982
rect 21086 41970 21138 41982
rect 23550 41970 23602 41982
rect 20626 41918 20638 41970
rect 20690 41918 20702 41970
rect 21298 41918 21310 41970
rect 21362 41918 21374 41970
rect 21858 41918 21870 41970
rect 21922 41918 21934 41970
rect 22194 41918 22206 41970
rect 22258 41918 22270 41970
rect 20414 41906 20466 41918
rect 21086 41906 21138 41918
rect 23550 41906 23602 41918
rect 23998 41970 24050 41982
rect 23998 41906 24050 41918
rect 24670 41970 24722 41982
rect 28018 41918 28030 41970
rect 28082 41918 28094 41970
rect 24670 41906 24722 41918
rect 7534 41858 7586 41870
rect 6962 41806 6974 41858
rect 7026 41806 7038 41858
rect 7534 41794 7586 41806
rect 9886 41858 9938 41870
rect 15822 41858 15874 41870
rect 13010 41806 13022 41858
rect 13074 41806 13086 41858
rect 15138 41806 15150 41858
rect 15202 41806 15214 41858
rect 25218 41806 25230 41858
rect 25282 41806 25294 41858
rect 27346 41806 27358 41858
rect 27410 41806 27422 41858
rect 9886 41794 9938 41806
rect 15822 41794 15874 41806
rect 22206 41746 22258 41758
rect 2706 41694 2718 41746
rect 2770 41694 2782 41746
rect 16258 41694 16270 41746
rect 16322 41694 16334 41746
rect 21634 41694 21646 41746
rect 21698 41694 21710 41746
rect 22866 41694 22878 41746
rect 22930 41743 22942 41746
rect 23314 41743 23326 41746
rect 22930 41697 23326 41743
rect 22930 41694 22942 41697
rect 23314 41694 23326 41697
rect 23378 41694 23390 41746
rect 22206 41682 22258 41694
rect 1344 41578 28560 41612
rect 1344 41526 4616 41578
rect 4668 41526 4720 41578
rect 4772 41526 4824 41578
rect 4876 41526 11420 41578
rect 11472 41526 11524 41578
rect 11576 41526 11628 41578
rect 11680 41526 18224 41578
rect 18276 41526 18328 41578
rect 18380 41526 18432 41578
rect 18484 41526 25028 41578
rect 25080 41526 25132 41578
rect 25184 41526 25236 41578
rect 25288 41526 28560 41578
rect 1344 41492 28560 41526
rect 2718 41410 2770 41422
rect 2718 41346 2770 41358
rect 3054 41410 3106 41422
rect 3266 41358 3278 41410
rect 3330 41407 3342 41410
rect 3938 41407 3950 41410
rect 3330 41361 3950 41407
rect 3330 41358 3342 41361
rect 3938 41358 3950 41361
rect 4002 41358 4014 41410
rect 22418 41358 22430 41410
rect 22482 41407 22494 41410
rect 22754 41407 22766 41410
rect 22482 41361 22766 41407
rect 22482 41358 22494 41361
rect 22754 41358 22766 41361
rect 22818 41358 22830 41410
rect 26338 41358 26350 41410
rect 26402 41358 26414 41410
rect 3054 41346 3106 41358
rect 3950 41298 4002 41310
rect 3950 41234 4002 41246
rect 4846 41298 4898 41310
rect 11790 41298 11842 41310
rect 10546 41246 10558 41298
rect 10610 41246 10622 41298
rect 4846 41234 4898 41246
rect 11790 41234 11842 41246
rect 14590 41298 14642 41310
rect 19518 41298 19570 41310
rect 15586 41246 15598 41298
rect 15650 41246 15662 41298
rect 17714 41246 17726 41298
rect 17778 41246 17790 41298
rect 14590 41234 14642 41246
rect 19518 41234 19570 41246
rect 20414 41298 20466 41310
rect 20414 41234 20466 41246
rect 21422 41298 21474 41310
rect 21422 41234 21474 41246
rect 22766 41298 22818 41310
rect 22766 41234 22818 41246
rect 23998 41298 24050 41310
rect 23998 41234 24050 41246
rect 24670 41298 24722 41310
rect 24670 41234 24722 41246
rect 25118 41298 25170 41310
rect 25118 41234 25170 41246
rect 27358 41298 27410 41310
rect 27358 41234 27410 41246
rect 28030 41298 28082 41310
rect 28030 41234 28082 41246
rect 5854 41186 5906 41198
rect 5854 41122 5906 41134
rect 6862 41186 6914 41198
rect 13582 41186 13634 41198
rect 7634 41134 7646 41186
rect 7698 41134 7710 41186
rect 6862 41122 6914 41134
rect 13582 41122 13634 41134
rect 14030 41186 14082 41198
rect 18846 41186 18898 41198
rect 14802 41134 14814 41186
rect 14866 41134 14878 41186
rect 14030 41122 14082 41134
rect 18846 41122 18898 41134
rect 19406 41186 19458 41198
rect 19954 41134 19966 41186
rect 20018 41134 20030 41186
rect 26338 41134 26350 41186
rect 26402 41134 26414 41186
rect 26674 41134 26686 41186
rect 26738 41134 26750 41186
rect 19406 41122 19458 41134
rect 6302 41074 6354 41086
rect 12238 41074 12290 41086
rect 8418 41022 8430 41074
rect 8482 41022 8494 41074
rect 6302 41010 6354 41022
rect 12238 41010 12290 41022
rect 13470 41074 13522 41086
rect 13470 41010 13522 41022
rect 13806 41074 13858 41086
rect 13806 41010 13858 41022
rect 18286 41074 18338 41086
rect 18286 41010 18338 41022
rect 18622 41074 18674 41086
rect 18622 41010 18674 41022
rect 26910 41074 26962 41086
rect 26910 41010 26962 41022
rect 2046 40962 2098 40974
rect 2046 40898 2098 40910
rect 2382 40962 2434 40974
rect 2382 40898 2434 40910
rect 2830 40962 2882 40974
rect 2830 40898 2882 40910
rect 3502 40962 3554 40974
rect 3502 40898 3554 40910
rect 4398 40962 4450 40974
rect 4398 40898 4450 40910
rect 6190 40962 6242 40974
rect 6190 40898 6242 40910
rect 7310 40962 7362 40974
rect 7310 40898 7362 40910
rect 11342 40962 11394 40974
rect 11342 40898 11394 40910
rect 12798 40962 12850 40974
rect 12798 40898 12850 40910
rect 18510 40962 18562 40974
rect 18510 40898 18562 40910
rect 19630 40962 19682 40974
rect 19630 40898 19682 40910
rect 21870 40962 21922 40974
rect 21870 40898 21922 40910
rect 22318 40962 22370 40974
rect 22318 40898 22370 40910
rect 23550 40962 23602 40974
rect 23550 40898 23602 40910
rect 25790 40962 25842 40974
rect 25790 40898 25842 40910
rect 26798 40962 26850 40974
rect 26798 40898 26850 40910
rect 1344 40794 28720 40828
rect 1344 40742 8018 40794
rect 8070 40742 8122 40794
rect 8174 40742 8226 40794
rect 8278 40742 14822 40794
rect 14874 40742 14926 40794
rect 14978 40742 15030 40794
rect 15082 40742 21626 40794
rect 21678 40742 21730 40794
rect 21782 40742 21834 40794
rect 21886 40742 28430 40794
rect 28482 40742 28534 40794
rect 28586 40742 28638 40794
rect 28690 40742 28720 40794
rect 1344 40708 28720 40742
rect 10334 40626 10386 40638
rect 2706 40574 2718 40626
rect 2770 40574 2782 40626
rect 8418 40574 8430 40626
rect 8482 40574 8494 40626
rect 10334 40562 10386 40574
rect 10782 40626 10834 40638
rect 13246 40626 13298 40638
rect 11554 40574 11566 40626
rect 11618 40574 11630 40626
rect 10782 40562 10834 40574
rect 13246 40562 13298 40574
rect 13582 40626 13634 40638
rect 13582 40562 13634 40574
rect 14030 40626 14082 40638
rect 14030 40562 14082 40574
rect 15150 40626 15202 40638
rect 15150 40562 15202 40574
rect 15598 40626 15650 40638
rect 15598 40562 15650 40574
rect 16046 40626 16098 40638
rect 16046 40562 16098 40574
rect 16718 40626 16770 40638
rect 16718 40562 16770 40574
rect 21086 40626 21138 40638
rect 21086 40562 21138 40574
rect 21534 40626 21586 40638
rect 21534 40562 21586 40574
rect 22430 40626 22482 40638
rect 22430 40562 22482 40574
rect 22878 40626 22930 40638
rect 22878 40562 22930 40574
rect 23326 40626 23378 40638
rect 23326 40562 23378 40574
rect 23886 40626 23938 40638
rect 23886 40562 23938 40574
rect 25342 40626 25394 40638
rect 25342 40562 25394 40574
rect 27470 40626 27522 40638
rect 27470 40562 27522 40574
rect 28142 40626 28194 40638
rect 28142 40562 28194 40574
rect 2046 40514 2098 40526
rect 2046 40450 2098 40462
rect 3166 40514 3218 40526
rect 3166 40450 3218 40462
rect 8206 40514 8258 40526
rect 8206 40450 8258 40462
rect 11118 40514 11170 40526
rect 21982 40514 22034 40526
rect 18498 40462 18510 40514
rect 18562 40462 18574 40514
rect 11118 40450 11170 40462
rect 21982 40450 22034 40462
rect 24110 40514 24162 40526
rect 24110 40450 24162 40462
rect 26350 40514 26402 40526
rect 26350 40450 26402 40462
rect 1710 40402 1762 40414
rect 24334 40402 24386 40414
rect 25790 40402 25842 40414
rect 2482 40350 2494 40402
rect 2546 40350 2558 40402
rect 2930 40350 2942 40402
rect 2994 40350 3006 40402
rect 3602 40350 3614 40402
rect 3666 40350 3678 40402
rect 4274 40350 4286 40402
rect 4338 40350 4350 40402
rect 8418 40350 8430 40402
rect 8482 40350 8494 40402
rect 8978 40350 8990 40402
rect 9042 40350 9054 40402
rect 9874 40350 9886 40402
rect 9938 40350 9950 40402
rect 11330 40350 11342 40402
rect 11394 40350 11406 40402
rect 11778 40350 11790 40402
rect 11842 40350 11854 40402
rect 12562 40350 12574 40402
rect 12626 40350 12638 40402
rect 17714 40350 17726 40402
rect 17778 40350 17790 40402
rect 24658 40350 24670 40402
rect 24722 40350 24734 40402
rect 1710 40338 1762 40350
rect 24334 40338 24386 40350
rect 25790 40338 25842 40350
rect 26798 40402 26850 40414
rect 26798 40338 26850 40350
rect 7870 40290 7922 40302
rect 5058 40238 5070 40290
rect 5122 40238 5134 40290
rect 7186 40238 7198 40290
rect 7250 40238 7262 40290
rect 7870 40226 7922 40238
rect 9550 40290 9602 40302
rect 9550 40226 9602 40238
rect 9662 40290 9714 40302
rect 9662 40226 9714 40238
rect 12238 40290 12290 40302
rect 12238 40226 12290 40238
rect 12350 40290 12402 40302
rect 12350 40226 12402 40238
rect 14478 40290 14530 40302
rect 24222 40290 24274 40302
rect 20626 40238 20638 40290
rect 20690 40238 20702 40290
rect 14478 40226 14530 40238
rect 24222 40226 24274 40238
rect 3726 40178 3778 40190
rect 2594 40126 2606 40178
rect 2658 40126 2670 40178
rect 8754 40126 8766 40178
rect 8818 40126 8830 40178
rect 11666 40126 11678 40178
rect 11730 40126 11742 40178
rect 3726 40114 3778 40126
rect 1344 40010 28560 40044
rect 1344 39958 4616 40010
rect 4668 39958 4720 40010
rect 4772 39958 4824 40010
rect 4876 39958 11420 40010
rect 11472 39958 11524 40010
rect 11576 39958 11628 40010
rect 11680 39958 18224 40010
rect 18276 39958 18328 40010
rect 18380 39958 18432 40010
rect 18484 39958 25028 40010
rect 25080 39958 25132 40010
rect 25184 39958 25236 40010
rect 25288 39958 28560 40010
rect 1344 39924 28560 39958
rect 5966 39842 6018 39854
rect 27358 39842 27410 39854
rect 7298 39790 7310 39842
rect 7362 39839 7374 39842
rect 7858 39839 7870 39842
rect 7362 39793 7870 39839
rect 7362 39790 7374 39793
rect 7858 39790 7870 39793
rect 7922 39790 7934 39842
rect 8754 39790 8766 39842
rect 8818 39839 8830 39842
rect 9650 39839 9662 39842
rect 8818 39793 9662 39839
rect 8818 39790 8830 39793
rect 9650 39790 9662 39793
rect 9714 39790 9726 39842
rect 13570 39790 13582 39842
rect 13634 39839 13646 39842
rect 14466 39839 14478 39842
rect 13634 39793 14478 39839
rect 13634 39790 13646 39793
rect 14466 39790 14478 39793
rect 14530 39790 14542 39842
rect 17826 39790 17838 39842
rect 17890 39839 17902 39842
rect 18722 39839 18734 39842
rect 17890 39793 18734 39839
rect 17890 39790 17902 39793
rect 18722 39790 18734 39793
rect 18786 39790 18798 39842
rect 19394 39790 19406 39842
rect 19458 39839 19470 39842
rect 19618 39839 19630 39842
rect 19458 39793 19630 39839
rect 19458 39790 19470 39793
rect 19618 39790 19630 39793
rect 19682 39790 19694 39842
rect 26786 39790 26798 39842
rect 26850 39790 26862 39842
rect 5966 39778 6018 39790
rect 27358 39778 27410 39790
rect 27694 39842 27746 39854
rect 27694 39778 27746 39790
rect 5070 39730 5122 39742
rect 2482 39678 2494 39730
rect 2546 39678 2558 39730
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 5070 39666 5122 39678
rect 7198 39730 7250 39742
rect 7198 39666 7250 39678
rect 8094 39730 8146 39742
rect 8094 39666 8146 39678
rect 8542 39730 8594 39742
rect 8542 39666 8594 39678
rect 8990 39730 9042 39742
rect 16046 39730 16098 39742
rect 10770 39678 10782 39730
rect 10834 39678 10846 39730
rect 12898 39678 12910 39730
rect 12962 39678 12974 39730
rect 8990 39666 9042 39678
rect 16046 39666 16098 39678
rect 16382 39730 16434 39742
rect 16382 39666 16434 39678
rect 19406 39730 19458 39742
rect 19406 39666 19458 39678
rect 20414 39730 20466 39742
rect 20414 39666 20466 39678
rect 22654 39730 22706 39742
rect 28142 39730 28194 39742
rect 22978 39678 22990 39730
rect 23042 39678 23054 39730
rect 22654 39666 22706 39678
rect 28142 39666 28194 39678
rect 6414 39618 6466 39630
rect 14142 39618 14194 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 5618 39566 5630 39618
rect 5682 39566 5694 39618
rect 6178 39566 6190 39618
rect 6242 39566 6254 39618
rect 9986 39566 9998 39618
rect 10050 39566 10062 39618
rect 6414 39554 6466 39566
rect 14142 39554 14194 39566
rect 15150 39618 15202 39630
rect 26238 39618 26290 39630
rect 25890 39566 25902 39618
rect 25954 39566 25966 39618
rect 26450 39566 26462 39618
rect 26514 39566 26526 39618
rect 26898 39566 26910 39618
rect 26962 39566 26974 39618
rect 15150 39554 15202 39566
rect 26238 39554 26290 39566
rect 14590 39506 14642 39518
rect 14590 39442 14642 39454
rect 14926 39506 14978 39518
rect 14926 39442 14978 39454
rect 15486 39506 15538 39518
rect 25106 39454 25118 39506
rect 25170 39454 25182 39506
rect 15486 39442 15538 39454
rect 5630 39394 5682 39406
rect 5630 39330 5682 39342
rect 7758 39394 7810 39406
rect 7758 39330 7810 39342
rect 9550 39394 9602 39406
rect 9550 39330 9602 39342
rect 13582 39394 13634 39406
rect 13582 39330 13634 39342
rect 15150 39394 15202 39406
rect 15150 39330 15202 39342
rect 16942 39394 16994 39406
rect 16942 39330 16994 39342
rect 17838 39394 17890 39406
rect 17838 39330 17890 39342
rect 18174 39394 18226 39406
rect 18174 39330 18226 39342
rect 18622 39394 18674 39406
rect 18622 39330 18674 39342
rect 19854 39394 19906 39406
rect 19854 39330 19906 39342
rect 20750 39394 20802 39406
rect 20750 39330 20802 39342
rect 21422 39394 21474 39406
rect 21422 39330 21474 39342
rect 21870 39394 21922 39406
rect 21870 39330 21922 39342
rect 27022 39394 27074 39406
rect 27022 39330 27074 39342
rect 27470 39394 27522 39406
rect 27470 39330 27522 39342
rect 1344 39226 28720 39260
rect 1344 39174 8018 39226
rect 8070 39174 8122 39226
rect 8174 39174 8226 39226
rect 8278 39174 14822 39226
rect 14874 39174 14926 39226
rect 14978 39174 15030 39226
rect 15082 39174 21626 39226
rect 21678 39174 21730 39226
rect 21782 39174 21834 39226
rect 21886 39174 28430 39226
rect 28482 39174 28534 39226
rect 28586 39174 28638 39226
rect 28690 39174 28720 39226
rect 1344 39140 28720 39174
rect 2270 39058 2322 39070
rect 2270 38994 2322 39006
rect 3390 39058 3442 39070
rect 3390 38994 3442 39006
rect 3950 39058 4002 39070
rect 3950 38994 4002 39006
rect 4398 39058 4450 39070
rect 4398 38994 4450 39006
rect 5518 39058 5570 39070
rect 5518 38994 5570 39006
rect 10110 39058 10162 39070
rect 10110 38994 10162 39006
rect 10894 39058 10946 39070
rect 10894 38994 10946 39006
rect 11342 39058 11394 39070
rect 11342 38994 11394 39006
rect 12798 39058 12850 39070
rect 12798 38994 12850 39006
rect 19630 39058 19682 39070
rect 19630 38994 19682 39006
rect 19966 39058 20018 39070
rect 19966 38994 20018 39006
rect 23998 39058 24050 39070
rect 23998 38994 24050 39006
rect 3502 38946 3554 38958
rect 3502 38882 3554 38894
rect 5070 38946 5122 38958
rect 18062 38946 18114 38958
rect 14690 38894 14702 38946
rect 14754 38894 14766 38946
rect 5070 38882 5122 38894
rect 18062 38882 18114 38894
rect 18846 38946 18898 38958
rect 18846 38882 18898 38894
rect 19854 38946 19906 38958
rect 19854 38882 19906 38894
rect 24110 38946 24162 38958
rect 24110 38882 24162 38894
rect 24334 38946 24386 38958
rect 27346 38894 27358 38946
rect 27410 38894 27422 38946
rect 24334 38882 24386 38894
rect 1822 38834 1874 38846
rect 1822 38770 1874 38782
rect 12350 38834 12402 38846
rect 18734 38834 18786 38846
rect 19742 38834 19794 38846
rect 23662 38834 23714 38846
rect 14018 38782 14030 38834
rect 14082 38782 14094 38834
rect 18498 38782 18510 38834
rect 18562 38782 18574 38834
rect 19394 38782 19406 38834
rect 19458 38782 19470 38834
rect 20626 38782 20638 38834
rect 20690 38782 20702 38834
rect 28018 38782 28030 38834
rect 28082 38782 28094 38834
rect 12350 38770 12402 38782
rect 18734 38770 18786 38782
rect 19742 38770 19794 38782
rect 23662 38770 23714 38782
rect 11678 38722 11730 38734
rect 17502 38722 17554 38734
rect 16818 38670 16830 38722
rect 16882 38670 16894 38722
rect 11678 38658 11730 38670
rect 17502 38658 17554 38670
rect 19070 38722 19122 38734
rect 21298 38670 21310 38722
rect 21362 38670 21374 38722
rect 23426 38670 23438 38722
rect 23490 38670 23502 38722
rect 25218 38670 25230 38722
rect 25282 38670 25294 38722
rect 19070 38658 19122 38670
rect 1344 38442 28560 38476
rect 1344 38390 4616 38442
rect 4668 38390 4720 38442
rect 4772 38390 4824 38442
rect 4876 38390 11420 38442
rect 11472 38390 11524 38442
rect 11576 38390 11628 38442
rect 11680 38390 18224 38442
rect 18276 38390 18328 38442
rect 18380 38390 18432 38442
rect 18484 38390 25028 38442
rect 25080 38390 25132 38442
rect 25184 38390 25236 38442
rect 25288 38390 28560 38442
rect 1344 38356 28560 38390
rect 2370 38222 2382 38274
rect 2434 38222 2446 38274
rect 11778 38222 11790 38274
rect 11842 38271 11854 38274
rect 12114 38271 12126 38274
rect 11842 38225 12126 38271
rect 11842 38222 11854 38225
rect 12114 38222 12126 38225
rect 12178 38222 12190 38274
rect 13682 38222 13694 38274
rect 13746 38271 13758 38274
rect 14018 38271 14030 38274
rect 13746 38225 14030 38271
rect 13746 38222 13758 38225
rect 14018 38222 14030 38225
rect 14082 38222 14094 38274
rect 21970 38222 21982 38274
rect 22034 38222 22046 38274
rect 23538 38222 23550 38274
rect 23602 38271 23614 38274
rect 24098 38271 24110 38274
rect 23602 38225 24110 38271
rect 23602 38222 23614 38225
rect 24098 38222 24110 38225
rect 24162 38222 24174 38274
rect 26450 38222 26462 38274
rect 26514 38271 26526 38274
rect 27234 38271 27246 38274
rect 26514 38225 27246 38271
rect 26514 38222 26526 38225
rect 27234 38222 27246 38225
rect 27298 38222 27310 38274
rect 11790 38162 11842 38174
rect 9090 38110 9102 38162
rect 9154 38110 9166 38162
rect 11790 38098 11842 38110
rect 13582 38162 13634 38174
rect 20190 38162 20242 38174
rect 16482 38110 16494 38162
rect 16546 38110 16558 38162
rect 13582 38098 13634 38110
rect 20190 38098 20242 38110
rect 20750 38162 20802 38174
rect 20750 38098 20802 38110
rect 21534 38162 21586 38174
rect 21534 38098 21586 38110
rect 24110 38162 24162 38174
rect 24110 38098 24162 38110
rect 25230 38162 25282 38174
rect 25230 38098 25282 38110
rect 25678 38162 25730 38174
rect 25678 38098 25730 38110
rect 27022 38162 27074 38174
rect 27022 38098 27074 38110
rect 27470 38162 27522 38174
rect 27470 38098 27522 38110
rect 3390 38050 3442 38062
rect 10558 38050 10610 38062
rect 21758 38050 21810 38062
rect 22766 38050 22818 38062
rect 2370 37998 2382 38050
rect 2434 37998 2446 38050
rect 6178 37998 6190 38050
rect 6242 37998 6254 38050
rect 10098 37998 10110 38050
rect 10162 37998 10174 38050
rect 10770 37998 10782 38050
rect 10834 37998 10846 38050
rect 15922 37998 15934 38050
rect 15986 37998 15998 38050
rect 22082 37998 22094 38050
rect 22146 37998 22158 38050
rect 3390 37986 3442 37998
rect 10558 37986 10610 37998
rect 21758 37986 21810 37998
rect 22766 37986 22818 37998
rect 23102 38050 23154 38062
rect 23102 37986 23154 37998
rect 23662 38050 23714 38062
rect 23662 37986 23714 37998
rect 2942 37938 2994 37950
rect 21422 37938 21474 37950
rect 2706 37886 2718 37938
rect 2770 37886 2782 37938
rect 6962 37886 6974 37938
rect 7026 37886 7038 37938
rect 2942 37874 2994 37886
rect 21422 37874 21474 37886
rect 3838 37826 3890 37838
rect 2482 37774 2494 37826
rect 2546 37774 2558 37826
rect 3838 37762 3890 37774
rect 5854 37826 5906 37838
rect 5854 37762 5906 37774
rect 10334 37826 10386 37838
rect 10334 37762 10386 37774
rect 10446 37826 10498 37838
rect 10446 37762 10498 37774
rect 11230 37826 11282 37838
rect 11230 37762 11282 37774
rect 12238 37826 12290 37838
rect 12238 37762 12290 37774
rect 12910 37826 12962 37838
rect 12910 37762 12962 37774
rect 14142 37826 14194 37838
rect 14142 37762 14194 37774
rect 22654 37826 22706 37838
rect 22654 37762 22706 37774
rect 22878 37826 22930 37838
rect 22878 37762 22930 37774
rect 22990 37826 23042 37838
rect 22990 37762 23042 37774
rect 24782 37826 24834 37838
rect 24782 37762 24834 37774
rect 26126 37826 26178 37838
rect 26126 37762 26178 37774
rect 26574 37826 26626 37838
rect 26574 37762 26626 37774
rect 28142 37826 28194 37838
rect 28142 37762 28194 37774
rect 1344 37658 28720 37692
rect 1344 37606 8018 37658
rect 8070 37606 8122 37658
rect 8174 37606 8226 37658
rect 8278 37606 14822 37658
rect 14874 37606 14926 37658
rect 14978 37606 15030 37658
rect 15082 37606 21626 37658
rect 21678 37606 21730 37658
rect 21782 37606 21834 37658
rect 21886 37606 28430 37658
rect 28482 37606 28534 37658
rect 28586 37606 28638 37658
rect 28690 37606 28720 37658
rect 1344 37572 28720 37606
rect 6414 37490 6466 37502
rect 6414 37426 6466 37438
rect 6862 37490 6914 37502
rect 6862 37426 6914 37438
rect 7310 37490 7362 37502
rect 7310 37426 7362 37438
rect 8206 37490 8258 37502
rect 8206 37426 8258 37438
rect 8430 37490 8482 37502
rect 8430 37426 8482 37438
rect 9662 37490 9714 37502
rect 9662 37426 9714 37438
rect 11454 37490 11506 37502
rect 11454 37426 11506 37438
rect 13582 37490 13634 37502
rect 13582 37426 13634 37438
rect 13918 37490 13970 37502
rect 13918 37426 13970 37438
rect 15262 37490 15314 37502
rect 15262 37426 15314 37438
rect 16046 37490 16098 37502
rect 16046 37426 16098 37438
rect 16830 37490 16882 37502
rect 16830 37426 16882 37438
rect 17502 37490 17554 37502
rect 17502 37426 17554 37438
rect 17614 37490 17666 37502
rect 17614 37426 17666 37438
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 18846 37490 18898 37502
rect 18846 37426 18898 37438
rect 19070 37490 19122 37502
rect 19070 37426 19122 37438
rect 19854 37490 19906 37502
rect 19854 37426 19906 37438
rect 20862 37490 20914 37502
rect 20862 37426 20914 37438
rect 22318 37490 22370 37502
rect 22318 37426 22370 37438
rect 22990 37490 23042 37502
rect 22990 37426 23042 37438
rect 23438 37490 23490 37502
rect 23438 37426 23490 37438
rect 25230 37490 25282 37502
rect 25230 37426 25282 37438
rect 25678 37490 25730 37502
rect 25678 37426 25730 37438
rect 27358 37490 27410 37502
rect 27358 37426 27410 37438
rect 7534 37378 7586 37390
rect 2482 37326 2494 37378
rect 2546 37326 2558 37378
rect 7534 37314 7586 37326
rect 7758 37378 7810 37390
rect 11006 37378 11058 37390
rect 10098 37326 10110 37378
rect 10162 37326 10174 37378
rect 7758 37314 7810 37326
rect 11006 37314 11058 37326
rect 11230 37378 11282 37390
rect 11230 37314 11282 37326
rect 11790 37378 11842 37390
rect 11790 37314 11842 37326
rect 20414 37378 20466 37390
rect 20414 37314 20466 37326
rect 23998 37378 24050 37390
rect 23998 37314 24050 37326
rect 24334 37378 24386 37390
rect 24334 37314 24386 37326
rect 7086 37266 7138 37278
rect 1810 37214 1822 37266
rect 1874 37214 1886 37266
rect 7086 37202 7138 37214
rect 8318 37266 8370 37278
rect 9998 37266 10050 37278
rect 8754 37214 8766 37266
rect 8818 37214 8830 37266
rect 8318 37202 8370 37214
rect 9998 37202 10050 37214
rect 10334 37266 10386 37278
rect 11454 37266 11506 37278
rect 10546 37214 10558 37266
rect 10610 37214 10622 37266
rect 10334 37202 10386 37214
rect 11454 37202 11506 37214
rect 12126 37266 12178 37278
rect 12126 37202 12178 37214
rect 12574 37266 12626 37278
rect 12574 37202 12626 37214
rect 12798 37266 12850 37278
rect 12798 37202 12850 37214
rect 14254 37266 14306 37278
rect 14254 37202 14306 37214
rect 14478 37266 14530 37278
rect 14478 37202 14530 37214
rect 14590 37266 14642 37278
rect 14590 37202 14642 37214
rect 15038 37266 15090 37278
rect 15038 37202 15090 37214
rect 17390 37266 17442 37278
rect 18958 37266 19010 37278
rect 17938 37214 17950 37266
rect 18002 37214 18014 37266
rect 17390 37202 17442 37214
rect 18958 37202 19010 37214
rect 19182 37266 19234 37278
rect 24558 37266 24610 37278
rect 19394 37214 19406 37266
rect 19458 37214 19470 37266
rect 22530 37214 22542 37266
rect 22594 37214 22606 37266
rect 19182 37202 19234 37214
rect 24558 37202 24610 37214
rect 25342 37266 25394 37278
rect 25342 37202 25394 37214
rect 25454 37266 25506 37278
rect 26898 37214 26910 37266
rect 26962 37214 26974 37266
rect 25454 37202 25506 37214
rect 5070 37154 5122 37166
rect 4610 37102 4622 37154
rect 4674 37102 4686 37154
rect 5070 37090 5122 37102
rect 5966 37154 6018 37166
rect 5966 37090 6018 37102
rect 12686 37154 12738 37166
rect 12686 37090 12738 37102
rect 15598 37154 15650 37166
rect 15598 37090 15650 37102
rect 21310 37154 21362 37166
rect 21310 37090 21362 37102
rect 21758 37154 21810 37166
rect 24110 37154 24162 37166
rect 21970 37102 21982 37154
rect 22034 37102 22046 37154
rect 21758 37090 21810 37102
rect 5854 37042 5906 37054
rect 21298 36990 21310 37042
rect 21362 37039 21374 37042
rect 21985 37039 22031 37102
rect 24110 37090 24162 37102
rect 26238 37154 26290 37166
rect 27918 37154 27970 37166
rect 26786 37102 26798 37154
rect 26850 37102 26862 37154
rect 26238 37090 26290 37102
rect 27918 37090 27970 37102
rect 21362 36993 22031 37039
rect 22206 37042 22258 37054
rect 21362 36990 21374 36993
rect 5854 36978 5906 36990
rect 22206 36978 22258 36990
rect 26574 37042 26626 37054
rect 26574 36978 26626 36990
rect 1344 36874 28560 36908
rect 1344 36822 4616 36874
rect 4668 36822 4720 36874
rect 4772 36822 4824 36874
rect 4876 36822 11420 36874
rect 11472 36822 11524 36874
rect 11576 36822 11628 36874
rect 11680 36822 18224 36874
rect 18276 36822 18328 36874
rect 18380 36822 18432 36874
rect 18484 36822 25028 36874
rect 25080 36822 25132 36874
rect 25184 36822 25236 36874
rect 25288 36822 28560 36874
rect 1344 36788 28560 36822
rect 3166 36706 3218 36718
rect 3166 36642 3218 36654
rect 6862 36706 6914 36718
rect 6862 36642 6914 36654
rect 14366 36706 14418 36718
rect 18610 36654 18622 36706
rect 18674 36703 18686 36706
rect 18674 36657 18783 36703
rect 18674 36654 18686 36657
rect 14366 36642 14418 36654
rect 2494 36594 2546 36606
rect 2494 36530 2546 36542
rect 3278 36594 3330 36606
rect 3278 36530 3330 36542
rect 3950 36594 4002 36606
rect 9326 36594 9378 36606
rect 18398 36594 18450 36606
rect 5058 36542 5070 36594
rect 5122 36542 5134 36594
rect 8642 36542 8654 36594
rect 8706 36542 8718 36594
rect 9986 36542 9998 36594
rect 10050 36542 10062 36594
rect 12114 36542 12126 36594
rect 12178 36542 12190 36594
rect 14578 36542 14590 36594
rect 14642 36542 14654 36594
rect 3950 36530 4002 36542
rect 9326 36530 9378 36542
rect 18398 36530 18450 36542
rect 1710 36482 1762 36494
rect 1710 36418 1762 36430
rect 4734 36482 4786 36494
rect 5966 36482 6018 36494
rect 5618 36430 5630 36482
rect 5682 36430 5694 36482
rect 4734 36418 4786 36430
rect 5966 36418 6018 36430
rect 6078 36482 6130 36494
rect 8430 36482 8482 36494
rect 13694 36482 13746 36494
rect 6738 36430 6750 36482
rect 6802 36430 6814 36482
rect 8194 36430 8206 36482
rect 8258 36430 8270 36482
rect 8866 36430 8878 36482
rect 8930 36430 8942 36482
rect 12898 36430 12910 36482
rect 12962 36430 12974 36482
rect 6078 36418 6130 36430
rect 8430 36418 8482 36430
rect 13694 36418 13746 36430
rect 13918 36482 13970 36494
rect 13918 36418 13970 36430
rect 14030 36482 14082 36494
rect 15150 36482 15202 36494
rect 14690 36430 14702 36482
rect 14754 36430 14766 36482
rect 14030 36418 14082 36430
rect 15150 36418 15202 36430
rect 15262 36482 15314 36494
rect 15262 36418 15314 36430
rect 15486 36482 15538 36494
rect 16494 36482 16546 36494
rect 15698 36430 15710 36482
rect 15762 36430 15774 36482
rect 15486 36418 15538 36430
rect 16494 36418 16546 36430
rect 4958 36370 5010 36382
rect 4958 36306 5010 36318
rect 6414 36370 6466 36382
rect 6414 36306 6466 36318
rect 13470 36370 13522 36382
rect 13470 36306 13522 36318
rect 16046 36370 16098 36382
rect 16046 36306 16098 36318
rect 16606 36370 16658 36382
rect 16606 36306 16658 36318
rect 17614 36370 17666 36382
rect 17614 36306 17666 36318
rect 2046 36258 2098 36270
rect 2046 36194 2098 36206
rect 4398 36258 4450 36270
rect 4398 36194 4450 36206
rect 5630 36258 5682 36270
rect 5630 36194 5682 36206
rect 8654 36258 8706 36270
rect 8654 36194 8706 36206
rect 15374 36258 15426 36270
rect 15374 36194 15426 36206
rect 16270 36258 16322 36270
rect 16270 36194 16322 36206
rect 16382 36258 16434 36270
rect 16382 36194 16434 36206
rect 17166 36258 17218 36270
rect 18737 36258 18783 36657
rect 26786 36654 26798 36706
rect 26850 36654 26862 36706
rect 19966 36594 20018 36606
rect 19966 36530 20018 36542
rect 22430 36594 22482 36606
rect 22430 36530 22482 36542
rect 22766 36594 22818 36606
rect 27806 36594 27858 36606
rect 24098 36542 24110 36594
rect 24162 36542 24174 36594
rect 26226 36542 26238 36594
rect 26290 36542 26302 36594
rect 22766 36530 22818 36542
rect 27806 36530 27858 36542
rect 18958 36482 19010 36494
rect 18958 36418 19010 36430
rect 21310 36482 21362 36494
rect 27022 36482 27074 36494
rect 23426 36430 23438 36482
rect 23490 36430 23502 36482
rect 26562 36430 26574 36482
rect 26626 36430 26638 36482
rect 21310 36418 21362 36430
rect 27022 36418 27074 36430
rect 27358 36482 27410 36494
rect 27358 36418 27410 36430
rect 19406 36370 19458 36382
rect 19406 36306 19458 36318
rect 21422 36370 21474 36382
rect 21422 36306 21474 36318
rect 21646 36370 21698 36382
rect 21646 36306 21698 36318
rect 21870 36370 21922 36382
rect 21870 36306 21922 36318
rect 19070 36258 19122 36270
rect 18722 36206 18734 36258
rect 18786 36206 18798 36258
rect 17166 36194 17218 36206
rect 19070 36194 19122 36206
rect 19182 36258 19234 36270
rect 19182 36194 19234 36206
rect 20414 36258 20466 36270
rect 20414 36194 20466 36206
rect 27246 36258 27298 36270
rect 27246 36194 27298 36206
rect 1344 36090 28720 36124
rect 1344 36038 8018 36090
rect 8070 36038 8122 36090
rect 8174 36038 8226 36090
rect 8278 36038 14822 36090
rect 14874 36038 14926 36090
rect 14978 36038 15030 36090
rect 15082 36038 21626 36090
rect 21678 36038 21730 36090
rect 21782 36038 21834 36090
rect 21886 36038 28430 36090
rect 28482 36038 28534 36090
rect 28586 36038 28638 36090
rect 28690 36038 28720 36090
rect 1344 36004 28720 36038
rect 3726 35922 3778 35934
rect 3726 35858 3778 35870
rect 7422 35922 7474 35934
rect 7422 35858 7474 35870
rect 8542 35922 8594 35934
rect 8542 35858 8594 35870
rect 8990 35922 9042 35934
rect 8990 35858 9042 35870
rect 10110 35922 10162 35934
rect 10110 35858 10162 35870
rect 12462 35922 12514 35934
rect 12462 35858 12514 35870
rect 16718 35922 16770 35934
rect 16718 35858 16770 35870
rect 9662 35810 9714 35822
rect 4834 35758 4846 35810
rect 4898 35758 4910 35810
rect 22978 35758 22990 35810
rect 23042 35758 23054 35810
rect 27346 35758 27358 35810
rect 27410 35758 27422 35810
rect 9662 35746 9714 35758
rect 12126 35698 12178 35710
rect 4050 35646 4062 35698
rect 4114 35646 4126 35698
rect 12126 35634 12178 35646
rect 12238 35698 12290 35710
rect 12238 35634 12290 35646
rect 12574 35698 12626 35710
rect 13346 35646 13358 35698
rect 13410 35646 13422 35698
rect 17378 35646 17390 35698
rect 17442 35646 17454 35698
rect 23762 35646 23774 35698
rect 23826 35646 23838 35698
rect 28018 35646 28030 35698
rect 28082 35646 28094 35698
rect 12574 35634 12626 35646
rect 1822 35586 1874 35598
rect 10782 35586 10834 35598
rect 6962 35534 6974 35586
rect 7026 35534 7038 35586
rect 1822 35522 1874 35534
rect 10782 35522 10834 35534
rect 11678 35586 11730 35598
rect 11678 35522 11730 35534
rect 12350 35586 12402 35598
rect 24222 35586 24274 35598
rect 14130 35534 14142 35586
rect 14194 35534 14206 35586
rect 16258 35534 16270 35586
rect 16322 35534 16334 35586
rect 18162 35534 18174 35586
rect 18226 35534 18238 35586
rect 20290 35534 20302 35586
rect 20354 35534 20366 35586
rect 20850 35534 20862 35586
rect 20914 35534 20926 35586
rect 12350 35522 12402 35534
rect 24222 35522 24274 35534
rect 24670 35586 24722 35598
rect 25218 35534 25230 35586
rect 25282 35534 25294 35586
rect 24670 35522 24722 35534
rect 1344 35306 28560 35340
rect 1344 35254 4616 35306
rect 4668 35254 4720 35306
rect 4772 35254 4824 35306
rect 4876 35254 11420 35306
rect 11472 35254 11524 35306
rect 11576 35254 11628 35306
rect 11680 35254 18224 35306
rect 18276 35254 18328 35306
rect 18380 35254 18432 35306
rect 18484 35254 25028 35306
rect 25080 35254 25132 35306
rect 25184 35254 25236 35306
rect 25288 35254 28560 35306
rect 1344 35220 28560 35254
rect 11678 35138 11730 35150
rect 14478 35138 14530 35150
rect 19182 35138 19234 35150
rect 13570 35086 13582 35138
rect 13634 35135 13646 35138
rect 13906 35135 13918 35138
rect 13634 35089 13918 35135
rect 13634 35086 13646 35089
rect 13906 35086 13918 35089
rect 13970 35086 13982 35138
rect 16370 35086 16382 35138
rect 16434 35086 16446 35138
rect 18610 35086 18622 35138
rect 18674 35135 18686 35138
rect 18946 35135 18958 35138
rect 18674 35089 18958 35135
rect 18674 35086 18686 35089
rect 18946 35086 18958 35089
rect 19010 35086 19022 35138
rect 24770 35086 24782 35138
rect 24834 35135 24846 35138
rect 25106 35135 25118 35138
rect 24834 35089 25118 35135
rect 24834 35086 24846 35089
rect 25106 35086 25118 35089
rect 25170 35086 25182 35138
rect 25890 35086 25902 35138
rect 25954 35135 25966 35138
rect 26562 35135 26574 35138
rect 25954 35089 26574 35135
rect 25954 35086 25966 35089
rect 26562 35086 26574 35089
rect 26626 35086 26638 35138
rect 11678 35074 11730 35086
rect 14478 35074 14530 35086
rect 19182 35074 19234 35086
rect 4846 35026 4898 35038
rect 12910 35026 12962 35038
rect 2930 34974 2942 35026
rect 2994 34974 3006 35026
rect 8642 34974 8654 35026
rect 8706 34974 8718 35026
rect 4846 34962 4898 34974
rect 12910 34962 12962 34974
rect 13582 35026 13634 35038
rect 13582 34962 13634 34974
rect 14814 35026 14866 35038
rect 14814 34962 14866 34974
rect 18062 35026 18114 35038
rect 18062 34962 18114 34974
rect 21534 35026 21586 35038
rect 21534 34962 21586 34974
rect 21982 35026 22034 35038
rect 21982 34962 22034 34974
rect 24670 35026 24722 35038
rect 24670 34962 24722 34974
rect 26238 35026 26290 35038
rect 26238 34962 26290 34974
rect 26574 35026 26626 35038
rect 26574 34962 26626 34974
rect 27134 35026 27186 35038
rect 27134 34962 27186 34974
rect 3502 34914 3554 34926
rect 8318 34914 8370 34926
rect 2818 34862 2830 34914
rect 2882 34862 2894 34914
rect 8082 34862 8094 34914
rect 8146 34862 8158 34914
rect 3502 34850 3554 34862
rect 8318 34850 8370 34862
rect 10110 34914 10162 34926
rect 10110 34850 10162 34862
rect 10670 34914 10722 34926
rect 14926 34914 14978 34926
rect 11330 34862 11342 34914
rect 11394 34862 11406 34914
rect 14130 34862 14142 34914
rect 14194 34862 14206 34914
rect 14690 34862 14702 34914
rect 14754 34862 14766 34914
rect 10670 34850 10722 34862
rect 14926 34850 14978 34862
rect 15934 34914 15986 34926
rect 15934 34850 15986 34862
rect 17950 34914 18002 34926
rect 17950 34850 18002 34862
rect 18174 34914 18226 34926
rect 18174 34850 18226 34862
rect 18510 34914 18562 34926
rect 20190 34914 20242 34926
rect 19618 34862 19630 34914
rect 19682 34862 19694 34914
rect 18510 34850 18562 34862
rect 20190 34850 20242 34862
rect 22542 34914 22594 34926
rect 22542 34850 22594 34862
rect 1710 34802 1762 34814
rect 1710 34738 1762 34750
rect 3390 34802 3442 34814
rect 3390 34738 3442 34750
rect 7758 34802 7810 34814
rect 7758 34738 7810 34750
rect 8654 34802 8706 34814
rect 8654 34738 8706 34750
rect 9550 34802 9602 34814
rect 9550 34738 9602 34750
rect 9774 34802 9826 34814
rect 9774 34738 9826 34750
rect 10334 34802 10386 34814
rect 11006 34802 11058 34814
rect 10770 34750 10782 34802
rect 10834 34750 10846 34802
rect 10334 34738 10386 34750
rect 11006 34738 11058 34750
rect 15710 34802 15762 34814
rect 15710 34738 15762 34750
rect 15822 34802 15874 34814
rect 15822 34738 15874 34750
rect 17614 34802 17666 34814
rect 20638 34802 20690 34814
rect 19730 34750 19742 34802
rect 19794 34750 19806 34802
rect 20066 34750 20078 34802
rect 20130 34750 20142 34802
rect 17614 34738 17666 34750
rect 20638 34738 20690 34750
rect 2046 34690 2098 34702
rect 2046 34626 2098 34638
rect 8542 34690 8594 34702
rect 8542 34626 8594 34638
rect 10110 34690 10162 34702
rect 10110 34626 10162 34638
rect 12462 34690 12514 34702
rect 12462 34626 12514 34638
rect 17054 34690 17106 34702
rect 17054 34626 17106 34638
rect 18958 34690 19010 34702
rect 18958 34626 19010 34638
rect 21870 34690 21922 34702
rect 21870 34626 21922 34638
rect 22094 34690 22146 34702
rect 22094 34626 22146 34638
rect 22878 34690 22930 34702
rect 22878 34626 22930 34638
rect 23326 34690 23378 34702
rect 23326 34626 23378 34638
rect 23886 34690 23938 34702
rect 23886 34626 23938 34638
rect 24222 34690 24274 34702
rect 24222 34626 24274 34638
rect 25118 34690 25170 34702
rect 25118 34626 25170 34638
rect 25678 34690 25730 34702
rect 25678 34626 25730 34638
rect 27694 34690 27746 34702
rect 27694 34626 27746 34638
rect 28142 34690 28194 34702
rect 28142 34626 28194 34638
rect 1344 34522 28720 34556
rect 1344 34470 8018 34522
rect 8070 34470 8122 34522
rect 8174 34470 8226 34522
rect 8278 34470 14822 34522
rect 14874 34470 14926 34522
rect 14978 34470 15030 34522
rect 15082 34470 21626 34522
rect 21678 34470 21730 34522
rect 21782 34470 21834 34522
rect 21886 34470 28430 34522
rect 28482 34470 28534 34522
rect 28586 34470 28638 34522
rect 28690 34470 28720 34522
rect 1344 34436 28720 34470
rect 6414 34354 6466 34366
rect 6414 34290 6466 34302
rect 7198 34354 7250 34366
rect 7198 34290 7250 34302
rect 8990 34354 9042 34366
rect 8990 34290 9042 34302
rect 12126 34354 12178 34366
rect 12126 34290 12178 34302
rect 13918 34354 13970 34366
rect 13918 34290 13970 34302
rect 15822 34354 15874 34366
rect 15822 34290 15874 34302
rect 18622 34354 18674 34366
rect 18622 34290 18674 34302
rect 19070 34354 19122 34366
rect 19070 34290 19122 34302
rect 19966 34354 20018 34366
rect 19966 34290 20018 34302
rect 20190 34354 20242 34366
rect 20190 34290 20242 34302
rect 20750 34354 20802 34366
rect 20750 34290 20802 34302
rect 21198 34354 21250 34366
rect 21198 34290 21250 34302
rect 21758 34354 21810 34366
rect 21758 34290 21810 34302
rect 22766 34354 22818 34366
rect 22766 34290 22818 34302
rect 23326 34354 23378 34366
rect 23326 34290 23378 34302
rect 25342 34354 25394 34366
rect 25342 34290 25394 34302
rect 26686 34354 26738 34366
rect 26686 34290 26738 34302
rect 27806 34354 27858 34366
rect 27806 34290 27858 34302
rect 27134 34242 27186 34254
rect 5730 34190 5742 34242
rect 5794 34190 5806 34242
rect 27134 34178 27186 34190
rect 27358 34242 27410 34254
rect 27358 34178 27410 34190
rect 5966 34130 6018 34142
rect 8094 34130 8146 34142
rect 1810 34078 1822 34130
rect 1874 34078 1886 34130
rect 5170 34078 5182 34130
rect 5234 34078 5246 34130
rect 7858 34078 7870 34130
rect 7922 34078 7934 34130
rect 5966 34066 6018 34078
rect 8094 34066 8146 34078
rect 8318 34130 8370 34142
rect 8318 34066 8370 34078
rect 8430 34130 8482 34142
rect 9774 34130 9826 34142
rect 9538 34078 9550 34130
rect 9602 34078 9614 34130
rect 8430 34066 8482 34078
rect 9774 34066 9826 34078
rect 9998 34130 10050 34142
rect 9998 34066 10050 34078
rect 10110 34130 10162 34142
rect 10110 34066 10162 34078
rect 10558 34130 10610 34142
rect 10558 34066 10610 34078
rect 10782 34130 10834 34142
rect 10782 34066 10834 34078
rect 11118 34130 11170 34142
rect 19854 34130 19906 34142
rect 19618 34078 19630 34130
rect 19682 34078 19694 34130
rect 11118 34066 11170 34078
rect 19854 34066 19906 34078
rect 20078 34130 20130 34142
rect 20078 34066 20130 34078
rect 25902 34130 25954 34142
rect 26114 34078 26126 34130
rect 26178 34078 26190 34130
rect 26450 34078 26462 34130
rect 26514 34078 26526 34130
rect 25902 34066 25954 34078
rect 5854 34018 5906 34030
rect 2482 33966 2494 34018
rect 2546 33966 2558 34018
rect 4610 33966 4622 34018
rect 4674 33966 4686 34018
rect 5854 33954 5906 33966
rect 6526 34018 6578 34030
rect 6526 33954 6578 33966
rect 7534 34018 7586 34030
rect 7534 33954 7586 33966
rect 8206 34018 8258 34030
rect 8206 33954 8258 33966
rect 9886 34018 9938 34030
rect 9886 33954 9938 33966
rect 10670 34018 10722 34030
rect 10670 33954 10722 33966
rect 11566 34018 11618 34030
rect 11566 33954 11618 33966
rect 12462 34018 12514 34030
rect 12462 33954 12514 33966
rect 15374 34018 15426 34030
rect 15374 33954 15426 33966
rect 18062 34018 18114 34030
rect 18062 33954 18114 33966
rect 22094 34018 22146 34030
rect 22094 33954 22146 33966
rect 23662 34018 23714 34030
rect 23662 33954 23714 33966
rect 24222 34018 24274 34030
rect 24222 33954 24274 33966
rect 24670 34018 24722 34030
rect 24670 33954 24722 33966
rect 27022 33906 27074 33918
rect 5394 33854 5406 33906
rect 5458 33854 5470 33906
rect 23986 33854 23998 33906
rect 24050 33903 24062 33906
rect 24658 33903 24670 33906
rect 24050 33857 24670 33903
rect 24050 33854 24062 33857
rect 24658 33854 24670 33857
rect 24722 33854 24734 33906
rect 26450 33854 26462 33906
rect 26514 33854 26526 33906
rect 27022 33842 27074 33854
rect 1344 33738 28560 33772
rect 1344 33686 4616 33738
rect 4668 33686 4720 33738
rect 4772 33686 4824 33738
rect 4876 33686 11420 33738
rect 11472 33686 11524 33738
rect 11576 33686 11628 33738
rect 11680 33686 18224 33738
rect 18276 33686 18328 33738
rect 18380 33686 18432 33738
rect 18484 33686 25028 33738
rect 25080 33686 25132 33738
rect 25184 33686 25236 33738
rect 25288 33686 28560 33738
rect 1344 33652 28560 33686
rect 3726 33570 3778 33582
rect 21422 33570 21474 33582
rect 8978 33518 8990 33570
rect 9042 33567 9054 33570
rect 9538 33567 9550 33570
rect 9042 33521 9550 33567
rect 9042 33518 9054 33521
rect 9538 33518 9550 33521
rect 9602 33518 9614 33570
rect 9762 33518 9774 33570
rect 9826 33567 9838 33570
rect 10098 33567 10110 33570
rect 9826 33521 10110 33567
rect 9826 33518 9838 33521
rect 10098 33518 10110 33521
rect 10162 33518 10174 33570
rect 3726 33506 3778 33518
rect 21422 33506 21474 33518
rect 2606 33458 2658 33470
rect 9102 33458 9154 33470
rect 3490 33406 3502 33458
rect 3554 33406 3566 33458
rect 6402 33406 6414 33458
rect 6466 33406 6478 33458
rect 8530 33406 8542 33458
rect 8594 33406 8606 33458
rect 2606 33394 2658 33406
rect 9102 33394 9154 33406
rect 9550 33458 9602 33470
rect 9550 33394 9602 33406
rect 10110 33458 10162 33470
rect 10110 33394 10162 33406
rect 12798 33458 12850 33470
rect 12798 33394 12850 33406
rect 14926 33458 14978 33470
rect 14926 33394 14978 33406
rect 18062 33458 18114 33470
rect 18062 33394 18114 33406
rect 24894 33458 24946 33470
rect 25218 33406 25230 33458
rect 25282 33406 25294 33458
rect 27346 33406 27358 33458
rect 27410 33406 27422 33458
rect 24894 33394 24946 33406
rect 10446 33346 10498 33358
rect 2370 33294 2382 33346
rect 2434 33294 2446 33346
rect 2818 33294 2830 33346
rect 2882 33294 2894 33346
rect 3378 33294 3390 33346
rect 3442 33294 3454 33346
rect 5730 33294 5742 33346
rect 5794 33294 5806 33346
rect 10446 33282 10498 33294
rect 11118 33346 11170 33358
rect 11118 33282 11170 33294
rect 12014 33346 12066 33358
rect 20078 33346 20130 33358
rect 12338 33294 12350 33346
rect 12402 33294 12414 33346
rect 15138 33294 15150 33346
rect 15202 33294 15214 33346
rect 12014 33282 12066 33294
rect 20078 33282 20130 33294
rect 20190 33346 20242 33358
rect 20190 33282 20242 33294
rect 21310 33346 21362 33358
rect 21310 33282 21362 33294
rect 22430 33346 22482 33358
rect 22430 33282 22482 33294
rect 22654 33346 22706 33358
rect 23986 33294 23998 33346
rect 24050 33294 24062 33346
rect 28018 33294 28030 33346
rect 28082 33294 28094 33346
rect 22654 33282 22706 33294
rect 3054 33234 3106 33246
rect 3054 33170 3106 33182
rect 10558 33234 10610 33246
rect 10558 33170 10610 33182
rect 10670 33234 10722 33246
rect 10670 33170 10722 33182
rect 11678 33234 11730 33246
rect 11678 33170 11730 33182
rect 14814 33234 14866 33246
rect 14814 33170 14866 33182
rect 15598 33234 15650 33246
rect 15598 33170 15650 33182
rect 19070 33234 19122 33246
rect 19070 33170 19122 33182
rect 20526 33234 20578 33246
rect 20526 33170 20578 33182
rect 22878 33234 22930 33246
rect 22878 33170 22930 33182
rect 4398 33122 4450 33134
rect 2594 33070 2606 33122
rect 2658 33070 2670 33122
rect 4398 33058 4450 33070
rect 4846 33122 4898 33134
rect 4846 33058 4898 33070
rect 11342 33122 11394 33134
rect 11342 33058 11394 33070
rect 11902 33122 11954 33134
rect 11902 33058 11954 33070
rect 12126 33122 12178 33134
rect 12126 33058 12178 33070
rect 13582 33122 13634 33134
rect 13582 33058 13634 33070
rect 18510 33122 18562 33134
rect 18510 33058 18562 33070
rect 19518 33122 19570 33134
rect 19518 33058 19570 33070
rect 19966 33122 20018 33134
rect 19966 33058 20018 33070
rect 20302 33122 20354 33134
rect 20302 33058 20354 33070
rect 21422 33122 21474 33134
rect 21422 33058 21474 33070
rect 22318 33122 22370 33134
rect 22318 33058 22370 33070
rect 22542 33122 22594 33134
rect 22542 33058 22594 33070
rect 23438 33122 23490 33134
rect 23438 33058 23490 33070
rect 23550 33122 23602 33134
rect 23550 33058 23602 33070
rect 23662 33122 23714 33134
rect 23662 33058 23714 33070
rect 24446 33122 24498 33134
rect 24446 33058 24498 33070
rect 1344 32954 28720 32988
rect 1344 32902 8018 32954
rect 8070 32902 8122 32954
rect 8174 32902 8226 32954
rect 8278 32902 14822 32954
rect 14874 32902 14926 32954
rect 14978 32902 15030 32954
rect 15082 32902 21626 32954
rect 21678 32902 21730 32954
rect 21782 32902 21834 32954
rect 21886 32902 28430 32954
rect 28482 32902 28534 32954
rect 28586 32902 28638 32954
rect 28690 32902 28720 32954
rect 1344 32868 28720 32902
rect 2606 32786 2658 32798
rect 2606 32722 2658 32734
rect 3054 32786 3106 32798
rect 3054 32722 3106 32734
rect 3502 32786 3554 32798
rect 3502 32722 3554 32734
rect 10446 32786 10498 32798
rect 10446 32722 10498 32734
rect 11006 32786 11058 32798
rect 11006 32722 11058 32734
rect 11454 32786 11506 32798
rect 11454 32722 11506 32734
rect 12574 32786 12626 32798
rect 12574 32722 12626 32734
rect 18734 32786 18786 32798
rect 18734 32722 18786 32734
rect 20190 32786 20242 32798
rect 20190 32722 20242 32734
rect 25678 32786 25730 32798
rect 25678 32722 25730 32734
rect 27134 32786 27186 32798
rect 27134 32722 27186 32734
rect 17390 32674 17442 32686
rect 17390 32610 17442 32622
rect 17726 32562 17778 32574
rect 12898 32510 12910 32562
rect 12962 32510 12974 32562
rect 17726 32498 17778 32510
rect 17838 32562 17890 32574
rect 18622 32562 18674 32574
rect 18386 32510 18398 32562
rect 18450 32510 18462 32562
rect 17838 32498 17890 32510
rect 18622 32498 18674 32510
rect 18846 32562 18898 32574
rect 19518 32562 19570 32574
rect 19058 32510 19070 32562
rect 19122 32510 19134 32562
rect 18846 32498 18898 32510
rect 19518 32498 19570 32510
rect 19966 32562 20018 32574
rect 19966 32498 20018 32510
rect 20078 32562 20130 32574
rect 20078 32498 20130 32510
rect 20302 32562 20354 32574
rect 26014 32562 26066 32574
rect 20514 32510 20526 32562
rect 20578 32510 20590 32562
rect 21858 32510 21870 32562
rect 21922 32510 21934 32562
rect 26338 32510 26350 32562
rect 26402 32510 26414 32562
rect 20302 32498 20354 32510
rect 26014 32498 26066 32510
rect 1822 32450 1874 32462
rect 1822 32386 1874 32398
rect 3950 32450 4002 32462
rect 3950 32386 4002 32398
rect 8766 32450 8818 32462
rect 8766 32386 8818 32398
rect 12126 32450 12178 32462
rect 16270 32450 16322 32462
rect 13682 32398 13694 32450
rect 13746 32398 13758 32450
rect 15810 32398 15822 32450
rect 15874 32398 15886 32450
rect 12126 32386 12178 32398
rect 16270 32386 16322 32398
rect 16830 32450 16882 32462
rect 16830 32386 16882 32398
rect 17502 32450 17554 32462
rect 17502 32386 17554 32398
rect 20974 32450 21026 32462
rect 20974 32386 21026 32398
rect 21422 32450 21474 32462
rect 27918 32450 27970 32462
rect 22530 32398 22542 32450
rect 22594 32398 22606 32450
rect 24658 32398 24670 32450
rect 24722 32398 24734 32450
rect 21422 32386 21474 32398
rect 27918 32386 27970 32398
rect 26350 32338 26402 32350
rect 3154 32286 3166 32338
rect 3218 32335 3230 32338
rect 3490 32335 3502 32338
rect 3218 32289 3502 32335
rect 3218 32286 3230 32289
rect 3490 32286 3502 32289
rect 3554 32335 3566 32338
rect 3938 32335 3950 32338
rect 3554 32289 3950 32335
rect 3554 32286 3566 32289
rect 3938 32286 3950 32289
rect 4002 32286 4014 32338
rect 26350 32274 26402 32286
rect 26686 32338 26738 32350
rect 26686 32274 26738 32286
rect 1344 32170 28560 32204
rect 1344 32118 4616 32170
rect 4668 32118 4720 32170
rect 4772 32118 4824 32170
rect 4876 32118 11420 32170
rect 11472 32118 11524 32170
rect 11576 32118 11628 32170
rect 11680 32118 18224 32170
rect 18276 32118 18328 32170
rect 18380 32118 18432 32170
rect 18484 32118 25028 32170
rect 25080 32118 25132 32170
rect 25184 32118 25236 32170
rect 25288 32118 28560 32170
rect 1344 32084 28560 32118
rect 2494 32002 2546 32014
rect 12798 32002 12850 32014
rect 11890 31950 11902 32002
rect 11954 31950 11966 32002
rect 2494 31938 2546 31950
rect 12798 31938 12850 31950
rect 19182 32002 19234 32014
rect 19182 31938 19234 31950
rect 3390 31890 3442 31902
rect 23102 31890 23154 31902
rect 9090 31838 9102 31890
rect 9154 31838 9166 31890
rect 9986 31838 9998 31890
rect 10050 31838 10062 31890
rect 12450 31838 12462 31890
rect 12514 31838 12526 31890
rect 3390 31826 3442 31838
rect 23102 31826 23154 31838
rect 24222 31890 24274 31902
rect 25218 31838 25230 31890
rect 25282 31838 25294 31890
rect 24222 31826 24274 31838
rect 5854 31778 5906 31790
rect 9774 31778 9826 31790
rect 20750 31778 20802 31790
rect 22990 31778 23042 31790
rect 2818 31726 2830 31778
rect 2882 31726 2894 31778
rect 4050 31726 4062 31778
rect 4114 31726 4126 31778
rect 4722 31726 4734 31778
rect 4786 31726 4798 31778
rect 6290 31726 6302 31778
rect 6354 31726 6366 31778
rect 10210 31726 10222 31778
rect 10274 31726 10286 31778
rect 11554 31726 11566 31778
rect 11618 31726 11630 31778
rect 12002 31726 12014 31778
rect 12066 31726 12078 31778
rect 17266 31726 17278 31778
rect 17330 31726 17342 31778
rect 19394 31726 19406 31778
rect 19458 31726 19470 31778
rect 20178 31726 20190 31778
rect 20242 31726 20254 31778
rect 21298 31726 21310 31778
rect 21362 31726 21374 31778
rect 5854 31714 5906 31726
rect 9774 31714 9826 31726
rect 20750 31714 20802 31726
rect 22990 31714 23042 31726
rect 23550 31778 23602 31790
rect 28018 31726 28030 31778
rect 28082 31726 28094 31778
rect 23550 31714 23602 31726
rect 1710 31666 1762 31678
rect 1710 31602 1762 31614
rect 2046 31666 2098 31678
rect 2046 31602 2098 31614
rect 5070 31666 5122 31678
rect 9550 31666 9602 31678
rect 6962 31614 6974 31666
rect 7026 31614 7038 31666
rect 5070 31602 5122 31614
rect 9550 31602 9602 31614
rect 11342 31666 11394 31678
rect 11342 31602 11394 31614
rect 12574 31666 12626 31678
rect 19518 31666 19570 31678
rect 22542 31666 22594 31678
rect 16706 31614 16718 31666
rect 16770 31614 16782 31666
rect 21522 31614 21534 31666
rect 21586 31614 21598 31666
rect 22194 31614 22206 31666
rect 22258 31614 22270 31666
rect 12574 31602 12626 31614
rect 19518 31602 19570 31614
rect 22542 31602 22594 31614
rect 23326 31666 23378 31678
rect 23326 31602 23378 31614
rect 24670 31666 24722 31678
rect 27346 31614 27358 31666
rect 27410 31614 27422 31666
rect 24670 31602 24722 31614
rect 2606 31554 2658 31566
rect 2606 31490 2658 31502
rect 3278 31554 3330 31566
rect 3278 31490 3330 31502
rect 4174 31554 4226 31566
rect 4174 31490 4226 31502
rect 9998 31554 10050 31566
rect 9998 31490 10050 31502
rect 11006 31554 11058 31566
rect 11006 31490 11058 31502
rect 11454 31554 11506 31566
rect 11454 31490 11506 31502
rect 1344 31386 28720 31420
rect 1344 31334 8018 31386
rect 8070 31334 8122 31386
rect 8174 31334 8226 31386
rect 8278 31334 14822 31386
rect 14874 31334 14926 31386
rect 14978 31334 15030 31386
rect 15082 31334 21626 31386
rect 21678 31334 21730 31386
rect 21782 31334 21834 31386
rect 21886 31334 28430 31386
rect 28482 31334 28534 31386
rect 28586 31334 28638 31386
rect 28690 31334 28720 31386
rect 1344 31300 28720 31334
rect 5070 31218 5122 31230
rect 5070 31154 5122 31166
rect 5742 31218 5794 31230
rect 5742 31154 5794 31166
rect 6302 31218 6354 31230
rect 6302 31154 6354 31166
rect 7086 31218 7138 31230
rect 7086 31154 7138 31166
rect 9886 31218 9938 31230
rect 9886 31154 9938 31166
rect 10222 31218 10274 31230
rect 10222 31154 10274 31166
rect 14142 31218 14194 31230
rect 14142 31154 14194 31166
rect 15934 31218 15986 31230
rect 15934 31154 15986 31166
rect 16046 31218 16098 31230
rect 16046 31154 16098 31166
rect 16494 31218 16546 31230
rect 16494 31154 16546 31166
rect 16942 31218 16994 31230
rect 16942 31154 16994 31166
rect 17950 31218 18002 31230
rect 17950 31154 18002 31166
rect 19070 31218 19122 31230
rect 19070 31154 19122 31166
rect 19518 31218 19570 31230
rect 24110 31218 24162 31230
rect 21634 31166 21646 31218
rect 21698 31166 21710 31218
rect 19518 31154 19570 31166
rect 24110 31154 24162 31166
rect 26686 31218 26738 31230
rect 26686 31154 26738 31166
rect 8206 31106 8258 31118
rect 15486 31106 15538 31118
rect 7186 31054 7198 31106
rect 7250 31054 7262 31106
rect 11330 31054 11342 31106
rect 11394 31054 11406 31106
rect 8206 31042 8258 31054
rect 15486 31042 15538 31054
rect 18174 31106 18226 31118
rect 18174 31042 18226 31054
rect 18734 31106 18786 31118
rect 18734 31042 18786 31054
rect 18846 31106 18898 31118
rect 22542 31106 22594 31118
rect 19842 31054 19854 31106
rect 19906 31054 19918 31106
rect 18846 31042 18898 31054
rect 22542 31042 22594 31054
rect 24334 31106 24386 31118
rect 26114 31054 26126 31106
rect 26178 31054 26190 31106
rect 24334 31042 24386 31054
rect 6974 30994 7026 31006
rect 14030 30994 14082 31006
rect 17838 30994 17890 31006
rect 1810 30942 1822 30994
rect 1874 30942 1886 30994
rect 7522 30942 7534 30994
rect 7586 30942 7598 30994
rect 8418 30942 8430 30994
rect 8482 30942 8494 30994
rect 10658 30942 10670 30994
rect 10722 30942 10734 30994
rect 14242 30942 14254 30994
rect 14306 30942 14318 30994
rect 14578 30942 14590 30994
rect 14642 30942 14654 30994
rect 15698 30942 15710 30994
rect 15762 30942 15774 30994
rect 17602 30942 17614 30994
rect 17666 30942 17678 30994
rect 6974 30930 7026 30942
rect 14030 30930 14082 30942
rect 17838 30930 17890 30942
rect 18062 30994 18114 31006
rect 18062 30930 18114 30942
rect 21534 30994 21586 31006
rect 21534 30930 21586 30942
rect 21982 30994 22034 31006
rect 25902 30994 25954 31006
rect 24658 30942 24670 30994
rect 24722 30942 24734 30994
rect 21982 30930 22034 30942
rect 25902 30930 25954 30942
rect 26350 30994 26402 31006
rect 26450 30942 26462 30994
rect 26514 30942 26526 30994
rect 26350 30930 26402 30942
rect 6638 30882 6690 30894
rect 2482 30830 2494 30882
rect 2546 30830 2558 30882
rect 4610 30830 4622 30882
rect 4674 30830 4686 30882
rect 6638 30818 6690 30830
rect 8094 30882 8146 30894
rect 8094 30818 8146 30830
rect 8878 30882 8930 30894
rect 24222 30882 24274 30894
rect 13458 30830 13470 30882
rect 13522 30830 13534 30882
rect 8878 30818 8930 30830
rect 24222 30818 24274 30830
rect 25342 30882 25394 30894
rect 25342 30818 25394 30830
rect 27134 30882 27186 30894
rect 27134 30818 27186 30830
rect 27582 30882 27634 30894
rect 27582 30818 27634 30830
rect 28142 30882 28194 30894
rect 28142 30818 28194 30830
rect 7522 30718 7534 30770
rect 7586 30718 7598 30770
rect 14578 30718 14590 30770
rect 14642 30718 14654 30770
rect 27234 30718 27246 30770
rect 27298 30767 27310 30770
rect 28130 30767 28142 30770
rect 27298 30721 28142 30767
rect 27298 30718 27310 30721
rect 28130 30718 28142 30721
rect 28194 30718 28206 30770
rect 1344 30602 28560 30636
rect 1344 30550 4616 30602
rect 4668 30550 4720 30602
rect 4772 30550 4824 30602
rect 4876 30550 11420 30602
rect 11472 30550 11524 30602
rect 11576 30550 11628 30602
rect 11680 30550 18224 30602
rect 18276 30550 18328 30602
rect 18380 30550 18432 30602
rect 18484 30550 25028 30602
rect 25080 30550 25132 30602
rect 25184 30550 25236 30602
rect 25288 30550 28560 30602
rect 1344 30516 28560 30550
rect 2606 30434 2658 30446
rect 4734 30434 4786 30446
rect 3490 30382 3502 30434
rect 3554 30431 3566 30434
rect 4050 30431 4062 30434
rect 3554 30385 4062 30431
rect 3554 30382 3566 30385
rect 4050 30382 4062 30385
rect 4114 30382 4126 30434
rect 2606 30370 2658 30382
rect 4734 30370 4786 30382
rect 5070 30434 5122 30446
rect 20638 30434 20690 30446
rect 5842 30382 5854 30434
rect 5906 30382 5918 30434
rect 18834 30382 18846 30434
rect 18898 30431 18910 30434
rect 19058 30431 19070 30434
rect 18898 30385 19070 30431
rect 18898 30382 18910 30385
rect 19058 30382 19070 30385
rect 19122 30382 19134 30434
rect 5070 30370 5122 30382
rect 20638 30370 20690 30382
rect 6862 30322 6914 30334
rect 6862 30258 6914 30270
rect 7646 30322 7698 30334
rect 7646 30258 7698 30270
rect 8318 30322 8370 30334
rect 8318 30258 8370 30270
rect 8430 30322 8482 30334
rect 11454 30322 11506 30334
rect 9762 30270 9774 30322
rect 9826 30270 9838 30322
rect 10882 30270 10894 30322
rect 10946 30270 10958 30322
rect 8430 30258 8482 30270
rect 11454 30258 11506 30270
rect 12574 30322 12626 30334
rect 12574 30258 12626 30270
rect 14814 30322 14866 30334
rect 21422 30322 21474 30334
rect 18386 30270 18398 30322
rect 18450 30270 18462 30322
rect 14814 30258 14866 30270
rect 21422 30258 21474 30270
rect 2046 30210 2098 30222
rect 6414 30210 6466 30222
rect 2258 30158 2270 30210
rect 2322 30158 2334 30210
rect 2818 30158 2830 30210
rect 2882 30158 2894 30210
rect 5058 30158 5070 30210
rect 5122 30158 5134 30210
rect 5618 30158 5630 30210
rect 5682 30158 5694 30210
rect 2046 30146 2098 30158
rect 6414 30146 6466 30158
rect 7198 30210 7250 30222
rect 9550 30210 9602 30222
rect 7410 30158 7422 30210
rect 7474 30158 7486 30210
rect 7858 30158 7870 30210
rect 7922 30158 7934 30210
rect 7198 30146 7250 30158
rect 9550 30146 9602 30158
rect 9886 30210 9938 30222
rect 10558 30210 10610 30222
rect 10322 30158 10334 30210
rect 10386 30158 10398 30210
rect 9886 30146 9938 30158
rect 10558 30146 10610 30158
rect 12014 30210 12066 30222
rect 18846 30210 18898 30222
rect 15586 30158 15598 30210
rect 15650 30158 15662 30210
rect 16258 30158 16270 30210
rect 16322 30158 16334 30210
rect 12014 30146 12066 30158
rect 18846 30146 18898 30158
rect 19854 30210 19906 30222
rect 19854 30146 19906 30158
rect 20750 30210 20802 30222
rect 23986 30158 23998 30210
rect 24050 30158 24062 30210
rect 20750 30146 20802 30158
rect 3054 30098 3106 30110
rect 9326 30098 9378 30110
rect 6178 30046 6190 30098
rect 6242 30046 6254 30098
rect 3054 30034 3106 30046
rect 9326 30034 9378 30046
rect 10894 30098 10946 30110
rect 10894 30034 10946 30046
rect 15150 30098 15202 30110
rect 27906 30046 27918 30098
rect 27970 30046 27982 30098
rect 15150 30034 15202 30046
rect 3614 29986 3666 29998
rect 2594 29934 2606 29986
rect 2658 29934 2670 29986
rect 3614 29922 3666 29934
rect 3950 29986 4002 29998
rect 3950 29922 4002 29934
rect 4398 29986 4450 29998
rect 4398 29922 4450 29934
rect 5630 29986 5682 29998
rect 5630 29922 5682 29934
rect 7310 29986 7362 29998
rect 7310 29922 7362 29934
rect 8542 29986 8594 29998
rect 8542 29922 8594 29934
rect 9774 29986 9826 29998
rect 9774 29922 9826 29934
rect 10782 29986 10834 29998
rect 10782 29922 10834 29934
rect 12910 29986 12962 29998
rect 12910 29922 12962 29934
rect 13806 29986 13858 29998
rect 13806 29922 13858 29934
rect 14142 29986 14194 29998
rect 14142 29922 14194 29934
rect 14590 29986 14642 29998
rect 14590 29922 14642 29934
rect 14702 29986 14754 29998
rect 14702 29922 14754 29934
rect 14926 29986 14978 29998
rect 14926 29922 14978 29934
rect 19294 29986 19346 29998
rect 19294 29922 19346 29934
rect 20190 29986 20242 29998
rect 20190 29922 20242 29934
rect 20638 29986 20690 29998
rect 20638 29922 20690 29934
rect 21870 29986 21922 29998
rect 21870 29922 21922 29934
rect 22542 29986 22594 29998
rect 22542 29922 22594 29934
rect 1344 29818 28720 29852
rect 1344 29766 8018 29818
rect 8070 29766 8122 29818
rect 8174 29766 8226 29818
rect 8278 29766 14822 29818
rect 14874 29766 14926 29818
rect 14978 29766 15030 29818
rect 15082 29766 21626 29818
rect 21678 29766 21730 29818
rect 21782 29766 21834 29818
rect 21886 29766 28430 29818
rect 28482 29766 28534 29818
rect 28586 29766 28638 29818
rect 28690 29766 28720 29818
rect 1344 29732 28720 29766
rect 11902 29650 11954 29662
rect 10546 29598 10558 29650
rect 10610 29598 10622 29650
rect 11902 29586 11954 29598
rect 12350 29650 12402 29662
rect 12350 29586 12402 29598
rect 16158 29650 16210 29662
rect 16158 29586 16210 29598
rect 17726 29650 17778 29662
rect 17726 29586 17778 29598
rect 17838 29650 17890 29662
rect 17838 29586 17890 29598
rect 2046 29538 2098 29550
rect 11230 29538 11282 29550
rect 21086 29538 21138 29550
rect 3602 29486 3614 29538
rect 3666 29486 3678 29538
rect 6850 29486 6862 29538
rect 6914 29486 6926 29538
rect 10322 29486 10334 29538
rect 10386 29486 10398 29538
rect 20178 29486 20190 29538
rect 20242 29486 20254 29538
rect 20402 29486 20414 29538
rect 20466 29486 20478 29538
rect 2046 29474 2098 29486
rect 11230 29474 11282 29486
rect 21086 29474 21138 29486
rect 1710 29426 1762 29438
rect 17950 29426 18002 29438
rect 2818 29374 2830 29426
rect 2882 29374 2894 29426
rect 6066 29374 6078 29426
rect 6130 29374 6142 29426
rect 10434 29374 10446 29426
rect 10498 29374 10510 29426
rect 10882 29374 10894 29426
rect 10946 29374 10958 29426
rect 12786 29374 12798 29426
rect 12850 29374 12862 29426
rect 17378 29374 17390 29426
rect 17442 29374 17454 29426
rect 18834 29374 18846 29426
rect 18898 29374 18910 29426
rect 19842 29374 19854 29426
rect 19906 29374 19918 29426
rect 24658 29374 24670 29426
rect 24722 29374 24734 29426
rect 28130 29374 28142 29426
rect 28194 29374 28206 29426
rect 1710 29362 1762 29374
rect 17950 29362 18002 29374
rect 2494 29314 2546 29326
rect 9662 29314 9714 29326
rect 16606 29314 16658 29326
rect 5730 29262 5742 29314
rect 5794 29262 5806 29314
rect 8978 29262 8990 29314
rect 9042 29262 9054 29314
rect 13570 29262 13582 29314
rect 13634 29262 13646 29314
rect 15698 29262 15710 29314
rect 15762 29262 15774 29314
rect 2494 29250 2546 29262
rect 9662 29250 9714 29262
rect 16606 29250 16658 29262
rect 19294 29314 19346 29326
rect 19294 29250 19346 29262
rect 21422 29314 21474 29326
rect 21746 29262 21758 29314
rect 21810 29262 21822 29314
rect 23874 29262 23886 29314
rect 23938 29262 23950 29314
rect 25218 29262 25230 29314
rect 25282 29262 25294 29314
rect 27346 29262 27358 29314
rect 27410 29262 27422 29314
rect 21422 29250 21474 29262
rect 18510 29202 18562 29214
rect 18510 29138 18562 29150
rect 18846 29202 18898 29214
rect 19058 29150 19070 29202
rect 19122 29199 19134 29202
rect 19618 29199 19630 29202
rect 19122 29153 19630 29199
rect 19122 29150 19134 29153
rect 19618 29150 19630 29153
rect 19682 29150 19694 29202
rect 18846 29138 18898 29150
rect 1344 29034 28560 29068
rect 1344 28982 4616 29034
rect 4668 28982 4720 29034
rect 4772 28982 4824 29034
rect 4876 28982 11420 29034
rect 11472 28982 11524 29034
rect 11576 28982 11628 29034
rect 11680 28982 18224 29034
rect 18276 28982 18328 29034
rect 18380 28982 18432 29034
rect 18484 28982 25028 29034
rect 25080 28982 25132 29034
rect 25184 28982 25236 29034
rect 25288 28982 28560 29034
rect 1344 28948 28560 28982
rect 3838 28866 3890 28878
rect 20414 28866 20466 28878
rect 2034 28814 2046 28866
rect 2098 28863 2110 28866
rect 2258 28863 2270 28866
rect 2098 28817 2270 28863
rect 2098 28814 2110 28817
rect 2258 28814 2270 28817
rect 2322 28814 2334 28866
rect 5954 28814 5966 28866
rect 6018 28863 6030 28866
rect 6402 28863 6414 28866
rect 6018 28817 6414 28863
rect 6018 28814 6030 28817
rect 6402 28814 6414 28817
rect 6466 28814 6478 28866
rect 3838 28802 3890 28814
rect 20414 28802 20466 28814
rect 2046 28754 2098 28766
rect 2046 28690 2098 28702
rect 2718 28754 2770 28766
rect 4286 28754 4338 28766
rect 3490 28702 3502 28754
rect 3554 28702 3566 28754
rect 2718 28690 2770 28702
rect 4286 28690 4338 28702
rect 5182 28754 5234 28766
rect 5182 28690 5234 28702
rect 5966 28754 6018 28766
rect 5966 28690 6018 28702
rect 6414 28754 6466 28766
rect 6414 28690 6466 28702
rect 6862 28754 6914 28766
rect 6862 28690 6914 28702
rect 7310 28754 7362 28766
rect 7310 28690 7362 28702
rect 12462 28754 12514 28766
rect 12462 28690 12514 28702
rect 12910 28754 12962 28766
rect 12910 28690 12962 28702
rect 13806 28754 13858 28766
rect 13806 28690 13858 28702
rect 14814 28754 14866 28766
rect 14814 28690 14866 28702
rect 15710 28754 15762 28766
rect 24670 28754 24722 28766
rect 19730 28702 19742 28754
rect 19794 28702 19806 28754
rect 21858 28702 21870 28754
rect 21922 28702 21934 28754
rect 15710 28690 15762 28702
rect 24670 28690 24722 28702
rect 27134 28754 27186 28766
rect 27134 28690 27186 28702
rect 27470 28754 27522 28766
rect 27470 28690 27522 28702
rect 4174 28642 4226 28654
rect 2370 28590 2382 28642
rect 2434 28590 2446 28642
rect 2930 28590 2942 28642
rect 2994 28590 3006 28642
rect 4174 28578 4226 28590
rect 11230 28642 11282 28654
rect 11230 28578 11282 28590
rect 14030 28642 14082 28654
rect 14030 28578 14082 28590
rect 14142 28642 14194 28654
rect 14926 28642 14978 28654
rect 16046 28642 16098 28654
rect 24222 28642 24274 28654
rect 14242 28590 14254 28642
rect 14306 28590 14318 28642
rect 15138 28590 15150 28642
rect 15202 28590 15214 28642
rect 16930 28590 16942 28642
rect 16994 28590 17006 28642
rect 20290 28590 20302 28642
rect 20354 28590 20366 28642
rect 23650 28590 23662 28642
rect 23714 28590 23726 28642
rect 14142 28578 14194 28590
rect 14926 28578 14978 28590
rect 16046 28578 16098 28590
rect 24222 28578 24274 28590
rect 24446 28642 24498 28654
rect 24446 28578 24498 28590
rect 24782 28642 24834 28654
rect 24782 28578 24834 28590
rect 25006 28642 25058 28654
rect 25006 28578 25058 28590
rect 25230 28642 25282 28654
rect 25230 28578 25282 28590
rect 25454 28642 25506 28654
rect 25454 28578 25506 28590
rect 25678 28642 25730 28654
rect 25678 28578 25730 28590
rect 26462 28642 26514 28654
rect 26462 28578 26514 28590
rect 3166 28530 3218 28542
rect 3166 28466 3218 28478
rect 3614 28530 3666 28542
rect 3614 28466 3666 28478
rect 13694 28530 13746 28542
rect 20750 28530 20802 28542
rect 17602 28478 17614 28530
rect 17666 28478 17678 28530
rect 13694 28466 13746 28478
rect 20750 28466 20802 28478
rect 26126 28530 26178 28542
rect 26126 28466 26178 28478
rect 26350 28530 26402 28542
rect 26350 28466 26402 28478
rect 2382 28418 2434 28430
rect 2382 28354 2434 28366
rect 11790 28418 11842 28430
rect 11790 28354 11842 28366
rect 20526 28418 20578 28430
rect 20526 28354 20578 28366
rect 26574 28418 26626 28430
rect 26574 28354 26626 28366
rect 28142 28418 28194 28430
rect 28142 28354 28194 28366
rect 1344 28250 28720 28284
rect 1344 28198 8018 28250
rect 8070 28198 8122 28250
rect 8174 28198 8226 28250
rect 8278 28198 14822 28250
rect 14874 28198 14926 28250
rect 14978 28198 15030 28250
rect 15082 28198 21626 28250
rect 21678 28198 21730 28250
rect 21782 28198 21834 28250
rect 21886 28198 28430 28250
rect 28482 28198 28534 28250
rect 28586 28198 28638 28250
rect 28690 28198 28720 28250
rect 1344 28164 28720 28198
rect 5070 28082 5122 28094
rect 5070 28018 5122 28030
rect 6638 28082 6690 28094
rect 6638 28018 6690 28030
rect 11454 28082 11506 28094
rect 11454 28018 11506 28030
rect 11566 28082 11618 28094
rect 11566 28018 11618 28030
rect 14254 28082 14306 28094
rect 14254 28018 14306 28030
rect 15710 28082 15762 28094
rect 15710 28018 15762 28030
rect 17726 28082 17778 28094
rect 17726 28018 17778 28030
rect 23998 28082 24050 28094
rect 23998 28018 24050 28030
rect 24670 28082 24722 28094
rect 24670 28018 24722 28030
rect 25678 28082 25730 28094
rect 25678 28018 25730 28030
rect 26686 28082 26738 28094
rect 26686 28018 26738 28030
rect 10222 27970 10274 27982
rect 2482 27918 2494 27970
rect 2546 27918 2558 27970
rect 10222 27906 10274 27918
rect 10446 27970 10498 27982
rect 10446 27906 10498 27918
rect 10782 27970 10834 27982
rect 10782 27906 10834 27918
rect 11006 27970 11058 27982
rect 25902 27970 25954 27982
rect 27134 27970 27186 27982
rect 17826 27918 17838 27970
rect 17890 27918 17902 27970
rect 26114 27918 26126 27970
rect 26178 27918 26190 27970
rect 11006 27906 11058 27918
rect 25902 27906 25954 27918
rect 27134 27906 27186 27918
rect 27358 27970 27410 27982
rect 27358 27906 27410 27918
rect 27806 27970 27858 27982
rect 27806 27906 27858 27918
rect 8990 27858 9042 27870
rect 1810 27806 1822 27858
rect 1874 27806 1886 27858
rect 8990 27794 9042 27806
rect 11342 27858 11394 27870
rect 11342 27794 11394 27806
rect 12014 27858 12066 27870
rect 17614 27858 17666 27870
rect 23102 27858 23154 27870
rect 14914 27806 14926 27858
rect 14978 27806 14990 27858
rect 18162 27806 18174 27858
rect 18226 27806 18238 27858
rect 19618 27806 19630 27858
rect 19682 27806 19694 27858
rect 22866 27806 22878 27858
rect 22930 27806 22942 27858
rect 12014 27794 12066 27806
rect 17614 27794 17666 27806
rect 23102 27794 23154 27806
rect 23326 27858 23378 27870
rect 23538 27806 23550 27858
rect 23602 27806 23614 27858
rect 26450 27806 26462 27858
rect 26514 27806 26526 27858
rect 23326 27794 23378 27806
rect 9662 27746 9714 27758
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 9662 27682 9714 27694
rect 10558 27746 10610 27758
rect 10558 27682 10610 27694
rect 12350 27746 12402 27758
rect 12350 27682 12402 27694
rect 12798 27746 12850 27758
rect 12798 27682 12850 27694
rect 15262 27746 15314 27758
rect 15262 27682 15314 27694
rect 16158 27746 16210 27758
rect 16158 27682 16210 27694
rect 16942 27746 16994 27758
rect 16942 27682 16994 27694
rect 18846 27746 18898 27758
rect 18846 27682 18898 27694
rect 19294 27746 19346 27758
rect 20402 27694 20414 27746
rect 20466 27694 20478 27746
rect 22530 27694 22542 27746
rect 22594 27694 22606 27746
rect 22978 27694 22990 27746
rect 23042 27694 23054 27746
rect 19294 27682 19346 27694
rect 14926 27634 14978 27646
rect 26350 27634 26402 27646
rect 18162 27582 18174 27634
rect 18226 27582 18238 27634
rect 14926 27570 14978 27582
rect 26350 27570 26402 27582
rect 27022 27634 27074 27646
rect 27022 27570 27074 27582
rect 1344 27466 28560 27500
rect 1344 27414 4616 27466
rect 4668 27414 4720 27466
rect 4772 27414 4824 27466
rect 4876 27414 11420 27466
rect 11472 27414 11524 27466
rect 11576 27414 11628 27466
rect 11680 27414 18224 27466
rect 18276 27414 18328 27466
rect 18380 27414 18432 27466
rect 18484 27414 25028 27466
rect 25080 27414 25132 27466
rect 25184 27414 25236 27466
rect 25288 27414 28560 27466
rect 1344 27380 28560 27414
rect 8542 27298 8594 27310
rect 17938 27246 17950 27298
rect 18002 27295 18014 27298
rect 18498 27295 18510 27298
rect 18002 27249 18510 27295
rect 18002 27246 18014 27249
rect 18498 27246 18510 27249
rect 18562 27246 18574 27298
rect 24658 27295 24670 27298
rect 24113 27249 24670 27295
rect 8542 27234 8594 27246
rect 2494 27186 2546 27198
rect 2494 27122 2546 27134
rect 3838 27186 3890 27198
rect 3838 27122 3890 27134
rect 4286 27186 4338 27198
rect 4286 27122 4338 27134
rect 5070 27186 5122 27198
rect 5070 27122 5122 27134
rect 5630 27186 5682 27198
rect 6414 27186 6466 27198
rect 7758 27186 7810 27198
rect 12910 27186 12962 27198
rect 16830 27186 16882 27198
rect 5954 27134 5966 27186
rect 6018 27134 6030 27186
rect 6850 27134 6862 27186
rect 6914 27134 6926 27186
rect 10322 27134 10334 27186
rect 10386 27134 10398 27186
rect 12450 27134 12462 27186
rect 12514 27134 12526 27186
rect 16370 27134 16382 27186
rect 16434 27134 16446 27186
rect 5630 27122 5682 27134
rect 6414 27122 6466 27134
rect 7758 27122 7810 27134
rect 12910 27122 12962 27134
rect 16830 27122 16882 27134
rect 19070 27186 19122 27198
rect 19070 27122 19122 27134
rect 20302 27186 20354 27198
rect 22306 27134 22318 27186
rect 22370 27134 22382 27186
rect 23986 27134 23998 27186
rect 24050 27183 24062 27186
rect 24113 27183 24159 27249
rect 24658 27246 24670 27249
rect 24722 27246 24734 27298
rect 24050 27137 24159 27183
rect 24446 27186 24498 27198
rect 24050 27134 24062 27137
rect 25218 27134 25230 27186
rect 25282 27134 25294 27186
rect 27346 27134 27358 27186
rect 27410 27134 27422 27186
rect 20302 27122 20354 27134
rect 24446 27122 24498 27134
rect 2942 27074 2994 27086
rect 18622 27074 18674 27086
rect 6738 27022 6750 27074
rect 6802 27022 6814 27074
rect 2942 27010 2994 27022
rect 8094 27018 8146 27030
rect 8306 27022 8318 27074
rect 8370 27022 8382 27074
rect 8866 27022 8878 27074
rect 8930 27022 8942 27074
rect 9650 27022 9662 27074
rect 9714 27022 9726 27074
rect 13570 27022 13582 27074
rect 13634 27022 13646 27074
rect 1710 26962 1762 26974
rect 1710 26898 1762 26910
rect 5854 26962 5906 26974
rect 18622 27010 18674 27022
rect 20414 27074 20466 27086
rect 23650 27022 23662 27074
rect 23714 27022 23726 27074
rect 28130 27022 28142 27074
rect 28194 27022 28206 27074
rect 20414 27010 20466 27022
rect 8094 26954 8146 26966
rect 18286 26962 18338 26974
rect 14242 26910 14254 26962
rect 14306 26910 14318 26962
rect 5854 26898 5906 26910
rect 18286 26898 18338 26910
rect 20190 26962 20242 26974
rect 20190 26898 20242 26910
rect 20750 26962 20802 26974
rect 20750 26898 20802 26910
rect 2046 26850 2098 26862
rect 2046 26786 2098 26798
rect 3390 26850 3442 26862
rect 3390 26786 3442 26798
rect 6302 26850 6354 26862
rect 6302 26786 6354 26798
rect 8206 26850 8258 26862
rect 8206 26786 8258 26798
rect 19854 26850 19906 26862
rect 19854 26786 19906 26798
rect 24894 26850 24946 26862
rect 24894 26786 24946 26798
rect 1344 26682 28720 26716
rect 1344 26630 8018 26682
rect 8070 26630 8122 26682
rect 8174 26630 8226 26682
rect 8278 26630 14822 26682
rect 14874 26630 14926 26682
rect 14978 26630 15030 26682
rect 15082 26630 21626 26682
rect 21678 26630 21730 26682
rect 21782 26630 21834 26682
rect 21886 26630 28430 26682
rect 28482 26630 28534 26682
rect 28586 26630 28638 26682
rect 28690 26630 28720 26682
rect 1344 26596 28720 26630
rect 2830 26514 2882 26526
rect 2830 26450 2882 26462
rect 9662 26514 9714 26526
rect 9662 26450 9714 26462
rect 12574 26514 12626 26526
rect 12574 26450 12626 26462
rect 13470 26514 13522 26526
rect 15262 26514 15314 26526
rect 14242 26462 14254 26514
rect 14306 26462 14318 26514
rect 13470 26450 13522 26462
rect 15262 26450 15314 26462
rect 15710 26514 15762 26526
rect 15710 26450 15762 26462
rect 16382 26514 16434 26526
rect 16382 26450 16434 26462
rect 20190 26514 20242 26526
rect 20190 26450 20242 26462
rect 21310 26514 21362 26526
rect 21310 26450 21362 26462
rect 21422 26514 21474 26526
rect 21422 26450 21474 26462
rect 21534 26514 21586 26526
rect 21534 26450 21586 26462
rect 23886 26514 23938 26526
rect 23886 26450 23938 26462
rect 24334 26514 24386 26526
rect 24334 26450 24386 26462
rect 25230 26514 25282 26526
rect 25230 26450 25282 26462
rect 26238 26514 26290 26526
rect 26238 26450 26290 26462
rect 26910 26514 26962 26526
rect 26910 26450 26962 26462
rect 27358 26514 27410 26526
rect 27358 26450 27410 26462
rect 13358 26402 13410 26414
rect 3378 26350 3390 26402
rect 3442 26350 3454 26402
rect 6066 26350 6078 26402
rect 6130 26350 6142 26402
rect 13358 26338 13410 26350
rect 14030 26402 14082 26414
rect 14030 26338 14082 26350
rect 17390 26402 17442 26414
rect 17390 26338 17442 26350
rect 19294 26402 19346 26414
rect 19294 26338 19346 26350
rect 19742 26402 19794 26414
rect 19742 26338 19794 26350
rect 10782 26290 10834 26302
rect 4946 26238 4958 26290
rect 5010 26238 5022 26290
rect 9874 26238 9886 26290
rect 9938 26238 9950 26290
rect 10782 26226 10834 26238
rect 12798 26290 12850 26302
rect 14366 26290 14418 26302
rect 21982 26290 22034 26302
rect 25454 26290 25506 26302
rect 13122 26238 13134 26290
rect 13186 26238 13198 26290
rect 14802 26238 14814 26290
rect 14866 26238 14878 26290
rect 17602 26238 17614 26290
rect 17666 26238 17678 26290
rect 18162 26238 18174 26290
rect 18226 26238 18238 26290
rect 18498 26238 18510 26290
rect 18562 26238 18574 26290
rect 22642 26238 22654 26290
rect 22706 26238 22718 26290
rect 12798 26226 12850 26238
rect 14366 26226 14418 26238
rect 21982 26226 22034 26238
rect 25454 26226 25506 26238
rect 25902 26290 25954 26302
rect 25902 26226 25954 26238
rect 10334 26178 10386 26190
rect 10334 26114 10386 26126
rect 12126 26178 12178 26190
rect 12126 26114 12178 26126
rect 16830 26178 16882 26190
rect 16830 26114 16882 26126
rect 17502 26178 17554 26190
rect 17502 26114 17554 26126
rect 20974 26178 21026 26190
rect 20974 26114 21026 26126
rect 22318 26178 22370 26190
rect 23438 26178 23490 26190
rect 22754 26126 22766 26178
rect 22818 26126 22830 26178
rect 22318 26114 22370 26126
rect 23438 26114 23490 26126
rect 25342 26178 25394 26190
rect 25342 26114 25394 26126
rect 28142 26178 28194 26190
rect 28142 26114 28194 26126
rect 9550 26066 9602 26078
rect 17838 26066 17890 26078
rect 14578 26014 14590 26066
rect 14642 26014 14654 26066
rect 15138 26014 15150 26066
rect 15202 26063 15214 26066
rect 15810 26063 15822 26066
rect 15202 26017 15822 26063
rect 15202 26014 15214 26017
rect 15810 26014 15822 26017
rect 15874 26014 15886 26066
rect 9550 26002 9602 26014
rect 17838 26002 17890 26014
rect 18510 26066 18562 26078
rect 18510 26002 18562 26014
rect 18846 26066 18898 26078
rect 18846 26002 18898 26014
rect 22990 26066 23042 26078
rect 22990 26002 23042 26014
rect 1344 25898 28560 25932
rect 1344 25846 4616 25898
rect 4668 25846 4720 25898
rect 4772 25846 4824 25898
rect 4876 25846 11420 25898
rect 11472 25846 11524 25898
rect 11576 25846 11628 25898
rect 11680 25846 18224 25898
rect 18276 25846 18328 25898
rect 18380 25846 18432 25898
rect 18484 25846 25028 25898
rect 25080 25846 25132 25898
rect 25184 25846 25236 25898
rect 25288 25846 28560 25898
rect 1344 25812 28560 25846
rect 2494 25730 2546 25742
rect 2494 25666 2546 25678
rect 5966 25730 6018 25742
rect 5966 25666 6018 25678
rect 2270 25618 2322 25630
rect 2270 25554 2322 25566
rect 5070 25618 5122 25630
rect 12910 25618 12962 25630
rect 7858 25566 7870 25618
rect 7922 25566 7934 25618
rect 9986 25566 9998 25618
rect 10050 25566 10062 25618
rect 5070 25554 5122 25566
rect 12910 25554 12962 25566
rect 13806 25618 13858 25630
rect 20190 25618 20242 25630
rect 16706 25566 16718 25618
rect 16770 25566 16782 25618
rect 18834 25566 18846 25618
rect 18898 25566 18910 25618
rect 13806 25554 13858 25566
rect 20190 25554 20242 25566
rect 20750 25618 20802 25630
rect 21634 25566 21646 25618
rect 21698 25566 21710 25618
rect 24882 25566 24894 25618
rect 24946 25566 24958 25618
rect 20750 25554 20802 25566
rect 4062 25506 4114 25518
rect 6414 25506 6466 25518
rect 14142 25506 14194 25518
rect 19294 25506 19346 25518
rect 3490 25454 3502 25506
rect 3554 25454 3566 25506
rect 5730 25454 5742 25506
rect 5794 25454 5806 25506
rect 6178 25454 6190 25506
rect 6242 25454 6254 25506
rect 7186 25454 7198 25506
rect 7250 25454 7262 25506
rect 16034 25454 16046 25506
rect 16098 25454 16110 25506
rect 24546 25454 24558 25506
rect 24610 25454 24622 25506
rect 27794 25454 27806 25506
rect 27858 25454 27870 25506
rect 4062 25442 4114 25454
rect 6414 25442 6466 25454
rect 14142 25442 14194 25454
rect 19294 25442 19346 25454
rect 2718 25394 2770 25406
rect 2718 25330 2770 25342
rect 4622 25394 4674 25406
rect 4622 25330 4674 25342
rect 14478 25394 14530 25406
rect 23762 25342 23774 25394
rect 23826 25342 23838 25394
rect 27010 25342 27022 25394
rect 27074 25342 27086 25394
rect 14478 25330 14530 25342
rect 2606 25282 2658 25294
rect 2606 25218 2658 25230
rect 5630 25282 5682 25294
rect 5630 25218 5682 25230
rect 10446 25282 10498 25294
rect 10446 25218 10498 25230
rect 14366 25282 14418 25294
rect 14366 25218 14418 25230
rect 14926 25282 14978 25294
rect 14926 25218 14978 25230
rect 15374 25282 15426 25294
rect 15374 25218 15426 25230
rect 19742 25282 19794 25294
rect 19742 25218 19794 25230
rect 1344 25114 28720 25148
rect 1344 25062 8018 25114
rect 8070 25062 8122 25114
rect 8174 25062 8226 25114
rect 8278 25062 14822 25114
rect 14874 25062 14926 25114
rect 14978 25062 15030 25114
rect 15082 25062 21626 25114
rect 21678 25062 21730 25114
rect 21782 25062 21834 25114
rect 21886 25062 28430 25114
rect 28482 25062 28534 25114
rect 28586 25062 28638 25114
rect 28690 25062 28720 25114
rect 1344 25028 28720 25062
rect 2382 24946 2434 24958
rect 2382 24882 2434 24894
rect 7758 24946 7810 24958
rect 7758 24882 7810 24894
rect 8990 24946 9042 24958
rect 8990 24882 9042 24894
rect 14254 24946 14306 24958
rect 14254 24882 14306 24894
rect 15150 24946 15202 24958
rect 15150 24882 15202 24894
rect 15710 24946 15762 24958
rect 15710 24882 15762 24894
rect 16942 24946 16994 24958
rect 20190 24946 20242 24958
rect 18722 24894 18734 24946
rect 18786 24894 18798 24946
rect 16942 24882 16994 24894
rect 20190 24882 20242 24894
rect 20974 24946 21026 24958
rect 20974 24882 21026 24894
rect 21198 24946 21250 24958
rect 21198 24882 21250 24894
rect 22990 24946 23042 24958
rect 22990 24882 23042 24894
rect 25678 24946 25730 24958
rect 25678 24882 25730 24894
rect 3614 24834 3666 24846
rect 16270 24834 16322 24846
rect 5170 24782 5182 24834
rect 5234 24782 5246 24834
rect 3614 24770 3666 24782
rect 16270 24770 16322 24782
rect 19630 24834 19682 24846
rect 19630 24770 19682 24782
rect 20078 24834 20130 24846
rect 20078 24770 20130 24782
rect 20414 24834 20466 24846
rect 20414 24770 20466 24782
rect 20862 24834 20914 24846
rect 20862 24770 20914 24782
rect 25454 24834 25506 24846
rect 25454 24770 25506 24782
rect 2046 24722 2098 24734
rect 3166 24722 3218 24734
rect 2370 24670 2382 24722
rect 2434 24670 2446 24722
rect 2930 24670 2942 24722
rect 2994 24670 3006 24722
rect 2046 24658 2098 24670
rect 3166 24658 3218 24670
rect 3502 24722 3554 24734
rect 3502 24658 3554 24670
rect 4062 24722 4114 24734
rect 13358 24722 13410 24734
rect 4498 24670 4510 24722
rect 4562 24670 4574 24722
rect 9650 24670 9662 24722
rect 9714 24670 9726 24722
rect 4062 24658 4114 24670
rect 13358 24658 13410 24670
rect 16158 24722 16210 24734
rect 22206 24722 22258 24734
rect 16594 24670 16606 24722
rect 16658 24670 16670 24722
rect 19842 24670 19854 24722
rect 19906 24670 19918 24722
rect 20626 24670 20638 24722
rect 20690 24670 20702 24722
rect 21410 24670 21422 24722
rect 21474 24670 21486 24722
rect 21634 24670 21646 24722
rect 21698 24670 21710 24722
rect 16158 24658 16210 24670
rect 22206 24658 22258 24670
rect 22542 24722 22594 24734
rect 25342 24722 25394 24734
rect 22866 24670 22878 24722
rect 22930 24670 22942 24722
rect 22542 24658 22594 24670
rect 25342 24658 25394 24670
rect 25902 24722 25954 24734
rect 25902 24658 25954 24670
rect 12910 24610 12962 24622
rect 7298 24558 7310 24610
rect 7362 24558 7374 24610
rect 10322 24558 10334 24610
rect 10386 24558 10398 24610
rect 12450 24558 12462 24610
rect 12514 24558 12526 24610
rect 12910 24546 12962 24558
rect 14702 24610 14754 24622
rect 14702 24546 14754 24558
rect 15934 24610 15986 24622
rect 15934 24546 15986 24558
rect 17614 24610 17666 24622
rect 17614 24546 17666 24558
rect 17950 24610 18002 24622
rect 17950 24546 18002 24558
rect 18398 24610 18450 24622
rect 18398 24546 18450 24558
rect 19294 24610 19346 24622
rect 19294 24546 19346 24558
rect 21534 24610 21586 24622
rect 21534 24546 21586 24558
rect 23438 24610 23490 24622
rect 23438 24546 23490 24558
rect 24222 24610 24274 24622
rect 24222 24546 24274 24558
rect 24670 24610 24722 24622
rect 24670 24546 24722 24558
rect 26238 24610 26290 24622
rect 26238 24546 26290 24558
rect 26910 24610 26962 24622
rect 26910 24546 26962 24558
rect 27358 24610 27410 24622
rect 27358 24546 27410 24558
rect 28142 24610 28194 24622
rect 28142 24546 28194 24558
rect 19070 24498 19122 24510
rect 2594 24446 2606 24498
rect 2658 24446 2670 24498
rect 14242 24446 14254 24498
rect 14306 24495 14318 24498
rect 14914 24495 14926 24498
rect 14306 24449 14926 24495
rect 14306 24446 14318 24449
rect 14914 24446 14926 24449
rect 14978 24446 14990 24498
rect 22754 24446 22766 24498
rect 22818 24446 22830 24498
rect 23090 24446 23102 24498
rect 23154 24495 23166 24498
rect 23426 24495 23438 24498
rect 23154 24449 23438 24495
rect 23154 24446 23166 24449
rect 23426 24446 23438 24449
rect 23490 24446 23502 24498
rect 19070 24434 19122 24446
rect 1344 24330 28560 24364
rect 1344 24278 4616 24330
rect 4668 24278 4720 24330
rect 4772 24278 4824 24330
rect 4876 24278 11420 24330
rect 11472 24278 11524 24330
rect 11576 24278 11628 24330
rect 11680 24278 18224 24330
rect 18276 24278 18328 24330
rect 18380 24278 18432 24330
rect 18484 24278 25028 24330
rect 25080 24278 25132 24330
rect 25184 24278 25236 24330
rect 25288 24278 28560 24330
rect 1344 24244 28560 24278
rect 15822 24162 15874 24174
rect 15822 24098 15874 24110
rect 16606 24162 16658 24174
rect 16606 24098 16658 24110
rect 16942 24162 16994 24174
rect 16942 24098 16994 24110
rect 18510 24162 18562 24174
rect 22082 24110 22094 24162
rect 22146 24159 22158 24162
rect 22866 24159 22878 24162
rect 22146 24113 22878 24159
rect 22146 24110 22158 24113
rect 22866 24110 22878 24113
rect 22930 24110 22942 24162
rect 18510 24098 18562 24110
rect 5742 24050 5794 24062
rect 2482 23998 2494 24050
rect 2546 23998 2558 24050
rect 4610 23998 4622 24050
rect 4674 23998 4686 24050
rect 8978 24024 8990 24076
rect 9042 24024 9054 24076
rect 9774 24050 9826 24062
rect 13470 24050 13522 24062
rect 20190 24050 20242 24062
rect 5742 23986 5794 23998
rect 12786 23998 12798 24050
rect 12850 23998 12862 24050
rect 14018 23998 14030 24050
rect 14082 23998 14094 24050
rect 19282 23998 19294 24050
rect 19346 23998 19358 24050
rect 9774 23986 9826 23998
rect 13470 23986 13522 23998
rect 20190 23986 20242 23998
rect 20638 24050 20690 24062
rect 20638 23986 20690 23998
rect 21422 24050 21474 24062
rect 21422 23986 21474 23998
rect 24558 24050 24610 24062
rect 24558 23986 24610 23998
rect 25342 24050 25394 24062
rect 25342 23986 25394 23998
rect 27246 24050 27298 24062
rect 27246 23986 27298 23998
rect 27694 24050 27746 24062
rect 27694 23986 27746 23998
rect 10110 23938 10162 23950
rect 1810 23886 1822 23938
rect 1874 23886 1886 23938
rect 6066 23886 6078 23938
rect 6130 23886 6142 23938
rect 10110 23874 10162 23886
rect 10446 23938 10498 23950
rect 10446 23874 10498 23886
rect 11230 23938 11282 23950
rect 11230 23874 11282 23886
rect 11566 23938 11618 23950
rect 11566 23874 11618 23886
rect 11790 23938 11842 23950
rect 11790 23874 11842 23886
rect 12350 23938 12402 23950
rect 12350 23874 12402 23886
rect 13694 23938 13746 23950
rect 13694 23874 13746 23886
rect 14478 23938 14530 23950
rect 14478 23874 14530 23886
rect 14926 23938 14978 23950
rect 19854 23938 19906 23950
rect 26350 23938 26402 23950
rect 16706 23886 16718 23938
rect 16770 23886 16782 23938
rect 26226 23886 26238 23938
rect 26290 23886 26302 23938
rect 14926 23874 14978 23886
rect 19854 23874 19906 23886
rect 26350 23874 26402 23886
rect 10670 23826 10722 23838
rect 6850 23774 6862 23826
rect 6914 23774 6926 23826
rect 10670 23762 10722 23774
rect 11678 23826 11730 23838
rect 11678 23762 11730 23774
rect 12014 23826 12066 23838
rect 12014 23762 12066 23774
rect 12686 23826 12738 23838
rect 12686 23762 12738 23774
rect 15150 23826 15202 23838
rect 15150 23762 15202 23774
rect 15710 23826 15762 23838
rect 15710 23762 15762 23774
rect 16270 23826 16322 23838
rect 16270 23762 16322 23774
rect 17502 23826 17554 23838
rect 17502 23762 17554 23774
rect 17950 23826 18002 23838
rect 17950 23762 18002 23774
rect 18398 23826 18450 23838
rect 26798 23826 26850 23838
rect 26562 23774 26574 23826
rect 26626 23774 26638 23826
rect 18398 23762 18450 23774
rect 26798 23762 26850 23774
rect 5070 23714 5122 23726
rect 5070 23650 5122 23662
rect 10334 23714 10386 23726
rect 10334 23650 10386 23662
rect 12910 23714 12962 23726
rect 12910 23650 12962 23662
rect 14702 23714 14754 23726
rect 14702 23650 14754 23662
rect 15822 23714 15874 23726
rect 15822 23650 15874 23662
rect 16494 23714 16546 23726
rect 16494 23650 16546 23662
rect 17054 23714 17106 23726
rect 17054 23650 17106 23662
rect 17278 23714 17330 23726
rect 17278 23650 17330 23662
rect 18174 23714 18226 23726
rect 18174 23650 18226 23662
rect 18846 23714 18898 23726
rect 18846 23650 18898 23662
rect 19294 23714 19346 23726
rect 19294 23650 19346 23662
rect 19518 23714 19570 23726
rect 19518 23650 19570 23662
rect 21870 23714 21922 23726
rect 21870 23650 21922 23662
rect 22318 23714 22370 23726
rect 22318 23650 22370 23662
rect 22766 23714 22818 23726
rect 22766 23650 22818 23662
rect 23214 23714 23266 23726
rect 23214 23650 23266 23662
rect 23998 23714 24050 23726
rect 23998 23650 24050 23662
rect 25006 23714 25058 23726
rect 25006 23650 25058 23662
rect 26686 23714 26738 23726
rect 26686 23650 26738 23662
rect 28142 23714 28194 23726
rect 28142 23650 28194 23662
rect 1344 23546 28720 23580
rect 1344 23494 8018 23546
rect 8070 23494 8122 23546
rect 8174 23494 8226 23546
rect 8278 23494 14822 23546
rect 14874 23494 14926 23546
rect 14978 23494 15030 23546
rect 15082 23494 21626 23546
rect 21678 23494 21730 23546
rect 21782 23494 21834 23546
rect 21886 23494 28430 23546
rect 28482 23494 28534 23546
rect 28586 23494 28638 23546
rect 28690 23494 28720 23546
rect 1344 23460 28720 23494
rect 2046 23378 2098 23390
rect 2046 23314 2098 23326
rect 3166 23378 3218 23390
rect 3166 23314 3218 23326
rect 4622 23378 4674 23390
rect 4622 23314 4674 23326
rect 6974 23378 7026 23390
rect 6974 23314 7026 23326
rect 10894 23378 10946 23390
rect 10894 23314 10946 23326
rect 12686 23378 12738 23390
rect 12686 23314 12738 23326
rect 12798 23378 12850 23390
rect 12798 23314 12850 23326
rect 13246 23378 13298 23390
rect 13246 23314 13298 23326
rect 17614 23378 17666 23390
rect 17614 23314 17666 23326
rect 20078 23378 20130 23390
rect 20078 23314 20130 23326
rect 23214 23378 23266 23390
rect 23214 23314 23266 23326
rect 23662 23378 23714 23390
rect 23662 23314 23714 23326
rect 3838 23266 3890 23278
rect 3838 23202 3890 23214
rect 6638 23266 6690 23278
rect 22430 23266 22482 23278
rect 23774 23266 23826 23278
rect 7522 23214 7534 23266
rect 7586 23214 7598 23266
rect 8642 23214 8654 23266
rect 8706 23263 8718 23266
rect 8866 23263 8878 23266
rect 8706 23217 8878 23263
rect 8706 23214 8718 23217
rect 8866 23214 8878 23217
rect 8930 23214 8942 23266
rect 14242 23214 14254 23266
rect 14306 23214 14318 23266
rect 22642 23214 22654 23266
rect 22706 23214 22718 23266
rect 6638 23202 6690 23214
rect 22430 23202 22482 23214
rect 23774 23202 23826 23214
rect 1710 23154 1762 23166
rect 1710 23090 1762 23102
rect 3390 23154 3442 23166
rect 7758 23154 7810 23166
rect 20526 23154 20578 23166
rect 23998 23154 24050 23166
rect 4498 23102 4510 23154
rect 4562 23102 4574 23154
rect 7186 23102 7198 23154
rect 7250 23102 7262 23154
rect 8530 23102 8542 23154
rect 8594 23102 8606 23154
rect 12226 23102 12238 23154
rect 12290 23102 12302 23154
rect 12450 23102 12462 23154
rect 12514 23102 12526 23154
rect 13570 23102 13582 23154
rect 13634 23102 13646 23154
rect 20738 23102 20750 23154
rect 20802 23102 20814 23154
rect 22978 23102 22990 23154
rect 23042 23102 23054 23154
rect 24210 23102 24222 23154
rect 24274 23102 24286 23154
rect 27346 23102 27358 23154
rect 27410 23102 27422 23154
rect 28018 23102 28030 23154
rect 28082 23102 28094 23154
rect 3390 23090 3442 23102
rect 7758 23090 7810 23102
rect 20526 23090 20578 23102
rect 23998 23090 24050 23102
rect 2718 23042 2770 23054
rect 2718 22978 2770 22990
rect 5518 23042 5570 23054
rect 5518 22978 5570 22990
rect 6190 23042 6242 23054
rect 6190 22978 6242 22990
rect 8318 23042 8370 23054
rect 8318 22978 8370 22990
rect 8990 23042 9042 23054
rect 8990 22978 9042 22990
rect 11902 23042 11954 23054
rect 16830 23042 16882 23054
rect 16370 22990 16382 23042
rect 16434 22990 16446 23042
rect 11902 22978 11954 22990
rect 16830 22978 16882 22990
rect 17950 23042 18002 23054
rect 17950 22978 18002 22990
rect 18622 23042 18674 23054
rect 18622 22978 18674 22990
rect 19070 23042 19122 23054
rect 19070 22978 19122 22990
rect 19518 23042 19570 23054
rect 19518 22978 19570 22990
rect 21198 23042 21250 23054
rect 21198 22978 21250 22990
rect 21870 23042 21922 23054
rect 21870 22978 21922 22990
rect 23886 23042 23938 23054
rect 23886 22978 23938 22990
rect 24670 23042 24722 23054
rect 25218 22990 25230 23042
rect 25282 22990 25294 23042
rect 24670 22978 24722 22990
rect 3054 22930 3106 22942
rect 3054 22866 3106 22878
rect 3726 22930 3778 22942
rect 3726 22866 3778 22878
rect 7310 22930 7362 22942
rect 7310 22866 7362 22878
rect 8206 22930 8258 22942
rect 20414 22930 20466 22942
rect 18610 22878 18622 22930
rect 18674 22927 18686 22930
rect 18946 22927 18958 22930
rect 18674 22881 18958 22927
rect 18674 22878 18686 22881
rect 18946 22878 18958 22881
rect 19010 22878 19022 22930
rect 21858 22878 21870 22930
rect 21922 22927 21934 22930
rect 22194 22927 22206 22930
rect 21922 22881 22206 22927
rect 21922 22878 21934 22881
rect 22194 22878 22206 22881
rect 22258 22878 22270 22930
rect 22978 22878 22990 22930
rect 23042 22878 23054 22930
rect 8206 22866 8258 22878
rect 20414 22866 20466 22878
rect 1344 22762 28560 22796
rect 1344 22710 4616 22762
rect 4668 22710 4720 22762
rect 4772 22710 4824 22762
rect 4876 22710 11420 22762
rect 11472 22710 11524 22762
rect 11576 22710 11628 22762
rect 11680 22710 18224 22762
rect 18276 22710 18328 22762
rect 18380 22710 18432 22762
rect 18484 22710 25028 22762
rect 25080 22710 25132 22762
rect 25184 22710 25236 22762
rect 25288 22710 28560 22762
rect 1344 22676 28560 22710
rect 20178 22542 20190 22594
rect 20242 22542 20254 22594
rect 8878 22482 8930 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 8878 22418 8930 22430
rect 10222 22482 10274 22494
rect 10222 22418 10274 22430
rect 11006 22482 11058 22494
rect 11006 22418 11058 22430
rect 13022 22482 13074 22494
rect 13022 22418 13074 22430
rect 13694 22482 13746 22494
rect 13694 22418 13746 22430
rect 15710 22482 15762 22494
rect 15710 22418 15762 22430
rect 16606 22482 16658 22494
rect 16606 22418 16658 22430
rect 18622 22482 18674 22494
rect 18622 22418 18674 22430
rect 21870 22482 21922 22494
rect 21870 22418 21922 22430
rect 22318 22482 22370 22494
rect 22318 22418 22370 22430
rect 24558 22482 24610 22494
rect 24558 22418 24610 22430
rect 25006 22482 25058 22494
rect 26898 22430 26910 22482
rect 26962 22430 26974 22482
rect 25006 22418 25058 22430
rect 15822 22370 15874 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 15822 22306 15874 22318
rect 17054 22370 17106 22382
rect 17054 22306 17106 22318
rect 19070 22370 19122 22382
rect 19842 22318 19854 22370
rect 19906 22318 19918 22370
rect 20290 22318 20302 22370
rect 20354 22318 20366 22370
rect 23202 22318 23214 22370
rect 23266 22318 23278 22370
rect 23650 22318 23662 22370
rect 23714 22318 23726 22370
rect 25218 22318 25230 22370
rect 25282 22318 25294 22370
rect 26002 22318 26014 22370
rect 26066 22318 26078 22370
rect 19070 22306 19122 22318
rect 10446 22258 10498 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 10446 22194 10498 22206
rect 16046 22258 16098 22270
rect 16046 22194 16098 22206
rect 19630 22258 19682 22270
rect 24894 22258 24946 22270
rect 23986 22206 23998 22258
rect 24050 22206 24062 22258
rect 19630 22194 19682 22206
rect 24894 22194 24946 22206
rect 5070 22146 5122 22158
rect 5070 22082 5122 22094
rect 7982 22146 8034 22158
rect 7982 22082 8034 22094
rect 10334 22146 10386 22158
rect 10334 22082 10386 22094
rect 15598 22146 15650 22158
rect 15598 22082 15650 22094
rect 17502 22146 17554 22158
rect 17502 22082 17554 22094
rect 18174 22146 18226 22158
rect 18174 22082 18226 22094
rect 19742 22146 19794 22158
rect 19742 22082 19794 22094
rect 21422 22146 21474 22158
rect 21422 22082 21474 22094
rect 22878 22146 22930 22158
rect 22978 22094 22990 22146
rect 23042 22094 23054 22146
rect 22878 22082 22930 22094
rect 1344 21978 28720 22012
rect 1344 21926 8018 21978
rect 8070 21926 8122 21978
rect 8174 21926 8226 21978
rect 8278 21926 14822 21978
rect 14874 21926 14926 21978
rect 14978 21926 15030 21978
rect 15082 21926 21626 21978
rect 21678 21926 21730 21978
rect 21782 21926 21834 21978
rect 21886 21926 28430 21978
rect 28482 21926 28534 21978
rect 28586 21926 28638 21978
rect 28690 21926 28720 21978
rect 1344 21892 28720 21926
rect 2718 21810 2770 21822
rect 2718 21746 2770 21758
rect 3950 21810 4002 21822
rect 3950 21746 4002 21758
rect 4398 21810 4450 21822
rect 4398 21746 4450 21758
rect 12910 21810 12962 21822
rect 12910 21746 12962 21758
rect 13358 21810 13410 21822
rect 13358 21746 13410 21758
rect 17950 21810 18002 21822
rect 17950 21746 18002 21758
rect 24334 21810 24386 21822
rect 24334 21746 24386 21758
rect 2046 21698 2098 21710
rect 8430 21698 8482 21710
rect 3266 21646 3278 21698
rect 3330 21646 3342 21698
rect 2046 21634 2098 21646
rect 8430 21634 8482 21646
rect 8654 21698 8706 21710
rect 8654 21634 8706 21646
rect 14478 21698 14530 21710
rect 24222 21698 24274 21710
rect 19730 21646 19742 21698
rect 19794 21646 19806 21698
rect 14478 21634 14530 21646
rect 24222 21634 24274 21646
rect 3054 21586 3106 21598
rect 1810 21534 1822 21586
rect 1874 21534 1886 21586
rect 2706 21534 2718 21586
rect 2770 21534 2782 21586
rect 3054 21522 3106 21534
rect 3502 21586 3554 21598
rect 17614 21586 17666 21598
rect 5058 21534 5070 21586
rect 5122 21534 5134 21586
rect 9650 21534 9662 21586
rect 9714 21534 9726 21586
rect 18946 21534 18958 21586
rect 19010 21534 19022 21586
rect 22754 21534 22766 21586
rect 22818 21534 22830 21586
rect 26002 21534 26014 21586
rect 26066 21534 26078 21586
rect 3502 21522 3554 21534
rect 17614 21522 17666 21534
rect 14254 21474 14306 21486
rect 5842 21422 5854 21474
rect 5906 21422 5918 21474
rect 7970 21422 7982 21474
rect 8034 21422 8046 21474
rect 10322 21422 10334 21474
rect 10386 21422 10398 21474
rect 12450 21422 12462 21474
rect 12514 21422 12526 21474
rect 14254 21410 14306 21422
rect 14366 21474 14418 21486
rect 14366 21410 14418 21422
rect 15038 21474 15090 21486
rect 15038 21410 15090 21422
rect 15486 21474 15538 21486
rect 15486 21410 15538 21422
rect 18398 21474 18450 21486
rect 21858 21422 21870 21474
rect 21922 21422 21934 21474
rect 23426 21422 23438 21474
rect 23490 21422 23502 21474
rect 27010 21422 27022 21474
rect 27074 21422 27086 21474
rect 18398 21410 18450 21422
rect 8318 21362 8370 21374
rect 8318 21298 8370 21310
rect 24446 21362 24498 21374
rect 24446 21298 24498 21310
rect 1344 21194 28560 21228
rect 1344 21142 4616 21194
rect 4668 21142 4720 21194
rect 4772 21142 4824 21194
rect 4876 21142 11420 21194
rect 11472 21142 11524 21194
rect 11576 21142 11628 21194
rect 11680 21142 18224 21194
rect 18276 21142 18328 21194
rect 18380 21142 18432 21194
rect 18484 21142 25028 21194
rect 25080 21142 25132 21194
rect 25184 21142 25236 21194
rect 25288 21142 28560 21194
rect 1344 21108 28560 21142
rect 3054 21026 3106 21038
rect 6862 21026 6914 21038
rect 11006 21026 11058 21038
rect 4274 21023 4286 21026
rect 3054 20962 3106 20974
rect 3841 20977 4286 21023
rect 1822 20914 1874 20926
rect 1822 20850 1874 20862
rect 2382 20914 2434 20926
rect 2382 20850 2434 20862
rect 3502 20802 3554 20814
rect 2706 20750 2718 20802
rect 2770 20750 2782 20802
rect 3602 20750 3614 20802
rect 3666 20799 3678 20802
rect 3841 20799 3887 20977
rect 4274 20974 4286 20977
rect 4338 21023 4350 21026
rect 4834 21023 4846 21026
rect 4338 20977 4846 21023
rect 4338 20974 4350 20977
rect 4834 20974 4846 20977
rect 4898 20974 4910 21026
rect 5842 20974 5854 21026
rect 5906 21023 5918 21026
rect 6402 21023 6414 21026
rect 5906 20977 6414 21023
rect 5906 20974 5918 20977
rect 6402 20974 6414 20977
rect 6466 20974 6478 21026
rect 9986 20974 9998 21026
rect 10050 20974 10062 21026
rect 6862 20962 6914 20974
rect 11006 20962 11058 20974
rect 11678 21026 11730 21038
rect 11678 20962 11730 20974
rect 12014 21026 12066 21038
rect 20078 21026 20130 21038
rect 27134 21026 27186 21038
rect 12226 20974 12238 21026
rect 12290 21023 12302 21026
rect 12450 21023 12462 21026
rect 12290 20977 12462 21023
rect 12290 20974 12302 20977
rect 12450 20974 12462 20977
rect 12514 20974 12526 21026
rect 14018 20974 14030 21026
rect 14082 20974 14094 21026
rect 19506 20974 19518 21026
rect 19570 20974 19582 21026
rect 26338 20974 26350 21026
rect 26402 20974 26414 21026
rect 12014 20962 12066 20974
rect 20078 20962 20130 20974
rect 27134 20962 27186 20974
rect 27470 21026 27522 21038
rect 27470 20962 27522 20974
rect 4846 20914 4898 20926
rect 4846 20850 4898 20862
rect 8206 20914 8258 20926
rect 8206 20850 8258 20862
rect 9102 20914 9154 20926
rect 9102 20850 9154 20862
rect 12462 20914 12514 20926
rect 12462 20850 12514 20862
rect 12910 20914 12962 20926
rect 12910 20850 12962 20862
rect 14926 20914 14978 20926
rect 18610 20862 18622 20914
rect 18674 20862 18686 20914
rect 23314 20862 23326 20914
rect 23378 20862 23390 20914
rect 25442 20862 25454 20914
rect 25506 20862 25518 20914
rect 14926 20850 14978 20862
rect 8654 20802 8706 20814
rect 3666 20753 3887 20799
rect 3666 20750 3678 20753
rect 6626 20750 6638 20802
rect 6690 20750 6702 20802
rect 3502 20738 3554 20750
rect 8654 20738 8706 20750
rect 9774 20802 9826 20814
rect 18958 20802 19010 20814
rect 26126 20802 26178 20814
rect 10210 20750 10222 20802
rect 10274 20750 10286 20802
rect 10770 20750 10782 20802
rect 10834 20750 10846 20802
rect 11330 20750 11342 20802
rect 11394 20750 11406 20802
rect 14242 20750 14254 20802
rect 14306 20750 14318 20802
rect 15810 20750 15822 20802
rect 15874 20750 15886 20802
rect 19170 20750 19182 20802
rect 19234 20750 19246 20802
rect 19506 20750 19518 20802
rect 19570 20750 19582 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 22642 20750 22654 20802
rect 22706 20750 22718 20802
rect 26338 20750 26350 20802
rect 26402 20750 26414 20802
rect 27122 20750 27134 20802
rect 27186 20750 27198 20802
rect 9774 20738 9826 20750
rect 18958 20738 19010 20750
rect 26126 20738 26178 20750
rect 6190 20690 6242 20702
rect 7310 20690 7362 20702
rect 7074 20638 7086 20690
rect 7138 20638 7150 20690
rect 6190 20626 6242 20638
rect 7310 20626 7362 20638
rect 7758 20690 7810 20702
rect 7758 20626 7810 20638
rect 9438 20690 9490 20702
rect 9438 20626 9490 20638
rect 10558 20690 10610 20702
rect 10558 20626 10610 20638
rect 11790 20690 11842 20702
rect 11790 20626 11842 20638
rect 13470 20690 13522 20702
rect 20414 20690 20466 20702
rect 13682 20638 13694 20690
rect 13746 20638 13758 20690
rect 16482 20638 16494 20690
rect 16546 20638 16558 20690
rect 13470 20626 13522 20638
rect 20414 20626 20466 20638
rect 25790 20690 25842 20702
rect 25790 20626 25842 20638
rect 2942 20578 2994 20590
rect 2942 20514 2994 20526
rect 3390 20578 3442 20590
rect 3390 20514 3442 20526
rect 3950 20578 4002 20590
rect 3950 20514 4002 20526
rect 4398 20578 4450 20590
rect 4398 20514 4450 20526
rect 5742 20578 5794 20590
rect 5742 20514 5794 20526
rect 6526 20578 6578 20590
rect 6526 20514 6578 20526
rect 10222 20578 10274 20590
rect 10222 20514 10274 20526
rect 10670 20578 10722 20590
rect 10670 20514 10722 20526
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 15374 20578 15426 20590
rect 15374 20514 15426 20526
rect 19070 20578 19122 20590
rect 19070 20514 19122 20526
rect 21422 20578 21474 20590
rect 21422 20514 21474 20526
rect 22094 20578 22146 20590
rect 22094 20514 22146 20526
rect 25902 20578 25954 20590
rect 25902 20514 25954 20526
rect 27918 20578 27970 20590
rect 27918 20514 27970 20526
rect 1344 20410 28720 20444
rect 1344 20358 8018 20410
rect 8070 20358 8122 20410
rect 8174 20358 8226 20410
rect 8278 20358 14822 20410
rect 14874 20358 14926 20410
rect 14978 20358 15030 20410
rect 15082 20358 21626 20410
rect 21678 20358 21730 20410
rect 21782 20358 21834 20410
rect 21886 20358 28430 20410
rect 28482 20358 28534 20410
rect 28586 20358 28638 20410
rect 28690 20358 28720 20410
rect 1344 20324 28720 20358
rect 2494 20242 2546 20254
rect 2494 20178 2546 20190
rect 7198 20242 7250 20254
rect 7198 20178 7250 20190
rect 10446 20242 10498 20254
rect 10446 20178 10498 20190
rect 11454 20242 11506 20254
rect 23102 20242 23154 20254
rect 11666 20190 11678 20242
rect 11730 20239 11742 20242
rect 11730 20193 11839 20239
rect 11730 20190 11742 20193
rect 11454 20178 11506 20190
rect 3278 20130 3330 20142
rect 3042 20078 3054 20130
rect 3106 20078 3118 20130
rect 3278 20066 3330 20078
rect 5406 20130 5458 20142
rect 5406 20066 5458 20078
rect 8878 20130 8930 20142
rect 8878 20066 8930 20078
rect 9998 20130 10050 20142
rect 9998 20066 10050 20078
rect 2830 20018 2882 20030
rect 2594 19966 2606 20018
rect 2658 19966 2670 20018
rect 3938 19966 3950 20018
rect 4002 19966 4014 20018
rect 2830 19954 2882 19966
rect 4958 19906 5010 19918
rect 4958 19842 5010 19854
rect 8318 19906 8370 19918
rect 8318 19842 8370 19854
rect 4498 19742 4510 19794
rect 4562 19742 4574 19794
rect 11793 19791 11839 20193
rect 16482 20190 16494 20242
rect 16546 20190 16558 20242
rect 23102 20178 23154 20190
rect 11902 20130 11954 20142
rect 15710 20130 15762 20142
rect 13010 20078 13022 20130
rect 13074 20078 13086 20130
rect 11902 20066 11954 20078
rect 15710 20066 15762 20078
rect 16046 20130 16098 20142
rect 16046 20066 16098 20078
rect 23662 20130 23714 20142
rect 23662 20066 23714 20078
rect 24670 20130 24722 20142
rect 26002 20078 26014 20130
rect 26066 20078 26078 20130
rect 24670 20066 24722 20078
rect 12338 19966 12350 20018
rect 12402 19966 12414 20018
rect 16258 19966 16270 20018
rect 16322 19966 16334 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 17602 19966 17614 20018
rect 17666 19966 17678 20018
rect 25330 19966 25342 20018
rect 25394 19966 25406 20018
rect 24110 19906 24162 19918
rect 15138 19854 15150 19906
rect 15202 19854 15214 19906
rect 19394 19854 19406 19906
rect 19458 19854 19470 19906
rect 28130 19854 28142 19906
rect 28194 19854 28206 19906
rect 24110 19842 24162 19854
rect 11890 19791 11902 19794
rect 11793 19745 11902 19791
rect 11890 19742 11902 19745
rect 11954 19742 11966 19794
rect 16594 19742 16606 19794
rect 16658 19742 16670 19794
rect 1344 19626 28560 19660
rect 1344 19574 4616 19626
rect 4668 19574 4720 19626
rect 4772 19574 4824 19626
rect 4876 19574 11420 19626
rect 11472 19574 11524 19626
rect 11576 19574 11628 19626
rect 11680 19574 18224 19626
rect 18276 19574 18328 19626
rect 18380 19574 18432 19626
rect 18484 19574 25028 19626
rect 25080 19574 25132 19626
rect 25184 19574 25236 19626
rect 25288 19574 28560 19626
rect 1344 19540 28560 19574
rect 18174 19458 18226 19470
rect 18174 19394 18226 19406
rect 8654 19346 8706 19358
rect 12462 19346 12514 19358
rect 2482 19294 2494 19346
rect 2546 19294 2558 19346
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 9762 19294 9774 19346
rect 9826 19294 9838 19346
rect 11890 19294 11902 19346
rect 11954 19294 11966 19346
rect 8654 19282 8706 19294
rect 12462 19282 12514 19294
rect 12910 19346 12962 19358
rect 17054 19346 17106 19358
rect 15362 19294 15374 19346
rect 15426 19294 15438 19346
rect 12910 19282 12962 19294
rect 17054 19282 17106 19294
rect 18286 19346 18338 19358
rect 18286 19282 18338 19294
rect 20526 19346 20578 19358
rect 20526 19282 20578 19294
rect 22654 19346 22706 19358
rect 27022 19346 27074 19358
rect 23090 19294 23102 19346
rect 23154 19294 23166 19346
rect 22654 19282 22706 19294
rect 27022 19282 27074 19294
rect 28030 19346 28082 19358
rect 28030 19282 28082 19294
rect 6078 19234 6130 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 6078 19170 6130 19182
rect 6414 19234 6466 19246
rect 6414 19170 6466 19182
rect 6638 19234 6690 19246
rect 6638 19170 6690 19182
rect 7758 19234 7810 19246
rect 7758 19170 7810 19182
rect 8206 19234 8258 19246
rect 13358 19234 13410 19246
rect 8978 19182 8990 19234
rect 9042 19182 9054 19234
rect 8206 19170 8258 19182
rect 13358 19170 13410 19182
rect 13806 19234 13858 19246
rect 13806 19170 13858 19182
rect 13918 19234 13970 19246
rect 16494 19234 16546 19246
rect 19518 19234 19570 19246
rect 14578 19182 14590 19234
rect 14642 19182 14654 19234
rect 16034 19182 16046 19234
rect 16098 19182 16110 19234
rect 18498 19182 18510 19234
rect 18562 19182 18574 19234
rect 13918 19170 13970 19182
rect 16494 19170 16546 19182
rect 19518 19170 19570 19182
rect 19742 19234 19794 19246
rect 21646 19234 21698 19246
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 19742 19170 19794 19182
rect 21646 19170 21698 19182
rect 21870 19234 21922 19246
rect 21870 19170 21922 19182
rect 22318 19234 22370 19246
rect 25890 19182 25902 19234
rect 25954 19182 25966 19234
rect 22318 19170 22370 19182
rect 6974 19122 7026 19134
rect 21758 19122 21810 19134
rect 15586 19070 15598 19122
rect 15650 19070 15662 19122
rect 25218 19070 25230 19122
rect 25282 19070 25294 19122
rect 6974 19058 7026 19070
rect 21758 19058 21810 19070
rect 5070 19010 5122 19022
rect 5070 18946 5122 18958
rect 6526 19010 6578 19022
rect 6526 18946 6578 18958
rect 7534 19010 7586 19022
rect 7534 18946 7586 18958
rect 7646 19010 7698 19022
rect 7646 18946 7698 18958
rect 13582 19010 13634 19022
rect 17502 19010 17554 19022
rect 14690 18958 14702 19010
rect 14754 18958 14766 19010
rect 13582 18946 13634 18958
rect 17502 18946 17554 18958
rect 18958 19010 19010 19022
rect 18958 18946 19010 18958
rect 19630 19010 19682 19022
rect 19630 18946 19682 18958
rect 26462 19010 26514 19022
rect 26462 18946 26514 18958
rect 27358 19010 27410 19022
rect 27358 18946 27410 18958
rect 1344 18842 28720 18876
rect 1344 18790 8018 18842
rect 8070 18790 8122 18842
rect 8174 18790 8226 18842
rect 8278 18790 14822 18842
rect 14874 18790 14926 18842
rect 14978 18790 15030 18842
rect 15082 18790 21626 18842
rect 21678 18790 21730 18842
rect 21782 18790 21834 18842
rect 21886 18790 28430 18842
rect 28482 18790 28534 18842
rect 28586 18790 28638 18842
rect 28690 18790 28720 18842
rect 1344 18756 28720 18790
rect 3278 18674 3330 18686
rect 3278 18610 3330 18622
rect 8990 18674 9042 18686
rect 8990 18610 9042 18622
rect 25342 18674 25394 18686
rect 25342 18610 25394 18622
rect 26126 18674 26178 18686
rect 26126 18610 26178 18622
rect 26350 18674 26402 18686
rect 26350 18610 26402 18622
rect 2046 18562 2098 18574
rect 5954 18510 5966 18562
rect 6018 18510 6030 18562
rect 2046 18498 2098 18510
rect 1710 18450 1762 18462
rect 1710 18386 1762 18398
rect 3726 18450 3778 18462
rect 8542 18450 8594 18462
rect 24670 18450 24722 18462
rect 5170 18398 5182 18450
rect 5234 18398 5246 18450
rect 11554 18398 11566 18450
rect 11618 18398 11630 18450
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 19170 18398 19182 18450
rect 19234 18398 19246 18450
rect 23986 18398 23998 18450
rect 24050 18398 24062 18450
rect 3726 18386 3778 18398
rect 8542 18386 8594 18398
rect 24670 18386 24722 18398
rect 25230 18450 25282 18462
rect 25230 18386 25282 18398
rect 25454 18450 25506 18462
rect 25454 18386 25506 18398
rect 25678 18450 25730 18462
rect 25678 18386 25730 18398
rect 26238 18450 26290 18462
rect 26238 18386 26290 18398
rect 26798 18450 26850 18462
rect 26798 18386 26850 18398
rect 28030 18450 28082 18462
rect 28030 18386 28082 18398
rect 2494 18338 2546 18350
rect 11230 18338 11282 18350
rect 17502 18338 17554 18350
rect 8082 18286 8094 18338
rect 8146 18286 8158 18338
rect 13570 18286 13582 18338
rect 13634 18286 13646 18338
rect 2494 18274 2546 18286
rect 11230 18274 11282 18286
rect 17502 18274 17554 18286
rect 17950 18338 18002 18350
rect 27134 18338 27186 18350
rect 21298 18286 21310 18338
rect 21362 18286 21374 18338
rect 22194 18286 22206 18338
rect 22258 18286 22270 18338
rect 17950 18274 18002 18286
rect 27134 18274 27186 18286
rect 27582 18338 27634 18350
rect 27582 18274 27634 18286
rect 27122 18174 27134 18226
rect 27186 18223 27198 18226
rect 27794 18223 27806 18226
rect 27186 18177 27806 18223
rect 27186 18174 27198 18177
rect 27794 18174 27806 18177
rect 27858 18174 27870 18226
rect 1344 18058 28560 18092
rect 1344 18006 4616 18058
rect 4668 18006 4720 18058
rect 4772 18006 4824 18058
rect 4876 18006 11420 18058
rect 11472 18006 11524 18058
rect 11576 18006 11628 18058
rect 11680 18006 18224 18058
rect 18276 18006 18328 18058
rect 18380 18006 18432 18058
rect 18484 18006 25028 18058
rect 25080 18006 25132 18058
rect 25184 18006 25236 18058
rect 25288 18006 28560 18058
rect 1344 17972 28560 18006
rect 2718 17890 2770 17902
rect 12674 17838 12686 17890
rect 12738 17887 12750 17890
rect 12898 17887 12910 17890
rect 12738 17841 12910 17887
rect 12738 17838 12750 17841
rect 12898 17838 12910 17841
rect 12962 17838 12974 17890
rect 2718 17826 2770 17838
rect 3502 17778 3554 17790
rect 8990 17778 9042 17790
rect 8530 17726 8542 17778
rect 8594 17726 8606 17778
rect 3502 17714 3554 17726
rect 8990 17714 9042 17726
rect 10110 17778 10162 17790
rect 10110 17714 10162 17726
rect 12910 17778 12962 17790
rect 12910 17714 12962 17726
rect 13918 17778 13970 17790
rect 16942 17778 16994 17790
rect 27582 17778 27634 17790
rect 15250 17726 15262 17778
rect 15314 17726 15326 17778
rect 20738 17726 20750 17778
rect 20802 17726 20814 17778
rect 21298 17726 21310 17778
rect 21362 17726 21374 17778
rect 25218 17726 25230 17778
rect 25282 17726 25294 17778
rect 13918 17714 13970 17726
rect 16942 17714 16994 17726
rect 27582 17714 27634 17726
rect 10446 17666 10498 17678
rect 4162 17614 4174 17666
rect 4226 17614 4238 17666
rect 5730 17614 5742 17666
rect 5794 17614 5806 17666
rect 10446 17602 10498 17614
rect 10782 17666 10834 17678
rect 10782 17602 10834 17614
rect 11006 17666 11058 17678
rect 11006 17602 11058 17614
rect 11566 17666 11618 17678
rect 11566 17602 11618 17614
rect 11678 17666 11730 17678
rect 14030 17666 14082 17678
rect 12002 17614 12014 17666
rect 12066 17614 12078 17666
rect 11678 17602 11730 17614
rect 14030 17602 14082 17614
rect 14926 17666 14978 17678
rect 15934 17666 15986 17678
rect 15362 17614 15374 17666
rect 15426 17614 15438 17666
rect 14926 17602 14978 17614
rect 15934 17602 15986 17614
rect 16494 17666 16546 17678
rect 16494 17602 16546 17614
rect 17054 17666 17106 17678
rect 17826 17614 17838 17666
rect 17890 17614 17902 17666
rect 24098 17614 24110 17666
rect 24162 17614 24174 17666
rect 26562 17614 26574 17666
rect 26626 17614 26638 17666
rect 17054 17602 17106 17614
rect 2942 17554 2994 17566
rect 13806 17554 13858 17566
rect 6402 17502 6414 17554
rect 6466 17502 6478 17554
rect 2942 17490 2994 17502
rect 13806 17490 13858 17502
rect 14702 17554 14754 17566
rect 14702 17490 14754 17502
rect 16270 17554 16322 17566
rect 18610 17502 18622 17554
rect 18674 17502 18686 17554
rect 23426 17502 23438 17554
rect 23490 17502 23502 17554
rect 16270 17490 16322 17502
rect 2830 17442 2882 17454
rect 2830 17378 2882 17390
rect 3390 17442 3442 17454
rect 9438 17442 9490 17454
rect 4722 17390 4734 17442
rect 4786 17390 4798 17442
rect 3390 17378 3442 17390
rect 9438 17378 9490 17390
rect 10558 17442 10610 17454
rect 10558 17378 10610 17390
rect 11454 17442 11506 17454
rect 11454 17378 11506 17390
rect 12462 17442 12514 17454
rect 12462 17378 12514 17390
rect 14254 17442 14306 17454
rect 14254 17378 14306 17390
rect 15150 17442 15202 17454
rect 15150 17378 15202 17390
rect 16046 17442 16098 17454
rect 16046 17378 16098 17390
rect 16830 17442 16882 17454
rect 16830 17378 16882 17390
rect 17278 17442 17330 17454
rect 17278 17378 17330 17390
rect 28030 17442 28082 17454
rect 28030 17378 28082 17390
rect 1344 17274 28720 17308
rect 1344 17222 8018 17274
rect 8070 17222 8122 17274
rect 8174 17222 8226 17274
rect 8278 17222 14822 17274
rect 14874 17222 14926 17274
rect 14978 17222 15030 17274
rect 15082 17222 21626 17274
rect 21678 17222 21730 17274
rect 21782 17222 21834 17274
rect 21886 17222 28430 17274
rect 28482 17222 28534 17274
rect 28586 17222 28638 17274
rect 28690 17222 28720 17274
rect 1344 17188 28720 17222
rect 5070 17106 5122 17118
rect 5070 17042 5122 17054
rect 6526 17106 6578 17118
rect 6526 17042 6578 17054
rect 7646 17106 7698 17118
rect 7646 17042 7698 17054
rect 7870 17106 7922 17118
rect 7870 17042 7922 17054
rect 8990 17106 9042 17118
rect 8990 17042 9042 17054
rect 9662 17106 9714 17118
rect 9662 17042 9714 17054
rect 10334 17106 10386 17118
rect 10334 17042 10386 17054
rect 11230 17106 11282 17118
rect 11230 17042 11282 17054
rect 11678 17106 11730 17118
rect 11678 17042 11730 17054
rect 15934 17106 15986 17118
rect 15934 17042 15986 17054
rect 16718 17106 16770 17118
rect 16718 17042 16770 17054
rect 18062 17106 18114 17118
rect 18062 17042 18114 17054
rect 18510 17106 18562 17118
rect 18510 17042 18562 17054
rect 18958 17106 19010 17118
rect 18958 17042 19010 17054
rect 20302 17106 20354 17118
rect 20302 17042 20354 17054
rect 20750 17106 20802 17118
rect 20750 17042 20802 17054
rect 21310 17106 21362 17118
rect 21310 17042 21362 17054
rect 23102 17106 23154 17118
rect 23102 17042 23154 17054
rect 23550 17106 23602 17118
rect 23550 17042 23602 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 24670 17106 24722 17118
rect 24670 17042 24722 17054
rect 6974 16994 7026 17006
rect 6974 16930 7026 16942
rect 7758 16994 7810 17006
rect 16270 16994 16322 17006
rect 12786 16942 12798 16994
rect 12850 16942 12862 16994
rect 7758 16930 7810 16942
rect 16270 16930 16322 16942
rect 18846 16994 18898 17006
rect 18846 16930 18898 16942
rect 19182 16994 19234 17006
rect 19182 16930 19234 16942
rect 19406 16994 19458 17006
rect 19406 16930 19458 16942
rect 21198 16994 21250 17006
rect 21198 16930 21250 16942
rect 22654 16994 22706 17006
rect 26338 16942 26350 16994
rect 26402 16942 26414 16994
rect 22654 16930 22706 16942
rect 6078 16882 6130 16894
rect 1810 16830 1822 16882
rect 1874 16830 1886 16882
rect 6078 16818 6130 16830
rect 6302 16882 6354 16894
rect 6302 16818 6354 16830
rect 6750 16882 6802 16894
rect 6750 16818 6802 16830
rect 8318 16882 8370 16894
rect 8318 16818 8370 16830
rect 10782 16882 10834 16894
rect 15374 16882 15426 16894
rect 12114 16830 12126 16882
rect 12178 16830 12190 16882
rect 10782 16818 10834 16830
rect 15374 16818 15426 16830
rect 17614 16882 17666 16894
rect 17614 16818 17666 16830
rect 21534 16882 21586 16894
rect 21534 16818 21586 16830
rect 21646 16882 21698 16894
rect 21646 16818 21698 16830
rect 22206 16882 22258 16894
rect 27570 16830 27582 16882
rect 27634 16830 27646 16882
rect 22206 16818 22258 16830
rect 5630 16770 5682 16782
rect 19854 16770 19906 16782
rect 2482 16718 2494 16770
rect 2546 16718 2558 16770
rect 4610 16718 4622 16770
rect 4674 16718 4686 16770
rect 5282 16718 5294 16770
rect 5346 16718 5358 16770
rect 14914 16718 14926 16770
rect 14978 16718 14990 16770
rect 5297 16655 5343 16718
rect 5630 16706 5682 16718
rect 19854 16706 19906 16718
rect 6066 16655 6078 16658
rect 5297 16609 6078 16655
rect 6066 16606 6078 16609
rect 6130 16606 6142 16658
rect 15250 16606 15262 16658
rect 15314 16655 15326 16658
rect 16482 16655 16494 16658
rect 15314 16609 16494 16655
rect 15314 16606 15326 16609
rect 16482 16606 16494 16609
rect 16546 16606 16558 16658
rect 17266 16606 17278 16658
rect 17330 16655 17342 16658
rect 17826 16655 17838 16658
rect 17330 16609 17838 16655
rect 17330 16606 17342 16609
rect 17826 16606 17838 16609
rect 17890 16606 17902 16658
rect 22194 16606 22206 16658
rect 22258 16655 22270 16658
rect 23202 16655 23214 16658
rect 22258 16609 23214 16655
rect 22258 16606 22270 16609
rect 23202 16606 23214 16609
rect 23266 16606 23278 16658
rect 1344 16490 28560 16524
rect 1344 16438 4616 16490
rect 4668 16438 4720 16490
rect 4772 16438 4824 16490
rect 4876 16438 11420 16490
rect 11472 16438 11524 16490
rect 11576 16438 11628 16490
rect 11680 16438 18224 16490
rect 18276 16438 18328 16490
rect 18380 16438 18432 16490
rect 18484 16438 25028 16490
rect 25080 16438 25132 16490
rect 25184 16438 25236 16490
rect 25288 16438 28560 16490
rect 1344 16404 28560 16438
rect 2830 16322 2882 16334
rect 13570 16270 13582 16322
rect 13634 16319 13646 16322
rect 14130 16319 14142 16322
rect 13634 16273 14142 16319
rect 13634 16270 13646 16273
rect 14130 16270 14142 16273
rect 14194 16270 14206 16322
rect 2830 16258 2882 16270
rect 14142 16210 14194 16222
rect 8866 16158 8878 16210
rect 8930 16158 8942 16210
rect 14142 16146 14194 16158
rect 14590 16210 14642 16222
rect 18398 16210 18450 16222
rect 15810 16158 15822 16210
rect 15874 16158 15886 16210
rect 17938 16158 17950 16210
rect 18002 16158 18014 16210
rect 14590 16146 14642 16158
rect 18398 16146 18450 16158
rect 20750 16210 20802 16222
rect 27022 16210 27074 16222
rect 24098 16158 24110 16210
rect 24162 16158 24174 16210
rect 20750 16146 20802 16158
rect 27022 16146 27074 16158
rect 27582 16210 27634 16222
rect 27582 16146 27634 16158
rect 28142 16210 28194 16222
rect 28142 16146 28194 16158
rect 12574 16098 12626 16110
rect 20302 16098 20354 16110
rect 1810 16046 1822 16098
rect 1874 16046 1886 16098
rect 2594 16046 2606 16098
rect 2658 16046 2670 16098
rect 3042 16046 3054 16098
rect 3106 16046 3118 16098
rect 8194 16046 8206 16098
rect 8258 16046 8270 16098
rect 15138 16046 15150 16098
rect 15202 16046 15214 16098
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 12574 16034 12626 16046
rect 20302 16034 20354 16046
rect 3278 15986 3330 15998
rect 3278 15922 3330 15934
rect 12798 15986 12850 15998
rect 12798 15922 12850 15934
rect 2046 15874 2098 15886
rect 2046 15810 2098 15822
rect 2494 15874 2546 15886
rect 2494 15810 2546 15822
rect 3726 15874 3778 15886
rect 3726 15810 3778 15822
rect 4174 15874 4226 15886
rect 4174 15810 4226 15822
rect 12350 15874 12402 15886
rect 12350 15810 12402 15822
rect 12462 15874 12514 15886
rect 12462 15810 12514 15822
rect 13694 15874 13746 15886
rect 13694 15810 13746 15822
rect 1344 15706 28720 15740
rect 1344 15654 8018 15706
rect 8070 15654 8122 15706
rect 8174 15654 8226 15706
rect 8278 15654 14822 15706
rect 14874 15654 14926 15706
rect 14978 15654 15030 15706
rect 15082 15654 21626 15706
rect 21678 15654 21730 15706
rect 21782 15654 21834 15706
rect 21886 15654 28430 15706
rect 28482 15654 28534 15706
rect 28586 15654 28638 15706
rect 28690 15654 28720 15706
rect 1344 15620 28720 15654
rect 1822 15538 1874 15550
rect 1822 15474 1874 15486
rect 3054 15538 3106 15550
rect 3054 15474 3106 15486
rect 3502 15538 3554 15550
rect 3502 15474 3554 15486
rect 6078 15538 6130 15550
rect 6078 15474 6130 15486
rect 6526 15538 6578 15550
rect 6526 15474 6578 15486
rect 7758 15538 7810 15550
rect 7758 15474 7810 15486
rect 8990 15538 9042 15550
rect 8990 15474 9042 15486
rect 13022 15538 13074 15550
rect 13022 15474 13074 15486
rect 13358 15538 13410 15550
rect 13358 15474 13410 15486
rect 13582 15538 13634 15550
rect 13582 15474 13634 15486
rect 13806 15538 13858 15550
rect 13806 15474 13858 15486
rect 15374 15538 15426 15550
rect 15374 15474 15426 15486
rect 15598 15538 15650 15550
rect 15598 15474 15650 15486
rect 16158 15538 16210 15550
rect 16158 15474 16210 15486
rect 18958 15538 19010 15550
rect 18958 15474 19010 15486
rect 20638 15538 20690 15550
rect 20638 15474 20690 15486
rect 21758 15538 21810 15550
rect 21758 15474 21810 15486
rect 22206 15538 22258 15550
rect 22206 15474 22258 15486
rect 24222 15538 24274 15550
rect 24222 15474 24274 15486
rect 24334 15538 24386 15550
rect 24334 15474 24386 15486
rect 7422 15426 7474 15438
rect 14254 15426 14306 15438
rect 10322 15374 10334 15426
rect 10386 15374 10398 15426
rect 7422 15362 7474 15374
rect 14254 15362 14306 15374
rect 19742 15426 19794 15438
rect 19742 15362 19794 15374
rect 23774 15426 23826 15438
rect 23774 15362 23826 15374
rect 6862 15314 6914 15326
rect 6862 15250 6914 15262
rect 7982 15314 8034 15326
rect 14478 15314 14530 15326
rect 8306 15262 8318 15314
rect 8370 15262 8382 15314
rect 9650 15262 9662 15314
rect 9714 15262 9726 15314
rect 7982 15250 8034 15262
rect 14478 15250 14530 15262
rect 14814 15314 14866 15326
rect 14814 15250 14866 15262
rect 15150 15314 15202 15326
rect 15150 15250 15202 15262
rect 15262 15314 15314 15326
rect 15262 15250 15314 15262
rect 16606 15314 16658 15326
rect 16606 15250 16658 15262
rect 18734 15314 18786 15326
rect 20190 15314 20242 15326
rect 19282 15262 19294 15314
rect 19346 15262 19358 15314
rect 18734 15250 18786 15262
rect 20190 15250 20242 15262
rect 21982 15314 22034 15326
rect 21982 15250 22034 15262
rect 22654 15314 22706 15326
rect 22654 15250 22706 15262
rect 23214 15314 23266 15326
rect 23214 15250 23266 15262
rect 23326 15314 23378 15326
rect 23326 15250 23378 15262
rect 23550 15314 23602 15326
rect 23550 15250 23602 15262
rect 24110 15314 24162 15326
rect 24658 15262 24670 15314
rect 24722 15262 24734 15314
rect 25778 15262 25790 15314
rect 25842 15262 25854 15314
rect 24110 15250 24162 15262
rect 3950 15202 4002 15214
rect 3950 15138 4002 15150
rect 4398 15202 4450 15214
rect 4398 15138 4450 15150
rect 5630 15202 5682 15214
rect 5630 15138 5682 15150
rect 7870 15202 7922 15214
rect 13470 15202 13522 15214
rect 12450 15150 12462 15202
rect 12514 15150 12526 15202
rect 7870 15138 7922 15150
rect 13470 15138 13522 15150
rect 14366 15202 14418 15214
rect 14366 15138 14418 15150
rect 18846 15202 18898 15214
rect 18846 15138 18898 15150
rect 21198 15202 21250 15214
rect 21198 15138 21250 15150
rect 22094 15202 22146 15214
rect 26338 15150 26350 15202
rect 26402 15150 26414 15202
rect 22094 15138 22146 15150
rect 3154 15038 3166 15090
rect 3218 15087 3230 15090
rect 3938 15087 3950 15090
rect 3218 15041 3950 15087
rect 3218 15038 3230 15041
rect 3938 15038 3950 15041
rect 4002 15038 4014 15090
rect 1344 14922 28560 14956
rect 1344 14870 4616 14922
rect 4668 14870 4720 14922
rect 4772 14870 4824 14922
rect 4876 14870 11420 14922
rect 11472 14870 11524 14922
rect 11576 14870 11628 14922
rect 11680 14870 18224 14922
rect 18276 14870 18328 14922
rect 18380 14870 18432 14922
rect 18484 14870 25028 14922
rect 25080 14870 25132 14922
rect 25184 14870 25236 14922
rect 25288 14870 28560 14922
rect 1344 14836 28560 14870
rect 2046 14642 2098 14654
rect 20750 14642 20802 14654
rect 9426 14590 9438 14642
rect 9490 14590 9502 14642
rect 12674 14590 12686 14642
rect 12738 14590 12750 14642
rect 14354 14590 14366 14642
rect 14418 14590 14430 14642
rect 16482 14590 16494 14642
rect 16546 14590 16558 14642
rect 19842 14590 19854 14642
rect 19906 14590 19918 14642
rect 2046 14578 2098 14590
rect 20750 14578 20802 14590
rect 22430 14642 22482 14654
rect 27022 14642 27074 14654
rect 23538 14590 23550 14642
rect 23602 14590 23614 14642
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 22430 14578 22482 14590
rect 27022 14578 27074 14590
rect 27806 14642 27858 14654
rect 27806 14578 27858 14590
rect 28142 14642 28194 14654
rect 28142 14578 28194 14590
rect 2606 14530 2658 14542
rect 5070 14530 5122 14542
rect 2258 14478 2270 14530
rect 2322 14478 2334 14530
rect 3602 14478 3614 14530
rect 3666 14478 3678 14530
rect 2606 14466 2658 14478
rect 5070 14466 5122 14478
rect 5518 14530 5570 14542
rect 5518 14466 5570 14478
rect 6190 14530 6242 14542
rect 21198 14530 21250 14542
rect 6626 14478 6638 14530
rect 6690 14478 6702 14530
rect 9874 14478 9886 14530
rect 9938 14478 9950 14530
rect 13682 14478 13694 14530
rect 13746 14478 13758 14530
rect 17042 14478 17054 14530
rect 17106 14478 17118 14530
rect 6190 14466 6242 14478
rect 21198 14466 21250 14478
rect 21534 14530 21586 14542
rect 21534 14466 21586 14478
rect 21870 14530 21922 14542
rect 22754 14478 22766 14530
rect 22818 14478 22830 14530
rect 21870 14466 21922 14478
rect 3054 14418 3106 14430
rect 2818 14366 2830 14418
rect 2882 14366 2894 14418
rect 3054 14354 3106 14366
rect 4622 14418 4674 14430
rect 4622 14354 4674 14366
rect 5966 14418 6018 14430
rect 7298 14366 7310 14418
rect 7362 14366 7374 14418
rect 10546 14366 10558 14418
rect 10610 14366 10622 14418
rect 17714 14366 17726 14418
rect 17778 14366 17790 14418
rect 5966 14354 6018 14366
rect 5742 14306 5794 14318
rect 2594 14254 2606 14306
rect 2658 14254 2670 14306
rect 4162 14254 4174 14306
rect 4226 14254 4238 14306
rect 5742 14242 5794 14254
rect 20302 14306 20354 14318
rect 20302 14242 20354 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 26126 14306 26178 14318
rect 26126 14242 26178 14254
rect 26574 14306 26626 14318
rect 26574 14242 26626 14254
rect 1344 14138 28720 14172
rect 1344 14086 8018 14138
rect 8070 14086 8122 14138
rect 8174 14086 8226 14138
rect 8278 14086 14822 14138
rect 14874 14086 14926 14138
rect 14978 14086 15030 14138
rect 15082 14086 21626 14138
rect 21678 14086 21730 14138
rect 21782 14086 21834 14138
rect 21886 14086 28430 14138
rect 28482 14086 28534 14138
rect 28586 14086 28638 14138
rect 28690 14086 28720 14138
rect 1344 14052 28720 14086
rect 2270 13970 2322 13982
rect 2270 13906 2322 13918
rect 3278 13970 3330 13982
rect 3278 13906 3330 13918
rect 8542 13970 8594 13982
rect 8542 13906 8594 13918
rect 9662 13970 9714 13982
rect 9662 13906 9714 13918
rect 10670 13970 10722 13982
rect 10670 13906 10722 13918
rect 11566 13970 11618 13982
rect 11566 13906 11618 13918
rect 15262 13970 15314 13982
rect 15262 13906 15314 13918
rect 15710 13970 15762 13982
rect 15710 13906 15762 13918
rect 18174 13970 18226 13982
rect 18174 13906 18226 13918
rect 25454 13970 25506 13982
rect 25454 13906 25506 13918
rect 26686 13970 26738 13982
rect 26686 13906 26738 13918
rect 27134 13970 27186 13982
rect 27134 13906 27186 13918
rect 2718 13858 2770 13870
rect 8766 13858 8818 13870
rect 5282 13806 5294 13858
rect 5346 13806 5358 13858
rect 2718 13794 2770 13806
rect 8766 13794 8818 13806
rect 8990 13858 9042 13870
rect 8990 13794 9042 13806
rect 11118 13858 11170 13870
rect 11118 13794 11170 13806
rect 18622 13858 18674 13870
rect 18622 13794 18674 13806
rect 19070 13858 19122 13870
rect 20962 13806 20974 13858
rect 21026 13806 21038 13858
rect 19070 13794 19122 13806
rect 8094 13746 8146 13758
rect 4498 13694 4510 13746
rect 4562 13694 4574 13746
rect 8094 13682 8146 13694
rect 8318 13746 8370 13758
rect 8318 13682 8370 13694
rect 9550 13746 9602 13758
rect 9550 13682 9602 13694
rect 9774 13746 9826 13758
rect 10446 13746 10498 13758
rect 10098 13694 10110 13746
rect 10162 13694 10174 13746
rect 9774 13682 9826 13694
rect 10446 13682 10498 13694
rect 10782 13746 10834 13758
rect 17950 13746 18002 13758
rect 12002 13694 12014 13746
rect 12066 13694 12078 13746
rect 10782 13682 10834 13694
rect 17950 13682 18002 13694
rect 18398 13746 18450 13758
rect 23550 13746 23602 13758
rect 20178 13694 20190 13746
rect 20242 13694 20254 13746
rect 18398 13682 18450 13694
rect 23550 13682 23602 13694
rect 2494 13634 2546 13646
rect 3390 13634 3442 13646
rect 2818 13582 2830 13634
rect 2882 13582 2894 13634
rect 2494 13570 2546 13582
rect 3390 13570 3442 13582
rect 4174 13634 4226 13646
rect 17726 13634 17778 13646
rect 24222 13634 24274 13646
rect 7410 13582 7422 13634
rect 7474 13582 7486 13634
rect 12674 13582 12686 13634
rect 12738 13582 12750 13634
rect 14802 13582 14814 13634
rect 14866 13582 14878 13634
rect 23090 13582 23102 13634
rect 23154 13582 23166 13634
rect 4174 13570 4226 13582
rect 17726 13570 17778 13582
rect 24222 13570 24274 13582
rect 24670 13634 24722 13646
rect 24670 13570 24722 13582
rect 25790 13634 25842 13646
rect 25790 13570 25842 13582
rect 26238 13634 26290 13646
rect 26238 13570 26290 13582
rect 1344 13354 28560 13388
rect 1344 13302 4616 13354
rect 4668 13302 4720 13354
rect 4772 13302 4824 13354
rect 4876 13302 11420 13354
rect 11472 13302 11524 13354
rect 11576 13302 11628 13354
rect 11680 13302 18224 13354
rect 18276 13302 18328 13354
rect 18380 13302 18432 13354
rect 18484 13302 25028 13354
rect 25080 13302 25132 13354
rect 25184 13302 25236 13354
rect 25288 13302 28560 13354
rect 1344 13268 28560 13302
rect 12002 13134 12014 13186
rect 12066 13183 12078 13186
rect 12674 13183 12686 13186
rect 12066 13137 12686 13183
rect 12066 13134 12078 13137
rect 12674 13134 12686 13137
rect 12738 13183 12750 13186
rect 13010 13183 13022 13186
rect 12738 13137 13022 13183
rect 12738 13134 12750 13137
rect 13010 13134 13022 13137
rect 13074 13134 13086 13186
rect 14354 13134 14366 13186
rect 14418 13183 14430 13186
rect 15026 13183 15038 13186
rect 14418 13137 15038 13183
rect 14418 13134 14430 13137
rect 15026 13134 15038 13137
rect 15090 13134 15102 13186
rect 26450 13134 26462 13186
rect 26514 13183 26526 13186
rect 27010 13183 27022 13186
rect 26514 13137 27022 13183
rect 26514 13134 26526 13137
rect 27010 13134 27022 13137
rect 27074 13134 27086 13186
rect 5070 13074 5122 13086
rect 2482 13022 2494 13074
rect 2546 13022 2558 13074
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 5070 13010 5122 13022
rect 8094 13074 8146 13086
rect 8094 13010 8146 13022
rect 10894 13074 10946 13086
rect 10894 13010 10946 13022
rect 11342 13074 11394 13086
rect 11342 13010 11394 13022
rect 12238 13074 12290 13086
rect 12238 13010 12290 13022
rect 12686 13074 12738 13086
rect 12686 13010 12738 13022
rect 14590 13074 14642 13086
rect 14590 13010 14642 13022
rect 14926 13074 14978 13086
rect 14926 13010 14978 13022
rect 17054 13074 17106 13086
rect 17054 13010 17106 13022
rect 22094 13074 22146 13086
rect 26238 13074 26290 13086
rect 24434 13022 24446 13074
rect 24498 13022 24510 13074
rect 22094 13010 22146 13022
rect 26238 13010 26290 13022
rect 27022 13074 27074 13086
rect 27022 13010 27074 13022
rect 5518 12962 5570 12974
rect 1810 12910 1822 12962
rect 1874 12910 1886 12962
rect 5518 12898 5570 12910
rect 6974 12962 7026 12974
rect 6974 12898 7026 12910
rect 7198 12962 7250 12974
rect 7198 12898 7250 12910
rect 13470 12962 13522 12974
rect 13470 12898 13522 12910
rect 13694 12962 13746 12974
rect 13694 12898 13746 12910
rect 14142 12962 14194 12974
rect 14142 12898 14194 12910
rect 17614 12962 17666 12974
rect 17614 12898 17666 12910
rect 18958 12962 19010 12974
rect 18958 12898 19010 12910
rect 19742 12962 19794 12974
rect 19742 12898 19794 12910
rect 22766 12962 22818 12974
rect 26574 12962 26626 12974
rect 23426 12910 23438 12962
rect 23490 12910 23502 12962
rect 22766 12898 22818 12910
rect 26574 12898 26626 12910
rect 5966 12850 6018 12862
rect 5966 12786 6018 12798
rect 6190 12850 6242 12862
rect 6190 12786 6242 12798
rect 7086 12850 7138 12862
rect 7086 12786 7138 12798
rect 10110 12850 10162 12862
rect 10110 12786 10162 12798
rect 17390 12850 17442 12862
rect 17390 12786 17442 12798
rect 17950 12850 18002 12862
rect 17950 12786 18002 12798
rect 18398 12850 18450 12862
rect 18398 12786 18450 12798
rect 5742 12738 5794 12750
rect 5742 12674 5794 12686
rect 6638 12738 6690 12750
rect 6638 12674 6690 12686
rect 7422 12738 7474 12750
rect 7422 12674 7474 12686
rect 8542 12738 8594 12750
rect 8542 12674 8594 12686
rect 9326 12738 9378 12750
rect 9326 12674 9378 12686
rect 9662 12738 9714 12750
rect 9662 12674 9714 12686
rect 9774 12738 9826 12750
rect 9774 12674 9826 12686
rect 9886 12738 9938 12750
rect 9886 12674 9938 12686
rect 11790 12738 11842 12750
rect 11790 12674 11842 12686
rect 13806 12738 13858 12750
rect 13806 12674 13858 12686
rect 17502 12738 17554 12750
rect 17502 12674 17554 12686
rect 18286 12738 18338 12750
rect 18286 12674 18338 12686
rect 18510 12738 18562 12750
rect 18510 12674 18562 12686
rect 19294 12738 19346 12750
rect 19294 12674 19346 12686
rect 20190 12738 20242 12750
rect 20190 12674 20242 12686
rect 1344 12570 28720 12604
rect 1344 12518 8018 12570
rect 8070 12518 8122 12570
rect 8174 12518 8226 12570
rect 8278 12518 14822 12570
rect 14874 12518 14926 12570
rect 14978 12518 15030 12570
rect 15082 12518 21626 12570
rect 21678 12518 21730 12570
rect 21782 12518 21834 12570
rect 21886 12518 28430 12570
rect 28482 12518 28534 12570
rect 28586 12518 28638 12570
rect 28690 12518 28720 12570
rect 1344 12484 28720 12518
rect 4062 12402 4114 12414
rect 4062 12338 4114 12350
rect 8206 12402 8258 12414
rect 8206 12338 8258 12350
rect 11454 12402 11506 12414
rect 11454 12338 11506 12350
rect 12014 12402 12066 12414
rect 12014 12338 12066 12350
rect 13246 12402 13298 12414
rect 13246 12338 13298 12350
rect 16382 12402 16434 12414
rect 16382 12338 16434 12350
rect 17726 12402 17778 12414
rect 17726 12338 17778 12350
rect 18174 12402 18226 12414
rect 20974 12402 21026 12414
rect 18946 12350 18958 12402
rect 19010 12350 19022 12402
rect 18174 12338 18226 12350
rect 20974 12338 21026 12350
rect 21758 12402 21810 12414
rect 21758 12338 21810 12350
rect 22990 12402 23042 12414
rect 22990 12338 23042 12350
rect 23550 12402 23602 12414
rect 23550 12338 23602 12350
rect 24110 12402 24162 12414
rect 24110 12338 24162 12350
rect 2382 12290 2434 12302
rect 2034 12238 2046 12290
rect 2098 12238 2110 12290
rect 2382 12226 2434 12238
rect 2606 12290 2658 12302
rect 10558 12290 10610 12302
rect 3378 12238 3390 12290
rect 3442 12238 3454 12290
rect 5170 12238 5182 12290
rect 5234 12238 5246 12290
rect 2606 12226 2658 12238
rect 10558 12226 10610 12238
rect 11006 12290 11058 12302
rect 19854 12290 19906 12302
rect 18722 12238 18734 12290
rect 18786 12238 18798 12290
rect 11006 12226 11058 12238
rect 19854 12226 19906 12238
rect 22206 12290 22258 12302
rect 22206 12226 22258 12238
rect 22542 12290 22594 12302
rect 22542 12226 22594 12238
rect 1710 12178 1762 12190
rect 1710 12114 1762 12126
rect 3054 12178 3106 12190
rect 8990 12178 9042 12190
rect 4498 12126 4510 12178
rect 4562 12126 4574 12178
rect 3054 12114 3106 12126
rect 8990 12114 9042 12126
rect 9662 12178 9714 12190
rect 9662 12114 9714 12126
rect 9774 12178 9826 12190
rect 9774 12114 9826 12126
rect 10222 12178 10274 12190
rect 22094 12178 22146 12190
rect 18610 12126 18622 12178
rect 18674 12126 18686 12178
rect 19506 12126 19518 12178
rect 19570 12126 19582 12178
rect 25218 12126 25230 12178
rect 25282 12126 25294 12178
rect 10222 12114 10274 12126
rect 22094 12114 22146 12126
rect 8542 12066 8594 12078
rect 2594 12014 2606 12066
rect 2658 12014 2670 12066
rect 7298 12014 7310 12066
rect 7362 12014 7374 12066
rect 8542 12002 8594 12014
rect 9998 12066 10050 12078
rect 9998 12002 10050 12014
rect 14366 12066 14418 12078
rect 14366 12002 14418 12014
rect 15262 12066 15314 12078
rect 15262 12002 15314 12014
rect 16830 12066 16882 12078
rect 16830 12002 16882 12014
rect 20526 12066 20578 12078
rect 20526 12002 20578 12014
rect 22430 12066 22482 12078
rect 22430 12002 22482 12014
rect 24670 12066 24722 12078
rect 27122 12014 27134 12066
rect 27186 12014 27198 12066
rect 24670 12002 24722 12014
rect 20402 11902 20414 11954
rect 20466 11951 20478 11954
rect 20850 11951 20862 11954
rect 20466 11905 20862 11951
rect 20466 11902 20478 11905
rect 20850 11902 20862 11905
rect 20914 11902 20926 11954
rect 22754 11902 22766 11954
rect 22818 11951 22830 11954
rect 23426 11951 23438 11954
rect 22818 11905 23438 11951
rect 22818 11902 22830 11905
rect 23426 11902 23438 11905
rect 23490 11902 23502 11954
rect 1344 11786 28560 11820
rect 1344 11734 4616 11786
rect 4668 11734 4720 11786
rect 4772 11734 4824 11786
rect 4876 11734 11420 11786
rect 11472 11734 11524 11786
rect 11576 11734 11628 11786
rect 11680 11734 18224 11786
rect 18276 11734 18328 11786
rect 18380 11734 18432 11786
rect 18484 11734 25028 11786
rect 25080 11734 25132 11786
rect 25184 11734 25236 11786
rect 25288 11734 28560 11786
rect 1344 11700 28560 11734
rect 2606 11618 2658 11630
rect 3938 11566 3950 11618
rect 4002 11566 4014 11618
rect 2606 11554 2658 11566
rect 7198 11506 7250 11518
rect 7198 11442 7250 11454
rect 7646 11506 7698 11518
rect 7858 11454 7870 11506
rect 7922 11454 7934 11506
rect 9986 11454 9998 11506
rect 10050 11454 10062 11506
rect 15810 11454 15822 11506
rect 15874 11454 15886 11506
rect 17042 11454 17054 11506
rect 17106 11454 17118 11506
rect 19170 11454 19182 11506
rect 19234 11454 19246 11506
rect 21298 11454 21310 11506
rect 21362 11454 21374 11506
rect 23426 11454 23438 11506
rect 23490 11454 23502 11506
rect 25778 11454 25790 11506
rect 25842 11454 25854 11506
rect 7646 11442 7698 11454
rect 3054 11394 3106 11406
rect 19630 11394 19682 11406
rect 2258 11342 2270 11394
rect 2322 11342 2334 11394
rect 3378 11342 3390 11394
rect 3442 11342 3454 11394
rect 10658 11342 10670 11394
rect 10722 11342 10734 11394
rect 14466 11342 14478 11394
rect 14530 11342 14542 11394
rect 15922 11342 15934 11394
rect 15986 11342 15998 11394
rect 16370 11342 16382 11394
rect 16434 11342 16446 11394
rect 3054 11330 3106 11342
rect 19630 11330 19682 11342
rect 20078 11394 20130 11406
rect 20078 11330 20130 11342
rect 20190 11394 20242 11406
rect 20190 11330 20242 11342
rect 20750 11394 20802 11406
rect 24098 11342 24110 11394
rect 24162 11342 24174 11394
rect 24658 11342 24670 11394
rect 24722 11342 24734 11394
rect 20750 11330 20802 11342
rect 4286 11282 4338 11294
rect 2818 11230 2830 11282
rect 2882 11230 2894 11282
rect 4286 11218 4338 11230
rect 4958 11282 5010 11294
rect 4958 11218 5010 11230
rect 5070 11282 5122 11294
rect 5070 11218 5122 11230
rect 6302 11282 6354 11294
rect 6302 11218 6354 11230
rect 6526 11282 6578 11294
rect 6526 11218 6578 11230
rect 11230 11282 11282 11294
rect 11230 11218 11282 11230
rect 12910 11282 12962 11294
rect 12910 11218 12962 11230
rect 13582 11282 13634 11294
rect 13582 11218 13634 11230
rect 13918 11282 13970 11294
rect 13918 11218 13970 11230
rect 14142 11282 14194 11294
rect 14142 11218 14194 11230
rect 14702 11282 14754 11294
rect 15810 11230 15822 11282
rect 15874 11230 15886 11282
rect 14702 11218 14754 11230
rect 2046 11170 2098 11182
rect 4398 11170 4450 11182
rect 2594 11118 2606 11170
rect 2658 11118 2670 11170
rect 2046 11106 2098 11118
rect 4398 11106 4450 11118
rect 4510 11170 4562 11182
rect 4510 11106 4562 11118
rect 5966 11170 6018 11182
rect 5966 11106 6018 11118
rect 6414 11170 6466 11182
rect 6414 11106 6466 11118
rect 12014 11170 12066 11182
rect 12014 11106 12066 11118
rect 12462 11170 12514 11182
rect 12462 11106 12514 11118
rect 13806 11170 13858 11182
rect 13806 11106 13858 11118
rect 19854 11170 19906 11182
rect 19854 11106 19906 11118
rect 1344 11002 28720 11036
rect 1344 10950 8018 11002
rect 8070 10950 8122 11002
rect 8174 10950 8226 11002
rect 8278 10950 14822 11002
rect 14874 10950 14926 11002
rect 14978 10950 15030 11002
rect 15082 10950 21626 11002
rect 21678 10950 21730 11002
rect 21782 10950 21834 11002
rect 21886 10950 28430 11002
rect 28482 10950 28534 11002
rect 28586 10950 28638 11002
rect 28690 10950 28720 11002
rect 1344 10916 28720 10950
rect 9886 10834 9938 10846
rect 8642 10782 8654 10834
rect 8706 10782 8718 10834
rect 9886 10770 9938 10782
rect 11678 10834 11730 10846
rect 11678 10770 11730 10782
rect 11902 10834 11954 10846
rect 11902 10770 11954 10782
rect 12126 10834 12178 10846
rect 12126 10770 12178 10782
rect 12798 10834 12850 10846
rect 12798 10770 12850 10782
rect 13582 10834 13634 10846
rect 13582 10770 13634 10782
rect 14590 10834 14642 10846
rect 14590 10770 14642 10782
rect 14702 10834 14754 10846
rect 14702 10770 14754 10782
rect 14926 10834 14978 10846
rect 14926 10770 14978 10782
rect 16382 10834 16434 10846
rect 18622 10834 18674 10846
rect 17938 10782 17950 10834
rect 18002 10782 18014 10834
rect 16382 10770 16434 10782
rect 18622 10770 18674 10782
rect 19630 10834 19682 10846
rect 22318 10834 22370 10846
rect 20290 10782 20302 10834
rect 20354 10782 20366 10834
rect 19630 10770 19682 10782
rect 22318 10770 22370 10782
rect 22430 10834 22482 10846
rect 22430 10770 22482 10782
rect 24110 10834 24162 10846
rect 24110 10770 24162 10782
rect 7758 10722 7810 10734
rect 2258 10670 2270 10722
rect 2322 10670 2334 10722
rect 7758 10658 7810 10670
rect 14030 10722 14082 10734
rect 14030 10658 14082 10670
rect 15710 10722 15762 10734
rect 15710 10658 15762 10670
rect 15934 10722 15986 10734
rect 21646 10722 21698 10734
rect 17602 10670 17614 10722
rect 17666 10670 17678 10722
rect 20850 10670 20862 10722
rect 20914 10670 20926 10722
rect 15934 10658 15986 10670
rect 21646 10658 21698 10670
rect 22654 10722 22706 10734
rect 22654 10658 22706 10670
rect 23214 10722 23266 10734
rect 23214 10658 23266 10670
rect 23662 10722 23714 10734
rect 23662 10658 23714 10670
rect 10222 10610 10274 10622
rect 7298 10558 7310 10610
rect 7362 10558 7374 10610
rect 8082 10558 8094 10610
rect 8146 10558 8158 10610
rect 10222 10546 10274 10558
rect 10446 10610 10498 10622
rect 10446 10546 10498 10558
rect 10782 10610 10834 10622
rect 10782 10546 10834 10558
rect 11118 10610 11170 10622
rect 11118 10546 11170 10558
rect 11790 10610 11842 10622
rect 11790 10546 11842 10558
rect 13806 10610 13858 10622
rect 13806 10546 13858 10558
rect 14478 10610 14530 10622
rect 14478 10546 14530 10558
rect 15262 10610 15314 10622
rect 15262 10546 15314 10558
rect 16270 10610 16322 10622
rect 16270 10546 16322 10558
rect 16494 10610 16546 10622
rect 21198 10610 21250 10622
rect 16818 10558 16830 10610
rect 16882 10558 16894 10610
rect 17378 10558 17390 10610
rect 17442 10558 17454 10610
rect 18498 10558 18510 10610
rect 18562 10558 18574 10610
rect 19954 10558 19966 10610
rect 20018 10558 20030 10610
rect 20290 10558 20302 10610
rect 20354 10558 20366 10610
rect 16494 10546 16546 10558
rect 21198 10546 21250 10558
rect 21310 10610 21362 10622
rect 21310 10546 21362 10558
rect 21422 10610 21474 10622
rect 21422 10546 21474 10558
rect 22206 10610 22258 10622
rect 25554 10558 25566 10610
rect 25618 10558 25630 10610
rect 22206 10546 22258 10558
rect 10670 10498 10722 10510
rect 10670 10434 10722 10446
rect 13358 10498 13410 10510
rect 13358 10434 13410 10446
rect 13694 10498 13746 10510
rect 13694 10434 13746 10446
rect 15486 10498 15538 10510
rect 15486 10434 15538 10446
rect 24558 10498 24610 10510
rect 26338 10446 26350 10498
rect 26402 10446 26414 10498
rect 24558 10434 24610 10446
rect 7646 10386 7698 10398
rect 7646 10322 7698 10334
rect 1344 10218 28560 10252
rect 1344 10166 4616 10218
rect 4668 10166 4720 10218
rect 4772 10166 4824 10218
rect 4876 10166 11420 10218
rect 11472 10166 11524 10218
rect 11576 10166 11628 10218
rect 11680 10166 18224 10218
rect 18276 10166 18328 10218
rect 18380 10166 18432 10218
rect 18484 10166 25028 10218
rect 25080 10166 25132 10218
rect 25184 10166 25236 10218
rect 25288 10166 28560 10218
rect 1344 10132 28560 10166
rect 2482 9886 2494 9938
rect 2546 9886 2558 9938
rect 4610 9886 4622 9938
rect 4674 9886 4686 9938
rect 8754 9886 8766 9938
rect 8818 9886 8830 9938
rect 10434 9886 10446 9938
rect 10498 9886 10510 9938
rect 12562 9886 12574 9938
rect 12626 9886 12638 9938
rect 14242 9886 14254 9938
rect 14306 9886 14318 9938
rect 16370 9886 16382 9938
rect 16434 9886 16446 9938
rect 18610 9886 18622 9938
rect 18674 9886 18686 9938
rect 20738 9912 20750 9964
rect 20802 9912 20814 9964
rect 21534 9938 21586 9950
rect 21534 9874 21586 9886
rect 21982 9938 22034 9950
rect 22978 9886 22990 9938
rect 23042 9886 23054 9938
rect 21982 9874 22034 9886
rect 16718 9826 16770 9838
rect 1810 9774 1822 9826
rect 1874 9774 1886 9826
rect 5954 9774 5966 9826
rect 6018 9774 6030 9826
rect 9762 9774 9774 9826
rect 9826 9774 9838 9826
rect 13458 9774 13470 9826
rect 13522 9774 13534 9826
rect 16718 9762 16770 9774
rect 17054 9826 17106 9838
rect 25566 9826 25618 9838
rect 17826 9774 17838 9826
rect 17890 9774 17902 9826
rect 24882 9774 24894 9826
rect 24946 9774 24958 9826
rect 17054 9762 17106 9774
rect 25566 9762 25618 9774
rect 26014 9826 26066 9838
rect 26014 9762 26066 9774
rect 17390 9714 17442 9726
rect 6626 9662 6638 9714
rect 6690 9662 6702 9714
rect 17390 9650 17442 9662
rect 5070 9602 5122 9614
rect 5070 9538 5122 9550
rect 9214 9602 9266 9614
rect 9214 9538 9266 9550
rect 17054 9602 17106 9614
rect 17054 9538 17106 9550
rect 1344 9434 28720 9468
rect 1344 9382 8018 9434
rect 8070 9382 8122 9434
rect 8174 9382 8226 9434
rect 8278 9382 14822 9434
rect 14874 9382 14926 9434
rect 14978 9382 15030 9434
rect 15082 9382 21626 9434
rect 21678 9382 21730 9434
rect 21782 9382 21834 9434
rect 21886 9382 28430 9434
rect 28482 9382 28534 9434
rect 28586 9382 28638 9434
rect 28690 9382 28720 9434
rect 1344 9348 28720 9382
rect 7534 9266 7586 9278
rect 6514 9214 6526 9266
rect 6578 9214 6590 9266
rect 7534 9202 7586 9214
rect 7870 9266 7922 9278
rect 7870 9202 7922 9214
rect 8878 9266 8930 9278
rect 8878 9202 8930 9214
rect 12462 9266 12514 9278
rect 12462 9202 12514 9214
rect 12798 9266 12850 9278
rect 12798 9202 12850 9214
rect 15038 9266 15090 9278
rect 15038 9202 15090 9214
rect 17614 9266 17666 9278
rect 17614 9202 17666 9214
rect 18062 9266 18114 9278
rect 18062 9202 18114 9214
rect 18174 9266 18226 9278
rect 18174 9202 18226 9214
rect 19070 9266 19122 9278
rect 19070 9202 19122 9214
rect 19518 9266 19570 9278
rect 19518 9202 19570 9214
rect 19966 9266 20018 9278
rect 19966 9202 20018 9214
rect 24222 9266 24274 9278
rect 24222 9202 24274 9214
rect 13134 9154 13186 9166
rect 2370 9102 2382 9154
rect 2434 9102 2446 9154
rect 3154 9102 3166 9154
rect 3218 9102 3230 9154
rect 4498 9102 4510 9154
rect 4562 9102 4574 9154
rect 6290 9102 6302 9154
rect 6354 9102 6366 9154
rect 13134 9090 13186 9102
rect 13694 9154 13746 9166
rect 13694 9090 13746 9102
rect 14142 9154 14194 9166
rect 14142 9090 14194 9102
rect 16830 9154 16882 9166
rect 16830 9090 16882 9102
rect 17950 9154 18002 9166
rect 17950 9090 18002 9102
rect 6078 9042 6130 9054
rect 4386 8990 4398 9042
rect 4450 8990 4462 9042
rect 6078 8978 6130 8990
rect 6526 9042 6578 9054
rect 13358 9042 13410 9054
rect 6626 8990 6638 9042
rect 6690 8990 6702 9042
rect 7746 8990 7758 9042
rect 7810 8990 7822 9042
rect 6526 8978 6578 8990
rect 13358 8978 13410 8990
rect 15486 9042 15538 9054
rect 15486 8978 15538 8990
rect 18622 9042 18674 9054
rect 18622 8978 18674 8990
rect 23438 9042 23490 9054
rect 23438 8978 23490 8990
rect 2158 8930 2210 8942
rect 2158 8866 2210 8878
rect 5518 8930 5570 8942
rect 5518 8866 5570 8878
rect 13246 8930 13298 8942
rect 13246 8866 13298 8878
rect 14702 8930 14754 8942
rect 14702 8866 14754 8878
rect 16158 8930 16210 8942
rect 16158 8866 16210 8878
rect 20974 8930 21026 8942
rect 20974 8866 21026 8878
rect 1344 8650 28560 8684
rect 1344 8598 4616 8650
rect 4668 8598 4720 8650
rect 4772 8598 4824 8650
rect 4876 8598 11420 8650
rect 11472 8598 11524 8650
rect 11576 8598 11628 8650
rect 11680 8598 18224 8650
rect 18276 8598 18328 8650
rect 18380 8598 18432 8650
rect 18484 8598 25028 8650
rect 25080 8598 25132 8650
rect 25184 8598 25236 8650
rect 25288 8598 28560 8650
rect 1344 8564 28560 8598
rect 6850 8430 6862 8482
rect 6914 8430 6926 8482
rect 16930 8430 16942 8482
rect 16994 8479 17006 8482
rect 17154 8479 17166 8482
rect 16994 8433 17166 8479
rect 16994 8430 17006 8433
rect 17154 8430 17166 8433
rect 17218 8430 17230 8482
rect 1822 8370 1874 8382
rect 7534 8370 7586 8382
rect 16942 8370 16994 8382
rect 5058 8318 5070 8370
rect 5122 8318 5134 8370
rect 14242 8318 14254 8370
rect 14306 8318 14318 8370
rect 16370 8318 16382 8370
rect 16434 8318 16446 8370
rect 1822 8306 1874 8318
rect 7534 8306 7586 8318
rect 16942 8306 16994 8318
rect 17390 8370 17442 8382
rect 17390 8306 17442 8318
rect 17838 8370 17890 8382
rect 17838 8306 17890 8318
rect 18174 8370 18226 8382
rect 18174 8306 18226 8318
rect 18846 8370 18898 8382
rect 18846 8306 18898 8318
rect 21422 8370 21474 8382
rect 22642 8318 22654 8370
rect 22706 8318 22718 8370
rect 21422 8306 21474 8318
rect 6638 8258 6690 8270
rect 19294 8258 19346 8270
rect 20638 8258 20690 8270
rect 2258 8206 2270 8258
rect 2322 8206 2334 8258
rect 6850 8206 6862 8258
rect 6914 8206 6926 8258
rect 13570 8206 13582 8258
rect 13634 8206 13646 8258
rect 20066 8206 20078 8258
rect 20130 8206 20142 8258
rect 6638 8194 6690 8206
rect 19294 8194 19346 8206
rect 20638 8194 20690 8206
rect 22094 8258 22146 8270
rect 22094 8194 22146 8206
rect 22318 8258 22370 8270
rect 24782 8258 24834 8270
rect 24546 8206 24558 8258
rect 24610 8206 24622 8258
rect 22318 8194 22370 8206
rect 24782 8194 24834 8206
rect 6302 8146 6354 8158
rect 2930 8094 2942 8146
rect 2994 8094 3006 8146
rect 6302 8082 6354 8094
rect 7422 8146 7474 8158
rect 7422 8082 7474 8094
rect 8094 8146 8146 8158
rect 8094 8082 8146 8094
rect 8206 8146 8258 8158
rect 20302 8146 20354 8158
rect 19730 8094 19742 8146
rect 19794 8094 19806 8146
rect 8206 8082 8258 8094
rect 20302 8082 20354 8094
rect 20750 8146 20802 8158
rect 20750 8082 20802 8094
rect 23998 8146 24050 8158
rect 23998 8082 24050 8094
rect 6078 8034 6130 8046
rect 7646 8034 7698 8046
rect 6738 7982 6750 8034
rect 6802 7982 6814 8034
rect 6078 7970 6130 7982
rect 7646 7970 7698 7982
rect 8654 8034 8706 8046
rect 8654 7970 8706 7982
rect 24446 8034 24498 8046
rect 24446 7970 24498 7982
rect 1344 7866 28720 7900
rect 1344 7814 8018 7866
rect 8070 7814 8122 7866
rect 8174 7814 8226 7866
rect 8278 7814 14822 7866
rect 14874 7814 14926 7866
rect 14978 7814 15030 7866
rect 15082 7814 21626 7866
rect 21678 7814 21730 7866
rect 21782 7814 21834 7866
rect 21886 7814 28430 7866
rect 28482 7814 28534 7866
rect 28586 7814 28638 7866
rect 28690 7814 28720 7866
rect 1344 7780 28720 7814
rect 2830 7698 2882 7710
rect 2034 7646 2046 7698
rect 2098 7646 2110 7698
rect 2830 7634 2882 7646
rect 3726 7698 3778 7710
rect 9662 7698 9714 7710
rect 5058 7646 5070 7698
rect 5122 7646 5134 7698
rect 3726 7634 3778 7646
rect 9662 7634 9714 7646
rect 13582 7698 13634 7710
rect 20626 7646 20638 7698
rect 20690 7646 20702 7698
rect 22754 7646 22766 7698
rect 22818 7646 22830 7698
rect 23202 7646 23214 7698
rect 23266 7646 23278 7698
rect 13582 7634 13634 7646
rect 5518 7586 5570 7598
rect 6850 7534 6862 7586
rect 6914 7534 6926 7586
rect 14690 7534 14702 7586
rect 14754 7534 14766 7586
rect 19842 7534 19854 7586
rect 19906 7534 19918 7586
rect 5518 7522 5570 7534
rect 1710 7474 1762 7486
rect 5182 7474 5234 7486
rect 21198 7474 21250 7486
rect 23662 7474 23714 7486
rect 3266 7422 3278 7474
rect 3330 7422 3342 7474
rect 4722 7422 4734 7474
rect 4786 7422 4798 7474
rect 6178 7422 6190 7474
rect 6242 7422 6254 7474
rect 13906 7422 13918 7474
rect 13970 7422 13982 7474
rect 20514 7422 20526 7474
rect 20578 7422 20590 7474
rect 22418 7422 22430 7474
rect 22482 7422 22494 7474
rect 1710 7410 1762 7422
rect 5182 7410 5234 7422
rect 21198 7410 21250 7422
rect 23662 7410 23714 7422
rect 23774 7474 23826 7486
rect 23774 7410 23826 7422
rect 23886 7474 23938 7486
rect 23886 7410 23938 7422
rect 19070 7362 19122 7374
rect 8978 7310 8990 7362
rect 9042 7310 9054 7362
rect 16818 7310 16830 7362
rect 16882 7310 16894 7362
rect 19070 7298 19122 7310
rect 4946 7198 4958 7250
rect 5010 7198 5022 7250
rect 1344 7082 28560 7116
rect 1344 7030 4616 7082
rect 4668 7030 4720 7082
rect 4772 7030 4824 7082
rect 4876 7030 11420 7082
rect 11472 7030 11524 7082
rect 11576 7030 11628 7082
rect 11680 7030 18224 7082
rect 18276 7030 18328 7082
rect 18380 7030 18432 7082
rect 18484 7030 25028 7082
rect 25080 7030 25132 7082
rect 25184 7030 25236 7082
rect 25288 7030 28560 7082
rect 1344 6996 28560 7030
rect 22430 6914 22482 6926
rect 5842 6862 5854 6914
rect 5906 6911 5918 6914
rect 6290 6911 6302 6914
rect 5906 6865 6302 6911
rect 5906 6862 5918 6865
rect 6290 6862 6302 6865
rect 6354 6911 6366 6914
rect 6626 6911 6638 6914
rect 6354 6865 6638 6911
rect 6354 6862 6366 6865
rect 6626 6862 6638 6865
rect 6690 6862 6702 6914
rect 22430 6850 22482 6862
rect 2494 6802 2546 6814
rect 2494 6738 2546 6750
rect 3390 6802 3442 6814
rect 3390 6738 3442 6750
rect 5854 6802 5906 6814
rect 5854 6738 5906 6750
rect 6638 6802 6690 6814
rect 24670 6802 24722 6814
rect 18946 6750 18958 6802
rect 19010 6750 19022 6802
rect 19506 6750 19518 6802
rect 19570 6750 19582 6802
rect 6638 6738 6690 6750
rect 24670 6738 24722 6750
rect 4734 6690 4786 6702
rect 4734 6626 4786 6638
rect 4846 6690 4898 6702
rect 4846 6626 4898 6638
rect 6190 6690 6242 6702
rect 21646 6690 21698 6702
rect 16146 6638 16158 6690
rect 16210 6638 16222 6690
rect 16818 6638 16830 6690
rect 16882 6638 16894 6690
rect 20066 6638 20078 6690
rect 20130 6638 20142 6690
rect 6190 6626 6242 6638
rect 21646 6626 21698 6638
rect 22094 6690 22146 6702
rect 24434 6638 24446 6690
rect 24498 6638 24510 6690
rect 22094 6626 22146 6638
rect 4398 6578 4450 6590
rect 21310 6578 21362 6590
rect 20514 6526 20526 6578
rect 20578 6526 20590 6578
rect 4398 6514 4450 6526
rect 21310 6514 21362 6526
rect 22542 6578 22594 6590
rect 22542 6514 22594 6526
rect 23886 6578 23938 6590
rect 23886 6514 23938 6526
rect 3838 6466 3890 6478
rect 24882 6414 24894 6466
rect 24946 6414 24958 6466
rect 3838 6402 3890 6414
rect 1344 6298 28720 6332
rect 1344 6246 8018 6298
rect 8070 6246 8122 6298
rect 8174 6246 8226 6298
rect 8278 6246 14822 6298
rect 14874 6246 14926 6298
rect 14978 6246 15030 6298
rect 15082 6246 21626 6298
rect 21678 6246 21730 6298
rect 21782 6246 21834 6298
rect 21886 6246 28430 6298
rect 28482 6246 28534 6298
rect 28586 6246 28638 6298
rect 28690 6246 28720 6298
rect 1344 6212 28720 6246
rect 5182 6130 5234 6142
rect 5182 6066 5234 6078
rect 5854 6130 5906 6142
rect 25454 6130 25506 6142
rect 18722 6078 18734 6130
rect 18786 6078 18798 6130
rect 21410 6078 21422 6130
rect 21474 6078 21486 6130
rect 5854 6066 5906 6078
rect 25454 6066 25506 6078
rect 26014 6018 26066 6030
rect 20066 5966 20078 6018
rect 20130 5966 20142 6018
rect 21858 5966 21870 6018
rect 21922 5966 21934 6018
rect 22530 5966 22542 6018
rect 22594 5966 22606 6018
rect 24210 5966 24222 6018
rect 24274 5966 24286 6018
rect 26014 5954 26066 5966
rect 22990 5906 23042 5918
rect 19842 5854 19854 5906
rect 19906 5854 19918 5906
rect 21746 5854 21758 5906
rect 21810 5854 21822 5906
rect 22990 5842 23042 5854
rect 23102 5906 23154 5918
rect 23102 5842 23154 5854
rect 23438 5906 23490 5918
rect 23438 5842 23490 5854
rect 23662 5906 23714 5918
rect 25902 5906 25954 5918
rect 23874 5854 23886 5906
rect 23938 5854 23950 5906
rect 23662 5842 23714 5854
rect 25902 5842 25954 5854
rect 25566 5794 25618 5806
rect 24098 5742 24110 5794
rect 24162 5742 24174 5794
rect 25566 5730 25618 5742
rect 1344 5514 28560 5548
rect 1344 5462 4616 5514
rect 4668 5462 4720 5514
rect 4772 5462 4824 5514
rect 4876 5462 11420 5514
rect 11472 5462 11524 5514
rect 11576 5462 11628 5514
rect 11680 5462 18224 5514
rect 18276 5462 18328 5514
rect 18380 5462 18432 5514
rect 18484 5462 25028 5514
rect 25080 5462 25132 5514
rect 25184 5462 25236 5514
rect 25288 5462 28560 5514
rect 1344 5428 28560 5462
rect 22530 5182 22542 5234
rect 22594 5182 22606 5234
rect 1710 5122 1762 5134
rect 1710 5058 1762 5070
rect 2494 5122 2546 5134
rect 2494 5058 2546 5070
rect 18734 5122 18786 5134
rect 18734 5058 18786 5070
rect 20638 5122 20690 5134
rect 25454 5122 25506 5134
rect 21522 5070 21534 5122
rect 21586 5070 21598 5122
rect 22978 5070 22990 5122
rect 23042 5070 23054 5122
rect 20638 5058 20690 5070
rect 25454 5058 25506 5070
rect 26910 5122 26962 5134
rect 26910 5058 26962 5070
rect 27358 5122 27410 5134
rect 27358 5058 27410 5070
rect 27806 5122 27858 5134
rect 27806 5058 27858 5070
rect 19742 5010 19794 5022
rect 2034 4958 2046 5010
rect 2098 4958 2110 5010
rect 19742 4946 19794 4958
rect 20414 5010 20466 5022
rect 23202 4958 23214 5010
rect 23266 4958 23278 5010
rect 23874 4958 23886 5010
rect 23938 4958 23950 5010
rect 20414 4946 20466 4958
rect 19070 4898 19122 4910
rect 19070 4834 19122 4846
rect 19854 4898 19906 4910
rect 19854 4834 19906 4846
rect 20078 4898 20130 4910
rect 20078 4834 20130 4846
rect 20526 4898 20578 4910
rect 20526 4834 20578 4846
rect 21310 4898 21362 4910
rect 21310 4834 21362 4846
rect 26014 4898 26066 4910
rect 26014 4834 26066 4846
rect 26462 4898 26514 4910
rect 26462 4834 26514 4846
rect 1344 4730 28720 4764
rect 1344 4678 8018 4730
rect 8070 4678 8122 4730
rect 8174 4678 8226 4730
rect 8278 4678 14822 4730
rect 14874 4678 14926 4730
rect 14978 4678 15030 4730
rect 15082 4678 21626 4730
rect 21678 4678 21730 4730
rect 21782 4678 21834 4730
rect 21886 4678 28430 4730
rect 28482 4678 28534 4730
rect 28586 4678 28638 4730
rect 28690 4678 28720 4730
rect 1344 4644 28720 4678
rect 19630 4562 19682 4574
rect 19630 4498 19682 4510
rect 22430 4562 22482 4574
rect 22430 4498 22482 4510
rect 11790 4450 11842 4462
rect 11790 4386 11842 4398
rect 18510 4450 18562 4462
rect 18510 4386 18562 4398
rect 18846 4450 18898 4462
rect 18846 4386 18898 4398
rect 19182 4450 19234 4462
rect 19182 4386 19234 4398
rect 20638 4450 20690 4462
rect 20638 4386 20690 4398
rect 22990 4450 23042 4462
rect 22990 4386 23042 4398
rect 25230 4450 25282 4462
rect 25230 4386 25282 4398
rect 11230 4338 11282 4350
rect 21534 4338 21586 4350
rect 24222 4338 24274 4350
rect 11554 4286 11566 4338
rect 11618 4286 11630 4338
rect 19394 4286 19406 4338
rect 19458 4286 19470 4338
rect 23426 4286 23438 4338
rect 23490 4286 23502 4338
rect 25330 4286 25342 4338
rect 25394 4286 25406 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 11230 4274 11282 4286
rect 21534 4274 21586 4286
rect 24222 4274 24274 4286
rect 10782 4226 10834 4238
rect 12238 4226 12290 4238
rect 11666 4174 11678 4226
rect 11730 4174 11742 4226
rect 10782 4162 10834 4174
rect 12238 4162 12290 4174
rect 17838 4226 17890 4238
rect 17838 4162 17890 4174
rect 18286 4226 18338 4238
rect 18286 4162 18338 4174
rect 21870 4226 21922 4238
rect 21870 4162 21922 4174
rect 23214 4226 23266 4238
rect 23214 4162 23266 4174
rect 24110 4226 24162 4238
rect 24110 4162 24162 4174
rect 24670 4226 24722 4238
rect 24670 4162 24722 4174
rect 26462 4226 26514 4238
rect 26462 4162 26514 4174
rect 26910 4226 26962 4238
rect 26910 4162 26962 4174
rect 27358 4226 27410 4238
rect 27358 4162 27410 4174
rect 27806 4226 27858 4238
rect 27806 4162 27858 4174
rect 19742 4114 19794 4126
rect 19742 4050 19794 4062
rect 24558 4114 24610 4126
rect 27010 4062 27022 4114
rect 27074 4111 27086 4114
rect 27794 4111 27806 4114
rect 27074 4065 27806 4111
rect 27074 4062 27086 4065
rect 27794 4062 27806 4065
rect 27858 4062 27870 4114
rect 24558 4050 24610 4062
rect 1344 3946 28560 3980
rect 1344 3894 4616 3946
rect 4668 3894 4720 3946
rect 4772 3894 4824 3946
rect 4876 3894 11420 3946
rect 11472 3894 11524 3946
rect 11576 3894 11628 3946
rect 11680 3894 18224 3946
rect 18276 3894 18328 3946
rect 18380 3894 18432 3946
rect 18484 3894 25028 3946
rect 25080 3894 25132 3946
rect 25184 3894 25236 3946
rect 25288 3894 28560 3946
rect 1344 3860 28560 3894
rect 20066 3726 20078 3778
rect 20130 3726 20142 3778
rect 22194 3726 22206 3778
rect 22258 3726 22270 3778
rect 13022 3666 13074 3678
rect 10994 3614 11006 3666
rect 11058 3614 11070 3666
rect 13022 3602 13074 3614
rect 21422 3666 21474 3678
rect 27918 3666 27970 3678
rect 21970 3614 21982 3666
rect 22034 3614 22046 3666
rect 21422 3602 21474 3614
rect 27918 3602 27970 3614
rect 17278 3554 17330 3566
rect 7634 3502 7646 3554
rect 7698 3502 7710 3554
rect 9650 3502 9662 3554
rect 9714 3502 9726 3554
rect 11778 3502 11790 3554
rect 11842 3502 11854 3554
rect 15138 3502 15150 3554
rect 15202 3502 15214 3554
rect 17278 3490 17330 3502
rect 19294 3554 19346 3566
rect 20302 3554 20354 3566
rect 23662 3554 23714 3566
rect 20066 3502 20078 3554
rect 20130 3502 20142 3554
rect 22306 3502 22318 3554
rect 22370 3502 22382 3554
rect 22642 3502 22654 3554
rect 22706 3502 22718 3554
rect 24098 3502 24110 3554
rect 24162 3502 24174 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 26114 3502 26126 3554
rect 26178 3502 26190 3554
rect 19294 3490 19346 3502
rect 20302 3490 20354 3502
rect 23662 3490 23714 3502
rect 5182 3442 5234 3454
rect 5182 3378 5234 3390
rect 5630 3442 5682 3454
rect 5630 3378 5682 3390
rect 5742 3442 5794 3454
rect 10222 3442 10274 3454
rect 16270 3442 16322 3454
rect 7746 3390 7758 3442
rect 7810 3390 7822 3442
rect 12114 3390 12126 3442
rect 12178 3390 12190 3442
rect 12338 3390 12350 3442
rect 12402 3390 12414 3442
rect 5742 3378 5794 3390
rect 10222 3378 10274 3390
rect 16270 3378 16322 3390
rect 17726 3442 17778 3454
rect 17726 3378 17778 3390
rect 19630 3442 19682 3454
rect 19630 3378 19682 3390
rect 23326 3442 23378 3454
rect 27470 3442 27522 3454
rect 25666 3390 25678 3442
rect 25730 3390 25742 3442
rect 27122 3390 27134 3442
rect 27186 3390 27198 3442
rect 23326 3378 23378 3390
rect 27470 3378 27522 3390
rect 4622 3330 4674 3342
rect 4622 3266 4674 3278
rect 5966 3330 6018 3342
rect 5966 3266 6018 3278
rect 6302 3330 6354 3342
rect 6302 3266 6354 3278
rect 6862 3330 6914 3342
rect 6862 3266 6914 3278
rect 7422 3330 7474 3342
rect 7422 3266 7474 3278
rect 13582 3330 13634 3342
rect 21310 3330 21362 3342
rect 18834 3278 18846 3330
rect 18898 3278 18910 3330
rect 13582 3266 13634 3278
rect 21310 3266 21362 3278
rect 1344 3162 28720 3196
rect 1344 3110 8018 3162
rect 8070 3110 8122 3162
rect 8174 3110 8226 3162
rect 8278 3110 14822 3162
rect 14874 3110 14926 3162
rect 14978 3110 15030 3162
rect 15082 3110 21626 3162
rect 21678 3110 21730 3162
rect 21782 3110 21834 3162
rect 21886 3110 28430 3162
rect 28482 3110 28534 3162
rect 28586 3110 28638 3162
rect 28690 3110 28720 3162
rect 1344 3076 28720 3110
rect 9102 2994 9154 3006
rect 12574 2994 12626 3006
rect 6178 2942 6190 2994
rect 6242 2942 6254 2994
rect 12002 2942 12014 2994
rect 12066 2942 12078 2994
rect 9102 2930 9154 2942
rect 12574 2930 12626 2942
rect 17502 2994 17554 3006
rect 24322 2942 24334 2994
rect 24386 2942 24398 2994
rect 25330 2942 25342 2994
rect 25394 2942 25406 2994
rect 17502 2930 17554 2942
rect 9998 2882 10050 2894
rect 26686 2882 26738 2894
rect 17938 2830 17950 2882
rect 18002 2830 18014 2882
rect 19506 2830 19518 2882
rect 19570 2830 19582 2882
rect 20738 2830 20750 2882
rect 20802 2830 20814 2882
rect 21634 2830 21646 2882
rect 21698 2830 21710 2882
rect 25442 2830 25454 2882
rect 25506 2830 25518 2882
rect 26114 2830 26126 2882
rect 26178 2830 26190 2882
rect 9998 2818 10050 2830
rect 26686 2818 26738 2830
rect 27358 2882 27410 2894
rect 27358 2818 27410 2830
rect 6190 2770 6242 2782
rect 9662 2770 9714 2782
rect 2930 2718 2942 2770
rect 2994 2718 3006 2770
rect 6290 2718 6302 2770
rect 6354 2718 6366 2770
rect 6190 2706 6242 2718
rect 9662 2706 9714 2718
rect 10558 2770 10610 2782
rect 10558 2706 10610 2718
rect 11678 2770 11730 2782
rect 11678 2706 11730 2718
rect 12686 2770 12738 2782
rect 12686 2706 12738 2718
rect 17390 2770 17442 2782
rect 17390 2706 17442 2718
rect 18398 2770 18450 2782
rect 22990 2770 23042 2782
rect 25342 2770 25394 2782
rect 18946 2718 18958 2770
rect 19010 2718 19022 2770
rect 21186 2718 21198 2770
rect 21250 2718 21262 2770
rect 24098 2718 24110 2770
rect 24162 2718 24174 2770
rect 24322 2718 24334 2770
rect 24386 2718 24398 2770
rect 18398 2706 18450 2718
rect 22990 2706 23042 2718
rect 25342 2706 25394 2718
rect 27022 2770 27074 2782
rect 27570 2718 27582 2770
rect 27634 2718 27646 2770
rect 27022 2706 27074 2718
rect 7758 2658 7810 2670
rect 4050 2606 4062 2658
rect 4114 2606 4126 2658
rect 5954 2606 5966 2658
rect 6018 2606 6030 2658
rect 7758 2594 7810 2606
rect 8206 2658 8258 2670
rect 8206 2594 8258 2606
rect 8654 2658 8706 2670
rect 8654 2594 8706 2606
rect 11118 2658 11170 2670
rect 11118 2594 11170 2606
rect 11454 2658 11506 2670
rect 11454 2594 11506 2606
rect 13694 2658 13746 2670
rect 13694 2594 13746 2606
rect 14142 2658 14194 2670
rect 14142 2594 14194 2606
rect 14814 2658 14866 2670
rect 14814 2594 14866 2606
rect 15486 2658 15538 2670
rect 15486 2594 15538 2606
rect 16270 2658 16322 2670
rect 16270 2594 16322 2606
rect 16718 2658 16770 2670
rect 28142 2658 28194 2670
rect 18610 2606 18622 2658
rect 18674 2606 18686 2658
rect 20850 2606 20862 2658
rect 20914 2606 20926 2658
rect 23762 2606 23774 2658
rect 23826 2606 23838 2658
rect 16718 2594 16770 2606
rect 28142 2594 28194 2606
rect 10446 2546 10498 2558
rect 10446 2482 10498 2494
rect 10782 2546 10834 2558
rect 10782 2482 10834 2494
rect 11006 2546 11058 2558
rect 11006 2482 11058 2494
rect 12574 2546 12626 2558
rect 12574 2482 12626 2494
rect 12910 2546 12962 2558
rect 12910 2482 12962 2494
rect 13134 2546 13186 2558
rect 13134 2482 13186 2494
rect 1344 2378 28560 2412
rect 1344 2326 4616 2378
rect 4668 2326 4720 2378
rect 4772 2326 4824 2378
rect 4876 2326 11420 2378
rect 11472 2326 11524 2378
rect 11576 2326 11628 2378
rect 11680 2326 18224 2378
rect 18276 2326 18328 2378
rect 18380 2326 18432 2378
rect 18484 2326 25028 2378
rect 25080 2326 25132 2378
rect 25184 2326 25236 2378
rect 25288 2326 28560 2378
rect 1344 2292 28560 2326
rect 20750 2098 20802 2110
rect 18946 2046 18958 2098
rect 19010 2046 19022 2098
rect 20750 2034 20802 2046
rect 20974 2098 21026 2110
rect 20974 2034 21026 2046
rect 21870 2098 21922 2110
rect 25454 2098 25506 2110
rect 22866 2046 22878 2098
rect 22930 2046 22942 2098
rect 24658 2046 24670 2098
rect 24722 2046 24734 2098
rect 21870 2034 21922 2046
rect 25454 2034 25506 2046
rect 26462 2098 26514 2110
rect 26462 2034 26514 2046
rect 1934 1986 1986 1998
rect 6078 1986 6130 1998
rect 11230 1986 11282 1998
rect 13470 1986 13522 1998
rect 14702 1986 14754 1998
rect 2706 1934 2718 1986
rect 2770 1934 2782 1986
rect 4050 1934 4062 1986
rect 4114 1934 4126 1986
rect 4722 1934 4734 1986
rect 4786 1934 4798 1986
rect 6514 1934 6526 1986
rect 6578 1934 6590 1986
rect 7186 1934 7198 1986
rect 7250 1934 7262 1986
rect 7858 1934 7870 1986
rect 7922 1934 7934 1986
rect 8530 1934 8542 1986
rect 8594 1934 8606 1986
rect 9650 1934 9662 1986
rect 9714 1934 9726 1986
rect 10322 1934 10334 1986
rect 10386 1934 10398 1986
rect 11666 1934 11678 1986
rect 11730 1934 11742 1986
rect 12338 1934 12350 1986
rect 12402 1934 12414 1986
rect 13906 1934 13918 1986
rect 13970 1934 13982 1986
rect 1934 1922 1986 1934
rect 6078 1922 6130 1934
rect 11230 1922 11282 1934
rect 13470 1922 13522 1934
rect 14702 1922 14754 1934
rect 17614 1986 17666 1998
rect 19854 1986 19906 1998
rect 18610 1934 18622 1986
rect 18674 1934 18686 1986
rect 17614 1922 17666 1934
rect 19854 1922 19906 1934
rect 20190 1986 20242 1998
rect 20190 1922 20242 1934
rect 21086 1986 21138 1998
rect 21086 1922 21138 1934
rect 22430 1986 22482 1998
rect 23998 1986 24050 1998
rect 23202 1934 23214 1986
rect 23266 1934 23278 1986
rect 24994 1934 25006 1986
rect 25058 1934 25070 1986
rect 25890 1934 25902 1986
rect 25954 1934 25966 1986
rect 26898 1934 26910 1986
rect 26962 1934 26974 1986
rect 27570 1934 27582 1986
rect 27634 1934 27646 1986
rect 22430 1922 22482 1934
rect 23998 1922 24050 1934
rect 2942 1874 2994 1886
rect 2942 1810 2994 1822
rect 3278 1874 3330 1886
rect 3278 1810 3330 1822
rect 3614 1874 3666 1886
rect 3614 1810 3666 1822
rect 4286 1874 4338 1886
rect 4286 1810 4338 1822
rect 4958 1874 5010 1886
rect 4958 1810 5010 1822
rect 5742 1874 5794 1886
rect 5742 1810 5794 1822
rect 6750 1874 6802 1886
rect 6750 1810 6802 1822
rect 7422 1874 7474 1886
rect 7422 1810 7474 1822
rect 8094 1874 8146 1886
rect 8094 1810 8146 1822
rect 8766 1874 8818 1886
rect 8766 1810 8818 1822
rect 9886 1874 9938 1886
rect 9886 1810 9938 1822
rect 10558 1874 10610 1886
rect 10558 1810 10610 1822
rect 11902 1874 11954 1886
rect 11902 1810 11954 1822
rect 12574 1874 12626 1886
rect 12574 1810 12626 1822
rect 13694 1874 13746 1886
rect 13694 1810 13746 1822
rect 14366 1874 14418 1886
rect 14366 1810 14418 1822
rect 15038 1874 15090 1886
rect 15038 1810 15090 1822
rect 15374 1874 15426 1886
rect 15374 1810 15426 1822
rect 15710 1874 15762 1886
rect 15710 1810 15762 1822
rect 16046 1874 16098 1886
rect 16046 1810 16098 1822
rect 16942 1874 16994 1886
rect 16942 1810 16994 1822
rect 17278 1874 17330 1886
rect 17278 1810 17330 1822
rect 17950 1874 18002 1886
rect 19294 1874 19346 1886
rect 18498 1822 18510 1874
rect 18562 1822 18574 1874
rect 17950 1810 18002 1822
rect 19294 1810 19346 1822
rect 19630 1874 19682 1886
rect 19630 1810 19682 1822
rect 20078 1874 20130 1886
rect 20078 1810 20130 1822
rect 23662 1874 23714 1886
rect 23662 1810 23714 1822
rect 27358 1874 27410 1886
rect 27358 1810 27410 1822
rect 2382 1762 2434 1774
rect 2382 1698 2434 1710
rect 10894 1762 10946 1774
rect 10894 1698 10946 1710
rect 1344 1594 28720 1628
rect 1344 1542 8018 1594
rect 8070 1542 8122 1594
rect 8174 1542 8226 1594
rect 8278 1542 14822 1594
rect 14874 1542 14926 1594
rect 14978 1542 15030 1594
rect 15082 1542 21626 1594
rect 21678 1542 21730 1594
rect 21782 1542 21834 1594
rect 21886 1542 28430 1594
rect 28482 1542 28534 1594
rect 28586 1542 28638 1594
rect 28690 1542 28720 1594
rect 1344 1508 28720 1542
<< via1 >>
rect 8542 118750 8594 118802
rect 9326 118750 9378 118802
rect 4616 118358 4668 118410
rect 4720 118358 4772 118410
rect 4824 118358 4876 118410
rect 11420 118358 11472 118410
rect 11524 118358 11576 118410
rect 11628 118358 11680 118410
rect 18224 118358 18276 118410
rect 18328 118358 18380 118410
rect 18432 118358 18484 118410
rect 25028 118358 25080 118410
rect 25132 118358 25184 118410
rect 25236 118358 25288 118410
rect 13806 117966 13858 118018
rect 14702 117966 14754 118018
rect 19406 117966 19458 118018
rect 20078 117966 20130 118018
rect 1710 117854 1762 117906
rect 3390 117854 3442 117906
rect 5518 117854 5570 117906
rect 6974 117854 7026 117906
rect 9326 117854 9378 117906
rect 10558 117854 10610 117906
rect 12350 117854 12402 117906
rect 13358 117854 13410 117906
rect 16046 117742 16098 117794
rect 16382 117742 16434 117794
rect 17838 117742 17890 117794
rect 20862 117742 20914 117794
rect 8018 117574 8070 117626
rect 8122 117574 8174 117626
rect 8226 117574 8278 117626
rect 14822 117574 14874 117626
rect 14926 117574 14978 117626
rect 15030 117574 15082 117626
rect 21626 117574 21678 117626
rect 21730 117574 21782 117626
rect 21834 117574 21886 117626
rect 28430 117574 28482 117626
rect 28534 117574 28586 117626
rect 28638 117574 28690 117626
rect 25678 117406 25730 117458
rect 13806 117182 13858 117234
rect 14702 117182 14754 117234
rect 17390 117182 17442 117234
rect 18398 117182 18450 117234
rect 20078 117182 20130 117234
rect 20750 117182 20802 117234
rect 25342 117182 25394 117234
rect 16046 117070 16098 117122
rect 16382 117070 16434 117122
rect 16830 117070 16882 117122
rect 22318 117070 22370 117122
rect 22654 117070 22706 117122
rect 24670 117070 24722 117122
rect 19518 116958 19570 117010
rect 4616 116790 4668 116842
rect 4720 116790 4772 116842
rect 4824 116790 4876 116842
rect 11420 116790 11472 116842
rect 11524 116790 11576 116842
rect 11628 116790 11680 116842
rect 18224 116790 18276 116842
rect 18328 116790 18380 116842
rect 18432 116790 18484 116842
rect 25028 116790 25080 116842
rect 25132 116790 25184 116842
rect 25236 116790 25288 116842
rect 16270 116510 16322 116562
rect 18622 116510 18674 116562
rect 19854 116510 19906 116562
rect 10782 116398 10834 116450
rect 11454 116398 11506 116450
rect 13918 116398 13970 116450
rect 14926 116398 14978 116450
rect 16718 116398 16770 116450
rect 17726 116398 17778 116450
rect 13022 116174 13074 116226
rect 13582 116174 13634 116226
rect 20302 116174 20354 116226
rect 20750 116174 20802 116226
rect 8018 116006 8070 116058
rect 8122 116006 8174 116058
rect 8226 116006 8278 116058
rect 14822 116006 14874 116058
rect 14926 116006 14978 116058
rect 15030 116006 15082 116058
rect 21626 116006 21678 116058
rect 21730 116006 21782 116058
rect 21834 116006 21886 116058
rect 28430 116006 28482 116058
rect 28534 116006 28586 116058
rect 28638 116006 28690 116058
rect 12686 115838 12738 115890
rect 16158 115838 16210 115890
rect 19742 115838 19794 115890
rect 1710 115726 1762 115778
rect 11230 115614 11282 115666
rect 12238 115614 12290 115666
rect 13470 115614 13522 115666
rect 14478 115614 14530 115666
rect 17502 115614 17554 115666
rect 18398 115614 18450 115666
rect 20078 115614 20130 115666
rect 20862 115614 20914 115666
rect 22318 115502 22370 115554
rect 22654 115502 22706 115554
rect 10110 115390 10162 115442
rect 15598 115390 15650 115442
rect 4616 115222 4668 115274
rect 4720 115222 4772 115274
rect 4824 115222 4876 115274
rect 11420 115222 11472 115274
rect 11524 115222 11576 115274
rect 11628 115222 11680 115274
rect 18224 115222 18276 115274
rect 18328 115222 18380 115274
rect 18432 115222 18484 115274
rect 25028 115222 25080 115274
rect 25132 115222 25184 115274
rect 25236 115222 25288 115274
rect 15710 114942 15762 114994
rect 19854 114942 19906 114994
rect 17278 114830 17330 114882
rect 18062 114830 18114 114882
rect 21422 114830 21474 114882
rect 22430 114830 22482 114882
rect 18510 114606 18562 114658
rect 23774 114606 23826 114658
rect 24110 114606 24162 114658
rect 8018 114438 8070 114490
rect 8122 114438 8174 114490
rect 8226 114438 8278 114490
rect 14822 114438 14874 114490
rect 14926 114438 14978 114490
rect 15030 114438 15082 114490
rect 21626 114438 21678 114490
rect 21730 114438 21782 114490
rect 21834 114438 21886 114490
rect 28430 114438 28482 114490
rect 28534 114438 28586 114490
rect 28638 114438 28690 114490
rect 11230 114046 11282 114098
rect 12126 114046 12178 114098
rect 13582 114046 13634 114098
rect 14590 114046 14642 114098
rect 17502 114046 17554 114098
rect 18174 114046 18226 114098
rect 20078 114046 20130 114098
rect 20862 114046 20914 114098
rect 16270 113934 16322 113986
rect 22654 113934 22706 113986
rect 10110 113822 10162 113874
rect 15710 113822 15762 113874
rect 19518 113822 19570 113874
rect 22094 113822 22146 113874
rect 4616 113654 4668 113706
rect 4720 113654 4772 113706
rect 4824 113654 4876 113706
rect 11420 113654 11472 113706
rect 11524 113654 11576 113706
rect 11628 113654 11680 113706
rect 18224 113654 18276 113706
rect 18328 113654 18380 113706
rect 18432 113654 18484 113706
rect 25028 113654 25080 113706
rect 25132 113654 25184 113706
rect 25236 113654 25288 113706
rect 22094 113486 22146 113538
rect 16382 113374 16434 113426
rect 7982 113262 8034 113314
rect 8878 113262 8930 113314
rect 10558 113262 10610 113314
rect 11230 113262 11282 113314
rect 18622 113262 18674 113314
rect 19294 113262 19346 113314
rect 23438 113262 23490 113314
rect 24110 113262 24162 113314
rect 25902 113262 25954 113314
rect 26686 113262 26738 113314
rect 10222 113038 10274 113090
rect 12798 113038 12850 113090
rect 13806 113038 13858 113090
rect 20862 113038 20914 113090
rect 21422 113038 21474 113090
rect 28254 113038 28306 113090
rect 8018 112870 8070 112922
rect 8122 112870 8174 112922
rect 8226 112870 8278 112922
rect 14822 112870 14874 112922
rect 14926 112870 14978 112922
rect 15030 112870 15082 112922
rect 21626 112870 21678 112922
rect 21730 112870 21782 112922
rect 21834 112870 21886 112922
rect 28430 112870 28482 112922
rect 28534 112870 28586 112922
rect 28638 112870 28690 112922
rect 28254 112702 28306 112754
rect 11454 112478 11506 112530
rect 12126 112478 12178 112530
rect 13918 112478 13970 112530
rect 14702 112478 14754 112530
rect 16606 112478 16658 112530
rect 19182 112478 19234 112530
rect 19966 112478 20018 112530
rect 22542 112478 22594 112530
rect 23438 112478 23490 112530
rect 24782 112478 24834 112530
rect 25902 112478 25954 112530
rect 26686 112478 26738 112530
rect 21534 112366 21586 112418
rect 21870 112366 21922 112418
rect 13470 112254 13522 112306
rect 16046 112254 16098 112306
rect 4616 112086 4668 112138
rect 4720 112086 4772 112138
rect 4824 112086 4876 112138
rect 11420 112086 11472 112138
rect 11524 112086 11576 112138
rect 11628 112086 11680 112138
rect 18224 112086 18276 112138
rect 18328 112086 18380 112138
rect 18432 112086 18484 112138
rect 25028 112086 25080 112138
rect 25132 112086 25184 112138
rect 25236 112086 25288 112138
rect 11678 111918 11730 111970
rect 16046 111918 16098 111970
rect 25230 111918 25282 111970
rect 28030 111806 28082 111858
rect 8318 111694 8370 111746
rect 9214 111694 9266 111746
rect 9550 111694 9602 111746
rect 10334 111694 10386 111746
rect 13918 111694 13970 111746
rect 14702 111694 14754 111746
rect 16718 111694 16770 111746
rect 17390 111694 17442 111746
rect 18958 111694 19010 111746
rect 19294 111694 19346 111746
rect 23214 111694 23266 111746
rect 24110 111694 24162 111746
rect 25790 111694 25842 111746
rect 26686 111694 26738 111746
rect 6862 111470 6914 111522
rect 12350 111470 12402 111522
rect 13694 111470 13746 111522
rect 8018 111302 8070 111354
rect 8122 111302 8174 111354
rect 8226 111302 8278 111354
rect 14822 111302 14874 111354
rect 14926 111302 14978 111354
rect 15030 111302 15082 111354
rect 21626 111302 21678 111354
rect 21730 111302 21782 111354
rect 21834 111302 21886 111354
rect 28430 111302 28482 111354
rect 28534 111302 28586 111354
rect 28638 111302 28690 111354
rect 28254 111134 28306 111186
rect 12686 111022 12738 111074
rect 9550 110910 9602 110962
rect 10334 110910 10386 110962
rect 12126 110910 12178 110962
rect 13918 110910 13970 110962
rect 14702 110910 14754 110962
rect 17502 110910 17554 110962
rect 18174 110910 18226 110962
rect 20078 110910 20130 110962
rect 20750 110910 20802 110962
rect 25902 110910 25954 110962
rect 26686 110910 26738 110962
rect 13134 110798 13186 110850
rect 13582 110798 13634 110850
rect 16606 110798 16658 110850
rect 22318 110798 22370 110850
rect 22654 110798 22706 110850
rect 11678 110686 11730 110738
rect 16046 110686 16098 110738
rect 19518 110686 19570 110738
rect 4616 110518 4668 110570
rect 4720 110518 4772 110570
rect 4824 110518 4876 110570
rect 11420 110518 11472 110570
rect 11524 110518 11576 110570
rect 11628 110518 11680 110570
rect 18224 110518 18276 110570
rect 18328 110518 18380 110570
rect 18432 110518 18484 110570
rect 25028 110518 25080 110570
rect 25132 110518 25184 110570
rect 25236 110518 25288 110570
rect 11006 110350 11058 110402
rect 12014 110350 12066 110402
rect 16046 110350 16098 110402
rect 11454 110238 11506 110290
rect 16606 110238 16658 110290
rect 19854 110238 19906 110290
rect 28254 110238 28306 110290
rect 8878 110126 8930 110178
rect 9662 110126 9714 110178
rect 11678 110126 11730 110178
rect 12686 110126 12738 110178
rect 12910 110126 12962 110178
rect 13918 110126 13970 110178
rect 14702 110126 14754 110178
rect 21422 110126 21474 110178
rect 22318 110126 22370 110178
rect 25902 110126 25954 110178
rect 26686 110126 26738 110178
rect 13470 110014 13522 110066
rect 23662 110014 23714 110066
rect 12350 109902 12402 109954
rect 13582 109902 13634 109954
rect 19406 109902 19458 109954
rect 20638 109902 20690 109954
rect 23998 109902 24050 109954
rect 8018 109734 8070 109786
rect 8122 109734 8174 109786
rect 8226 109734 8278 109786
rect 14822 109734 14874 109786
rect 14926 109734 14978 109786
rect 15030 109734 15082 109786
rect 21626 109734 21678 109786
rect 21730 109734 21782 109786
rect 21834 109734 21886 109786
rect 28430 109734 28482 109786
rect 28534 109734 28586 109786
rect 28638 109734 28690 109786
rect 21422 109566 21474 109618
rect 28254 109566 28306 109618
rect 12126 109454 12178 109506
rect 14254 109454 14306 109506
rect 20526 109454 20578 109506
rect 10782 109342 10834 109394
rect 11678 109342 11730 109394
rect 12350 109342 12402 109394
rect 13582 109342 13634 109394
rect 15374 109342 15426 109394
rect 15822 109342 15874 109394
rect 16718 109342 16770 109394
rect 19518 109342 19570 109394
rect 21310 109342 21362 109394
rect 25902 109342 25954 109394
rect 26686 109342 26738 109394
rect 13022 109230 13074 109282
rect 16158 109230 16210 109282
rect 18174 109230 18226 109282
rect 18958 109230 19010 109282
rect 19966 109230 20018 109282
rect 22430 109230 22482 109282
rect 9662 109118 9714 109170
rect 4616 108950 4668 109002
rect 4720 108950 4772 109002
rect 4824 108950 4876 109002
rect 11420 108950 11472 109002
rect 11524 108950 11576 109002
rect 11628 108950 11680 109002
rect 18224 108950 18276 109002
rect 18328 108950 18380 109002
rect 18432 108950 18484 109002
rect 25028 108950 25080 109002
rect 25132 108950 25184 109002
rect 25236 108950 25288 109002
rect 9662 108782 9714 108834
rect 12798 108782 12850 108834
rect 14254 108782 14306 108834
rect 16942 108782 16994 108834
rect 21310 108782 21362 108834
rect 8990 108670 9042 108722
rect 14030 108670 14082 108722
rect 15038 108670 15090 108722
rect 17390 108670 17442 108722
rect 18734 108670 18786 108722
rect 20414 108670 20466 108722
rect 10782 108558 10834 108610
rect 11678 108558 11730 108610
rect 12574 108558 12626 108610
rect 12798 108558 12850 108610
rect 13694 108558 13746 108610
rect 14926 108558 14978 108610
rect 16942 108558 16994 108610
rect 17838 108558 17890 108610
rect 18510 108558 18562 108610
rect 19854 108558 19906 108610
rect 22318 108558 22370 108610
rect 23102 108558 23154 108610
rect 24894 108558 24946 108610
rect 25678 108558 25730 108610
rect 9214 108446 9266 108498
rect 16046 108446 16098 108498
rect 16606 108446 16658 108498
rect 18174 108446 18226 108498
rect 19182 108446 19234 108498
rect 20750 108446 20802 108498
rect 21422 108446 21474 108498
rect 15710 108334 15762 108386
rect 17278 108334 17330 108386
rect 17502 108334 17554 108386
rect 19070 108334 19122 108386
rect 21870 108334 21922 108386
rect 24670 108334 24722 108386
rect 27246 108334 27298 108386
rect 8018 108166 8070 108218
rect 8122 108166 8174 108218
rect 8226 108166 8278 108218
rect 14822 108166 14874 108218
rect 14926 108166 14978 108218
rect 15030 108166 15082 108218
rect 21626 108166 21678 108218
rect 21730 108166 21782 108218
rect 21834 108166 21886 108218
rect 28430 108166 28482 108218
rect 28534 108166 28586 108218
rect 28638 108166 28690 108218
rect 14478 107998 14530 108050
rect 20526 107998 20578 108050
rect 21086 107998 21138 108050
rect 28254 107998 28306 108050
rect 13134 107886 13186 107938
rect 17390 107886 17442 107938
rect 10782 107774 10834 107826
rect 11678 107774 11730 107826
rect 12126 107774 12178 107826
rect 12350 107774 12402 107826
rect 12686 107774 12738 107826
rect 13582 107774 13634 107826
rect 16046 107774 16098 107826
rect 16718 107774 16770 107826
rect 17726 107774 17778 107826
rect 18174 107774 18226 107826
rect 19182 107774 19234 107826
rect 20750 107774 20802 107826
rect 22318 107774 22370 107826
rect 23102 107774 23154 107826
rect 25902 107774 25954 107826
rect 26686 107774 26738 107826
rect 8990 107662 9042 107714
rect 12238 107662 12290 107714
rect 14030 107662 14082 107714
rect 21534 107662 21586 107714
rect 9662 107550 9714 107602
rect 24334 107550 24386 107602
rect 4616 107382 4668 107434
rect 4720 107382 4772 107434
rect 4824 107382 4876 107434
rect 11420 107382 11472 107434
rect 11524 107382 11576 107434
rect 11628 107382 11680 107434
rect 18224 107382 18276 107434
rect 18328 107382 18380 107434
rect 18432 107382 18484 107434
rect 25028 107382 25080 107434
rect 25132 107382 25184 107434
rect 25236 107382 25288 107434
rect 8542 107214 8594 107266
rect 8990 107214 9042 107266
rect 9438 107214 9490 107266
rect 9886 107214 9938 107266
rect 14926 107214 14978 107266
rect 21534 107214 21586 107266
rect 9438 107102 9490 107154
rect 9886 107102 9938 107154
rect 14254 107102 14306 107154
rect 20078 107102 20130 107154
rect 25006 107102 25058 107154
rect 28254 107102 28306 107154
rect 11454 106990 11506 107042
rect 12462 106990 12514 107042
rect 13582 106990 13634 107042
rect 14590 106990 14642 107042
rect 15486 106990 15538 107042
rect 16158 106990 16210 107042
rect 18174 106990 18226 107042
rect 19182 106990 19234 107042
rect 21310 106990 21362 107042
rect 22318 106990 22370 107042
rect 23102 106990 23154 107042
rect 25902 106990 25954 107042
rect 26686 106990 26738 107042
rect 13470 106878 13522 106930
rect 7534 106766 7586 106818
rect 8094 106766 8146 106818
rect 8542 106766 8594 106818
rect 9102 106766 9154 106818
rect 10110 106766 10162 106818
rect 13022 106766 13074 106818
rect 17726 106766 17778 106818
rect 21870 106766 21922 106818
rect 24670 106766 24722 106818
rect 8018 106598 8070 106650
rect 8122 106598 8174 106650
rect 8226 106598 8278 106650
rect 14822 106598 14874 106650
rect 14926 106598 14978 106650
rect 15030 106598 15082 106650
rect 21626 106598 21678 106650
rect 21730 106598 21782 106650
rect 21834 106598 21886 106650
rect 28430 106598 28482 106650
rect 28534 106598 28586 106650
rect 28638 106598 28690 106650
rect 9886 106430 9938 106482
rect 16830 106430 16882 106482
rect 19854 106430 19906 106482
rect 21310 106430 21362 106482
rect 22766 106430 22818 106482
rect 28254 106430 28306 106482
rect 3166 106318 3218 106370
rect 9102 106318 9154 106370
rect 9774 106318 9826 106370
rect 21870 106318 21922 106370
rect 6078 106206 6130 106258
rect 8094 106206 8146 106258
rect 15486 106206 15538 106258
rect 15934 106206 15986 106258
rect 17502 106206 17554 106258
rect 18286 106206 18338 106258
rect 22206 106206 22258 106258
rect 25342 106206 25394 106258
rect 25902 106206 25954 106258
rect 26686 106206 26738 106258
rect 3278 106094 3330 106146
rect 3838 106094 3890 106146
rect 4734 106094 4786 106146
rect 5294 106094 5346 106146
rect 5742 106094 5794 106146
rect 6302 106094 6354 106146
rect 7310 106094 7362 106146
rect 7646 106094 7698 106146
rect 8542 106094 8594 106146
rect 11230 106094 11282 106146
rect 16270 106094 16322 106146
rect 20190 106094 20242 106146
rect 23326 106094 23378 106146
rect 23774 106094 23826 106146
rect 3390 105982 3442 106034
rect 6414 105982 6466 106034
rect 7310 105982 7362 106034
rect 8318 105982 8370 106034
rect 8542 105982 8594 106034
rect 9102 105982 9154 106034
rect 15822 105982 15874 106034
rect 16494 105982 16546 106034
rect 23438 105982 23490 106034
rect 23998 105982 24050 106034
rect 24334 105982 24386 106034
rect 4616 105814 4668 105866
rect 4720 105814 4772 105866
rect 4824 105814 4876 105866
rect 11420 105814 11472 105866
rect 11524 105814 11576 105866
rect 11628 105814 11680 105866
rect 18224 105814 18276 105866
rect 18328 105814 18380 105866
rect 18432 105814 18484 105866
rect 25028 105814 25080 105866
rect 25132 105814 25184 105866
rect 25236 105814 25288 105866
rect 9662 105646 9714 105698
rect 19966 105646 20018 105698
rect 22542 105646 22594 105698
rect 1710 105534 1762 105586
rect 3838 105534 3890 105586
rect 5630 105534 5682 105586
rect 7758 105534 7810 105586
rect 16382 105534 16434 105586
rect 22206 105534 22258 105586
rect 26238 105534 26290 105586
rect 4510 105422 4562 105474
rect 8542 105422 8594 105474
rect 10782 105422 10834 105474
rect 11678 105422 11730 105474
rect 12686 105422 12738 105474
rect 13806 105422 13858 105474
rect 14030 105422 14082 105474
rect 14590 105422 14642 105474
rect 20302 105422 20354 105474
rect 20526 105422 20578 105474
rect 22542 105422 22594 105474
rect 23214 105422 23266 105474
rect 24446 105422 24498 105474
rect 25006 105422 25058 105474
rect 8878 105310 8930 105362
rect 21310 105310 21362 105362
rect 21534 105310 21586 105362
rect 23886 105310 23938 105362
rect 5182 105198 5234 105250
rect 8990 105198 9042 105250
rect 12462 105198 12514 105250
rect 12798 105198 12850 105250
rect 12910 105198 12962 105250
rect 13470 105198 13522 105250
rect 21422 105198 21474 105250
rect 25342 105198 25394 105250
rect 25678 105198 25730 105250
rect 26686 105198 26738 105250
rect 8018 105030 8070 105082
rect 8122 105030 8174 105082
rect 8226 105030 8278 105082
rect 14822 105030 14874 105082
rect 14926 105030 14978 105082
rect 15030 105030 15082 105082
rect 21626 105030 21678 105082
rect 21730 105030 21782 105082
rect 21834 105030 21886 105082
rect 28430 105030 28482 105082
rect 28534 105030 28586 105082
rect 28638 105030 28690 105082
rect 3838 104862 3890 104914
rect 3950 104862 4002 104914
rect 4062 104862 4114 104914
rect 6750 104862 6802 104914
rect 7982 104862 8034 104914
rect 8094 104862 8146 104914
rect 28030 104862 28082 104914
rect 4286 104750 4338 104802
rect 7310 104750 7362 104802
rect 7534 104750 7586 104802
rect 8318 104750 8370 104802
rect 8990 104750 9042 104802
rect 10446 104750 10498 104802
rect 19070 104750 19122 104802
rect 25230 104750 25282 104802
rect 3726 104638 3778 104690
rect 5182 104638 5234 104690
rect 6526 104638 6578 104690
rect 6638 104638 6690 104690
rect 6862 104638 6914 104690
rect 7086 104638 7138 104690
rect 7646 104638 7698 104690
rect 7870 104638 7922 104690
rect 8654 104638 8706 104690
rect 9662 104638 9714 104690
rect 11230 104638 11282 104690
rect 11790 104638 11842 104690
rect 18174 104638 18226 104690
rect 19406 104638 19458 104690
rect 25678 104638 25730 104690
rect 26686 104638 26738 104690
rect 2830 104526 2882 104578
rect 3278 104526 3330 104578
rect 4734 104526 4786 104578
rect 5630 104526 5682 104578
rect 6078 104526 6130 104578
rect 15486 104526 15538 104578
rect 17614 104526 17666 104578
rect 18510 104526 18562 104578
rect 22206 104526 22258 104578
rect 2942 104414 2994 104466
rect 3390 104414 3442 104466
rect 4616 104246 4668 104298
rect 4720 104246 4772 104298
rect 4824 104246 4876 104298
rect 11420 104246 11472 104298
rect 11524 104246 11576 104298
rect 11628 104246 11680 104298
rect 18224 104246 18276 104298
rect 18328 104246 18380 104298
rect 18432 104246 18484 104298
rect 25028 104246 25080 104298
rect 25132 104246 25184 104298
rect 25236 104246 25288 104298
rect 14702 104078 14754 104130
rect 27582 104078 27634 104130
rect 1710 103966 1762 104018
rect 5854 103966 5906 104018
rect 11230 103966 11282 104018
rect 12350 103966 12402 104018
rect 13582 103966 13634 104018
rect 23662 103966 23714 104018
rect 24670 103966 24722 104018
rect 26014 103966 26066 104018
rect 4510 103854 4562 103906
rect 8654 103854 8706 103906
rect 9886 103854 9938 103906
rect 10670 103854 10722 103906
rect 10894 103854 10946 103906
rect 12126 103854 12178 103906
rect 12238 103854 12290 103906
rect 13918 103854 13970 103906
rect 15038 103854 15090 103906
rect 15486 103854 15538 103906
rect 21422 103854 21474 103906
rect 22318 103854 22370 103906
rect 24446 103854 24498 103906
rect 24894 103854 24946 103906
rect 27694 103854 27746 103906
rect 3838 103742 3890 103794
rect 7982 103742 8034 103794
rect 9326 103742 9378 103794
rect 9662 103742 9714 103794
rect 11118 103742 11170 103794
rect 13806 103742 13858 103794
rect 17502 103742 17554 103794
rect 26910 103742 26962 103794
rect 5070 103630 5122 103682
rect 9214 103630 9266 103682
rect 10222 103630 10274 103682
rect 11342 103630 11394 103682
rect 13022 103630 13074 103682
rect 14142 103630 14194 103682
rect 14366 103630 14418 103682
rect 14814 103630 14866 103682
rect 24110 103630 24162 103682
rect 8018 103462 8070 103514
rect 8122 103462 8174 103514
rect 8226 103462 8278 103514
rect 14822 103462 14874 103514
rect 14926 103462 14978 103514
rect 15030 103462 15082 103514
rect 21626 103462 21678 103514
rect 21730 103462 21782 103514
rect 21834 103462 21886 103514
rect 28430 103462 28482 103514
rect 28534 103462 28586 103514
rect 28638 103462 28690 103514
rect 4286 103294 4338 103346
rect 5294 103294 5346 103346
rect 6974 103294 7026 103346
rect 7086 103294 7138 103346
rect 7870 103294 7922 103346
rect 8990 103294 9042 103346
rect 9550 103294 9602 103346
rect 17502 103294 17554 103346
rect 18398 103294 18450 103346
rect 22878 103294 22930 103346
rect 23326 103294 23378 103346
rect 23662 103294 23714 103346
rect 23998 103294 24050 103346
rect 3502 103182 3554 103234
rect 3726 103182 3778 103234
rect 4062 103182 4114 103234
rect 7198 103182 7250 103234
rect 7758 103182 7810 103234
rect 18286 103182 18338 103234
rect 2606 103070 2658 103122
rect 3278 103070 3330 103122
rect 3950 103070 4002 103122
rect 4398 103070 4450 103122
rect 7646 103070 7698 103122
rect 8094 103070 8146 103122
rect 8318 103070 8370 103122
rect 8766 103070 8818 103122
rect 9774 103070 9826 103122
rect 9998 103070 10050 103122
rect 10222 103070 10274 103122
rect 10670 103070 10722 103122
rect 10894 103070 10946 103122
rect 11790 103070 11842 103122
rect 12126 103070 12178 103122
rect 12574 103070 12626 103122
rect 13134 103070 13186 103122
rect 14030 103070 14082 103122
rect 14926 103070 14978 103122
rect 16158 103070 16210 103122
rect 17278 103070 17330 103122
rect 17726 103070 17778 103122
rect 17950 103070 18002 103122
rect 18846 103070 18898 103122
rect 22206 103070 22258 103122
rect 24222 103070 24274 103122
rect 2158 102958 2210 103010
rect 2942 102958 2994 103010
rect 5630 102958 5682 103010
rect 6078 102958 6130 103010
rect 6526 102958 6578 103010
rect 8878 102958 8930 103010
rect 10782 102958 10834 103010
rect 12238 102958 12290 103010
rect 14254 102958 14306 103010
rect 19518 102958 19570 103010
rect 21646 102958 21698 103010
rect 21982 102958 22034 103010
rect 22542 102958 22594 103010
rect 22990 102958 23042 103010
rect 25342 102958 25394 103010
rect 5070 102846 5122 102898
rect 6078 102846 6130 102898
rect 9438 102846 9490 102898
rect 12686 102846 12738 102898
rect 4616 102678 4668 102730
rect 4720 102678 4772 102730
rect 4824 102678 4876 102730
rect 11420 102678 11472 102730
rect 11524 102678 11576 102730
rect 11628 102678 11680 102730
rect 18224 102678 18276 102730
rect 18328 102678 18380 102730
rect 18432 102678 18484 102730
rect 25028 102678 25080 102730
rect 25132 102678 25184 102730
rect 25236 102678 25288 102730
rect 4174 102510 4226 102562
rect 5070 102510 5122 102562
rect 8318 102510 8370 102562
rect 12238 102510 12290 102562
rect 22542 102510 22594 102562
rect 5966 102398 6018 102450
rect 8654 102398 8706 102450
rect 11118 102398 11170 102450
rect 16830 102398 16882 102450
rect 20190 102398 20242 102450
rect 20638 102398 20690 102450
rect 20750 102398 20802 102450
rect 22766 102398 22818 102450
rect 23662 102398 23714 102450
rect 24222 102398 24274 102450
rect 24782 102398 24834 102450
rect 3390 102286 3442 102338
rect 7646 102286 7698 102338
rect 8878 102286 8930 102338
rect 9214 102286 9266 102338
rect 9550 102286 9602 102338
rect 10110 102286 10162 102338
rect 12350 102286 12402 102338
rect 12574 102286 12626 102338
rect 12798 102286 12850 102338
rect 13806 102286 13858 102338
rect 14254 102286 14306 102338
rect 20414 102286 20466 102338
rect 21534 102286 21586 102338
rect 21870 102286 21922 102338
rect 23214 102286 23266 102338
rect 23998 102286 24050 102338
rect 9662 102174 9714 102226
rect 13470 102174 13522 102226
rect 13582 102174 13634 102226
rect 19742 102174 19794 102226
rect 19966 102174 20018 102226
rect 24334 102174 24386 102226
rect 2606 102062 2658 102114
rect 3054 102062 3106 102114
rect 3502 102062 3554 102114
rect 3726 102062 3778 102114
rect 4286 102062 4338 102114
rect 4734 102062 4786 102114
rect 5070 102062 5122 102114
rect 6526 102062 6578 102114
rect 6862 102062 6914 102114
rect 7310 102062 7362 102114
rect 7758 102062 7810 102114
rect 9774 102062 9826 102114
rect 12238 102062 12290 102114
rect 21310 102062 21362 102114
rect 21422 102062 21474 102114
rect 22206 102062 22258 102114
rect 8018 101894 8070 101946
rect 8122 101894 8174 101946
rect 8226 101894 8278 101946
rect 14822 101894 14874 101946
rect 14926 101894 14978 101946
rect 15030 101894 15082 101946
rect 21626 101894 21678 101946
rect 21730 101894 21782 101946
rect 21834 101894 21886 101946
rect 28430 101894 28482 101946
rect 28534 101894 28586 101946
rect 28638 101894 28690 101946
rect 17502 101726 17554 101778
rect 9886 101614 9938 101666
rect 19406 101614 19458 101666
rect 24558 101614 24610 101666
rect 4510 101502 4562 101554
rect 5854 101502 5906 101554
rect 10222 101502 10274 101554
rect 11118 101502 11170 101554
rect 12238 101502 12290 101554
rect 22206 101502 22258 101554
rect 23326 101502 23378 101554
rect 23662 101502 23714 101554
rect 23886 101502 23938 101554
rect 1710 101390 1762 101442
rect 3838 101390 3890 101442
rect 5182 101390 5234 101442
rect 5630 101390 5682 101442
rect 6638 101390 6690 101442
rect 8766 101390 8818 101442
rect 10670 101390 10722 101442
rect 14254 101390 14306 101442
rect 23550 101390 23602 101442
rect 25342 101390 25394 101442
rect 24334 101278 24386 101330
rect 24670 101278 24722 101330
rect 4616 101110 4668 101162
rect 4720 101110 4772 101162
rect 4824 101110 4876 101162
rect 11420 101110 11472 101162
rect 11524 101110 11576 101162
rect 11628 101110 11680 101162
rect 18224 101110 18276 101162
rect 18328 101110 18380 101162
rect 18432 101110 18484 101162
rect 25028 101110 25080 101162
rect 25132 101110 25184 101162
rect 25236 101110 25288 101162
rect 3726 100830 3778 100882
rect 6302 100830 6354 100882
rect 7422 100830 7474 100882
rect 10670 100830 10722 100882
rect 12574 100830 12626 100882
rect 21310 100830 21362 100882
rect 24558 100830 24610 100882
rect 3278 100718 3330 100770
rect 3502 100718 3554 100770
rect 3950 100718 4002 100770
rect 5742 100718 5794 100770
rect 7310 100718 7362 100770
rect 9326 100718 9378 100770
rect 10446 100718 10498 100770
rect 12910 100718 12962 100770
rect 13470 100718 13522 100770
rect 19742 100718 19794 100770
rect 20078 100718 20130 100770
rect 24222 100718 24274 100770
rect 27358 100718 27410 100770
rect 2606 100606 2658 100658
rect 4846 100606 4898 100658
rect 6414 100606 6466 100658
rect 7758 100606 7810 100658
rect 9550 100606 9602 100658
rect 15486 100606 15538 100658
rect 20302 100606 20354 100658
rect 23438 100606 23490 100658
rect 26686 100606 26738 100658
rect 2158 100494 2210 100546
rect 3054 100494 3106 100546
rect 4510 100494 4562 100546
rect 4958 100494 5010 100546
rect 5182 100494 5234 100546
rect 6190 100494 6242 100546
rect 7422 100494 7474 100546
rect 20750 100494 20802 100546
rect 8018 100326 8070 100378
rect 8122 100326 8174 100378
rect 8226 100326 8278 100378
rect 14822 100326 14874 100378
rect 14926 100326 14978 100378
rect 15030 100326 15082 100378
rect 21626 100326 21678 100378
rect 21730 100326 21782 100378
rect 21834 100326 21886 100378
rect 28430 100326 28482 100378
rect 28534 100326 28586 100378
rect 28638 100326 28690 100378
rect 4286 100158 4338 100210
rect 8766 100158 8818 100210
rect 8990 100158 9042 100210
rect 23438 100158 23490 100210
rect 23550 100158 23602 100210
rect 25230 100158 25282 100210
rect 25342 100158 25394 100210
rect 3502 100046 3554 100098
rect 5294 100046 5346 100098
rect 8542 100046 8594 100098
rect 11118 100046 11170 100098
rect 21198 100046 21250 100098
rect 25678 100046 25730 100098
rect 2942 99934 2994 99986
rect 3166 99934 3218 99986
rect 4622 99934 4674 99986
rect 10110 99934 10162 99986
rect 11790 99934 11842 99986
rect 18286 99934 18338 99986
rect 22878 99934 22930 99986
rect 23326 99934 23378 99986
rect 24110 99934 24162 99986
rect 25454 99934 25506 99986
rect 2158 99822 2210 99874
rect 2606 99822 2658 99874
rect 2830 99822 2882 99874
rect 3390 99822 3442 99874
rect 2158 99710 2210 99762
rect 7422 99822 7474 99874
rect 8206 99822 8258 99874
rect 8878 99822 8930 99874
rect 10782 99822 10834 99874
rect 13582 99822 13634 99874
rect 23886 99822 23938 99874
rect 26238 99822 26290 99874
rect 26686 99822 26738 99874
rect 24446 99710 24498 99762
rect 4616 99542 4668 99594
rect 4720 99542 4772 99594
rect 4824 99542 4876 99594
rect 11420 99542 11472 99594
rect 11524 99542 11576 99594
rect 11628 99542 11680 99594
rect 18224 99542 18276 99594
rect 18328 99542 18380 99594
rect 18432 99542 18484 99594
rect 25028 99542 25080 99594
rect 25132 99542 25184 99594
rect 25236 99542 25288 99594
rect 22318 99374 22370 99426
rect 1710 99262 1762 99314
rect 3838 99262 3890 99314
rect 5182 99262 5234 99314
rect 11790 99262 11842 99314
rect 15486 99262 15538 99314
rect 20638 99262 20690 99314
rect 24894 99262 24946 99314
rect 4622 99150 4674 99202
rect 5854 99150 5906 99202
rect 6078 99150 6130 99202
rect 6302 99150 6354 99202
rect 6638 99150 6690 99202
rect 6750 99150 6802 99202
rect 7422 99150 7474 99202
rect 7646 99150 7698 99202
rect 14254 99150 14306 99202
rect 19182 99150 19234 99202
rect 19854 99150 19906 99202
rect 20190 99150 20242 99202
rect 21534 99150 21586 99202
rect 21758 99150 21810 99202
rect 21870 99150 21922 99202
rect 22878 99150 22930 99202
rect 6526 99038 6578 99090
rect 7086 99038 7138 99090
rect 6862 98926 6914 98978
rect 19070 98926 19122 98978
rect 19294 98926 19346 98978
rect 19518 98926 19570 98978
rect 20078 98926 20130 98978
rect 8018 98758 8070 98810
rect 8122 98758 8174 98810
rect 8226 98758 8278 98810
rect 14822 98758 14874 98810
rect 14926 98758 14978 98810
rect 15030 98758 15082 98810
rect 21626 98758 21678 98810
rect 21730 98758 21782 98810
rect 21834 98758 21886 98810
rect 28430 98758 28482 98810
rect 28534 98758 28586 98810
rect 28638 98758 28690 98810
rect 2830 98590 2882 98642
rect 3054 98590 3106 98642
rect 3278 98590 3330 98642
rect 4398 98590 4450 98642
rect 10894 98590 10946 98642
rect 18062 98590 18114 98642
rect 18174 98590 18226 98642
rect 18734 98590 18786 98642
rect 18846 98590 18898 98642
rect 21870 98590 21922 98642
rect 22766 98590 22818 98642
rect 23886 98590 23938 98642
rect 4062 98478 4114 98530
rect 6638 98478 6690 98530
rect 9886 98478 9938 98530
rect 11790 98478 11842 98530
rect 17838 98478 17890 98530
rect 17950 98478 18002 98530
rect 20862 98478 20914 98530
rect 21198 98478 21250 98530
rect 24446 98478 24498 98530
rect 3390 98366 3442 98418
rect 5182 98366 5234 98418
rect 5966 98366 6018 98418
rect 9550 98366 9602 98418
rect 9774 98366 9826 98418
rect 10110 98366 10162 98418
rect 10334 98366 10386 98418
rect 10782 98366 10834 98418
rect 15598 98366 15650 98418
rect 18286 98366 18338 98418
rect 18622 98366 18674 98418
rect 19182 98366 19234 98418
rect 20190 98366 20242 98418
rect 23998 98366 24050 98418
rect 24558 98366 24610 98418
rect 28030 98366 28082 98418
rect 2382 98254 2434 98306
rect 4846 98254 4898 98306
rect 5406 98254 5458 98306
rect 8766 98254 8818 98306
rect 19742 98254 19794 98306
rect 22318 98254 22370 98306
rect 23550 98254 23602 98306
rect 25230 98254 25282 98306
rect 27358 98254 27410 98306
rect 5518 98142 5570 98194
rect 20526 98142 20578 98194
rect 21870 98142 21922 98194
rect 22318 98142 22370 98194
rect 23886 98142 23938 98194
rect 24446 98142 24498 98194
rect 4616 97974 4668 98026
rect 4720 97974 4772 98026
rect 4824 97974 4876 98026
rect 11420 97974 11472 98026
rect 11524 97974 11576 98026
rect 11628 97974 11680 98026
rect 18224 97974 18276 98026
rect 18328 97974 18380 98026
rect 18432 97974 18484 98026
rect 25028 97974 25080 98026
rect 25132 97974 25184 98026
rect 25236 97974 25288 98026
rect 15150 97806 15202 97858
rect 23438 97806 23490 97858
rect 25342 97806 25394 97858
rect 3278 97694 3330 97746
rect 4622 97694 4674 97746
rect 17726 97694 17778 97746
rect 21870 97694 21922 97746
rect 22542 97694 22594 97746
rect 24446 97694 24498 97746
rect 25454 97694 25506 97746
rect 3838 97582 3890 97634
rect 5742 97582 5794 97634
rect 5854 97582 5906 97634
rect 6078 97582 6130 97634
rect 6190 97582 6242 97634
rect 6750 97582 6802 97634
rect 6862 97582 6914 97634
rect 7870 97582 7922 97634
rect 14702 97582 14754 97634
rect 15038 97582 15090 97634
rect 15934 97582 15986 97634
rect 16606 97582 16658 97634
rect 17502 97582 17554 97634
rect 19294 97582 19346 97634
rect 20078 97582 20130 97634
rect 23102 97582 23154 97634
rect 23550 97582 23602 97634
rect 24222 97582 24274 97634
rect 25678 97582 25730 97634
rect 27358 97582 27410 97634
rect 5070 97470 5122 97522
rect 7198 97470 7250 97522
rect 10446 97470 10498 97522
rect 14142 97470 14194 97522
rect 16718 97470 16770 97522
rect 17390 97470 17442 97522
rect 18958 97470 19010 97522
rect 19966 97470 20018 97522
rect 21422 97470 21474 97522
rect 22878 97470 22930 97522
rect 24894 97470 24946 97522
rect 26686 97470 26738 97522
rect 26798 97470 26850 97522
rect 2830 97358 2882 97410
rect 4174 97358 4226 97410
rect 6974 97358 7026 97410
rect 13806 97358 13858 97410
rect 14030 97358 14082 97410
rect 14254 97358 14306 97410
rect 17726 97358 17778 97410
rect 17950 97358 18002 97410
rect 18398 97358 18450 97410
rect 20638 97358 20690 97410
rect 23326 97358 23378 97410
rect 27022 97358 27074 97410
rect 8018 97190 8070 97242
rect 8122 97190 8174 97242
rect 8226 97190 8278 97242
rect 14822 97190 14874 97242
rect 14926 97190 14978 97242
rect 15030 97190 15082 97242
rect 21626 97190 21678 97242
rect 21730 97190 21782 97242
rect 21834 97190 21886 97242
rect 28430 97190 28482 97242
rect 28534 97190 28586 97242
rect 28638 97190 28690 97242
rect 7534 97022 7586 97074
rect 8878 97022 8930 97074
rect 13806 97022 13858 97074
rect 18174 97022 18226 97074
rect 18510 97022 18562 97074
rect 23550 97022 23602 97074
rect 2270 96910 2322 96962
rect 2718 96910 2770 96962
rect 6302 96910 6354 96962
rect 11902 96910 11954 96962
rect 13470 96910 13522 96962
rect 13694 96910 13746 96962
rect 14030 96910 14082 96962
rect 15710 96910 15762 96962
rect 17950 96910 18002 96962
rect 20190 96910 20242 96962
rect 20862 96910 20914 96962
rect 21310 96910 21362 96962
rect 22654 96910 22706 96962
rect 27358 96910 27410 96962
rect 1934 96798 1986 96850
rect 2158 96798 2210 96850
rect 2494 96798 2546 96850
rect 2942 96798 2994 96850
rect 3278 96798 3330 96850
rect 6974 96798 7026 96850
rect 8542 96798 8594 96850
rect 8766 96798 8818 96850
rect 9102 96798 9154 96850
rect 10894 96798 10946 96850
rect 11790 96798 11842 96850
rect 12350 96798 12402 96850
rect 14366 96798 14418 96850
rect 15150 96798 15202 96850
rect 16494 96798 16546 96850
rect 17390 96798 17442 96850
rect 17726 96798 17778 96850
rect 18846 96798 18898 96850
rect 22094 96798 22146 96850
rect 28030 96798 28082 96850
rect 3166 96686 3218 96738
rect 4174 96686 4226 96738
rect 8094 96686 8146 96738
rect 10222 96686 10274 96738
rect 12014 96686 12066 96738
rect 13134 96686 13186 96738
rect 15038 96686 15090 96738
rect 16270 96686 16322 96738
rect 16830 96686 16882 96738
rect 17838 96686 17890 96738
rect 19070 96686 19122 96738
rect 19630 96686 19682 96738
rect 23886 96686 23938 96738
rect 25230 96686 25282 96738
rect 7870 96574 7922 96626
rect 20526 96574 20578 96626
rect 4616 96406 4668 96458
rect 4720 96406 4772 96458
rect 4824 96406 4876 96458
rect 11420 96406 11472 96458
rect 11524 96406 11576 96458
rect 11628 96406 11680 96458
rect 18224 96406 18276 96458
rect 18328 96406 18380 96458
rect 18432 96406 18484 96458
rect 25028 96406 25080 96458
rect 25132 96406 25184 96458
rect 25236 96406 25288 96458
rect 18286 96238 18338 96290
rect 18622 96238 18674 96290
rect 19518 96238 19570 96290
rect 21870 96238 21922 96290
rect 22094 96238 22146 96290
rect 22766 96238 22818 96290
rect 1710 96126 1762 96178
rect 3838 96126 3890 96178
rect 6638 96126 6690 96178
rect 12126 96126 12178 96178
rect 14702 96126 14754 96178
rect 16718 96126 16770 96178
rect 24334 96126 24386 96178
rect 4622 96014 4674 96066
rect 11230 96014 11282 96066
rect 12014 96014 12066 96066
rect 14030 96014 14082 96066
rect 14814 96014 14866 96066
rect 15934 96014 15986 96066
rect 16382 96014 16434 96066
rect 17502 96014 17554 96066
rect 18062 96014 18114 96066
rect 19854 96014 19906 96066
rect 22318 96014 22370 96066
rect 23662 96014 23714 96066
rect 25230 96014 25282 96066
rect 25902 96014 25954 96066
rect 6078 95902 6130 95954
rect 12126 95902 12178 95954
rect 15374 95902 15426 95954
rect 17614 95902 17666 95954
rect 18846 95902 18898 95954
rect 20078 95902 20130 95954
rect 20638 95902 20690 95954
rect 21646 95902 21698 95954
rect 23214 95902 23266 95954
rect 25342 95902 25394 95954
rect 5070 95790 5122 95842
rect 13694 95790 13746 95842
rect 15710 95790 15762 95842
rect 15822 95790 15874 95842
rect 17726 95790 17778 95842
rect 23326 95790 23378 95842
rect 25454 95790 25506 95842
rect 26238 95790 26290 95842
rect 8018 95622 8070 95674
rect 8122 95622 8174 95674
rect 8226 95622 8278 95674
rect 14822 95622 14874 95674
rect 14926 95622 14978 95674
rect 15030 95622 15082 95674
rect 21626 95622 21678 95674
rect 21730 95622 21782 95674
rect 21834 95622 21886 95674
rect 28430 95622 28482 95674
rect 28534 95622 28586 95674
rect 28638 95622 28690 95674
rect 2382 95454 2434 95506
rect 3278 95454 3330 95506
rect 6526 95454 6578 95506
rect 13246 95454 13298 95506
rect 15598 95454 15650 95506
rect 16830 95454 16882 95506
rect 18622 95454 18674 95506
rect 20526 95454 20578 95506
rect 24110 95454 24162 95506
rect 24446 95454 24498 95506
rect 2830 95342 2882 95394
rect 5966 95342 6018 95394
rect 6862 95342 6914 95394
rect 9662 95342 9714 95394
rect 10222 95342 10274 95394
rect 13918 95342 13970 95394
rect 15038 95342 15090 95394
rect 15934 95342 15986 95394
rect 16270 95342 16322 95394
rect 18174 95342 18226 95394
rect 18846 95342 18898 95394
rect 20078 95342 20130 95394
rect 24558 95342 24610 95394
rect 25454 95342 25506 95394
rect 5854 95230 5906 95282
rect 6078 95230 6130 95282
rect 7198 95230 7250 95282
rect 8542 95230 8594 95282
rect 9550 95230 9602 95282
rect 10334 95230 10386 95282
rect 10558 95230 10610 95282
rect 10782 95230 10834 95282
rect 11006 95230 11058 95282
rect 12014 95230 12066 95282
rect 12350 95230 12402 95282
rect 13582 95230 13634 95282
rect 14030 95230 14082 95282
rect 14478 95230 14530 95282
rect 14702 95230 14754 95282
rect 15374 95230 15426 95282
rect 15598 95230 15650 95282
rect 16382 95230 16434 95282
rect 17614 95230 17666 95282
rect 18398 95230 18450 95282
rect 19070 95230 19122 95282
rect 24222 95230 24274 95282
rect 25342 95230 25394 95282
rect 25678 95230 25730 95282
rect 26014 95230 26066 95282
rect 3726 95118 3778 95170
rect 4062 95118 4114 95170
rect 4510 95118 4562 95170
rect 4958 95118 5010 95170
rect 5406 95118 5458 95170
rect 6974 95118 7026 95170
rect 7646 95118 7698 95170
rect 8094 95118 8146 95170
rect 8990 95118 9042 95170
rect 13694 95118 13746 95170
rect 14590 95118 14642 95170
rect 17502 95118 17554 95170
rect 4398 95006 4450 95058
rect 4958 95006 5010 95058
rect 5406 95006 5458 95058
rect 9662 95006 9714 95058
rect 11790 95006 11842 95058
rect 19518 95006 19570 95058
rect 19854 95006 19906 95058
rect 4616 94838 4668 94890
rect 4720 94838 4772 94890
rect 4824 94838 4876 94890
rect 11420 94838 11472 94890
rect 11524 94838 11576 94890
rect 11628 94838 11680 94890
rect 18224 94838 18276 94890
rect 18328 94838 18380 94890
rect 18432 94838 18484 94890
rect 25028 94838 25080 94890
rect 25132 94838 25184 94890
rect 25236 94838 25288 94890
rect 6414 94670 6466 94722
rect 14142 94670 14194 94722
rect 3054 94558 3106 94610
rect 3390 94558 3442 94610
rect 4622 94558 4674 94610
rect 5070 94558 5122 94610
rect 5742 94558 5794 94610
rect 6638 94558 6690 94610
rect 9774 94558 9826 94610
rect 11230 94558 11282 94610
rect 12462 94558 12514 94610
rect 14366 94558 14418 94610
rect 16606 94558 16658 94610
rect 19630 94558 19682 94610
rect 25790 94558 25842 94610
rect 3726 94446 3778 94498
rect 3950 94446 4002 94498
rect 10446 94446 10498 94498
rect 11118 94446 11170 94498
rect 11342 94446 11394 94498
rect 11678 94446 11730 94498
rect 12798 94446 12850 94498
rect 13694 94446 13746 94498
rect 15598 94446 15650 94498
rect 16158 94446 16210 94498
rect 16382 94446 16434 94498
rect 16942 94446 16994 94498
rect 18734 94446 18786 94498
rect 19070 94446 19122 94498
rect 21198 94446 21250 94498
rect 21646 94446 21698 94498
rect 25006 94446 25058 94498
rect 13918 94334 13970 94386
rect 14590 94334 14642 94386
rect 14926 94334 14978 94386
rect 15038 94334 15090 94386
rect 16718 94334 16770 94386
rect 17390 94334 17442 94386
rect 17614 94334 17666 94386
rect 18062 94334 18114 94386
rect 18174 94334 18226 94386
rect 18286 94334 18338 94386
rect 19182 94334 19234 94386
rect 21870 94334 21922 94386
rect 2494 94222 2546 94274
rect 3390 94222 3442 94274
rect 3502 94222 3554 94274
rect 6078 94222 6130 94274
rect 7086 94222 7138 94274
rect 7534 94222 7586 94274
rect 14030 94222 14082 94274
rect 15262 94222 15314 94274
rect 15710 94222 15762 94274
rect 17166 94222 17218 94274
rect 17950 94222 18002 94274
rect 21422 94222 21474 94274
rect 22430 94222 22482 94274
rect 28030 94222 28082 94274
rect 8018 94054 8070 94106
rect 8122 94054 8174 94106
rect 8226 94054 8278 94106
rect 14822 94054 14874 94106
rect 14926 94054 14978 94106
rect 15030 94054 15082 94106
rect 21626 94054 21678 94106
rect 21730 94054 21782 94106
rect 21834 94054 21886 94106
rect 28430 94054 28482 94106
rect 28534 94054 28586 94106
rect 28638 94054 28690 94106
rect 4062 93886 4114 93938
rect 8654 93886 8706 93938
rect 11118 93886 11170 93938
rect 12350 93886 12402 93938
rect 12798 93886 12850 93938
rect 13918 93886 13970 93938
rect 14366 93886 14418 93938
rect 15262 93886 15314 93938
rect 16270 93886 16322 93938
rect 16382 93886 16434 93938
rect 20974 93886 21026 93938
rect 22318 93886 22370 93938
rect 26910 93886 26962 93938
rect 2494 93774 2546 93826
rect 2942 93774 2994 93826
rect 3166 93774 3218 93826
rect 9886 93774 9938 93826
rect 10334 93774 10386 93826
rect 10782 93774 10834 93826
rect 15150 93774 15202 93826
rect 15486 93774 15538 93826
rect 19070 93774 19122 93826
rect 4846 93662 4898 93714
rect 8430 93662 8482 93714
rect 8654 93662 8706 93714
rect 8990 93662 9042 93714
rect 9550 93662 9602 93714
rect 12126 93662 12178 93714
rect 12462 93662 12514 93714
rect 13134 93662 13186 93714
rect 14254 93662 14306 93714
rect 14590 93662 14642 93714
rect 14814 93662 14866 93714
rect 15710 93662 15762 93714
rect 16046 93662 16098 93714
rect 16158 93662 16210 93714
rect 17614 93662 17666 93714
rect 18510 93662 18562 93714
rect 20302 93662 20354 93714
rect 20526 93662 20578 93714
rect 22542 93662 22594 93714
rect 27134 93662 27186 93714
rect 3054 93550 3106 93602
rect 4510 93550 4562 93602
rect 5518 93550 5570 93602
rect 7646 93550 7698 93602
rect 13358 93550 13410 93602
rect 19182 93550 19234 93602
rect 23102 93550 23154 93602
rect 27806 93550 27858 93602
rect 4616 93270 4668 93322
rect 4720 93270 4772 93322
rect 4824 93270 4876 93322
rect 11420 93270 11472 93322
rect 11524 93270 11576 93322
rect 11628 93270 11680 93322
rect 18224 93270 18276 93322
rect 18328 93270 18380 93322
rect 18432 93270 18484 93322
rect 25028 93270 25080 93322
rect 25132 93270 25184 93322
rect 25236 93270 25288 93322
rect 11566 93102 11618 93154
rect 14926 93102 14978 93154
rect 22318 93102 22370 93154
rect 1710 92990 1762 93042
rect 3838 92990 3890 93042
rect 5182 92990 5234 93042
rect 6190 92990 6242 93042
rect 9214 92990 9266 93042
rect 11342 92990 11394 93042
rect 15598 92990 15650 93042
rect 17502 92990 17554 93042
rect 19966 92990 20018 93042
rect 21646 92990 21698 93042
rect 22878 92990 22930 93042
rect 25790 92990 25842 93042
rect 4622 92878 4674 92930
rect 6078 92878 6130 92930
rect 6302 92878 6354 92930
rect 6974 92878 7026 92930
rect 7758 92878 7810 92930
rect 8430 92878 8482 92930
rect 12238 92878 12290 92930
rect 13694 92878 13746 92930
rect 14590 92878 14642 92930
rect 16494 92878 16546 92930
rect 17614 92878 17666 92930
rect 19742 92878 19794 92930
rect 21422 92878 21474 92930
rect 21758 92878 21810 92930
rect 21982 92878 22034 92930
rect 22654 92878 22706 92930
rect 23662 92878 23714 92930
rect 26238 92878 26290 92930
rect 26350 92878 26402 92930
rect 26574 92878 26626 92930
rect 11678 92766 11730 92818
rect 13918 92766 13970 92818
rect 14030 92766 14082 92818
rect 14366 92766 14418 92818
rect 15934 92766 15986 92818
rect 16606 92766 16658 92818
rect 16942 92766 16994 92818
rect 19966 92766 20018 92818
rect 20414 92766 20466 92818
rect 23326 92766 23378 92818
rect 23998 92766 24050 92818
rect 24110 92766 24162 92818
rect 25454 92766 25506 92818
rect 27134 92766 27186 92818
rect 5854 92654 5906 92706
rect 7534 92654 7586 92706
rect 8094 92654 8146 92706
rect 11902 92654 11954 92706
rect 12686 92654 12738 92706
rect 19406 92654 19458 92706
rect 20190 92654 20242 92706
rect 21534 92654 21586 92706
rect 23438 92654 23490 92706
rect 23774 92654 23826 92706
rect 25678 92654 25730 92706
rect 26238 92654 26290 92706
rect 27022 92654 27074 92706
rect 8018 92486 8070 92538
rect 8122 92486 8174 92538
rect 8226 92486 8278 92538
rect 14822 92486 14874 92538
rect 14926 92486 14978 92538
rect 15030 92486 15082 92538
rect 21626 92486 21678 92538
rect 21730 92486 21782 92538
rect 21834 92486 21886 92538
rect 28430 92486 28482 92538
rect 28534 92486 28586 92538
rect 28638 92486 28690 92538
rect 10222 92318 10274 92370
rect 10334 92318 10386 92370
rect 10558 92318 10610 92370
rect 16830 92318 16882 92370
rect 17726 92318 17778 92370
rect 18510 92318 18562 92370
rect 20414 92318 20466 92370
rect 21310 92318 21362 92370
rect 22430 92318 22482 92370
rect 23998 92318 24050 92370
rect 2494 92206 2546 92258
rect 3278 92206 3330 92258
rect 6750 92206 6802 92258
rect 9774 92206 9826 92258
rect 20302 92206 20354 92258
rect 20638 92206 20690 92258
rect 22318 92206 22370 92258
rect 23102 92206 23154 92258
rect 23550 92206 23602 92258
rect 24110 92206 24162 92258
rect 25230 92206 25282 92258
rect 25454 92206 25506 92258
rect 26798 92206 26850 92258
rect 3054 92094 3106 92146
rect 3390 92094 3442 92146
rect 5070 92094 5122 92146
rect 10110 92094 10162 92146
rect 11006 92094 11058 92146
rect 17502 92094 17554 92146
rect 17838 92094 17890 92146
rect 17950 92094 18002 92146
rect 20750 92094 20802 92146
rect 21982 92094 22034 92146
rect 22542 92094 22594 92146
rect 22878 92094 22930 92146
rect 23326 92094 23378 92146
rect 23886 92094 23938 92146
rect 24334 92094 24386 92146
rect 24670 92094 24722 92146
rect 25790 92094 25842 92146
rect 26238 92094 26290 92146
rect 26462 92094 26514 92146
rect 27358 92094 27410 92146
rect 27582 92094 27634 92146
rect 28030 92094 28082 92146
rect 2830 91982 2882 92034
rect 13470 91982 13522 92034
rect 18958 91982 19010 92034
rect 25678 91982 25730 92034
rect 26686 91982 26738 92034
rect 27470 91982 27522 92034
rect 23438 91870 23490 91922
rect 27022 91870 27074 91922
rect 4616 91702 4668 91754
rect 4720 91702 4772 91754
rect 4824 91702 4876 91754
rect 11420 91702 11472 91754
rect 11524 91702 11576 91754
rect 11628 91702 11680 91754
rect 18224 91702 18276 91754
rect 18328 91702 18380 91754
rect 18432 91702 18484 91754
rect 25028 91702 25080 91754
rect 25132 91702 25184 91754
rect 25236 91702 25288 91754
rect 5742 91534 5794 91586
rect 22878 91534 22930 91586
rect 26126 91534 26178 91586
rect 26350 91534 26402 91586
rect 26462 91534 26514 91586
rect 27246 91534 27298 91586
rect 2494 91422 2546 91474
rect 4622 91422 4674 91474
rect 6078 91422 6130 91474
rect 10782 91422 10834 91474
rect 12686 91422 12738 91474
rect 14590 91422 14642 91474
rect 17278 91422 17330 91474
rect 18062 91422 18114 91474
rect 18958 91422 19010 91474
rect 22990 91422 23042 91474
rect 28142 91422 28194 91474
rect 1822 91310 1874 91362
rect 6526 91310 6578 91362
rect 7310 91310 7362 91362
rect 7982 91310 8034 91362
rect 12798 91310 12850 91362
rect 15486 91310 15538 91362
rect 16046 91310 16098 91362
rect 18510 91310 18562 91362
rect 18846 91310 18898 91362
rect 19182 91310 19234 91362
rect 19406 91310 19458 91362
rect 22206 91310 22258 91362
rect 22318 91310 22370 91362
rect 23550 91310 23602 91362
rect 25566 91310 25618 91362
rect 26910 91310 26962 91362
rect 8654 91198 8706 91250
rect 12910 91198 12962 91250
rect 13582 91198 13634 91250
rect 13694 91198 13746 91250
rect 14254 91198 14306 91250
rect 16382 91198 16434 91250
rect 16830 91198 16882 91250
rect 18062 91198 18114 91250
rect 22094 91198 22146 91250
rect 22542 91198 22594 91250
rect 23774 91198 23826 91250
rect 23998 91198 24050 91250
rect 24222 91198 24274 91250
rect 24334 91198 24386 91250
rect 25118 91198 25170 91250
rect 25678 91198 25730 91250
rect 26014 91198 26066 91250
rect 5070 91086 5122 91138
rect 6974 91086 7026 91138
rect 7198 91086 7250 91138
rect 11454 91086 11506 91138
rect 12014 91086 12066 91138
rect 13358 91086 13410 91138
rect 17950 91086 18002 91138
rect 18286 91086 18338 91138
rect 23214 91086 23266 91138
rect 23326 91086 23378 91138
rect 25230 91086 25282 91138
rect 27134 91086 27186 91138
rect 8018 90918 8070 90970
rect 8122 90918 8174 90970
rect 8226 90918 8278 90970
rect 14822 90918 14874 90970
rect 14926 90918 14978 90970
rect 15030 90918 15082 90970
rect 21626 90918 21678 90970
rect 21730 90918 21782 90970
rect 21834 90918 21886 90970
rect 28430 90918 28482 90970
rect 28534 90918 28586 90970
rect 28638 90918 28690 90970
rect 4734 90750 4786 90802
rect 8654 90750 8706 90802
rect 11454 90750 11506 90802
rect 15710 90750 15762 90802
rect 19406 90750 19458 90802
rect 19966 90750 20018 90802
rect 22766 90750 22818 90802
rect 4510 90638 4562 90690
rect 5294 90638 5346 90690
rect 5742 90638 5794 90690
rect 7534 90638 7586 90690
rect 8430 90638 8482 90690
rect 8766 90638 8818 90690
rect 9662 90638 9714 90690
rect 10558 90638 10610 90690
rect 10894 90638 10946 90690
rect 11902 90638 11954 90690
rect 14030 90638 14082 90690
rect 14702 90638 14754 90690
rect 14926 90638 14978 90690
rect 20078 90638 20130 90690
rect 21870 90638 21922 90690
rect 22878 90638 22930 90690
rect 23438 90638 23490 90690
rect 23550 90638 23602 90690
rect 6414 90526 6466 90578
rect 6974 90526 7026 90578
rect 7086 90526 7138 90578
rect 7422 90526 7474 90578
rect 7758 90526 7810 90578
rect 8990 90526 9042 90578
rect 9774 90526 9826 90578
rect 9886 90526 9938 90578
rect 10334 90526 10386 90578
rect 11118 90526 11170 90578
rect 11678 90526 11730 90578
rect 12686 90526 12738 90578
rect 13470 90526 13522 90578
rect 15150 90526 15202 90578
rect 15374 90526 15426 90578
rect 15598 90526 15650 90578
rect 19742 90526 19794 90578
rect 20190 90526 20242 90578
rect 20414 90526 20466 90578
rect 20638 90526 20690 90578
rect 21086 90526 21138 90578
rect 21310 90526 21362 90578
rect 21646 90526 21698 90578
rect 21982 90526 22034 90578
rect 22542 90526 22594 90578
rect 27022 90526 27074 90578
rect 27582 90526 27634 90578
rect 8094 90414 8146 90466
rect 10670 90414 10722 90466
rect 11566 90414 11618 90466
rect 12350 90414 12402 90466
rect 12910 90414 12962 90466
rect 13358 90414 13410 90466
rect 16270 90414 16322 90466
rect 16606 90414 16658 90466
rect 17614 90414 17666 90466
rect 17950 90414 18002 90466
rect 18398 90414 18450 90466
rect 20862 90414 20914 90466
rect 28030 90414 28082 90466
rect 17950 90302 18002 90354
rect 18398 90302 18450 90354
rect 23438 90302 23490 90354
rect 27134 90302 27186 90354
rect 4616 90134 4668 90186
rect 4720 90134 4772 90186
rect 4824 90134 4876 90186
rect 11420 90134 11472 90186
rect 11524 90134 11576 90186
rect 11628 90134 11680 90186
rect 18224 90134 18276 90186
rect 18328 90134 18380 90186
rect 18432 90134 18484 90186
rect 25028 90134 25080 90186
rect 25132 90134 25184 90186
rect 25236 90134 25288 90186
rect 18846 89966 18898 90018
rect 23214 89966 23266 90018
rect 4846 89854 4898 89906
rect 5854 89854 5906 89906
rect 7982 89854 8034 89906
rect 9550 89854 9602 89906
rect 9998 89854 10050 89906
rect 12462 89854 12514 89906
rect 13918 89854 13970 89906
rect 15038 89854 15090 89906
rect 15486 89854 15538 89906
rect 8654 89742 8706 89794
rect 10782 89742 10834 89794
rect 13582 89742 13634 89794
rect 13806 89742 13858 89794
rect 14590 89742 14642 89794
rect 15262 89742 15314 89794
rect 15710 89742 15762 89794
rect 16606 89742 16658 89794
rect 17726 89742 17778 89794
rect 19630 89742 19682 89794
rect 20190 89742 20242 89794
rect 21758 89742 21810 89794
rect 22542 89742 22594 89794
rect 22878 89742 22930 89794
rect 24222 89742 24274 89794
rect 24558 89742 24610 89794
rect 26126 89742 26178 89794
rect 27022 89742 27074 89794
rect 14030 89630 14082 89682
rect 14814 89630 14866 89682
rect 15822 89630 15874 89682
rect 16270 89630 16322 89682
rect 19966 89630 20018 89682
rect 21870 89630 21922 89682
rect 22766 89630 22818 89682
rect 23326 89630 23378 89682
rect 23998 89630 24050 89682
rect 24894 89630 24946 89682
rect 27246 89630 27298 89682
rect 18062 89518 18114 89570
rect 19294 89518 19346 89570
rect 19742 89518 19794 89570
rect 21982 89518 22034 89570
rect 22206 89518 22258 89570
rect 24110 89518 24162 89570
rect 26014 89518 26066 89570
rect 8018 89350 8070 89402
rect 8122 89350 8174 89402
rect 8226 89350 8278 89402
rect 14822 89350 14874 89402
rect 14926 89350 14978 89402
rect 15030 89350 15082 89402
rect 21626 89350 21678 89402
rect 21730 89350 21782 89402
rect 21834 89350 21886 89402
rect 28430 89350 28482 89402
rect 28534 89350 28586 89402
rect 28638 89350 28690 89402
rect 18622 89182 18674 89234
rect 18846 89182 18898 89234
rect 21646 89182 21698 89234
rect 22430 89182 22482 89234
rect 15710 89070 15762 89122
rect 15822 89070 15874 89122
rect 23326 89070 23378 89122
rect 25566 89070 25618 89122
rect 27134 89070 27186 89122
rect 4622 88958 4674 89010
rect 5070 88958 5122 89010
rect 6862 88958 6914 89010
rect 7198 88958 7250 89010
rect 7758 88958 7810 89010
rect 15934 89014 15986 89066
rect 8654 88958 8706 89010
rect 10110 88958 10162 89010
rect 16382 88958 16434 89010
rect 16830 88958 16882 89010
rect 17502 88958 17554 89010
rect 17950 88958 18002 89010
rect 18174 88958 18226 89010
rect 18734 88958 18786 89010
rect 18958 88958 19010 89010
rect 19182 88958 19234 89010
rect 21422 88958 21474 89010
rect 22094 88958 22146 89010
rect 23550 88958 23602 89010
rect 25118 88958 25170 89010
rect 25342 88958 25394 89010
rect 25790 88958 25842 89010
rect 26350 88958 26402 89010
rect 28142 88958 28194 89010
rect 1710 88846 1762 88898
rect 3838 88846 3890 88898
rect 8094 88846 8146 88898
rect 9102 88846 9154 88898
rect 13358 88846 13410 88898
rect 17726 88846 17778 88898
rect 19630 88846 19682 88898
rect 21534 88846 21586 88898
rect 24558 88846 24610 88898
rect 26238 88846 26290 88898
rect 27134 88846 27186 88898
rect 7086 88734 7138 88786
rect 8206 88734 8258 88786
rect 19406 88734 19458 88786
rect 19742 88734 19794 88786
rect 22766 88734 22818 88786
rect 23998 88734 24050 88786
rect 24334 88734 24386 88786
rect 4616 88566 4668 88618
rect 4720 88566 4772 88618
rect 4824 88566 4876 88618
rect 11420 88566 11472 88618
rect 11524 88566 11576 88618
rect 11628 88566 11680 88618
rect 18224 88566 18276 88618
rect 18328 88566 18380 88618
rect 18432 88566 18484 88618
rect 25028 88566 25080 88618
rect 25132 88566 25184 88618
rect 25236 88566 25288 88618
rect 5630 88398 5682 88450
rect 6638 88398 6690 88450
rect 6862 88398 6914 88450
rect 7758 88398 7810 88450
rect 22654 88398 22706 88450
rect 22990 88398 23042 88450
rect 24782 88398 24834 88450
rect 5742 88286 5794 88338
rect 6190 88286 6242 88338
rect 6638 88286 6690 88338
rect 7198 88286 7250 88338
rect 8094 88286 8146 88338
rect 10782 88286 10834 88338
rect 12910 88286 12962 88338
rect 16830 88286 16882 88338
rect 19742 88286 19794 88338
rect 20078 88286 20130 88338
rect 20526 88286 20578 88338
rect 23214 88286 23266 88338
rect 8206 88174 8258 88226
rect 8542 88174 8594 88226
rect 9102 88174 9154 88226
rect 9550 88174 9602 88226
rect 10110 88174 10162 88226
rect 13470 88174 13522 88226
rect 18286 88174 18338 88226
rect 19294 88174 19346 88226
rect 20750 88174 20802 88226
rect 24558 88174 24610 88226
rect 25006 88174 25058 88226
rect 26462 88174 26514 88226
rect 26798 88174 26850 88226
rect 1710 88062 1762 88114
rect 2494 88062 2546 88114
rect 2830 88062 2882 88114
rect 7758 88062 7810 88114
rect 7982 88062 8034 88114
rect 9214 88062 9266 88114
rect 17726 88062 17778 88114
rect 18062 88062 18114 88114
rect 18510 88062 18562 88114
rect 18622 88062 18674 88114
rect 19182 88062 19234 88114
rect 19854 88062 19906 88114
rect 20414 88062 20466 88114
rect 2046 87950 2098 88002
rect 3390 87950 3442 88002
rect 8990 87950 9042 88002
rect 8018 87782 8070 87834
rect 8122 87782 8174 87834
rect 8226 87782 8278 87834
rect 14822 87782 14874 87834
rect 14926 87782 14978 87834
rect 15030 87782 15082 87834
rect 21626 87782 21678 87834
rect 21730 87782 21782 87834
rect 21834 87782 21886 87834
rect 28430 87782 28482 87834
rect 28534 87782 28586 87834
rect 28638 87782 28690 87834
rect 1822 87614 1874 87666
rect 15150 87614 15202 87666
rect 16606 87614 16658 87666
rect 17502 87614 17554 87666
rect 18846 87614 18898 87666
rect 19966 87614 20018 87666
rect 26126 87614 26178 87666
rect 27582 87614 27634 87666
rect 4734 87502 4786 87554
rect 6862 87502 6914 87554
rect 13806 87502 13858 87554
rect 15262 87502 15314 87554
rect 15822 87502 15874 87554
rect 24670 87502 24722 87554
rect 5406 87390 5458 87442
rect 5630 87390 5682 87442
rect 6078 87390 6130 87442
rect 9550 87390 9602 87442
rect 14030 87390 14082 87442
rect 14478 87390 14530 87442
rect 14702 87390 14754 87442
rect 14926 87390 14978 87442
rect 18398 87390 18450 87442
rect 24110 87390 24162 87442
rect 25790 87390 25842 87442
rect 27134 87390 27186 87442
rect 27358 87390 27410 87442
rect 4510 87278 4562 87330
rect 8990 87278 9042 87330
rect 13246 87278 13298 87330
rect 13918 87278 13970 87330
rect 15934 87278 15986 87330
rect 16046 87278 16098 87330
rect 16718 87278 16770 87330
rect 17838 87278 17890 87330
rect 19518 87278 19570 87330
rect 20302 87278 20354 87330
rect 20862 87278 20914 87330
rect 21310 87278 21362 87330
rect 21758 87278 21810 87330
rect 24334 87278 24386 87330
rect 25566 87278 25618 87330
rect 27470 87278 27522 87330
rect 28142 87278 28194 87330
rect 16382 87166 16434 87218
rect 18062 87166 18114 87218
rect 20862 87166 20914 87218
rect 21758 87166 21810 87218
rect 26686 87166 26738 87218
rect 26910 87166 26962 87218
rect 4616 86998 4668 87050
rect 4720 86998 4772 87050
rect 4824 86998 4876 87050
rect 11420 86998 11472 87050
rect 11524 86998 11576 87050
rect 11628 86998 11680 87050
rect 18224 86998 18276 87050
rect 18328 86998 18380 87050
rect 18432 86998 18484 87050
rect 25028 86998 25080 87050
rect 25132 86998 25184 87050
rect 25236 86998 25288 87050
rect 4510 86830 4562 86882
rect 7086 86830 7138 86882
rect 7870 86830 7922 86882
rect 18958 86830 19010 86882
rect 19742 86830 19794 86882
rect 23998 86830 24050 86882
rect 4734 86718 4786 86770
rect 6078 86718 6130 86770
rect 6526 86718 6578 86770
rect 7086 86718 7138 86770
rect 7870 86718 7922 86770
rect 8430 86718 8482 86770
rect 16494 86718 16546 86770
rect 24110 86718 24162 86770
rect 7534 86606 7586 86658
rect 8990 86606 9042 86658
rect 10110 86606 10162 86658
rect 12238 86606 12290 86658
rect 12574 86606 12626 86658
rect 15038 86606 15090 86658
rect 15710 86606 15762 86658
rect 17278 86606 17330 86658
rect 19182 86606 19234 86658
rect 21310 86606 21362 86658
rect 21870 86606 21922 86658
rect 25006 86606 25058 86658
rect 26014 86606 26066 86658
rect 27246 86606 27298 86658
rect 27918 86606 27970 86658
rect 3838 86494 3890 86546
rect 8654 86494 8706 86546
rect 9214 86494 9266 86546
rect 10894 86494 10946 86546
rect 11230 86494 11282 86546
rect 16382 86494 16434 86546
rect 19518 86494 19570 86546
rect 20078 86494 20130 86546
rect 21982 86494 22034 86546
rect 22878 86494 22930 86546
rect 3502 86382 3554 86434
rect 4174 86382 4226 86434
rect 8766 86382 8818 86434
rect 9550 86382 9602 86434
rect 9662 86382 9714 86434
rect 9774 86382 9826 86434
rect 10782 86382 10834 86434
rect 11006 86382 11058 86434
rect 12014 86382 12066 86434
rect 12126 86382 12178 86434
rect 15038 86382 15090 86434
rect 18846 86382 18898 86434
rect 20190 86382 20242 86434
rect 20414 86382 20466 86434
rect 20750 86382 20802 86434
rect 21534 86382 21586 86434
rect 8018 86214 8070 86266
rect 8122 86214 8174 86266
rect 8226 86214 8278 86266
rect 14822 86214 14874 86266
rect 14926 86214 14978 86266
rect 15030 86214 15082 86266
rect 21626 86214 21678 86266
rect 21730 86214 21782 86266
rect 21834 86214 21886 86266
rect 28430 86214 28482 86266
rect 28534 86214 28586 86266
rect 28638 86214 28690 86266
rect 7310 86046 7362 86098
rect 15262 86046 15314 86098
rect 24446 86046 24498 86098
rect 25678 86046 25730 86098
rect 25790 86046 25842 86098
rect 2046 85934 2098 85986
rect 3726 85934 3778 85986
rect 8094 85934 8146 85986
rect 8654 85934 8706 85986
rect 10782 85934 10834 85986
rect 15934 85934 15986 85986
rect 16158 85934 16210 85986
rect 16382 85934 16434 85986
rect 22990 85934 23042 85986
rect 23886 85934 23938 85986
rect 26462 85934 26514 85986
rect 27806 85934 27858 85986
rect 1710 85822 1762 85874
rect 3054 85822 3106 85874
rect 7758 85822 7810 85874
rect 8318 85822 8370 85874
rect 13470 85822 13522 85874
rect 19406 85822 19458 85874
rect 25454 85822 25506 85874
rect 26350 85822 26402 85874
rect 27246 85822 27298 85874
rect 2494 85710 2546 85762
rect 5854 85710 5906 85762
rect 6974 85710 7026 85762
rect 8206 85710 8258 85762
rect 17838 85710 17890 85762
rect 24558 85710 24610 85762
rect 24670 85710 24722 85762
rect 7198 85598 7250 85650
rect 7870 85598 7922 85650
rect 16718 85598 16770 85650
rect 23998 85598 24050 85650
rect 27470 85598 27522 85650
rect 27694 85598 27746 85650
rect 4616 85430 4668 85482
rect 4720 85430 4772 85482
rect 4824 85430 4876 85482
rect 11420 85430 11472 85482
rect 11524 85430 11576 85482
rect 11628 85430 11680 85482
rect 18224 85430 18276 85482
rect 18328 85430 18380 85482
rect 18432 85430 18484 85482
rect 25028 85430 25080 85482
rect 25132 85430 25184 85482
rect 25236 85430 25288 85482
rect 17390 85262 17442 85314
rect 18174 85262 18226 85314
rect 19182 85262 19234 85314
rect 20638 85262 20690 85314
rect 22990 85262 23042 85314
rect 23326 85262 23378 85314
rect 24670 85262 24722 85314
rect 25118 85262 25170 85314
rect 25454 85262 25506 85314
rect 3950 85150 4002 85202
rect 7198 85150 7250 85202
rect 9326 85150 9378 85202
rect 14478 85150 14530 85202
rect 16606 85150 16658 85202
rect 17614 85150 17666 85202
rect 21982 85150 22034 85202
rect 23326 85150 23378 85202
rect 24222 85150 24274 85202
rect 26574 85150 26626 85202
rect 3054 85038 3106 85090
rect 6526 85038 6578 85090
rect 9662 85038 9714 85090
rect 12574 85038 12626 85090
rect 13806 85038 13858 85090
rect 17950 85038 18002 85090
rect 18622 85038 18674 85090
rect 22318 85038 22370 85090
rect 25678 85038 25730 85090
rect 26238 85038 26290 85090
rect 27022 85038 27074 85090
rect 11454 84926 11506 84978
rect 12798 84926 12850 84978
rect 12910 84926 12962 84978
rect 17166 84926 17218 84978
rect 17614 84926 17666 84978
rect 20750 84926 20802 84978
rect 21310 84926 21362 84978
rect 22766 84926 22818 84978
rect 24782 84926 24834 84978
rect 27134 84926 27186 84978
rect 27358 84926 27410 84978
rect 27470 84926 27522 84978
rect 27918 84926 27970 84978
rect 6078 84814 6130 84866
rect 20638 84814 20690 84866
rect 21422 84814 21474 84866
rect 23662 84814 23714 84866
rect 24670 84814 24722 84866
rect 27694 84814 27746 84866
rect 8018 84646 8070 84698
rect 8122 84646 8174 84698
rect 8226 84646 8278 84698
rect 14822 84646 14874 84698
rect 14926 84646 14978 84698
rect 15030 84646 15082 84698
rect 21626 84646 21678 84698
rect 21730 84646 21782 84698
rect 21834 84646 21886 84698
rect 28430 84646 28482 84698
rect 28534 84646 28586 84698
rect 28638 84646 28690 84698
rect 5742 84478 5794 84530
rect 8990 84478 9042 84530
rect 14030 84478 14082 84530
rect 19854 84478 19906 84530
rect 19966 84478 20018 84530
rect 10222 84366 10274 84418
rect 11790 84366 11842 84418
rect 15374 84366 15426 84418
rect 20078 84366 20130 84418
rect 20190 84366 20242 84418
rect 22878 84366 22930 84418
rect 26238 84366 26290 84418
rect 26574 84366 26626 84418
rect 10670 84254 10722 84306
rect 11118 84254 11170 84306
rect 14478 84254 14530 84306
rect 17614 84254 17666 84306
rect 19742 84254 19794 84306
rect 20862 84254 20914 84306
rect 21086 84254 21138 84306
rect 21758 84254 21810 84306
rect 22542 84254 22594 84306
rect 23774 84254 23826 84306
rect 24446 84254 24498 84306
rect 25566 84254 25618 84306
rect 26126 84254 26178 84306
rect 27134 84254 27186 84306
rect 27470 84254 27522 84306
rect 27582 84254 27634 84306
rect 2494 84142 2546 84194
rect 5406 84142 5458 84194
rect 9774 84142 9826 84194
rect 16830 84142 16882 84194
rect 18622 84142 18674 84194
rect 21422 84142 21474 84194
rect 22654 84142 22706 84194
rect 23550 84142 23602 84194
rect 26686 84142 26738 84194
rect 28030 84142 28082 84194
rect 26910 84030 26962 84082
rect 28030 84030 28082 84082
rect 28254 84030 28306 84082
rect 4616 83862 4668 83914
rect 4720 83862 4772 83914
rect 4824 83862 4876 83914
rect 11420 83862 11472 83914
rect 11524 83862 11576 83914
rect 11628 83862 11680 83914
rect 18224 83862 18276 83914
rect 18328 83862 18380 83914
rect 18432 83862 18484 83914
rect 25028 83862 25080 83914
rect 25132 83862 25184 83914
rect 25236 83862 25288 83914
rect 7422 83694 7474 83746
rect 7758 83694 7810 83746
rect 26350 83694 26402 83746
rect 27470 83694 27522 83746
rect 12350 83582 12402 83634
rect 15598 83582 15650 83634
rect 18398 83582 18450 83634
rect 18958 83582 19010 83634
rect 19518 83582 19570 83634
rect 20302 83582 20354 83634
rect 21534 83582 21586 83634
rect 22654 83582 22706 83634
rect 24334 83582 24386 83634
rect 5742 83470 5794 83522
rect 5966 83470 6018 83522
rect 9550 83470 9602 83522
rect 14478 83470 14530 83522
rect 14590 83470 14642 83522
rect 14926 83470 14978 83522
rect 18062 83470 18114 83522
rect 19294 83470 19346 83522
rect 20750 83470 20802 83522
rect 21982 83470 22034 83522
rect 22766 83470 22818 83522
rect 23662 83470 23714 83522
rect 24446 83470 24498 83522
rect 26014 83470 26066 83522
rect 1710 83358 1762 83410
rect 3278 83358 3330 83410
rect 6190 83358 6242 83410
rect 6414 83358 6466 83410
rect 6862 83358 6914 83410
rect 10222 83358 10274 83410
rect 12910 83358 12962 83410
rect 14814 83358 14866 83410
rect 17838 83358 17890 83410
rect 18846 83358 18898 83410
rect 21310 83358 21362 83410
rect 23438 83358 23490 83410
rect 24558 83358 24610 83410
rect 25790 83358 25842 83410
rect 27134 83358 27186 83410
rect 2046 83246 2098 83298
rect 2830 83246 2882 83298
rect 3838 83246 3890 83298
rect 4174 83246 4226 83298
rect 4622 83246 4674 83298
rect 5070 83246 5122 83298
rect 5630 83246 5682 83298
rect 6750 83246 6802 83298
rect 7310 83246 7362 83298
rect 7758 83246 7810 83298
rect 12574 83246 12626 83298
rect 12798 83246 12850 83298
rect 13918 83246 13970 83298
rect 15934 83246 15986 83298
rect 16382 83246 16434 83298
rect 17166 83246 17218 83298
rect 17614 83246 17666 83298
rect 21534 83246 21586 83298
rect 26798 83246 26850 83298
rect 27358 83246 27410 83298
rect 28030 83246 28082 83298
rect 8018 83078 8070 83130
rect 8122 83078 8174 83130
rect 8226 83078 8278 83130
rect 14822 83078 14874 83130
rect 14926 83078 14978 83130
rect 15030 83078 15082 83130
rect 21626 83078 21678 83130
rect 21730 83078 21782 83130
rect 21834 83078 21886 83130
rect 28430 83078 28482 83130
rect 28534 83078 28586 83130
rect 28638 83078 28690 83130
rect 7422 82910 7474 82962
rect 9886 82910 9938 82962
rect 10334 82910 10386 82962
rect 10782 82910 10834 82962
rect 11118 82910 11170 82962
rect 11230 82910 11282 82962
rect 11566 82910 11618 82962
rect 16606 82910 16658 82962
rect 17502 82910 17554 82962
rect 19966 82910 20018 82962
rect 23550 82910 23602 82962
rect 25454 82910 25506 82962
rect 4846 82798 4898 82850
rect 16382 82798 16434 82850
rect 21086 82798 21138 82850
rect 22094 82798 22146 82850
rect 24222 82798 24274 82850
rect 26238 82798 26290 82850
rect 27470 82798 27522 82850
rect 2270 82686 2322 82738
rect 2606 82686 2658 82738
rect 3054 82686 3106 82738
rect 3390 82686 3442 82738
rect 4062 82686 4114 82738
rect 11342 82686 11394 82738
rect 12350 82686 12402 82738
rect 15598 82686 15650 82738
rect 15822 82686 15874 82738
rect 16270 82686 16322 82738
rect 16718 82686 16770 82738
rect 20302 82686 20354 82738
rect 20526 82686 20578 82738
rect 22542 82686 22594 82738
rect 23438 82686 23490 82738
rect 25454 82686 25506 82738
rect 26126 82686 26178 82738
rect 27022 82686 27074 82738
rect 27246 82686 27298 82738
rect 2382 82574 2434 82626
rect 6974 82574 7026 82626
rect 7422 82574 7474 82626
rect 8094 82574 8146 82626
rect 13470 82574 13522 82626
rect 15710 82574 15762 82626
rect 18062 82574 18114 82626
rect 18510 82574 18562 82626
rect 18958 82574 19010 82626
rect 19406 82574 19458 82626
rect 19854 82574 19906 82626
rect 26350 82574 26402 82626
rect 27134 82574 27186 82626
rect 28030 82574 28082 82626
rect 2830 82462 2882 82514
rect 3390 82462 3442 82514
rect 3726 82462 3778 82514
rect 7646 82462 7698 82514
rect 18062 82462 18114 82514
rect 18958 82462 19010 82514
rect 4616 82294 4668 82346
rect 4720 82294 4772 82346
rect 4824 82294 4876 82346
rect 11420 82294 11472 82346
rect 11524 82294 11576 82346
rect 11628 82294 11680 82346
rect 18224 82294 18276 82346
rect 18328 82294 18380 82346
rect 18432 82294 18484 82346
rect 25028 82294 25080 82346
rect 25132 82294 25184 82346
rect 25236 82294 25288 82346
rect 5966 82126 6018 82178
rect 10222 82126 10274 82178
rect 11230 82126 11282 82178
rect 21982 82126 22034 82178
rect 25230 82126 25282 82178
rect 26014 82126 26066 82178
rect 27694 82126 27746 82178
rect 2494 82014 2546 82066
rect 4622 82014 4674 82066
rect 4958 82014 5010 82066
rect 9326 82014 9378 82066
rect 9662 82014 9714 82066
rect 10222 82014 10274 82066
rect 15598 82014 15650 82066
rect 17726 82014 17778 82066
rect 18398 82014 18450 82066
rect 26574 82014 26626 82066
rect 27246 82014 27298 82066
rect 24782 81958 24834 82010
rect 1822 81902 1874 81954
rect 5966 81902 6018 81954
rect 6526 81902 6578 81954
rect 14814 81902 14866 81954
rect 20190 81902 20242 81954
rect 21310 81902 21362 81954
rect 21534 81902 21586 81954
rect 23214 81902 23266 81954
rect 24446 81902 24498 81954
rect 25454 81902 25506 81954
rect 26238 81902 26290 81954
rect 27470 81902 27522 81954
rect 5630 81790 5682 81842
rect 7198 81790 7250 81842
rect 20526 81790 20578 81842
rect 24670 81790 24722 81842
rect 5070 81678 5122 81730
rect 9774 81678 9826 81730
rect 10670 81678 10722 81730
rect 11118 81678 11170 81730
rect 11566 81678 11618 81730
rect 12014 81678 12066 81730
rect 12462 81678 12514 81730
rect 13022 81678 13074 81730
rect 13582 81678 13634 81730
rect 14030 81678 14082 81730
rect 14478 81678 14530 81730
rect 18846 81678 18898 81730
rect 19294 81678 19346 81730
rect 19742 81678 19794 81730
rect 20638 81678 20690 81730
rect 20750 81678 20802 81730
rect 28142 81678 28194 81730
rect 8018 81510 8070 81562
rect 8122 81510 8174 81562
rect 8226 81510 8278 81562
rect 14822 81510 14874 81562
rect 14926 81510 14978 81562
rect 15030 81510 15082 81562
rect 21626 81510 21678 81562
rect 21730 81510 21782 81562
rect 21834 81510 21886 81562
rect 28430 81510 28482 81562
rect 28534 81510 28586 81562
rect 28638 81510 28690 81562
rect 7198 81342 7250 81394
rect 10222 81342 10274 81394
rect 11902 81342 11954 81394
rect 17502 81342 17554 81394
rect 17838 81342 17890 81394
rect 19294 81342 19346 81394
rect 22878 81342 22930 81394
rect 23438 81342 23490 81394
rect 23662 81342 23714 81394
rect 23774 81342 23826 81394
rect 24558 81342 24610 81394
rect 26126 81342 26178 81394
rect 16606 81230 16658 81282
rect 16830 81230 16882 81282
rect 18398 81230 18450 81282
rect 18510 81230 18562 81282
rect 19966 81230 20018 81282
rect 22654 81230 22706 81282
rect 23886 81230 23938 81282
rect 24446 81230 24498 81282
rect 26350 81230 26402 81282
rect 3054 81118 3106 81170
rect 6974 81118 7026 81170
rect 7310 81118 7362 81170
rect 7422 81118 7474 81170
rect 7758 81118 7810 81170
rect 10558 81118 10610 81170
rect 10782 81118 10834 81170
rect 12238 81118 12290 81170
rect 17726 81118 17778 81170
rect 17950 81118 18002 81170
rect 18174 81118 18226 81170
rect 19406 81118 19458 81170
rect 20750 81118 20802 81170
rect 21646 81118 21698 81170
rect 22542 81118 22594 81170
rect 22990 81118 23042 81170
rect 26910 81118 26962 81170
rect 27134 81118 27186 81170
rect 28142 81118 28194 81170
rect 4846 81006 4898 81058
rect 5742 81006 5794 81058
rect 6190 81006 6242 81058
rect 6638 81006 6690 81058
rect 14030 81006 14082 81058
rect 20526 81006 20578 81058
rect 25230 81006 25282 81058
rect 28030 81006 28082 81058
rect 11006 80894 11058 80946
rect 11118 80894 11170 80946
rect 16494 80894 16546 80946
rect 19294 80894 19346 80946
rect 24558 80894 24610 80946
rect 25454 80894 25506 80946
rect 25678 80894 25730 80946
rect 26462 80894 26514 80946
rect 4616 80726 4668 80778
rect 4720 80726 4772 80778
rect 4824 80726 4876 80778
rect 11420 80726 11472 80778
rect 11524 80726 11576 80778
rect 11628 80726 11680 80778
rect 18224 80726 18276 80778
rect 18328 80726 18380 80778
rect 18432 80726 18484 80778
rect 25028 80726 25080 80778
rect 25132 80726 25184 80778
rect 25236 80726 25288 80778
rect 20190 80558 20242 80610
rect 21646 80558 21698 80610
rect 24110 80558 24162 80610
rect 24558 80558 24610 80610
rect 26238 80558 26290 80610
rect 26574 80558 26626 80610
rect 27246 80558 27298 80610
rect 27582 80558 27634 80610
rect 2830 80446 2882 80498
rect 4062 80446 4114 80498
rect 7086 80446 7138 80498
rect 10110 80446 10162 80498
rect 12238 80446 12290 80498
rect 16494 80446 16546 80498
rect 17502 80446 17554 80498
rect 18286 80446 18338 80498
rect 23438 80446 23490 80498
rect 27022 80446 27074 80498
rect 28030 80446 28082 80498
rect 3054 80334 3106 80386
rect 6078 80334 6130 80386
rect 9438 80334 9490 80386
rect 13582 80334 13634 80386
rect 17390 80334 17442 80386
rect 17838 80334 17890 80386
rect 18062 80334 18114 80386
rect 18846 80334 18898 80386
rect 19294 80334 19346 80386
rect 19966 80334 20018 80386
rect 21310 80334 21362 80386
rect 22094 80334 22146 80386
rect 24446 80334 24498 80386
rect 25230 80334 25282 80386
rect 25566 80334 25618 80386
rect 25902 80334 25954 80386
rect 5742 80222 5794 80274
rect 14366 80222 14418 80274
rect 20526 80222 20578 80274
rect 22430 80222 22482 80274
rect 23102 80222 23154 80274
rect 23998 80222 24050 80274
rect 26462 80222 26514 80274
rect 1710 80110 1762 80162
rect 2046 80110 2098 80162
rect 5070 80110 5122 80162
rect 5854 80110 5906 80162
rect 6526 80110 6578 80162
rect 13022 80110 13074 80162
rect 21534 80110 21586 80162
rect 23326 80110 23378 80162
rect 25006 80110 25058 80162
rect 25566 80110 25618 80162
rect 8018 79942 8070 79994
rect 8122 79942 8174 79994
rect 8226 79942 8278 79994
rect 14822 79942 14874 79994
rect 14926 79942 14978 79994
rect 15030 79942 15082 79994
rect 21626 79942 21678 79994
rect 21730 79942 21782 79994
rect 21834 79942 21886 79994
rect 28430 79942 28482 79994
rect 28534 79942 28586 79994
rect 28638 79942 28690 79994
rect 2494 79774 2546 79826
rect 17726 79774 17778 79826
rect 24670 79774 24722 79826
rect 26238 79774 26290 79826
rect 26686 79774 26738 79826
rect 27134 79774 27186 79826
rect 28030 79774 28082 79826
rect 12686 79662 12738 79714
rect 14814 79662 14866 79714
rect 15822 79662 15874 79714
rect 17614 79662 17666 79714
rect 19518 79662 19570 79714
rect 3278 79550 3330 79602
rect 4510 79550 4562 79602
rect 7758 79550 7810 79602
rect 10110 79550 10162 79602
rect 10334 79550 10386 79602
rect 11678 79550 11730 79602
rect 14926 79550 14978 79602
rect 16382 79550 16434 79602
rect 17950 79550 18002 79602
rect 18174 79550 18226 79602
rect 19070 79550 19122 79602
rect 19742 79550 19794 79602
rect 21086 79550 21138 79602
rect 21534 79550 21586 79602
rect 21870 79550 21922 79602
rect 23774 79550 23826 79602
rect 24222 79550 24274 79602
rect 25790 79550 25842 79602
rect 4062 79438 4114 79490
rect 5294 79438 5346 79490
rect 7422 79438 7474 79490
rect 8318 79438 8370 79490
rect 9102 79438 9154 79490
rect 10558 79438 10610 79490
rect 13134 79438 13186 79490
rect 19182 79438 19234 79490
rect 19966 79438 20018 79490
rect 22654 79438 22706 79490
rect 23326 79438 23378 79490
rect 25454 79438 25506 79490
rect 27582 79438 27634 79490
rect 3614 79326 3666 79378
rect 7870 79326 7922 79378
rect 10670 79326 10722 79378
rect 27358 79326 27410 79378
rect 28030 79326 28082 79378
rect 4616 79158 4668 79210
rect 4720 79158 4772 79210
rect 4824 79158 4876 79210
rect 11420 79158 11472 79210
rect 11524 79158 11576 79210
rect 11628 79158 11680 79210
rect 18224 79158 18276 79210
rect 18328 79158 18380 79210
rect 18432 79158 18484 79210
rect 25028 79158 25080 79210
rect 25132 79158 25184 79210
rect 25236 79158 25288 79210
rect 5854 78990 5906 79042
rect 14254 78990 14306 79042
rect 18958 78990 19010 79042
rect 19742 78990 19794 79042
rect 25342 78990 25394 79042
rect 25566 78990 25618 79042
rect 4622 78878 4674 78930
rect 11230 78878 11282 78930
rect 12014 78878 12066 78930
rect 17726 78878 17778 78930
rect 19070 78878 19122 78930
rect 21422 78878 21474 78930
rect 24222 78878 24274 78930
rect 26462 78878 26514 78930
rect 26910 78878 26962 78930
rect 27358 78878 27410 78930
rect 28142 78878 28194 78930
rect 1822 78766 1874 78818
rect 5854 78766 5906 78818
rect 6190 78766 6242 78818
rect 8430 78766 8482 78818
rect 12126 78766 12178 78818
rect 12238 78766 12290 78818
rect 13694 78766 13746 78818
rect 13918 78766 13970 78818
rect 14254 78766 14306 78818
rect 14814 78766 14866 78818
rect 18062 78766 18114 78818
rect 19294 78766 19346 78818
rect 20190 78766 20242 78818
rect 23774 78766 23826 78818
rect 2494 78654 2546 78706
rect 6414 78654 6466 78706
rect 9102 78654 9154 78706
rect 15598 78654 15650 78706
rect 19630 78654 19682 78706
rect 19742 78654 19794 78706
rect 20526 78654 20578 78706
rect 21310 78654 21362 78706
rect 22542 78654 22594 78706
rect 23326 78654 23378 78706
rect 5070 78542 5122 78594
rect 5630 78542 5682 78594
rect 6862 78542 6914 78594
rect 7870 78542 7922 78594
rect 13022 78542 13074 78594
rect 14478 78542 14530 78594
rect 18622 78542 18674 78594
rect 21534 78542 21586 78594
rect 22094 78542 22146 78594
rect 22654 78542 22706 78594
rect 22766 78542 22818 78594
rect 24670 78542 24722 78594
rect 25118 78542 25170 78594
rect 25678 78542 25730 78594
rect 26126 78542 26178 78594
rect 8018 78374 8070 78426
rect 8122 78374 8174 78426
rect 8226 78374 8278 78426
rect 14822 78374 14874 78426
rect 14926 78374 14978 78426
rect 15030 78374 15082 78426
rect 21626 78374 21678 78426
rect 21730 78374 21782 78426
rect 21834 78374 21886 78426
rect 28430 78374 28482 78426
rect 28534 78374 28586 78426
rect 28638 78374 28690 78426
rect 2382 78206 2434 78258
rect 4846 78206 4898 78258
rect 5294 78206 5346 78258
rect 6414 78206 6466 78258
rect 8990 78206 9042 78258
rect 11006 78206 11058 78258
rect 17502 78206 17554 78258
rect 2046 78094 2098 78146
rect 3166 78094 3218 78146
rect 18846 78094 18898 78146
rect 20190 78094 20242 78146
rect 1710 77982 1762 78034
rect 2606 77982 2658 78034
rect 2942 77982 2994 78034
rect 3502 77982 3554 78034
rect 3726 77982 3778 78034
rect 3614 77870 3666 77922
rect 2718 77758 2770 77810
rect 7870 77982 7922 78034
rect 8206 77982 8258 78034
rect 8542 77982 8594 78034
rect 8766 77982 8818 78034
rect 9886 77982 9938 78034
rect 13022 77982 13074 78034
rect 17390 77982 17442 78034
rect 17614 77982 17666 78034
rect 17950 77982 18002 78034
rect 18510 77982 18562 78034
rect 19742 77982 19794 78034
rect 21870 77982 21922 78034
rect 25342 77982 25394 78034
rect 4062 77870 4114 77922
rect 6078 77870 6130 77922
rect 6974 77870 7026 77922
rect 7422 77870 7474 77922
rect 13582 77870 13634 77922
rect 19294 77870 19346 77922
rect 20638 77870 20690 77922
rect 21086 77870 21138 77922
rect 22542 77870 22594 77922
rect 24670 77870 24722 77922
rect 26014 77870 26066 77922
rect 28142 77870 28194 77922
rect 4062 77758 4114 77810
rect 7422 77758 7474 77810
rect 7982 77758 8034 77810
rect 8766 77758 8818 77810
rect 17838 77758 17890 77810
rect 18510 77758 18562 77810
rect 20638 77758 20690 77810
rect 21422 77758 21474 77810
rect 4616 77590 4668 77642
rect 4720 77590 4772 77642
rect 4824 77590 4876 77642
rect 11420 77590 11472 77642
rect 11524 77590 11576 77642
rect 11628 77590 11680 77642
rect 18224 77590 18276 77642
rect 18328 77590 18380 77642
rect 18432 77590 18484 77642
rect 25028 77590 25080 77642
rect 25132 77590 25184 77642
rect 25236 77590 25288 77642
rect 20414 77422 20466 77474
rect 22542 77422 22594 77474
rect 2718 77310 2770 77362
rect 8542 77310 8594 77362
rect 12910 77310 12962 77362
rect 21422 77310 21474 77362
rect 23214 77310 23266 77362
rect 25230 77310 25282 77362
rect 3502 77198 3554 77250
rect 5630 77198 5682 77250
rect 9662 77198 9714 77250
rect 10110 77198 10162 77250
rect 15038 77198 15090 77250
rect 21982 77198 22034 77250
rect 22542 77198 22594 77250
rect 24446 77198 24498 77250
rect 28030 77198 28082 77250
rect 2494 77086 2546 77138
rect 2718 77086 2770 77138
rect 6414 77086 6466 77138
rect 10782 77086 10834 77138
rect 13582 77086 13634 77138
rect 18398 77086 18450 77138
rect 22206 77086 22258 77138
rect 23662 77086 23714 77138
rect 24334 77086 24386 77138
rect 24670 77086 24722 77138
rect 24894 77086 24946 77138
rect 27358 77086 27410 77138
rect 2158 76974 2210 77026
rect 4062 76974 4114 77026
rect 4734 76974 4786 77026
rect 5070 76974 5122 77026
rect 9326 76974 9378 77026
rect 13694 76974 13746 77026
rect 19966 76974 20018 77026
rect 20526 76974 20578 77026
rect 20638 76974 20690 77026
rect 22430 76974 22482 77026
rect 23102 76974 23154 77026
rect 8018 76806 8070 76858
rect 8122 76806 8174 76858
rect 8226 76806 8278 76858
rect 14822 76806 14874 76858
rect 14926 76806 14978 76858
rect 15030 76806 15082 76858
rect 21626 76806 21678 76858
rect 21730 76806 21782 76858
rect 21834 76806 21886 76858
rect 28430 76806 28482 76858
rect 28534 76806 28586 76858
rect 28638 76806 28690 76858
rect 6638 76638 6690 76690
rect 11118 76638 11170 76690
rect 11230 76638 11282 76690
rect 11902 76638 11954 76690
rect 13134 76638 13186 76690
rect 17502 76638 17554 76690
rect 22206 76638 22258 76690
rect 22654 76638 22706 76690
rect 24446 76638 24498 76690
rect 25342 76638 25394 76690
rect 26238 76638 26290 76690
rect 26910 76638 26962 76690
rect 27022 76638 27074 76690
rect 28142 76638 28194 76690
rect 2830 76526 2882 76578
rect 10446 76526 10498 76578
rect 15262 76526 15314 76578
rect 18174 76526 18226 76578
rect 27358 76526 27410 76578
rect 3726 76414 3778 76466
rect 5294 76414 5346 76466
rect 6526 76414 6578 76466
rect 6862 76414 6914 76466
rect 7086 76414 7138 76466
rect 7982 76414 8034 76466
rect 9774 76414 9826 76466
rect 10110 76414 10162 76466
rect 10670 76414 10722 76466
rect 11790 76414 11842 76466
rect 12126 76414 12178 76466
rect 12350 76414 12402 76466
rect 14030 76414 14082 76466
rect 16494 76414 16546 76466
rect 18958 76414 19010 76466
rect 25902 76414 25954 76466
rect 26350 76414 26402 76466
rect 26462 76414 26514 76466
rect 27134 76414 27186 76466
rect 1822 76302 1874 76354
rect 2270 76302 2322 76354
rect 2718 76302 2770 76354
rect 4622 76302 4674 76354
rect 5742 76302 5794 76354
rect 6302 76302 6354 76354
rect 7758 76302 7810 76354
rect 8542 76302 8594 76354
rect 8990 76302 9042 76354
rect 10222 76302 10274 76354
rect 19630 76302 19682 76354
rect 21758 76302 21810 76354
rect 23214 76302 23266 76354
rect 23550 76302 23602 76354
rect 24110 76302 24162 76354
rect 2606 76190 2658 76242
rect 7086 76190 7138 76242
rect 7646 76190 7698 76242
rect 11006 76190 11058 76242
rect 18062 76190 18114 76242
rect 21982 76190 22034 76242
rect 22878 76190 22930 76242
rect 24446 76190 24498 76242
rect 4616 76022 4668 76074
rect 4720 76022 4772 76074
rect 4824 76022 4876 76074
rect 11420 76022 11472 76074
rect 11524 76022 11576 76074
rect 11628 76022 11680 76074
rect 18224 76022 18276 76074
rect 18328 76022 18380 76074
rect 18432 76022 18484 76074
rect 25028 76022 25080 76074
rect 25132 76022 25184 76074
rect 25236 76022 25288 76074
rect 18286 75854 18338 75906
rect 20190 75854 20242 75906
rect 21870 75854 21922 75906
rect 22094 75854 22146 75906
rect 4622 75742 4674 75794
rect 8542 75742 8594 75794
rect 9774 75742 9826 75794
rect 11902 75742 11954 75794
rect 12462 75742 12514 75794
rect 16382 75742 16434 75794
rect 16830 75742 16882 75794
rect 19182 75742 19234 75794
rect 19742 75742 19794 75794
rect 21422 75742 21474 75794
rect 21870 75742 21922 75794
rect 22318 75742 22370 75794
rect 25678 75742 25730 75794
rect 26462 75742 26514 75794
rect 27358 75742 27410 75794
rect 1710 75630 1762 75682
rect 4958 75630 5010 75682
rect 5070 75630 5122 75682
rect 5630 75630 5682 75682
rect 9102 75630 9154 75682
rect 12574 75630 12626 75682
rect 12910 75630 12962 75682
rect 13582 75630 13634 75682
rect 18286 75630 18338 75682
rect 19966 75630 20018 75682
rect 20190 75630 20242 75682
rect 22878 75630 22930 75682
rect 27022 75630 27074 75682
rect 2494 75518 2546 75570
rect 6414 75518 6466 75570
rect 14254 75518 14306 75570
rect 17726 75518 17778 75570
rect 17950 75518 18002 75570
rect 19630 75518 19682 75570
rect 23550 75518 23602 75570
rect 12350 75406 12402 75458
rect 17278 75406 17330 75458
rect 18174 75406 18226 75458
rect 21310 75406 21362 75458
rect 26350 75406 26402 75458
rect 26574 75406 26626 75458
rect 27806 75406 27858 75458
rect 8018 75238 8070 75290
rect 8122 75238 8174 75290
rect 8226 75238 8278 75290
rect 14822 75238 14874 75290
rect 14926 75238 14978 75290
rect 15030 75238 15082 75290
rect 21626 75238 21678 75290
rect 21730 75238 21782 75290
rect 21834 75238 21886 75290
rect 28430 75238 28482 75290
rect 28534 75238 28586 75290
rect 28638 75238 28690 75290
rect 2382 75070 2434 75122
rect 4846 75070 4898 75122
rect 6414 75070 6466 75122
rect 6974 75070 7026 75122
rect 7534 75070 7586 75122
rect 7982 75070 8034 75122
rect 8542 75070 8594 75122
rect 8766 75070 8818 75122
rect 9774 75070 9826 75122
rect 9998 75070 10050 75122
rect 11006 75070 11058 75122
rect 11230 75070 11282 75122
rect 11342 75070 11394 75122
rect 12350 75070 12402 75122
rect 14254 75070 14306 75122
rect 15150 75070 15202 75122
rect 15934 75070 15986 75122
rect 20750 75070 20802 75122
rect 23774 75070 23826 75122
rect 24670 75070 24722 75122
rect 26686 75070 26738 75122
rect 28142 75070 28194 75122
rect 2046 74958 2098 75010
rect 2942 74958 2994 75010
rect 3166 74958 3218 75010
rect 5630 74958 5682 75010
rect 10222 74958 10274 75010
rect 13582 74958 13634 75010
rect 18174 74958 18226 75010
rect 1710 74846 1762 74898
rect 2494 74846 2546 74898
rect 2718 74846 2770 74898
rect 3614 74846 3666 74898
rect 5966 74846 6018 74898
rect 6078 74846 6130 74898
rect 6190 74846 6242 74898
rect 6862 74846 6914 74898
rect 8430 74846 8482 74898
rect 8990 74846 9042 74898
rect 9550 74846 9602 74898
rect 11454 74846 11506 74898
rect 11790 74846 11842 74898
rect 13246 74846 13298 74898
rect 14030 74846 14082 74898
rect 14254 74846 14306 74898
rect 14590 74846 14642 74898
rect 14926 74846 14978 74898
rect 15038 74846 15090 74898
rect 15598 74846 15650 74898
rect 16382 74846 16434 74898
rect 16830 74846 16882 74898
rect 17502 74846 17554 74898
rect 21982 74846 22034 74898
rect 4174 74734 4226 74786
rect 5294 74734 5346 74786
rect 10334 74734 10386 74786
rect 12798 74734 12850 74786
rect 20302 74734 20354 74786
rect 21310 74734 21362 74786
rect 22542 74734 22594 74786
rect 22990 74734 23042 74786
rect 23326 74734 23378 74786
rect 24222 74734 24274 74786
rect 25790 74734 25842 74786
rect 26126 74734 26178 74786
rect 27134 74734 27186 74786
rect 27582 74734 27634 74786
rect 6750 74622 6802 74674
rect 8878 74622 8930 74674
rect 12574 74622 12626 74674
rect 13358 74622 13410 74674
rect 13694 74622 13746 74674
rect 15710 74622 15762 74674
rect 16270 74622 16322 74674
rect 22206 74622 22258 74674
rect 23326 74622 23378 74674
rect 25902 74622 25954 74674
rect 26686 74622 26738 74674
rect 27134 74622 27186 74674
rect 27582 74622 27634 74674
rect 4616 74454 4668 74506
rect 4720 74454 4772 74506
rect 4824 74454 4876 74506
rect 11420 74454 11472 74506
rect 11524 74454 11576 74506
rect 11628 74454 11680 74506
rect 18224 74454 18276 74506
rect 18328 74454 18380 74506
rect 18432 74454 18484 74506
rect 25028 74454 25080 74506
rect 25132 74454 25184 74506
rect 25236 74454 25288 74506
rect 9102 74286 9154 74338
rect 10110 74286 10162 74338
rect 12574 74286 12626 74338
rect 18622 74286 18674 74338
rect 19294 74286 19346 74338
rect 20302 74286 20354 74338
rect 2270 74174 2322 74226
rect 5742 74174 5794 74226
rect 8654 74174 8706 74226
rect 9102 74174 9154 74226
rect 9998 74174 10050 74226
rect 10446 74174 10498 74226
rect 12126 74174 12178 74226
rect 12462 74174 12514 74226
rect 14030 74174 14082 74226
rect 17278 74174 17330 74226
rect 18734 74174 18786 74226
rect 24222 74174 24274 74226
rect 3614 74062 3666 74114
rect 15598 74062 15650 74114
rect 18958 74062 19010 74114
rect 19854 74062 19906 74114
rect 20302 74062 20354 74114
rect 21422 74062 21474 74114
rect 24782 74062 24834 74114
rect 25902 74062 25954 74114
rect 26238 74062 26290 74114
rect 26574 74062 26626 74114
rect 27022 74062 27074 74114
rect 27918 74062 27970 74114
rect 7198 73950 7250 74002
rect 10894 73950 10946 74002
rect 11678 73950 11730 74002
rect 14926 73950 14978 74002
rect 16046 73950 16098 74002
rect 19518 73950 19570 74002
rect 20750 73950 20802 74002
rect 22094 73950 22146 74002
rect 25006 73950 25058 74002
rect 25678 73950 25730 74002
rect 27134 73950 27186 74002
rect 27358 73950 27410 74002
rect 1822 73838 1874 73890
rect 2942 73838 2994 73890
rect 4062 73838 4114 73890
rect 4846 73838 4898 73890
rect 6750 73838 6802 73890
rect 9550 73838 9602 73890
rect 13582 73838 13634 73890
rect 14590 73838 14642 73890
rect 14814 73838 14866 73890
rect 15598 73838 15650 73890
rect 24558 73838 24610 73890
rect 24670 73838 24722 73890
rect 25566 73838 25618 73890
rect 26126 73838 26178 73890
rect 26910 73838 26962 73890
rect 8018 73670 8070 73722
rect 8122 73670 8174 73722
rect 8226 73670 8278 73722
rect 14822 73670 14874 73722
rect 14926 73670 14978 73722
rect 15030 73670 15082 73722
rect 21626 73670 21678 73722
rect 21730 73670 21782 73722
rect 21834 73670 21886 73722
rect 28430 73670 28482 73722
rect 28534 73670 28586 73722
rect 28638 73670 28690 73722
rect 8990 73502 9042 73554
rect 9662 73502 9714 73554
rect 10110 73502 10162 73554
rect 20302 73502 20354 73554
rect 21870 73502 21922 73554
rect 23550 73502 23602 73554
rect 2046 73390 2098 73442
rect 14030 73390 14082 73442
rect 18062 73390 18114 73442
rect 19294 73390 19346 73442
rect 20750 73390 20802 73442
rect 23998 73390 24050 73442
rect 26014 73390 26066 73442
rect 1710 73278 1762 73330
rect 2718 73278 2770 73330
rect 3166 73278 3218 73330
rect 4958 73278 5010 73330
rect 13134 73278 13186 73330
rect 13358 73278 13410 73330
rect 13694 73278 13746 73330
rect 13806 73278 13858 73330
rect 15934 73278 15986 73330
rect 17502 73278 17554 73330
rect 17950 73278 18002 73330
rect 18286 73278 18338 73330
rect 21086 73278 21138 73330
rect 21310 73278 21362 73330
rect 21870 73278 21922 73330
rect 22542 73278 22594 73330
rect 23438 73278 23490 73330
rect 23774 73278 23826 73330
rect 25342 73278 25394 73330
rect 3502 73166 3554 73218
rect 4174 73166 4226 73218
rect 4622 73166 4674 73218
rect 5742 73166 5794 73218
rect 7870 73166 7922 73218
rect 8318 73166 8370 73218
rect 13918 73166 13970 73218
rect 14590 73166 14642 73218
rect 15150 73166 15202 73218
rect 16382 73166 16434 73218
rect 16718 73166 16770 73218
rect 18734 73166 18786 73218
rect 19854 73166 19906 73218
rect 22318 73166 22370 73218
rect 22990 73166 23042 73218
rect 24446 73166 24498 73218
rect 28142 73166 28194 73218
rect 2382 73054 2434 73106
rect 2718 73054 2770 73106
rect 17278 73054 17330 73106
rect 19406 73054 19458 73106
rect 21646 73054 21698 73106
rect 22206 73054 22258 73106
rect 24334 73054 24386 73106
rect 4616 72886 4668 72938
rect 4720 72886 4772 72938
rect 4824 72886 4876 72938
rect 11420 72886 11472 72938
rect 11524 72886 11576 72938
rect 11628 72886 11680 72938
rect 18224 72886 18276 72938
rect 18328 72886 18380 72938
rect 18432 72886 18484 72938
rect 25028 72886 25080 72938
rect 25132 72886 25184 72938
rect 25236 72886 25288 72938
rect 8430 72718 8482 72770
rect 13694 72718 13746 72770
rect 14254 72718 14306 72770
rect 4622 72606 4674 72658
rect 5854 72606 5906 72658
rect 6190 72606 6242 72658
rect 6974 72606 7026 72658
rect 7982 72606 8034 72658
rect 12238 72606 12290 72658
rect 12910 72606 12962 72658
rect 13918 72606 13970 72658
rect 17838 72606 17890 72658
rect 18958 72606 19010 72658
rect 21422 72606 21474 72658
rect 27694 72606 27746 72658
rect 1822 72494 1874 72546
rect 6078 72494 6130 72546
rect 6302 72494 6354 72546
rect 7198 72494 7250 72546
rect 8318 72494 8370 72546
rect 8542 72494 8594 72546
rect 8766 72494 8818 72546
rect 8990 72494 9042 72546
rect 9326 72494 9378 72546
rect 13582 72494 13634 72546
rect 14142 72494 14194 72546
rect 15598 72494 15650 72546
rect 16382 72494 16434 72546
rect 18622 72494 18674 72546
rect 19182 72494 19234 72546
rect 22318 72494 22370 72546
rect 22430 72494 22482 72546
rect 22990 72494 23042 72546
rect 23214 72494 23266 72546
rect 23438 72494 23490 72546
rect 25678 72494 25730 72546
rect 2494 72382 2546 72434
rect 5070 72382 5122 72434
rect 5742 72382 5794 72434
rect 6862 72382 6914 72434
rect 10110 72382 10162 72434
rect 15262 72382 15314 72434
rect 16270 72382 16322 72434
rect 18510 72382 18562 72434
rect 21870 72382 21922 72434
rect 22094 72382 22146 72434
rect 19518 72270 19570 72322
rect 20190 72270 20242 72322
rect 20638 72270 20690 72322
rect 22206 72270 22258 72322
rect 23326 72270 23378 72322
rect 23550 72270 23602 72322
rect 24110 72270 24162 72322
rect 24558 72270 24610 72322
rect 25006 72270 25058 72322
rect 8018 72102 8070 72154
rect 8122 72102 8174 72154
rect 8226 72102 8278 72154
rect 14822 72102 14874 72154
rect 14926 72102 14978 72154
rect 15030 72102 15082 72154
rect 21626 72102 21678 72154
rect 21730 72102 21782 72154
rect 21834 72102 21886 72154
rect 28430 72102 28482 72154
rect 28534 72102 28586 72154
rect 28638 72102 28690 72154
rect 2494 71934 2546 71986
rect 7646 71934 7698 71986
rect 8542 71934 8594 71986
rect 8878 71934 8930 71986
rect 10558 71934 10610 71986
rect 11678 71934 11730 71986
rect 12462 71934 12514 71986
rect 12910 71934 12962 71986
rect 14366 71934 14418 71986
rect 15150 71934 15202 71986
rect 18846 71934 18898 71986
rect 23550 71934 23602 71986
rect 24558 71934 24610 71986
rect 26462 71934 26514 71986
rect 27470 71934 27522 71986
rect 28142 71934 28194 71986
rect 2270 71822 2322 71874
rect 10446 71822 10498 71874
rect 11006 71822 11058 71874
rect 11566 71822 11618 71874
rect 14254 71822 14306 71874
rect 16382 71822 16434 71874
rect 19406 71822 19458 71874
rect 21982 71822 22034 71874
rect 2606 71710 2658 71762
rect 2718 71710 2770 71762
rect 3054 71710 3106 71762
rect 3390 71710 3442 71762
rect 4398 71710 4450 71762
rect 5070 71710 5122 71762
rect 8766 71710 8818 71762
rect 8990 71710 9042 71762
rect 9550 71710 9602 71762
rect 9774 71710 9826 71762
rect 10222 71710 10274 71762
rect 10782 71710 10834 71762
rect 11454 71710 11506 71762
rect 12126 71710 12178 71762
rect 15710 71710 15762 71762
rect 15934 71710 15986 71762
rect 16158 71710 16210 71762
rect 17502 71710 17554 71762
rect 17950 71710 18002 71762
rect 18062 71710 18114 71762
rect 19070 71710 19122 71762
rect 20414 71710 20466 71762
rect 22654 71710 22706 71762
rect 23438 71710 23490 71762
rect 23774 71710 23826 71762
rect 23998 71710 24050 71762
rect 24334 71710 24386 71762
rect 26686 71710 26738 71762
rect 27134 71710 27186 71762
rect 3502 71598 3554 71650
rect 3950 71598 4002 71650
rect 7198 71598 7250 71650
rect 8094 71598 8146 71650
rect 9662 71598 9714 71650
rect 16270 71598 16322 71650
rect 18286 71598 18338 71650
rect 23662 71598 23714 71650
rect 25342 71598 25394 71650
rect 26014 71598 26066 71650
rect 26574 71598 26626 71650
rect 7534 71486 7586 71538
rect 8094 71486 8146 71538
rect 13470 71486 13522 71538
rect 13582 71486 13634 71538
rect 13806 71486 13858 71538
rect 13918 71486 13970 71538
rect 15486 71486 15538 71538
rect 17278 71486 17330 71538
rect 24670 71486 24722 71538
rect 4616 71318 4668 71370
rect 4720 71318 4772 71370
rect 4824 71318 4876 71370
rect 11420 71318 11472 71370
rect 11524 71318 11576 71370
rect 11628 71318 11680 71370
rect 18224 71318 18276 71370
rect 18328 71318 18380 71370
rect 18432 71318 18484 71370
rect 25028 71318 25080 71370
rect 25132 71318 25184 71370
rect 25236 71318 25288 71370
rect 3502 71150 3554 71202
rect 3950 71150 4002 71202
rect 7310 71150 7362 71202
rect 8094 71150 8146 71202
rect 8430 71150 8482 71202
rect 14926 71150 14978 71202
rect 15150 71150 15202 71202
rect 5742 71038 5794 71090
rect 8318 71038 8370 71090
rect 8878 71038 8930 71090
rect 9550 71038 9602 71090
rect 13582 71038 13634 71090
rect 14254 71038 14306 71090
rect 15374 71038 15426 71090
rect 18846 71038 18898 71090
rect 22206 71038 22258 71090
rect 24334 71038 24386 71090
rect 28142 71038 28194 71090
rect 1822 70926 1874 70978
rect 3502 70926 3554 70978
rect 6078 70926 6130 70978
rect 6190 70926 6242 70978
rect 6862 70926 6914 70978
rect 7086 70926 7138 70978
rect 9998 70926 10050 70978
rect 11230 70926 11282 70978
rect 13806 70926 13858 70978
rect 14030 70926 14082 70978
rect 14478 70926 14530 70978
rect 16830 70926 16882 70978
rect 17278 70926 17330 70978
rect 19294 70926 19346 70978
rect 20190 70926 20242 70978
rect 21534 70926 21586 70978
rect 25342 70926 25394 70978
rect 4622 70814 4674 70866
rect 5630 70814 5682 70866
rect 5854 70814 5906 70866
rect 6750 70814 6802 70866
rect 14254 70814 14306 70866
rect 16270 70814 16322 70866
rect 17950 70814 18002 70866
rect 18398 70814 18450 70866
rect 20750 70814 20802 70866
rect 26014 70814 26066 70866
rect 2046 70702 2098 70754
rect 2606 70702 2658 70754
rect 3054 70702 3106 70754
rect 3950 70702 4002 70754
rect 5182 70702 5234 70754
rect 7534 70702 7586 70754
rect 7982 70702 8034 70754
rect 9438 70702 9490 70754
rect 9662 70702 9714 70754
rect 10446 70702 10498 70754
rect 12462 70702 12514 70754
rect 12910 70702 12962 70754
rect 15598 70702 15650 70754
rect 15710 70702 15762 70754
rect 15822 70702 15874 70754
rect 17838 70702 17890 70754
rect 18286 70702 18338 70754
rect 19518 70702 19570 70754
rect 19630 70702 19682 70754
rect 24782 70702 24834 70754
rect 8018 70534 8070 70586
rect 8122 70534 8174 70586
rect 8226 70534 8278 70586
rect 14822 70534 14874 70586
rect 14926 70534 14978 70586
rect 15030 70534 15082 70586
rect 21626 70534 21678 70586
rect 21730 70534 21782 70586
rect 21834 70534 21886 70586
rect 28430 70534 28482 70586
rect 28534 70534 28586 70586
rect 28638 70534 28690 70586
rect 2270 70366 2322 70418
rect 9774 70366 9826 70418
rect 10222 70366 10274 70418
rect 10894 70366 10946 70418
rect 11342 70366 11394 70418
rect 13022 70366 13074 70418
rect 21310 70366 21362 70418
rect 25678 70366 25730 70418
rect 26126 70366 26178 70418
rect 27918 70366 27970 70418
rect 9550 70254 9602 70306
rect 15038 70254 15090 70306
rect 15934 70254 15986 70306
rect 26350 70254 26402 70306
rect 26574 70254 26626 70306
rect 27022 70254 27074 70306
rect 2718 70142 2770 70194
rect 7870 70142 7922 70194
rect 9998 70142 10050 70194
rect 10222 70142 10274 70194
rect 12238 70142 12290 70194
rect 12462 70142 12514 70194
rect 12910 70142 12962 70194
rect 13134 70142 13186 70194
rect 15262 70142 15314 70194
rect 15598 70142 15650 70194
rect 17390 70142 17442 70194
rect 22094 70142 22146 70194
rect 25902 70142 25954 70194
rect 3054 70030 3106 70082
rect 5070 70030 5122 70082
rect 11902 70030 11954 70082
rect 12686 70030 12738 70082
rect 14254 70030 14306 70082
rect 18174 70030 18226 70082
rect 20302 70030 20354 70082
rect 20750 70030 20802 70082
rect 21758 70030 21810 70082
rect 23886 70030 23938 70082
rect 27470 70030 27522 70082
rect 2046 69918 2098 69970
rect 2382 69918 2434 69970
rect 26910 69918 26962 69970
rect 4616 69750 4668 69802
rect 4720 69750 4772 69802
rect 4824 69750 4876 69802
rect 11420 69750 11472 69802
rect 11524 69750 11576 69802
rect 11628 69750 11680 69802
rect 18224 69750 18276 69802
rect 18328 69750 18380 69802
rect 18432 69750 18484 69802
rect 25028 69750 25080 69802
rect 25132 69750 25184 69802
rect 25236 69750 25288 69802
rect 8318 69582 8370 69634
rect 11790 69582 11842 69634
rect 12350 69582 12402 69634
rect 12686 69582 12738 69634
rect 4622 69470 4674 69522
rect 13358 69470 13410 69522
rect 16494 69470 16546 69522
rect 19406 69470 19458 69522
rect 21646 69470 21698 69522
rect 21982 69470 22034 69522
rect 23550 69470 23602 69522
rect 25342 69470 25394 69522
rect 25790 69470 25842 69522
rect 1710 69358 1762 69410
rect 8206 69358 8258 69410
rect 8766 69358 8818 69410
rect 13470 69358 13522 69410
rect 14030 69358 14082 69410
rect 14814 69358 14866 69410
rect 15822 69358 15874 69410
rect 16270 69358 16322 69410
rect 18286 69358 18338 69410
rect 18958 69358 19010 69410
rect 19518 69358 19570 69410
rect 19854 69358 19906 69410
rect 22318 69358 22370 69410
rect 26686 69358 26738 69410
rect 27582 69358 27634 69410
rect 2494 69246 2546 69298
rect 9326 69246 9378 69298
rect 12574 69246 12626 69298
rect 15262 69246 15314 69298
rect 16830 69246 16882 69298
rect 18734 69246 18786 69298
rect 26350 69246 26402 69298
rect 26910 69246 26962 69298
rect 27246 69246 27298 69298
rect 27806 69246 27858 69298
rect 5070 69134 5122 69186
rect 7870 69134 7922 69186
rect 9214 69134 9266 69186
rect 9438 69134 9490 69186
rect 10446 69134 10498 69186
rect 11790 69134 11842 69186
rect 12238 69134 12290 69186
rect 13694 69134 13746 69186
rect 13918 69134 13970 69186
rect 17390 69134 17442 69186
rect 17838 69134 17890 69186
rect 18622 69134 18674 69186
rect 19294 69134 19346 69186
rect 20414 69134 20466 69186
rect 20750 69134 20802 69186
rect 26574 69134 26626 69186
rect 27582 69134 27634 69186
rect 8018 68966 8070 69018
rect 8122 68966 8174 69018
rect 8226 68966 8278 69018
rect 14822 68966 14874 69018
rect 14926 68966 14978 69018
rect 15030 68966 15082 69018
rect 21626 68966 21678 69018
rect 21730 68966 21782 69018
rect 21834 68966 21886 69018
rect 28430 68966 28482 69018
rect 28534 68966 28586 69018
rect 28638 68966 28690 69018
rect 2606 68798 2658 68850
rect 8430 68798 8482 68850
rect 8990 68798 9042 68850
rect 14926 68798 14978 68850
rect 15374 68798 15426 68850
rect 16830 68798 16882 68850
rect 19406 68798 19458 68850
rect 20302 68798 20354 68850
rect 20750 68798 20802 68850
rect 3054 68686 3106 68738
rect 12798 68686 12850 68738
rect 17838 68686 17890 68738
rect 27358 68686 27410 68738
rect 2494 68574 2546 68626
rect 2830 68574 2882 68626
rect 3390 68574 3442 68626
rect 4846 68574 4898 68626
rect 9550 68574 9602 68626
rect 14030 68574 14082 68626
rect 17390 68574 17442 68626
rect 17614 68574 17666 68626
rect 22318 68574 22370 68626
rect 28142 68574 28194 68626
rect 3502 68462 3554 68514
rect 3950 68462 4002 68514
rect 4398 68462 4450 68514
rect 5518 68462 5570 68514
rect 7646 68462 7698 68514
rect 8318 68462 8370 68514
rect 10334 68462 10386 68514
rect 12462 68462 12514 68514
rect 14254 68462 14306 68514
rect 17502 68462 17554 68514
rect 18510 68462 18562 68514
rect 18958 68462 19010 68514
rect 19854 68462 19906 68514
rect 21198 68462 21250 68514
rect 21758 68462 21810 68514
rect 24222 68462 24274 68514
rect 25230 68462 25282 68514
rect 2494 68350 2546 68402
rect 3950 68350 4002 68402
rect 4510 68350 4562 68402
rect 19294 68350 19346 68402
rect 19966 68350 20018 68402
rect 21198 68350 21250 68402
rect 4616 68182 4668 68234
rect 4720 68182 4772 68234
rect 4824 68182 4876 68234
rect 11420 68182 11472 68234
rect 11524 68182 11576 68234
rect 11628 68182 11680 68234
rect 18224 68182 18276 68234
rect 18328 68182 18380 68234
rect 18432 68182 18484 68234
rect 25028 68182 25080 68234
rect 25132 68182 25184 68234
rect 25236 68182 25288 68234
rect 3278 67902 3330 67954
rect 6078 67902 6130 67954
rect 7758 67902 7810 67954
rect 10446 67902 10498 67954
rect 12910 67902 12962 67954
rect 13470 67902 13522 67954
rect 16046 67902 16098 67954
rect 21646 67902 21698 67954
rect 24222 67902 24274 67954
rect 27022 67902 27074 67954
rect 28142 67902 28194 67954
rect 10222 67790 10274 67842
rect 10894 67790 10946 67842
rect 11566 67790 11618 67842
rect 11678 67790 11730 67842
rect 12014 67790 12066 67842
rect 13694 67790 13746 67842
rect 18958 67790 19010 67842
rect 19294 67790 19346 67842
rect 20190 67790 20242 67842
rect 21870 67790 21922 67842
rect 22878 67790 22930 67842
rect 26014 67790 26066 67842
rect 5182 67678 5234 67730
rect 5966 67678 6018 67730
rect 6302 67678 6354 67730
rect 6526 67678 6578 67730
rect 10670 67678 10722 67730
rect 14030 67678 14082 67730
rect 18174 67678 18226 67730
rect 20526 67678 20578 67730
rect 21534 67678 21586 67730
rect 23214 67678 23266 67730
rect 27358 67678 27410 67730
rect 1822 67566 1874 67618
rect 7086 67566 7138 67618
rect 9662 67566 9714 67618
rect 9998 67566 10050 67618
rect 11454 67566 11506 67618
rect 12462 67566 12514 67618
rect 14478 67566 14530 67618
rect 19406 67566 19458 67618
rect 19630 67566 19682 67618
rect 22318 67566 22370 67618
rect 22990 67566 23042 67618
rect 23102 67566 23154 67618
rect 23326 67566 23378 67618
rect 26910 67566 26962 67618
rect 27134 67566 27186 67618
rect 8018 67398 8070 67450
rect 8122 67398 8174 67450
rect 8226 67398 8278 67450
rect 14822 67398 14874 67450
rect 14926 67398 14978 67450
rect 15030 67398 15082 67450
rect 21626 67398 21678 67450
rect 21730 67398 21782 67450
rect 21834 67398 21886 67450
rect 28430 67398 28482 67450
rect 28534 67398 28586 67450
rect 28638 67398 28690 67450
rect 8094 67230 8146 67282
rect 11342 67230 11394 67282
rect 13134 67230 13186 67282
rect 14030 67230 14082 67282
rect 17838 67230 17890 67282
rect 18734 67230 18786 67282
rect 2046 67118 2098 67170
rect 15822 67118 15874 67170
rect 16718 67118 16770 67170
rect 17950 67118 18002 67170
rect 19406 67118 19458 67170
rect 24446 67118 24498 67170
rect 24558 67118 24610 67170
rect 24670 67118 24722 67170
rect 27358 67118 27410 67170
rect 1710 67006 1762 67058
rect 2718 67006 2770 67058
rect 3054 67006 3106 67058
rect 4734 67006 4786 67058
rect 7870 67006 7922 67058
rect 8430 67006 8482 67058
rect 8878 67006 8930 67058
rect 11566 67006 11618 67058
rect 12014 67006 12066 67058
rect 12574 67006 12626 67058
rect 16158 67006 16210 67058
rect 17502 67006 17554 67058
rect 17614 67006 17666 67058
rect 18398 67006 18450 67058
rect 19070 67006 19122 67058
rect 19518 67006 19570 67058
rect 19630 67006 19682 67058
rect 20190 67006 20242 67058
rect 23998 67006 24050 67058
rect 28142 67006 28194 67058
rect 3838 66894 3890 66946
rect 5406 66894 5458 66946
rect 7534 66894 7586 66946
rect 7982 66894 8034 66946
rect 8430 66894 8482 66946
rect 8766 66894 8818 66946
rect 9662 66894 9714 66946
rect 11006 66894 11058 66946
rect 11454 66894 11506 66946
rect 13582 66894 13634 66946
rect 15262 66894 15314 66946
rect 20862 66894 20914 66946
rect 22990 66894 23042 66946
rect 23438 66894 23490 66946
rect 25230 66894 25282 66946
rect 2382 66782 2434 66834
rect 2718 66782 2770 66834
rect 3166 66782 3218 66834
rect 10782 66782 10834 66834
rect 11118 66782 11170 66834
rect 12798 66782 12850 66834
rect 15486 66782 15538 66834
rect 16382 66782 16434 66834
rect 4616 66614 4668 66666
rect 4720 66614 4772 66666
rect 4824 66614 4876 66666
rect 11420 66614 11472 66666
rect 11524 66614 11576 66666
rect 11628 66614 11680 66666
rect 18224 66614 18276 66666
rect 18328 66614 18380 66666
rect 18432 66614 18484 66666
rect 25028 66614 25080 66666
rect 25132 66614 25184 66666
rect 25236 66614 25288 66666
rect 21534 66446 21586 66498
rect 4622 66334 4674 66386
rect 5966 66334 6018 66386
rect 9550 66334 9602 66386
rect 12910 66334 12962 66386
rect 16382 66334 16434 66386
rect 17838 66334 17890 66386
rect 27918 66334 27970 66386
rect 1710 66222 1762 66274
rect 6078 66222 6130 66274
rect 6414 66222 6466 66274
rect 8318 66222 8370 66274
rect 13470 66222 13522 66274
rect 14254 66222 14306 66274
rect 17502 66222 17554 66274
rect 18510 66222 18562 66274
rect 21534 66222 21586 66274
rect 22878 66222 22930 66274
rect 2494 66110 2546 66162
rect 5182 66110 5234 66162
rect 5854 66110 5906 66162
rect 16830 66110 16882 66162
rect 17614 66110 17666 66162
rect 21870 66110 21922 66162
rect 22094 66110 22146 66162
rect 22542 66110 22594 66162
rect 6862 65998 6914 66050
rect 18846 65998 18898 66050
rect 19406 65998 19458 66050
rect 19966 65998 20018 66050
rect 20750 65998 20802 66050
rect 21310 65998 21362 66050
rect 8018 65830 8070 65882
rect 8122 65830 8174 65882
rect 8226 65830 8278 65882
rect 14822 65830 14874 65882
rect 14926 65830 14978 65882
rect 15030 65830 15082 65882
rect 21626 65830 21678 65882
rect 21730 65830 21782 65882
rect 21834 65830 21886 65882
rect 28430 65830 28482 65882
rect 28534 65830 28586 65882
rect 28638 65830 28690 65882
rect 2606 65662 2658 65714
rect 3390 65662 3442 65714
rect 7534 65662 7586 65714
rect 13582 65662 13634 65714
rect 14702 65662 14754 65714
rect 15934 65662 15986 65714
rect 23326 65662 23378 65714
rect 2830 65550 2882 65602
rect 3054 65550 3106 65602
rect 4398 65550 4450 65602
rect 13470 65550 13522 65602
rect 14478 65550 14530 65602
rect 17950 65550 18002 65602
rect 18062 65550 18114 65602
rect 18734 65550 18786 65602
rect 23102 65550 23154 65602
rect 2494 65438 2546 65490
rect 2606 65438 2658 65490
rect 7310 65438 7362 65490
rect 7422 65438 7474 65490
rect 7982 65438 8034 65490
rect 9662 65438 9714 65490
rect 13806 65438 13858 65490
rect 14030 65438 14082 65490
rect 14590 65438 14642 65490
rect 15150 65438 15202 65490
rect 17278 65438 17330 65490
rect 17502 65438 17554 65490
rect 21422 65438 21474 65490
rect 22878 65438 22930 65490
rect 23550 65438 23602 65490
rect 23998 65438 24050 65490
rect 24446 65438 24498 65490
rect 25342 65438 25394 65490
rect 25790 65438 25842 65490
rect 26126 65438 26178 65490
rect 26350 65438 26402 65490
rect 26910 65438 26962 65490
rect 27806 65438 27858 65490
rect 3502 65326 3554 65378
rect 3950 65326 4002 65378
rect 4846 65326 4898 65378
rect 8318 65326 8370 65378
rect 8766 65326 8818 65378
rect 10334 65326 10386 65378
rect 12462 65326 12514 65378
rect 13134 65326 13186 65378
rect 15486 65326 15538 65378
rect 16382 65326 16434 65378
rect 16942 65326 16994 65378
rect 18286 65326 18338 65378
rect 19406 65326 19458 65378
rect 19966 65326 20018 65378
rect 20974 65326 21026 65378
rect 21870 65326 21922 65378
rect 22318 65326 22370 65378
rect 23214 65326 23266 65378
rect 25902 65326 25954 65378
rect 27358 65326 27410 65378
rect 15486 65214 15538 65266
rect 16158 65214 16210 65266
rect 16830 65214 16882 65266
rect 20974 65214 21026 65266
rect 22094 65214 22146 65266
rect 4616 65046 4668 65098
rect 4720 65046 4772 65098
rect 4824 65046 4876 65098
rect 11420 65046 11472 65098
rect 11524 65046 11576 65098
rect 11628 65046 11680 65098
rect 18224 65046 18276 65098
rect 18328 65046 18380 65098
rect 18432 65046 18484 65098
rect 25028 65046 25080 65098
rect 25132 65046 25184 65098
rect 25236 65046 25288 65098
rect 3726 64878 3778 64930
rect 3950 64878 4002 64930
rect 12350 64878 12402 64930
rect 13022 64878 13074 64930
rect 16942 64878 16994 64930
rect 17166 64878 17218 64930
rect 17502 64878 17554 64930
rect 8542 64766 8594 64818
rect 8990 64766 9042 64818
rect 10334 64766 10386 64818
rect 18846 64766 18898 64818
rect 24222 64766 24274 64818
rect 24670 64766 24722 64818
rect 26014 64766 26066 64818
rect 28142 64766 28194 64818
rect 4174 64654 4226 64706
rect 5742 64654 5794 64706
rect 10446 64654 10498 64706
rect 10782 64654 10834 64706
rect 16942 64654 16994 64706
rect 20414 64654 20466 64706
rect 20526 64654 20578 64706
rect 21310 64654 21362 64706
rect 25342 64654 25394 64706
rect 1710 64542 1762 64594
rect 3054 64542 3106 64594
rect 4622 64542 4674 64594
rect 6414 64542 6466 64594
rect 10222 64542 10274 64594
rect 11230 64542 11282 64594
rect 19182 64542 19234 64594
rect 19966 64542 20018 64594
rect 20190 64542 20242 64594
rect 22094 64542 22146 64594
rect 2046 64430 2098 64482
rect 2830 64430 2882 64482
rect 2942 64430 2994 64482
rect 3726 64430 3778 64482
rect 9886 64430 9938 64482
rect 12686 64430 12738 64482
rect 13582 64430 13634 64482
rect 14254 64430 14306 64482
rect 17390 64430 17442 64482
rect 18958 64430 19010 64482
rect 19630 64430 19682 64482
rect 20750 64430 20802 64482
rect 8018 64262 8070 64314
rect 8122 64262 8174 64314
rect 8226 64262 8278 64314
rect 14822 64262 14874 64314
rect 14926 64262 14978 64314
rect 15030 64262 15082 64314
rect 21626 64262 21678 64314
rect 21730 64262 21782 64314
rect 21834 64262 21886 64314
rect 28430 64262 28482 64314
rect 28534 64262 28586 64314
rect 28638 64262 28690 64314
rect 2494 64094 2546 64146
rect 6302 64094 6354 64146
rect 7646 64094 7698 64146
rect 13582 64094 13634 64146
rect 20974 64094 21026 64146
rect 21870 64094 21922 64146
rect 24670 64094 24722 64146
rect 25566 64094 25618 64146
rect 25678 64094 25730 64146
rect 27022 64094 27074 64146
rect 3278 63982 3330 64034
rect 22430 63982 22482 64034
rect 26126 63982 26178 64034
rect 26350 63982 26402 64034
rect 27470 63982 27522 64034
rect 28030 63982 28082 64034
rect 1822 63870 1874 63922
rect 2718 63870 2770 63922
rect 2830 63870 2882 63922
rect 3054 63870 3106 63922
rect 3950 63870 4002 63922
rect 4510 63870 4562 63922
rect 5742 63870 5794 63922
rect 6078 63870 6130 63922
rect 6302 63870 6354 63922
rect 6638 63870 6690 63922
rect 7422 63870 7474 63922
rect 8094 63870 8146 63922
rect 8430 63870 8482 63922
rect 10110 63870 10162 63922
rect 13918 63870 13970 63922
rect 20414 63870 20466 63922
rect 21758 63870 21810 63922
rect 23102 63870 23154 63922
rect 23550 63870 23602 63922
rect 23774 63870 23826 63922
rect 24222 63870 24274 63922
rect 25118 63870 25170 63922
rect 25790 63870 25842 63922
rect 26798 63870 26850 63922
rect 27246 63870 27298 63922
rect 7086 63758 7138 63810
rect 7534 63758 7586 63810
rect 8878 63758 8930 63810
rect 9550 63758 9602 63810
rect 10894 63758 10946 63810
rect 13022 63758 13074 63810
rect 14702 63758 14754 63810
rect 16830 63758 16882 63810
rect 17614 63758 17666 63810
rect 19742 63758 19794 63810
rect 22878 63758 22930 63810
rect 23662 63758 23714 63810
rect 26574 63758 26626 63810
rect 27134 63758 27186 63810
rect 9662 63646 9714 63698
rect 21086 63646 21138 63698
rect 21422 63646 21474 63698
rect 21646 63646 21698 63698
rect 23998 63646 24050 63698
rect 24670 63646 24722 63698
rect 4616 63478 4668 63530
rect 4720 63478 4772 63530
rect 4824 63478 4876 63530
rect 11420 63478 11472 63530
rect 11524 63478 11576 63530
rect 11628 63478 11680 63530
rect 18224 63478 18276 63530
rect 18328 63478 18380 63530
rect 18432 63478 18484 63530
rect 25028 63478 25080 63530
rect 25132 63478 25184 63530
rect 25236 63478 25288 63530
rect 17614 63310 17666 63362
rect 18174 63310 18226 63362
rect 18846 63310 18898 63362
rect 19294 63310 19346 63362
rect 19742 63310 19794 63362
rect 2494 63198 2546 63250
rect 4622 63198 4674 63250
rect 5070 63198 5122 63250
rect 9662 63198 9714 63250
rect 11342 63198 11394 63250
rect 14478 63198 14530 63250
rect 14926 63198 14978 63250
rect 15374 63198 15426 63250
rect 16270 63198 16322 63250
rect 17726 63198 17778 63250
rect 23998 63198 24050 63250
rect 27022 63198 27074 63250
rect 27470 63198 27522 63250
rect 28142 63198 28194 63250
rect 1710 63086 1762 63138
rect 6750 63086 6802 63138
rect 10222 63086 10274 63138
rect 10558 63086 10610 63138
rect 11566 63086 11618 63138
rect 11790 63086 11842 63138
rect 12462 63086 12514 63138
rect 13470 63086 13522 63138
rect 15262 63086 15314 63138
rect 15486 63086 15538 63138
rect 15822 63086 15874 63138
rect 16158 63086 16210 63138
rect 16382 63086 16434 63138
rect 17166 63086 17218 63138
rect 19182 63086 19234 63138
rect 19630 63086 19682 63138
rect 20078 63086 20130 63138
rect 21422 63086 21474 63138
rect 7534 62974 7586 63026
rect 11230 62974 11282 63026
rect 12350 62974 12402 63026
rect 16606 62974 16658 63026
rect 18398 62974 18450 63026
rect 18622 62974 18674 63026
rect 9998 62862 10050 62914
rect 10110 62862 10162 62914
rect 12238 62862 12290 62914
rect 12686 62862 12738 62914
rect 13582 62862 13634 62914
rect 14030 62862 14082 62914
rect 19182 62862 19234 62914
rect 20526 62862 20578 62914
rect 8018 62694 8070 62746
rect 8122 62694 8174 62746
rect 8226 62694 8278 62746
rect 14822 62694 14874 62746
rect 14926 62694 14978 62746
rect 15030 62694 15082 62746
rect 21626 62694 21678 62746
rect 21730 62694 21782 62746
rect 21834 62694 21886 62746
rect 28430 62694 28482 62746
rect 28534 62694 28586 62746
rect 28638 62694 28690 62746
rect 3502 62526 3554 62578
rect 7870 62526 7922 62578
rect 8766 62526 8818 62578
rect 9886 62526 9938 62578
rect 10558 62526 10610 62578
rect 11006 62526 11058 62578
rect 11454 62526 11506 62578
rect 12014 62526 12066 62578
rect 12462 62526 12514 62578
rect 13022 62526 13074 62578
rect 13582 62526 13634 62578
rect 19294 62526 19346 62578
rect 19742 62526 19794 62578
rect 20190 62526 20242 62578
rect 20638 62526 20690 62578
rect 24670 62526 24722 62578
rect 3614 62414 3666 62466
rect 8318 62414 8370 62466
rect 14478 62414 14530 62466
rect 16270 62414 16322 62466
rect 17502 62414 17554 62466
rect 18622 62414 18674 62466
rect 27358 62414 27410 62466
rect 7758 62302 7810 62354
rect 8094 62302 8146 62354
rect 14366 62302 14418 62354
rect 14702 62302 14754 62354
rect 15374 62302 15426 62354
rect 16830 62302 16882 62354
rect 17614 62302 17666 62354
rect 18286 62302 18338 62354
rect 21310 62302 21362 62354
rect 28030 62302 28082 62354
rect 2494 62190 2546 62242
rect 6638 62190 6690 62242
rect 7422 62190 7474 62242
rect 15822 62190 15874 62242
rect 17502 62190 17554 62242
rect 22094 62190 22146 62242
rect 24222 62190 24274 62242
rect 25230 62190 25282 62242
rect 15374 62078 15426 62130
rect 16046 62078 16098 62130
rect 4616 61910 4668 61962
rect 4720 61910 4772 61962
rect 4824 61910 4876 61962
rect 11420 61910 11472 61962
rect 11524 61910 11576 61962
rect 11628 61910 11680 61962
rect 18224 61910 18276 61962
rect 18328 61910 18380 61962
rect 18432 61910 18484 61962
rect 25028 61910 25080 61962
rect 25132 61910 25184 61962
rect 25236 61910 25288 61962
rect 14478 61742 14530 61794
rect 2830 61630 2882 61682
rect 3502 61630 3554 61682
rect 4622 61630 4674 61682
rect 5070 61630 5122 61682
rect 7982 61630 8034 61682
rect 11790 61630 11842 61682
rect 12686 61630 12738 61682
rect 13582 61630 13634 61682
rect 17838 61630 17890 61682
rect 21422 61630 21474 61682
rect 22430 61630 22482 61682
rect 26910 61630 26962 61682
rect 3278 61518 3330 61570
rect 5966 61518 6018 61570
rect 6078 61518 6130 61570
rect 6190 61518 6242 61570
rect 6862 61518 6914 61570
rect 7086 61518 7138 61570
rect 8990 61518 9042 61570
rect 12350 61518 12402 61570
rect 14142 61518 14194 61570
rect 14926 61518 14978 61570
rect 15262 61518 15314 61570
rect 16046 61518 16098 61570
rect 16830 61518 16882 61570
rect 17278 61518 17330 61570
rect 20750 61518 20802 61570
rect 22654 61518 22706 61570
rect 22878 61518 22930 61570
rect 23326 61518 23378 61570
rect 23998 61518 24050 61570
rect 24222 61518 24274 61570
rect 24670 61518 24722 61570
rect 25678 61518 25730 61570
rect 1710 61406 1762 61458
rect 2046 61406 2098 61458
rect 5630 61406 5682 61458
rect 6750 61406 6802 61458
rect 9662 61406 9714 61458
rect 12126 61406 12178 61458
rect 13918 61406 13970 61458
rect 16158 61406 16210 61458
rect 19966 61406 20018 61458
rect 22318 61406 22370 61458
rect 4174 61294 4226 61346
rect 5742 61294 5794 61346
rect 7534 61294 7586 61346
rect 12574 61294 12626 61346
rect 12686 61294 12738 61346
rect 17390 61294 17442 61346
rect 21982 61294 22034 61346
rect 24334 61294 24386 61346
rect 24446 61294 24498 61346
rect 25118 61294 25170 61346
rect 8018 61126 8070 61178
rect 8122 61126 8174 61178
rect 8226 61126 8278 61178
rect 14822 61126 14874 61178
rect 14926 61126 14978 61178
rect 15030 61126 15082 61178
rect 21626 61126 21678 61178
rect 21730 61126 21782 61178
rect 21834 61126 21886 61178
rect 28430 61126 28482 61178
rect 28534 61126 28586 61178
rect 28638 61126 28690 61178
rect 2046 60958 2098 61010
rect 2606 60958 2658 61010
rect 10334 60958 10386 61010
rect 19966 60958 20018 61010
rect 20414 60958 20466 61010
rect 25454 60958 25506 61010
rect 27582 60958 27634 61010
rect 3054 60846 3106 60898
rect 5070 60846 5122 60898
rect 11454 60846 11506 60898
rect 13806 60846 13858 60898
rect 14926 60846 14978 60898
rect 17614 60846 17666 60898
rect 19182 60846 19234 60898
rect 19406 60846 19458 60898
rect 2382 60734 2434 60786
rect 2830 60734 2882 60786
rect 3390 60734 3442 60786
rect 4398 60734 4450 60786
rect 7870 60734 7922 60786
rect 8318 60734 8370 60786
rect 10110 60734 10162 60786
rect 10334 60734 10386 60786
rect 10670 60734 10722 60786
rect 12462 60734 12514 60786
rect 14142 60734 14194 60786
rect 16382 60734 16434 60786
rect 17390 60734 17442 60786
rect 17950 60734 18002 60786
rect 18622 60734 18674 60786
rect 19742 60734 19794 60786
rect 21870 60734 21922 60786
rect 26574 60734 26626 60786
rect 26798 60734 26850 60786
rect 27246 60734 27298 60786
rect 3726 60622 3778 60674
rect 7198 60622 7250 60674
rect 7646 60622 7698 60674
rect 8990 60622 9042 60674
rect 9774 60622 9826 60674
rect 10894 60622 10946 60674
rect 11118 60622 11170 60674
rect 12350 60622 12402 60674
rect 13918 60622 13970 60674
rect 22430 60622 22482 60674
rect 24334 60622 24386 60674
rect 26238 60622 26290 60674
rect 26686 60622 26738 60674
rect 2606 60510 2658 60562
rect 3390 60510 3442 60562
rect 7534 60510 7586 60562
rect 17278 60510 17330 60562
rect 19630 60510 19682 60562
rect 20302 60510 20354 60562
rect 20638 60510 20690 60562
rect 4616 60342 4668 60394
rect 4720 60342 4772 60394
rect 4824 60342 4876 60394
rect 11420 60342 11472 60394
rect 11524 60342 11576 60394
rect 11628 60342 11680 60394
rect 18224 60342 18276 60394
rect 18328 60342 18380 60394
rect 18432 60342 18484 60394
rect 25028 60342 25080 60394
rect 25132 60342 25184 60394
rect 25236 60342 25288 60394
rect 14366 60174 14418 60226
rect 19518 60174 19570 60226
rect 20078 60174 20130 60226
rect 20414 60174 20466 60226
rect 2494 60062 2546 60114
rect 4622 60062 4674 60114
rect 8542 60062 8594 60114
rect 8990 60062 9042 60114
rect 11342 60062 11394 60114
rect 12910 60062 12962 60114
rect 21646 60062 21698 60114
rect 28142 60062 28194 60114
rect 1822 59950 1874 60002
rect 5742 59950 5794 60002
rect 11454 59950 11506 60002
rect 11902 59950 11954 60002
rect 13470 59950 13522 60002
rect 13806 59950 13858 60002
rect 14254 59950 14306 60002
rect 14590 59950 14642 60002
rect 16382 59950 16434 60002
rect 16942 59950 16994 60002
rect 18958 59950 19010 60002
rect 19518 59950 19570 60002
rect 20078 59950 20130 60002
rect 24558 59950 24610 60002
rect 25342 59950 25394 60002
rect 6414 59838 6466 59890
rect 14814 59838 14866 59890
rect 17390 59838 17442 59890
rect 19182 59838 19234 59890
rect 23774 59838 23826 59890
rect 26014 59838 26066 59890
rect 5070 59726 5122 59778
rect 10446 59726 10498 59778
rect 10894 59726 10946 59778
rect 11230 59726 11282 59778
rect 12462 59726 12514 59778
rect 13582 59726 13634 59778
rect 14030 59726 14082 59778
rect 18510 59726 18562 59778
rect 19070 59726 19122 59778
rect 8018 59558 8070 59610
rect 8122 59558 8174 59610
rect 8226 59558 8278 59610
rect 14822 59558 14874 59610
rect 14926 59558 14978 59610
rect 15030 59558 15082 59610
rect 21626 59558 21678 59610
rect 21730 59558 21782 59610
rect 21834 59558 21886 59610
rect 28430 59558 28482 59610
rect 28534 59558 28586 59610
rect 28638 59558 28690 59610
rect 3166 59390 3218 59442
rect 5742 59390 5794 59442
rect 6638 59390 6690 59442
rect 9886 59390 9938 59442
rect 13806 59390 13858 59442
rect 22766 59390 22818 59442
rect 23662 59390 23714 59442
rect 26014 59390 26066 59442
rect 28142 59390 28194 59442
rect 2046 59278 2098 59330
rect 3278 59278 3330 59330
rect 14478 59278 14530 59330
rect 14814 59278 14866 59330
rect 15822 59278 15874 59330
rect 20302 59278 20354 59330
rect 22878 59278 22930 59330
rect 25902 59278 25954 59330
rect 26462 59278 26514 59330
rect 26910 59278 26962 59330
rect 27358 59278 27410 59330
rect 1710 59166 1762 59218
rect 6526 59166 6578 59218
rect 6750 59166 6802 59218
rect 7310 59166 7362 59218
rect 7758 59166 7810 59218
rect 9774 59166 9826 59218
rect 10446 59166 10498 59218
rect 14142 59166 14194 59218
rect 15486 59166 15538 59218
rect 16606 59166 16658 59218
rect 16830 59166 16882 59218
rect 21086 59166 21138 59218
rect 22542 59166 22594 59218
rect 22990 59166 23042 59218
rect 23438 59166 23490 59218
rect 23550 59166 23602 59218
rect 23998 59166 24050 59218
rect 26238 59166 26290 59218
rect 2494 59054 2546 59106
rect 3726 59054 3778 59106
rect 6190 59054 6242 59106
rect 11230 59054 11282 59106
rect 13358 59054 13410 59106
rect 17502 59054 17554 59106
rect 18174 59054 18226 59106
rect 21534 59054 21586 59106
rect 21982 59054 22034 59106
rect 24446 59054 24498 59106
rect 25342 59054 25394 59106
rect 7086 58942 7138 58994
rect 7422 58942 7474 58994
rect 7646 58942 7698 58994
rect 9886 58942 9938 58994
rect 15710 58942 15762 58994
rect 17502 58942 17554 58994
rect 17838 58942 17890 58994
rect 4616 58774 4668 58826
rect 4720 58774 4772 58826
rect 4824 58774 4876 58826
rect 11420 58774 11472 58826
rect 11524 58774 11576 58826
rect 11628 58774 11680 58826
rect 18224 58774 18276 58826
rect 18328 58774 18380 58826
rect 18432 58774 18484 58826
rect 25028 58774 25080 58826
rect 25132 58774 25184 58826
rect 25236 58774 25288 58826
rect 2942 58606 2994 58658
rect 3726 58606 3778 58658
rect 10110 58606 10162 58658
rect 10334 58606 10386 58658
rect 11790 58606 11842 58658
rect 14590 58606 14642 58658
rect 14926 58606 14978 58658
rect 4622 58494 4674 58546
rect 6078 58494 6130 58546
rect 10558 58494 10610 58546
rect 11454 58494 11506 58546
rect 12686 58494 12738 58546
rect 14926 58494 14978 58546
rect 15598 58494 15650 58546
rect 22542 58606 22594 58658
rect 23326 58606 23378 58658
rect 16158 58494 16210 58546
rect 19406 58494 19458 58546
rect 20638 58494 20690 58546
rect 22206 58494 22258 58546
rect 23326 58494 23378 58546
rect 23774 58494 23826 58546
rect 28142 58494 28194 58546
rect 2830 58382 2882 58434
rect 5630 58382 5682 58434
rect 12014 58382 12066 58434
rect 12910 58382 12962 58434
rect 16382 58382 16434 58434
rect 18398 58382 18450 58434
rect 25342 58382 25394 58434
rect 3166 58270 3218 58322
rect 3390 58270 3442 58322
rect 4062 58270 4114 58322
rect 9214 58270 9266 58322
rect 11342 58270 11394 58322
rect 11566 58270 11618 58322
rect 12574 58270 12626 58322
rect 14030 58270 14082 58322
rect 16494 58270 16546 58322
rect 19518 58270 19570 58322
rect 26014 58270 26066 58322
rect 2270 58158 2322 58210
rect 2606 58158 2658 58210
rect 3838 58158 3890 58210
rect 9662 58158 9714 58210
rect 10110 58158 10162 58210
rect 11006 58158 11058 58210
rect 13582 58158 13634 58210
rect 14478 58158 14530 58210
rect 21422 58158 21474 58210
rect 21870 58158 21922 58210
rect 22318 58158 22370 58210
rect 22766 58158 22818 58210
rect 24446 58158 24498 58210
rect 24894 58158 24946 58210
rect 8018 57990 8070 58042
rect 8122 57990 8174 58042
rect 8226 57990 8278 58042
rect 14822 57990 14874 58042
rect 14926 57990 14978 58042
rect 15030 57990 15082 58042
rect 21626 57990 21678 58042
rect 21730 57990 21782 58042
rect 21834 57990 21886 58042
rect 28430 57990 28482 58042
rect 28534 57990 28586 58042
rect 28638 57990 28690 58042
rect 5070 57822 5122 57874
rect 5966 57822 6018 57874
rect 7086 57822 7138 57874
rect 7534 57822 7586 57874
rect 8094 57822 8146 57874
rect 8542 57822 8594 57874
rect 8990 57822 9042 57874
rect 9550 57822 9602 57874
rect 13022 57822 13074 57874
rect 13470 57822 13522 57874
rect 17502 57822 17554 57874
rect 24222 57822 24274 57874
rect 26014 57822 26066 57874
rect 27246 57822 27298 57874
rect 27806 57822 27858 57874
rect 2494 57710 2546 57762
rect 6302 57710 6354 57762
rect 15486 57710 15538 57762
rect 17950 57710 18002 57762
rect 19966 57710 20018 57762
rect 21646 57710 21698 57762
rect 22878 57710 22930 57762
rect 23886 57710 23938 57762
rect 25902 57710 25954 57762
rect 26238 57710 26290 57762
rect 1822 57598 1874 57650
rect 6638 57598 6690 57650
rect 9774 57598 9826 57650
rect 10110 57598 10162 57650
rect 10670 57598 10722 57650
rect 11902 57598 11954 57650
rect 12238 57598 12290 57650
rect 12462 57598 12514 57650
rect 15150 57598 15202 57650
rect 15598 57598 15650 57650
rect 17390 57598 17442 57650
rect 21198 57598 21250 57650
rect 23214 57598 23266 57650
rect 23438 57598 23490 57650
rect 23774 57598 23826 57650
rect 23998 57598 24050 57650
rect 26462 57598 26514 57650
rect 26798 57598 26850 57650
rect 26910 57598 26962 57650
rect 27022 57598 27074 57650
rect 4622 57486 4674 57538
rect 6414 57486 6466 57538
rect 9662 57486 9714 57538
rect 11118 57486 11170 57538
rect 11566 57486 11618 57538
rect 12014 57486 12066 57538
rect 13918 57486 13970 57538
rect 14590 57486 14642 57538
rect 16830 57486 16882 57538
rect 22542 57486 22594 57538
rect 22990 57486 23042 57538
rect 25342 57486 25394 57538
rect 6862 57374 6914 57426
rect 7198 57374 7250 57426
rect 8094 57374 8146 57426
rect 11006 57374 11058 57426
rect 11566 57374 11618 57426
rect 4616 57206 4668 57258
rect 4720 57206 4772 57258
rect 4824 57206 4876 57258
rect 11420 57206 11472 57258
rect 11524 57206 11576 57258
rect 11628 57206 11680 57258
rect 18224 57206 18276 57258
rect 18328 57206 18380 57258
rect 18432 57206 18484 57258
rect 25028 57206 25080 57258
rect 25132 57206 25184 57258
rect 25236 57206 25288 57258
rect 3502 57038 3554 57090
rect 6190 57038 6242 57090
rect 20190 57038 20242 57090
rect 5070 56926 5122 56978
rect 9662 56926 9714 56978
rect 10782 56926 10834 56978
rect 12910 56926 12962 56978
rect 13582 56926 13634 56978
rect 14590 56926 14642 56978
rect 22654 56926 22706 56978
rect 24782 56926 24834 56978
rect 25566 56926 25618 56978
rect 27694 56926 27746 56978
rect 28142 56926 28194 56978
rect 5630 56814 5682 56866
rect 6190 56814 6242 56866
rect 6862 56814 6914 56866
rect 10110 56814 10162 56866
rect 13470 56814 13522 56866
rect 14142 56814 14194 56866
rect 16606 56814 16658 56866
rect 17054 56814 17106 56866
rect 21982 56814 22034 56866
rect 3614 56702 3666 56754
rect 4062 56702 4114 56754
rect 5854 56702 5906 56754
rect 7534 56702 7586 56754
rect 15598 56702 15650 56754
rect 18174 56702 18226 56754
rect 19518 56702 19570 56754
rect 21422 56702 21474 56754
rect 26910 56702 26962 56754
rect 5742 56590 5794 56642
rect 13694 56590 13746 56642
rect 15038 56590 15090 56642
rect 18958 56590 19010 56642
rect 19070 56590 19122 56642
rect 19294 56590 19346 56642
rect 19966 56590 20018 56642
rect 20078 56590 20130 56642
rect 20638 56590 20690 56642
rect 26014 56590 26066 56642
rect 26462 56590 26514 56642
rect 8018 56422 8070 56474
rect 8122 56422 8174 56474
rect 8226 56422 8278 56474
rect 14822 56422 14874 56474
rect 14926 56422 14978 56474
rect 15030 56422 15082 56474
rect 21626 56422 21678 56474
rect 21730 56422 21782 56474
rect 21834 56422 21886 56474
rect 28430 56422 28482 56474
rect 28534 56422 28586 56474
rect 28638 56422 28690 56474
rect 8430 56254 8482 56306
rect 11790 56254 11842 56306
rect 11902 56254 11954 56306
rect 13134 56254 13186 56306
rect 17838 56254 17890 56306
rect 23438 56254 23490 56306
rect 2046 56142 2098 56194
rect 3614 56142 3666 56194
rect 3838 56142 3890 56194
rect 5294 56142 5346 56194
rect 8654 56142 8706 56194
rect 8878 56142 8930 56194
rect 10222 56142 10274 56194
rect 11230 56142 11282 56194
rect 12238 56142 12290 56194
rect 13582 56142 13634 56194
rect 15038 56142 15090 56194
rect 15598 56142 15650 56194
rect 23886 56142 23938 56194
rect 1710 56030 1762 56082
rect 4174 56030 4226 56082
rect 4622 56030 4674 56082
rect 8318 56030 8370 56082
rect 9774 56030 9826 56082
rect 9998 56030 10050 56082
rect 10446 56030 10498 56082
rect 10894 56030 10946 56082
rect 11678 56030 11730 56082
rect 12014 56030 12066 56082
rect 12574 56030 12626 56082
rect 12798 56030 12850 56082
rect 12910 56030 12962 56082
rect 13022 56030 13074 56082
rect 13694 56030 13746 56082
rect 14478 56030 14530 56082
rect 14814 56030 14866 56082
rect 15486 56030 15538 56082
rect 16158 56030 16210 56082
rect 16606 56030 16658 56082
rect 17950 56030 18002 56082
rect 18286 56030 18338 56082
rect 19518 56030 19570 56082
rect 23326 56030 23378 56082
rect 23662 56030 23714 56082
rect 25342 56030 25394 56082
rect 2494 55918 2546 55970
rect 3950 55918 4002 55970
rect 7422 55918 7474 55970
rect 8094 55918 8146 55970
rect 10334 55918 10386 55970
rect 16942 55918 16994 55970
rect 17614 55918 17666 55970
rect 19070 55918 19122 55970
rect 20190 55918 20242 55970
rect 22318 55918 22370 55970
rect 22766 55918 22818 55970
rect 23438 55918 23490 55970
rect 24334 55918 24386 55970
rect 26014 55918 26066 55970
rect 28142 55918 28194 55970
rect 10894 55806 10946 55858
rect 4616 55638 4668 55690
rect 4720 55638 4772 55690
rect 4824 55638 4876 55690
rect 11420 55638 11472 55690
rect 11524 55638 11576 55690
rect 11628 55638 11680 55690
rect 18224 55638 18276 55690
rect 18328 55638 18380 55690
rect 18432 55638 18484 55690
rect 25028 55638 25080 55690
rect 25132 55638 25184 55690
rect 25236 55638 25288 55690
rect 10222 55470 10274 55522
rect 11678 55470 11730 55522
rect 12462 55470 12514 55522
rect 13022 55470 13074 55522
rect 13582 55470 13634 55522
rect 4622 55358 4674 55410
rect 6638 55358 6690 55410
rect 7198 55358 7250 55410
rect 7982 55358 8034 55410
rect 8878 55358 8930 55410
rect 9438 55358 9490 55410
rect 12574 55358 12626 55410
rect 20302 55470 20354 55522
rect 14254 55358 14306 55410
rect 21422 55358 21474 55410
rect 23214 55358 23266 55410
rect 1822 55246 1874 55298
rect 14366 55246 14418 55298
rect 20078 55246 20130 55298
rect 21310 55246 21362 55298
rect 21870 55246 21922 55298
rect 22318 55246 22370 55298
rect 22878 55246 22930 55298
rect 25118 55246 25170 55298
rect 25566 55246 25618 55298
rect 26350 55246 26402 55298
rect 26798 55246 26850 55298
rect 27358 55246 27410 55298
rect 27694 55246 27746 55298
rect 2494 55134 2546 55186
rect 11230 55134 11282 55186
rect 11566 55134 11618 55186
rect 12014 55134 12066 55186
rect 17166 55134 17218 55186
rect 20526 55134 20578 55186
rect 20750 55134 20802 55186
rect 21646 55134 21698 55186
rect 25790 55134 25842 55186
rect 27246 55134 27298 55186
rect 5070 55022 5122 55074
rect 6078 55022 6130 55074
rect 7646 55022 7698 55074
rect 8430 55022 8482 55074
rect 9886 55022 9938 55074
rect 10222 55022 10274 55074
rect 10670 55022 10722 55074
rect 12910 55022 12962 55074
rect 13582 55022 13634 55074
rect 14030 55022 14082 55074
rect 19966 55022 20018 55074
rect 22206 55022 22258 55074
rect 22430 55022 22482 55074
rect 23662 55022 23714 55074
rect 24110 55022 24162 55074
rect 24558 55022 24610 55074
rect 25454 55022 25506 55074
rect 26238 55022 26290 55074
rect 26462 55022 26514 55074
rect 26574 55022 26626 55074
rect 27134 55022 27186 55074
rect 28142 55022 28194 55074
rect 8018 54854 8070 54906
rect 8122 54854 8174 54906
rect 8226 54854 8278 54906
rect 14822 54854 14874 54906
rect 14926 54854 14978 54906
rect 15030 54854 15082 54906
rect 21626 54854 21678 54906
rect 21730 54854 21782 54906
rect 21834 54854 21886 54906
rect 28430 54854 28482 54906
rect 28534 54854 28586 54906
rect 28638 54854 28690 54906
rect 2942 54686 2994 54738
rect 5294 54686 5346 54738
rect 5742 54686 5794 54738
rect 15374 54686 15426 54738
rect 22878 54686 22930 54738
rect 24222 54686 24274 54738
rect 24670 54686 24722 54738
rect 25790 54686 25842 54738
rect 2606 54574 2658 54626
rect 2830 54574 2882 54626
rect 3054 54574 3106 54626
rect 4398 54574 4450 54626
rect 12798 54574 12850 54626
rect 15822 54574 15874 54626
rect 19518 54574 19570 54626
rect 2158 54462 2210 54514
rect 3390 54462 3442 54514
rect 7310 54462 7362 54514
rect 9662 54462 9714 54514
rect 10334 54462 10386 54514
rect 13134 54462 13186 54514
rect 15262 54462 15314 54514
rect 20190 54462 20242 54514
rect 20974 54462 21026 54514
rect 21198 54462 21250 54514
rect 4958 54350 5010 54402
rect 6190 54350 6242 54402
rect 6638 54350 6690 54402
rect 6974 54350 7026 54402
rect 7086 54350 7138 54402
rect 8206 54350 8258 54402
rect 8542 54350 8594 54402
rect 9102 54350 9154 54402
rect 12462 54350 12514 54402
rect 13246 54350 13298 54402
rect 15038 54350 15090 54402
rect 17390 54350 17442 54402
rect 21982 54350 22034 54402
rect 22430 54350 22482 54402
rect 23326 54350 23378 54402
rect 23774 54350 23826 54402
rect 25342 54350 25394 54402
rect 26238 54350 26290 54402
rect 26686 54350 26738 54402
rect 27134 54350 27186 54402
rect 27582 54350 27634 54402
rect 28030 54350 28082 54402
rect 3278 54238 3330 54290
rect 5070 54238 5122 54290
rect 5630 54238 5682 54290
rect 21534 54238 21586 54290
rect 22766 54238 22818 54290
rect 24558 54238 24610 54290
rect 25118 54238 25170 54290
rect 25454 54238 25506 54290
rect 25790 54238 25842 54290
rect 26686 54238 26738 54290
rect 28142 54238 28194 54290
rect 4616 54070 4668 54122
rect 4720 54070 4772 54122
rect 4824 54070 4876 54122
rect 11420 54070 11472 54122
rect 11524 54070 11576 54122
rect 11628 54070 11680 54122
rect 18224 54070 18276 54122
rect 18328 54070 18380 54122
rect 18432 54070 18484 54122
rect 25028 54070 25080 54122
rect 25132 54070 25184 54122
rect 25236 54070 25288 54122
rect 18734 53902 18786 53954
rect 19070 53902 19122 53954
rect 3390 53790 3442 53842
rect 4734 53790 4786 53842
rect 8542 53790 8594 53842
rect 10222 53790 10274 53842
rect 10670 53790 10722 53842
rect 11790 53790 11842 53842
rect 12910 53790 12962 53842
rect 13918 53790 13970 53842
rect 16494 53790 16546 53842
rect 21646 53790 21698 53842
rect 24110 53790 24162 53842
rect 2494 53678 2546 53730
rect 3838 53678 3890 53730
rect 4398 53678 4450 53730
rect 4622 53678 4674 53730
rect 5630 53678 5682 53730
rect 8766 53678 8818 53730
rect 9102 53678 9154 53730
rect 10782 53678 10834 53730
rect 11118 53678 11170 53730
rect 11902 53678 11954 53730
rect 12574 53678 12626 53730
rect 16270 53678 16322 53730
rect 18398 53678 18450 53730
rect 19630 53678 19682 53730
rect 20078 53678 20130 53730
rect 20302 53678 20354 53730
rect 20638 53678 20690 53730
rect 21534 53678 21586 53730
rect 21758 53678 21810 53730
rect 23102 53678 23154 53730
rect 23326 53678 23378 53730
rect 25790 53678 25842 53730
rect 26350 53678 26402 53730
rect 26798 53678 26850 53730
rect 27246 53678 27298 53730
rect 1710 53566 1762 53618
rect 2830 53566 2882 53618
rect 4174 53566 4226 53618
rect 6414 53566 6466 53618
rect 9438 53566 9490 53618
rect 10558 53566 10610 53618
rect 15262 53566 15314 53618
rect 18510 53566 18562 53618
rect 20526 53566 20578 53618
rect 22206 53566 22258 53618
rect 22766 53566 22818 53618
rect 23774 53566 23826 53618
rect 23998 53566 24050 53618
rect 26126 53566 26178 53618
rect 26686 53566 26738 53618
rect 27694 53566 27746 53618
rect 2046 53454 2098 53506
rect 4734 53454 4786 53506
rect 8990 53454 9042 53506
rect 11678 53454 11730 53506
rect 12126 53454 12178 53506
rect 12798 53454 12850 53506
rect 14366 53454 14418 53506
rect 18958 53454 19010 53506
rect 19406 53454 19458 53506
rect 21982 53454 22034 53506
rect 22990 53454 23042 53506
rect 24222 53454 24274 53506
rect 24670 53454 24722 53506
rect 25118 53454 25170 53506
rect 26014 53454 26066 53506
rect 26910 53454 26962 53506
rect 28142 53454 28194 53506
rect 8018 53286 8070 53338
rect 8122 53286 8174 53338
rect 8226 53286 8278 53338
rect 14822 53286 14874 53338
rect 14926 53286 14978 53338
rect 15030 53286 15082 53338
rect 21626 53286 21678 53338
rect 21730 53286 21782 53338
rect 21834 53286 21886 53338
rect 28430 53286 28482 53338
rect 28534 53286 28586 53338
rect 28638 53286 28690 53338
rect 2494 53118 2546 53170
rect 3278 53118 3330 53170
rect 3838 53118 3890 53170
rect 4286 53118 4338 53170
rect 4510 53118 4562 53170
rect 4622 53118 4674 53170
rect 5294 53118 5346 53170
rect 5518 53118 5570 53170
rect 5630 53118 5682 53170
rect 6414 53118 6466 53170
rect 8654 53118 8706 53170
rect 9102 53118 9154 53170
rect 9774 53118 9826 53170
rect 11230 53118 11282 53170
rect 19742 53118 19794 53170
rect 21310 53118 21362 53170
rect 6078 53006 6130 53058
rect 6302 53006 6354 53058
rect 9662 53006 9714 53058
rect 11902 53006 11954 53058
rect 12126 53006 12178 53058
rect 13694 53006 13746 53058
rect 15710 53006 15762 53058
rect 17950 53006 18002 53058
rect 20526 53006 20578 53058
rect 20638 53006 20690 53058
rect 23886 53006 23938 53058
rect 26014 53006 26066 53058
rect 4062 52894 4114 52946
rect 5070 52894 5122 52946
rect 6638 52894 6690 52946
rect 9886 52894 9938 52946
rect 10222 52894 10274 52946
rect 12574 52894 12626 52946
rect 14814 52894 14866 52946
rect 15150 52894 15202 52946
rect 17390 52894 17442 52946
rect 20302 52894 20354 52946
rect 21086 52894 21138 52946
rect 24558 52894 24610 52946
rect 25230 52894 25282 52946
rect 2158 52782 2210 52834
rect 2606 52782 2658 52834
rect 4622 52782 4674 52834
rect 5630 52782 5682 52834
rect 7646 52782 7698 52834
rect 8094 52782 8146 52834
rect 10894 52782 10946 52834
rect 12798 52782 12850 52834
rect 13582 52782 13634 52834
rect 19182 52782 19234 52834
rect 21758 52782 21810 52834
rect 28142 52782 28194 52834
rect 2718 52670 2770 52722
rect 6638 52670 6690 52722
rect 8206 52670 8258 52722
rect 8990 52670 9042 52722
rect 10446 52670 10498 52722
rect 11342 52670 11394 52722
rect 4616 52502 4668 52554
rect 4720 52502 4772 52554
rect 4824 52502 4876 52554
rect 11420 52502 11472 52554
rect 11524 52502 11576 52554
rect 11628 52502 11680 52554
rect 18224 52502 18276 52554
rect 18328 52502 18380 52554
rect 18432 52502 18484 52554
rect 25028 52502 25080 52554
rect 25132 52502 25184 52554
rect 25236 52502 25288 52554
rect 5966 52334 6018 52386
rect 6526 52334 6578 52386
rect 10670 52334 10722 52386
rect 11006 52334 11058 52386
rect 20750 52334 20802 52386
rect 21870 52334 21922 52386
rect 2830 52222 2882 52274
rect 3390 52222 3442 52274
rect 5854 52222 5906 52274
rect 6750 52222 6802 52274
rect 7086 52222 7138 52274
rect 8206 52222 8258 52274
rect 10334 52222 10386 52274
rect 11230 52222 11282 52274
rect 13022 52222 13074 52274
rect 14142 52222 14194 52274
rect 19742 52222 19794 52274
rect 23886 52222 23938 52274
rect 24334 52222 24386 52274
rect 24782 52222 24834 52274
rect 26238 52222 26290 52274
rect 27470 52222 27522 52274
rect 2494 52110 2546 52162
rect 3726 52110 3778 52162
rect 4174 52110 4226 52162
rect 4286 52110 4338 52162
rect 4734 52110 4786 52162
rect 7534 52110 7586 52162
rect 12014 52110 12066 52162
rect 12126 52110 12178 52162
rect 14030 52110 14082 52162
rect 15598 52110 15650 52162
rect 17614 52110 17666 52162
rect 19966 52110 20018 52162
rect 20078 52110 20130 52162
rect 20526 52110 20578 52162
rect 21534 52110 21586 52162
rect 21870 52110 21922 52162
rect 22430 52110 22482 52162
rect 22766 52110 22818 52162
rect 22990 52110 23042 52162
rect 25230 52110 25282 52162
rect 26350 52110 26402 52162
rect 26798 52110 26850 52162
rect 27134 52110 27186 52162
rect 2270 51998 2322 52050
rect 6190 51998 6242 52050
rect 12350 51998 12402 52050
rect 15038 51998 15090 52050
rect 16718 51998 16770 52050
rect 18174 51998 18226 52050
rect 21310 51998 21362 52050
rect 26238 51998 26290 52050
rect 26574 51998 26626 52050
rect 27582 51998 27634 52050
rect 27806 51998 27858 52050
rect 4398 51886 4450 51938
rect 4510 51886 4562 51938
rect 17726 51886 17778 51938
rect 21646 51886 21698 51938
rect 23438 51886 23490 51938
rect 25678 51886 25730 51938
rect 27358 51886 27410 51938
rect 8018 51718 8070 51770
rect 8122 51718 8174 51770
rect 8226 51718 8278 51770
rect 14822 51718 14874 51770
rect 14926 51718 14978 51770
rect 15030 51718 15082 51770
rect 21626 51718 21678 51770
rect 21730 51718 21782 51770
rect 21834 51718 21886 51770
rect 28430 51718 28482 51770
rect 28534 51718 28586 51770
rect 28638 51718 28690 51770
rect 2494 51550 2546 51602
rect 4734 51550 4786 51602
rect 5630 51550 5682 51602
rect 7310 51550 7362 51602
rect 7758 51550 7810 51602
rect 8990 51550 9042 51602
rect 16830 51550 16882 51602
rect 17502 51550 17554 51602
rect 19406 51550 19458 51602
rect 19742 51550 19794 51602
rect 23214 51550 23266 51602
rect 24334 51550 24386 51602
rect 27694 51550 27746 51602
rect 4062 51438 4114 51490
rect 5182 51438 5234 51490
rect 5854 51438 5906 51490
rect 10110 51438 10162 51490
rect 18622 51438 18674 51490
rect 18734 51438 18786 51490
rect 20862 51438 20914 51490
rect 23326 51438 23378 51490
rect 25790 51438 25842 51490
rect 26238 51438 26290 51490
rect 3614 51326 3666 51378
rect 6190 51326 6242 51378
rect 6414 51326 6466 51378
rect 8430 51326 8482 51378
rect 8766 51326 8818 51378
rect 13470 51326 13522 51378
rect 16158 51326 16210 51378
rect 16270 51326 16322 51378
rect 18398 51326 18450 51378
rect 19182 51326 19234 51378
rect 20190 51326 20242 51378
rect 23550 51326 23602 51378
rect 23886 51326 23938 51378
rect 24110 51326 24162 51378
rect 26462 51326 26514 51378
rect 26798 51326 26850 51378
rect 2046 51214 2098 51266
rect 3950 51214 4002 51266
rect 5966 51214 6018 51266
rect 8206 51214 8258 51266
rect 8878 51214 8930 51266
rect 15374 51214 15426 51266
rect 17950 51214 18002 51266
rect 22990 51214 23042 51266
rect 25342 51214 25394 51266
rect 26350 51214 26402 51266
rect 27246 51214 27298 51266
rect 28142 51214 28194 51266
rect 2382 51102 2434 51154
rect 2718 51102 2770 51154
rect 3838 51102 3890 51154
rect 15934 51102 15986 51154
rect 24446 51102 24498 51154
rect 27358 51102 27410 51154
rect 28030 51102 28082 51154
rect 4616 50934 4668 50986
rect 4720 50934 4772 50986
rect 4824 50934 4876 50986
rect 11420 50934 11472 50986
rect 11524 50934 11576 50986
rect 11628 50934 11680 50986
rect 18224 50934 18276 50986
rect 18328 50934 18380 50986
rect 18432 50934 18484 50986
rect 25028 50934 25080 50986
rect 25132 50934 25184 50986
rect 25236 50934 25288 50986
rect 20190 50766 20242 50818
rect 20750 50766 20802 50818
rect 22318 50766 22370 50818
rect 4622 50654 4674 50706
rect 5182 50654 5234 50706
rect 6526 50654 6578 50706
rect 10222 50654 10274 50706
rect 10670 50654 10722 50706
rect 11118 50654 11170 50706
rect 19630 50654 19682 50706
rect 24334 50654 24386 50706
rect 27806 50654 27858 50706
rect 1822 50542 1874 50594
rect 6190 50542 6242 50594
rect 6414 50542 6466 50594
rect 6638 50542 6690 50594
rect 7310 50542 7362 50594
rect 11454 50542 11506 50594
rect 12686 50542 12738 50594
rect 13582 50542 13634 50594
rect 15374 50542 15426 50594
rect 17390 50542 17442 50594
rect 21422 50542 21474 50594
rect 24894 50542 24946 50594
rect 12462 50486 12514 50538
rect 2494 50430 2546 50482
rect 6862 50430 6914 50482
rect 8094 50430 8146 50482
rect 11566 50430 11618 50482
rect 13022 50430 13074 50482
rect 14814 50430 14866 50482
rect 15038 50430 15090 50482
rect 16494 50430 16546 50482
rect 19182 50430 19234 50482
rect 25678 50430 25730 50482
rect 15598 50318 15650 50370
rect 20078 50318 20130 50370
rect 20526 50318 20578 50370
rect 8018 50150 8070 50202
rect 8122 50150 8174 50202
rect 8226 50150 8278 50202
rect 14822 50150 14874 50202
rect 14926 50150 14978 50202
rect 15030 50150 15082 50202
rect 21626 50150 21678 50202
rect 21730 50150 21782 50202
rect 21834 50150 21886 50202
rect 28430 50150 28482 50202
rect 28534 50150 28586 50202
rect 28638 50150 28690 50202
rect 3166 49982 3218 50034
rect 8094 49982 8146 50034
rect 8542 49982 8594 50034
rect 9998 49982 10050 50034
rect 11006 49982 11058 50034
rect 16718 49982 16770 50034
rect 25678 49982 25730 50034
rect 2046 49870 2098 49922
rect 2830 49870 2882 49922
rect 5294 49870 5346 49922
rect 9550 49870 9602 49922
rect 10558 49870 10610 49922
rect 12238 49870 12290 49922
rect 13582 49870 13634 49922
rect 16830 49870 16882 49922
rect 18510 49870 18562 49922
rect 19966 49870 20018 49922
rect 26126 49870 26178 49922
rect 1710 49758 1762 49810
rect 3166 49758 3218 49810
rect 3390 49758 3442 49810
rect 4622 49758 4674 49810
rect 8430 49758 8482 49810
rect 8654 49758 8706 49810
rect 8878 49758 8930 49810
rect 9774 49758 9826 49810
rect 10110 49758 10162 49810
rect 10782 49758 10834 49810
rect 11230 49758 11282 49810
rect 12462 49758 12514 49810
rect 12686 49758 12738 49810
rect 13022 49758 13074 49810
rect 15150 49758 15202 49810
rect 18958 49758 19010 49810
rect 19518 49758 19570 49810
rect 21870 49758 21922 49810
rect 25566 49758 25618 49810
rect 25902 49758 25954 49810
rect 2494 49646 2546 49698
rect 4174 49646 4226 49698
rect 7422 49646 7474 49698
rect 9886 49646 9938 49698
rect 11006 49646 11058 49698
rect 19742 49646 19794 49698
rect 22542 49646 22594 49698
rect 24670 49646 24722 49698
rect 26574 49646 26626 49698
rect 27022 49646 27074 49698
rect 27470 49646 27522 49698
rect 27918 49646 27970 49698
rect 3390 49534 3442 49586
rect 11902 49534 11954 49586
rect 26910 49534 26962 49586
rect 27918 49534 27970 49586
rect 4616 49366 4668 49418
rect 4720 49366 4772 49418
rect 4824 49366 4876 49418
rect 11420 49366 11472 49418
rect 11524 49366 11576 49418
rect 11628 49366 11680 49418
rect 18224 49366 18276 49418
rect 18328 49366 18380 49418
rect 18432 49366 18484 49418
rect 25028 49366 25080 49418
rect 25132 49366 25184 49418
rect 25236 49366 25288 49418
rect 7422 49198 7474 49250
rect 8206 49198 8258 49250
rect 13582 49198 13634 49250
rect 23886 49198 23938 49250
rect 25230 49198 25282 49250
rect 1822 49086 1874 49138
rect 2606 49086 2658 49138
rect 5630 49086 5682 49138
rect 6526 49086 6578 49138
rect 6862 49086 6914 49138
rect 7422 49086 7474 49138
rect 7870 49086 7922 49138
rect 8206 49086 8258 49138
rect 8654 49086 8706 49138
rect 9102 49086 9154 49138
rect 9550 49086 9602 49138
rect 10894 49086 10946 49138
rect 11342 49086 11394 49138
rect 15374 49086 15426 49138
rect 21422 49086 21474 49138
rect 23438 49086 23490 49138
rect 27134 49086 27186 49138
rect 27582 49086 27634 49138
rect 3614 48974 3666 49026
rect 3950 48974 4002 49026
rect 11790 48974 11842 49026
rect 12126 48974 12178 49026
rect 12350 48974 12402 49026
rect 13918 48974 13970 49026
rect 14142 48974 14194 49026
rect 15934 48974 15986 49026
rect 18622 48974 18674 49026
rect 18958 48974 19010 49026
rect 21870 48974 21922 49026
rect 23662 48974 23714 49026
rect 24110 48974 24162 49026
rect 24670 48974 24722 49026
rect 25230 48974 25282 49026
rect 26014 48974 26066 49026
rect 26350 48974 26402 49026
rect 12574 48862 12626 48914
rect 14366 48862 14418 48914
rect 14590 48862 14642 48914
rect 14926 48862 14978 48914
rect 17054 48862 17106 48914
rect 18846 48862 18898 48914
rect 20638 48862 20690 48914
rect 23326 48862 23378 48914
rect 24446 48862 24498 48914
rect 24894 48862 24946 48914
rect 25566 48862 25618 48914
rect 26686 48862 26738 48914
rect 2942 48750 2994 48802
rect 4062 48750 4114 48802
rect 4174 48750 4226 48802
rect 4958 48750 5010 48802
rect 5742 48750 5794 48802
rect 9998 48750 10050 48802
rect 10558 48750 10610 48802
rect 24334 48750 24386 48802
rect 26238 48750 26290 48802
rect 28030 48750 28082 48802
rect 8018 48582 8070 48634
rect 8122 48582 8174 48634
rect 8226 48582 8278 48634
rect 14822 48582 14874 48634
rect 14926 48582 14978 48634
rect 15030 48582 15082 48634
rect 21626 48582 21678 48634
rect 21730 48582 21782 48634
rect 21834 48582 21886 48634
rect 28430 48582 28482 48634
rect 28534 48582 28586 48634
rect 28638 48582 28690 48634
rect 6190 48414 6242 48466
rect 7534 48414 7586 48466
rect 9550 48414 9602 48466
rect 9998 48414 10050 48466
rect 11790 48414 11842 48466
rect 12238 48414 12290 48466
rect 12686 48414 12738 48466
rect 16606 48414 16658 48466
rect 5854 48302 5906 48354
rect 11342 48302 11394 48354
rect 14142 48302 14194 48354
rect 16830 48302 16882 48354
rect 17502 48302 17554 48354
rect 20526 48302 20578 48354
rect 22094 48302 22146 48354
rect 26014 48302 26066 48354
rect 1822 48190 1874 48242
rect 5294 48190 5346 48242
rect 8318 48190 8370 48242
rect 8542 48190 8594 48242
rect 8878 48190 8930 48242
rect 9774 48190 9826 48242
rect 14590 48190 14642 48242
rect 15038 48190 15090 48242
rect 17390 48190 17442 48242
rect 19518 48190 19570 48242
rect 21646 48190 21698 48242
rect 25342 48190 25394 48242
rect 2494 48078 2546 48130
rect 4622 48078 4674 48130
rect 6638 48078 6690 48130
rect 7086 48078 7138 48130
rect 8094 48078 8146 48130
rect 8430 48078 8482 48130
rect 9662 48078 9714 48130
rect 10782 48078 10834 48130
rect 19966 48078 20018 48130
rect 23326 48078 23378 48130
rect 23438 48078 23490 48130
rect 24558 48078 24610 48130
rect 28142 48078 28194 48130
rect 4958 47966 5010 48018
rect 5294 47966 5346 48018
rect 6078 47966 6130 48018
rect 6638 47966 6690 48018
rect 11790 47966 11842 48018
rect 12126 47966 12178 48018
rect 4616 47798 4668 47850
rect 4720 47798 4772 47850
rect 4824 47798 4876 47850
rect 11420 47798 11472 47850
rect 11524 47798 11576 47850
rect 11628 47798 11680 47850
rect 18224 47798 18276 47850
rect 18328 47798 18380 47850
rect 18432 47798 18484 47850
rect 25028 47798 25080 47850
rect 25132 47798 25184 47850
rect 25236 47798 25288 47850
rect 3502 47630 3554 47682
rect 11006 47630 11058 47682
rect 11566 47630 11618 47682
rect 20862 47630 20914 47682
rect 21310 47630 21362 47682
rect 2494 47518 2546 47570
rect 3054 47518 3106 47570
rect 4286 47518 4338 47570
rect 4734 47518 4786 47570
rect 7422 47518 7474 47570
rect 9550 47518 9602 47570
rect 10334 47518 10386 47570
rect 11230 47518 11282 47570
rect 11566 47518 11618 47570
rect 12462 47518 12514 47570
rect 19518 47518 19570 47570
rect 20078 47518 20130 47570
rect 21646 47518 21698 47570
rect 26350 47518 26402 47570
rect 26798 47518 26850 47570
rect 27246 47518 27298 47570
rect 28030 47630 28082 47682
rect 27694 47518 27746 47570
rect 28142 47518 28194 47570
rect 2942 47406 2994 47458
rect 3166 47406 3218 47458
rect 3502 47406 3554 47458
rect 5742 47406 5794 47458
rect 6750 47406 6802 47458
rect 10222 47406 10274 47458
rect 10558 47406 10610 47458
rect 13918 47406 13970 47458
rect 14142 47406 14194 47458
rect 14702 47406 14754 47458
rect 15262 47406 15314 47458
rect 18958 47406 19010 47458
rect 21870 47406 21922 47458
rect 23550 47406 23602 47458
rect 26686 47406 26738 47458
rect 1710 47294 1762 47346
rect 9998 47294 10050 47346
rect 10446 47294 10498 47346
rect 14366 47294 14418 47346
rect 16382 47294 16434 47346
rect 17054 47294 17106 47346
rect 18398 47294 18450 47346
rect 20302 47294 20354 47346
rect 22318 47294 22370 47346
rect 22766 47294 22818 47346
rect 24222 47294 24274 47346
rect 26910 47294 26962 47346
rect 2046 47182 2098 47234
rect 5854 47182 5906 47234
rect 12014 47182 12066 47234
rect 12910 47182 12962 47234
rect 13582 47182 13634 47234
rect 20526 47182 20578 47234
rect 20750 47182 20802 47234
rect 27134 47182 27186 47234
rect 8018 47014 8070 47066
rect 8122 47014 8174 47066
rect 8226 47014 8278 47066
rect 14822 47014 14874 47066
rect 14926 47014 14978 47066
rect 15030 47014 15082 47066
rect 21626 47014 21678 47066
rect 21730 47014 21782 47066
rect 21834 47014 21886 47066
rect 28430 47014 28482 47066
rect 28534 47014 28586 47066
rect 28638 47014 28690 47066
rect 4062 46846 4114 46898
rect 5070 46846 5122 46898
rect 9998 46846 10050 46898
rect 13918 46846 13970 46898
rect 15262 46846 15314 46898
rect 18958 46846 19010 46898
rect 21646 46846 21698 46898
rect 22878 46846 22930 46898
rect 24222 46846 24274 46898
rect 25454 46846 25506 46898
rect 26686 46846 26738 46898
rect 27134 46846 27186 46898
rect 28142 46846 28194 46898
rect 2046 46734 2098 46786
rect 4846 46734 4898 46786
rect 16270 46734 16322 46786
rect 17950 46734 18002 46786
rect 22094 46734 22146 46786
rect 1710 46622 1762 46674
rect 5518 46622 5570 46674
rect 10334 46622 10386 46674
rect 15038 46622 15090 46674
rect 15262 46622 15314 46674
rect 17390 46622 17442 46674
rect 20302 46622 20354 46674
rect 20526 46622 20578 46674
rect 20862 46622 20914 46674
rect 21198 46622 21250 46674
rect 21422 46622 21474 46674
rect 23102 46622 23154 46674
rect 23326 46622 23378 46674
rect 23886 46622 23938 46674
rect 24334 46622 24386 46674
rect 24558 46622 24610 46674
rect 25230 46622 25282 46674
rect 25342 46622 25394 46674
rect 25790 46622 25842 46674
rect 2718 46510 2770 46562
rect 3166 46510 3218 46562
rect 3614 46510 3666 46562
rect 4510 46510 4562 46562
rect 6302 46510 6354 46562
rect 8430 46510 8482 46562
rect 8990 46510 9042 46562
rect 11118 46510 11170 46562
rect 13246 46510 13298 46562
rect 19182 46510 19234 46562
rect 20414 46510 20466 46562
rect 21534 46510 21586 46562
rect 23214 46510 23266 46562
rect 26238 46510 26290 46562
rect 27582 46510 27634 46562
rect 5182 46398 5234 46450
rect 4616 46230 4668 46282
rect 4720 46230 4772 46282
rect 4824 46230 4876 46282
rect 11420 46230 11472 46282
rect 11524 46230 11576 46282
rect 11628 46230 11680 46282
rect 18224 46230 18276 46282
rect 18328 46230 18380 46282
rect 18432 46230 18484 46282
rect 25028 46230 25080 46282
rect 25132 46230 25184 46282
rect 25236 46230 25288 46282
rect 9438 46062 9490 46114
rect 9998 46062 10050 46114
rect 10334 46062 10386 46114
rect 10782 46062 10834 46114
rect 4622 45950 4674 46002
rect 6862 45950 6914 46002
rect 8990 45950 9042 46002
rect 10334 45950 10386 46002
rect 10782 45950 10834 46002
rect 24222 45950 24274 46002
rect 25118 45950 25170 46002
rect 26574 45950 26626 46002
rect 1822 45838 1874 45890
rect 7310 45838 7362 45890
rect 7870 45838 7922 45890
rect 7982 45838 8034 45890
rect 8318 45838 8370 45890
rect 9438 45838 9490 45890
rect 11230 45838 11282 45890
rect 14366 45838 14418 45890
rect 15822 45838 15874 45890
rect 17838 45838 17890 45890
rect 18286 45838 18338 45890
rect 21310 45838 21362 45890
rect 27806 45838 27858 45890
rect 2494 45726 2546 45778
rect 6414 45726 6466 45778
rect 6750 45726 6802 45778
rect 7086 45726 7138 45778
rect 11118 45726 11170 45778
rect 11454 45726 11506 45778
rect 11678 45726 11730 45778
rect 12238 45726 12290 45778
rect 16270 45726 16322 45778
rect 19294 45726 19346 45778
rect 22094 45726 22146 45778
rect 5182 45614 5234 45666
rect 6078 45614 6130 45666
rect 7758 45614 7810 45666
rect 9886 45614 9938 45666
rect 12126 45614 12178 45666
rect 12350 45614 12402 45666
rect 12574 45614 12626 45666
rect 13806 45614 13858 45666
rect 14702 45614 14754 45666
rect 17166 45614 17218 45666
rect 20414 45614 20466 45666
rect 24670 45614 24722 45666
rect 8018 45446 8070 45498
rect 8122 45446 8174 45498
rect 8226 45446 8278 45498
rect 14822 45446 14874 45498
rect 14926 45446 14978 45498
rect 15030 45446 15082 45498
rect 21626 45446 21678 45498
rect 21730 45446 21782 45498
rect 21834 45446 21886 45498
rect 28430 45446 28482 45498
rect 28534 45446 28586 45498
rect 28638 45446 28690 45498
rect 2606 45278 2658 45330
rect 4286 45278 4338 45330
rect 5182 45278 5234 45330
rect 5742 45278 5794 45330
rect 11454 45278 11506 45330
rect 11902 45278 11954 45330
rect 12798 45278 12850 45330
rect 15934 45278 15986 45330
rect 17502 45278 17554 45330
rect 22206 45278 22258 45330
rect 23214 45278 23266 45330
rect 23662 45278 23714 45330
rect 23998 45278 24050 45330
rect 7646 45166 7698 45218
rect 9550 45166 9602 45218
rect 13918 45166 13970 45218
rect 14030 45166 14082 45218
rect 14366 45166 14418 45218
rect 14814 45166 14866 45218
rect 15486 45166 15538 45218
rect 16830 45166 16882 45218
rect 22094 45166 22146 45218
rect 22430 45166 22482 45218
rect 22654 45166 22706 45218
rect 2270 45054 2322 45106
rect 2830 45054 2882 45106
rect 3054 45054 3106 45106
rect 3502 45054 3554 45106
rect 9102 45054 9154 45106
rect 9774 45054 9826 45106
rect 9998 45054 10050 45106
rect 10110 45054 10162 45106
rect 13470 45054 13522 45106
rect 13694 45054 13746 45106
rect 15262 45054 15314 45106
rect 16158 45054 16210 45106
rect 16382 45054 16434 45106
rect 16606 45054 16658 45106
rect 21198 45054 21250 45106
rect 28142 45054 28194 45106
rect 2046 44942 2098 44994
rect 3390 44942 3442 44994
rect 4846 44942 4898 44994
rect 6190 44942 6242 44994
rect 6750 44942 6802 44994
rect 7198 44942 7250 44994
rect 7982 44942 8034 44994
rect 8542 44942 8594 44994
rect 9886 44942 9938 44994
rect 11006 44942 11058 44994
rect 12350 44942 12402 44994
rect 13246 44942 13298 44994
rect 16270 44942 16322 44994
rect 17950 44942 18002 44994
rect 18398 44942 18450 44994
rect 20526 44942 20578 44994
rect 21758 44942 21810 44994
rect 24446 44942 24498 44994
rect 25230 44942 25282 44994
rect 27358 44942 27410 44994
rect 2494 44830 2546 44882
rect 6190 44830 6242 44882
rect 7758 44830 7810 44882
rect 8542 44830 8594 44882
rect 8878 44830 8930 44882
rect 11902 44830 11954 44882
rect 12350 44830 12402 44882
rect 13246 44830 13298 44882
rect 4616 44662 4668 44714
rect 4720 44662 4772 44714
rect 4824 44662 4876 44714
rect 11420 44662 11472 44714
rect 11524 44662 11576 44714
rect 11628 44662 11680 44714
rect 18224 44662 18276 44714
rect 18328 44662 18380 44714
rect 18432 44662 18484 44714
rect 25028 44662 25080 44714
rect 25132 44662 25184 44714
rect 25236 44662 25288 44714
rect 2270 44494 2322 44546
rect 3166 44494 3218 44546
rect 6190 44494 6242 44546
rect 9438 44494 9490 44546
rect 9998 44494 10050 44546
rect 2494 44382 2546 44434
rect 3726 44382 3778 44434
rect 8430 44382 8482 44434
rect 9662 44382 9714 44434
rect 10110 44382 10162 44434
rect 15262 44382 15314 44434
rect 26798 44382 26850 44434
rect 6414 44270 6466 44322
rect 6750 44270 6802 44322
rect 6862 44270 6914 44322
rect 7758 44270 7810 44322
rect 8654 44270 8706 44322
rect 10446 44270 10498 44322
rect 10670 44270 10722 44322
rect 12238 44270 12290 44322
rect 12574 44270 12626 44322
rect 13470 44270 13522 44322
rect 13582 44270 13634 44322
rect 14702 44270 14754 44322
rect 14926 44270 14978 44322
rect 15374 44270 15426 44322
rect 17502 44270 17554 44322
rect 19630 44270 19682 44322
rect 20190 44270 20242 44322
rect 20414 44270 20466 44322
rect 21422 44270 21474 44322
rect 23774 44270 23826 44322
rect 3390 44158 3442 44210
rect 4510 44158 4562 44210
rect 5630 44158 5682 44210
rect 5854 44158 5906 44210
rect 7870 44158 7922 44210
rect 8990 44158 9042 44210
rect 12014 44158 12066 44210
rect 15822 44158 15874 44210
rect 19518 44158 19570 44210
rect 19966 44158 20018 44210
rect 21198 44158 21250 44210
rect 21758 44158 21810 44210
rect 22318 44158 22370 44210
rect 2158 44046 2210 44098
rect 3054 44046 3106 44098
rect 3838 44046 3890 44098
rect 4398 44046 4450 44098
rect 5182 44046 5234 44098
rect 5742 44046 5794 44098
rect 6974 44046 7026 44098
rect 10782 44046 10834 44098
rect 10894 44046 10946 44098
rect 11006 44046 11058 44098
rect 11790 44046 11842 44098
rect 12126 44046 12178 44098
rect 13694 44046 13746 44098
rect 13918 44046 13970 44098
rect 15150 44046 15202 44098
rect 16046 44046 16098 44098
rect 20190 44046 20242 44098
rect 8018 43878 8070 43930
rect 8122 43878 8174 43930
rect 8226 43878 8278 43930
rect 14822 43878 14874 43930
rect 14926 43878 14978 43930
rect 15030 43878 15082 43930
rect 21626 43878 21678 43930
rect 21730 43878 21782 43930
rect 21834 43878 21886 43930
rect 28430 43878 28482 43930
rect 28534 43878 28586 43930
rect 28638 43878 28690 43930
rect 2158 43710 2210 43762
rect 19182 43710 19234 43762
rect 20190 43710 20242 43762
rect 22094 43710 22146 43762
rect 23438 43710 23490 43762
rect 25790 43710 25842 43762
rect 26462 43710 26514 43762
rect 2494 43598 2546 43650
rect 5406 43598 5458 43650
rect 10110 43598 10162 43650
rect 10446 43598 10498 43650
rect 11006 43598 11058 43650
rect 12126 43598 12178 43650
rect 17614 43598 17666 43650
rect 18846 43598 18898 43650
rect 19406 43598 19458 43650
rect 21310 43598 21362 43650
rect 23102 43598 23154 43650
rect 27358 43598 27410 43650
rect 28142 43598 28194 43650
rect 2830 43486 2882 43538
rect 4846 43486 4898 43538
rect 10782 43486 10834 43538
rect 11342 43486 11394 43538
rect 15038 43486 15090 43538
rect 15598 43486 15650 43538
rect 15934 43486 15986 43538
rect 16158 43486 16210 43538
rect 16830 43486 16882 43538
rect 17838 43486 17890 43538
rect 18510 43486 18562 43538
rect 19294 43486 19346 43538
rect 19742 43486 19794 43538
rect 23998 43486 24050 43538
rect 24222 43486 24274 43538
rect 24558 43486 24610 43538
rect 26238 43486 26290 43538
rect 26574 43486 26626 43538
rect 26798 43486 26850 43538
rect 27134 43486 27186 43538
rect 27246 43486 27298 43538
rect 27806 43486 27858 43538
rect 2606 43374 2658 43426
rect 9662 43374 9714 43426
rect 9998 43374 10050 43426
rect 14254 43374 14306 43426
rect 15710 43374 15762 43426
rect 16606 43374 16658 43426
rect 18174 43374 18226 43426
rect 20638 43374 20690 43426
rect 21646 43374 21698 43426
rect 22542 43374 22594 43426
rect 24110 43374 24162 43426
rect 16494 43262 16546 43314
rect 19966 43262 20018 43314
rect 20862 43262 20914 43314
rect 22318 43262 22370 43314
rect 23438 43262 23490 43314
rect 25566 43262 25618 43314
rect 25902 43262 25954 43314
rect 4616 43094 4668 43146
rect 4720 43094 4772 43146
rect 4824 43094 4876 43146
rect 11420 43094 11472 43146
rect 11524 43094 11576 43146
rect 11628 43094 11680 43146
rect 18224 43094 18276 43146
rect 18328 43094 18380 43146
rect 18432 43094 18484 43146
rect 25028 43094 25080 43146
rect 25132 43094 25184 43146
rect 25236 43094 25288 43146
rect 19294 42926 19346 42978
rect 4622 42814 4674 42866
rect 5070 42814 5122 42866
rect 6078 42814 6130 42866
rect 7198 42814 7250 42866
rect 9326 42814 9378 42866
rect 10782 42814 10834 42866
rect 12014 42814 12066 42866
rect 12910 42814 12962 42866
rect 13918 42814 13970 42866
rect 15822 42814 15874 42866
rect 17950 42814 18002 42866
rect 18622 42814 18674 42866
rect 21310 42814 21362 42866
rect 24558 42814 24610 42866
rect 27918 42814 27970 42866
rect 1822 42702 1874 42754
rect 6526 42702 6578 42754
rect 9662 42702 9714 42754
rect 15150 42702 15202 42754
rect 19518 42702 19570 42754
rect 20078 42702 20130 42754
rect 20302 42702 20354 42754
rect 20750 42702 20802 42754
rect 24110 42702 24162 42754
rect 27470 42702 27522 42754
rect 2494 42590 2546 42642
rect 9998 42590 10050 42642
rect 10446 42590 10498 42642
rect 14590 42590 14642 42642
rect 18286 42590 18338 42642
rect 18846 42590 18898 42642
rect 19966 42590 20018 42642
rect 23438 42590 23490 42642
rect 26686 42590 26738 42642
rect 9886 42478 9938 42530
rect 10670 42478 10722 42530
rect 10894 42478 10946 42530
rect 11006 42478 11058 42530
rect 11566 42478 11618 42530
rect 12462 42478 12514 42530
rect 14142 42478 14194 42530
rect 14254 42478 14306 42530
rect 14366 42478 14418 42530
rect 18510 42478 18562 42530
rect 18734 42478 18786 42530
rect 8018 42310 8070 42362
rect 8122 42310 8174 42362
rect 8226 42310 8278 42362
rect 14822 42310 14874 42362
rect 14926 42310 14978 42362
rect 15030 42310 15082 42362
rect 21626 42310 21678 42362
rect 21730 42310 21782 42362
rect 21834 42310 21886 42362
rect 28430 42310 28482 42362
rect 28534 42310 28586 42362
rect 28638 42310 28690 42362
rect 2494 42142 2546 42194
rect 8542 42142 8594 42194
rect 11230 42142 11282 42194
rect 19182 42142 19234 42194
rect 21870 42142 21922 42194
rect 23102 42142 23154 42194
rect 23886 42142 23938 42194
rect 2046 42030 2098 42082
rect 3054 42030 3106 42082
rect 3278 42030 3330 42082
rect 10558 42030 10610 42082
rect 11678 42030 11730 42082
rect 15710 42030 15762 42082
rect 19294 42030 19346 42082
rect 19406 42030 19458 42082
rect 22542 42030 22594 42082
rect 24222 42030 24274 42082
rect 1710 41918 1762 41970
rect 2718 41918 2770 41970
rect 3726 41918 3778 41970
rect 4174 41918 4226 41970
rect 4846 41918 4898 41970
rect 7758 41918 7810 41970
rect 8094 41918 8146 41970
rect 8206 41918 8258 41970
rect 8542 41918 8594 41970
rect 8990 41918 9042 41970
rect 10222 41918 10274 41970
rect 10334 41918 10386 41970
rect 10782 41918 10834 41970
rect 12350 41918 12402 41970
rect 15934 41918 15986 41970
rect 16494 41918 16546 41970
rect 17502 41918 17554 41970
rect 17614 41918 17666 41970
rect 17726 41918 17778 41970
rect 18174 41918 18226 41970
rect 18398 41918 18450 41970
rect 19070 41918 19122 41970
rect 19630 41918 19682 41970
rect 20078 41918 20130 41970
rect 20190 41918 20242 41970
rect 20302 41918 20354 41970
rect 20414 41918 20466 41970
rect 20638 41918 20690 41970
rect 21086 41918 21138 41970
rect 21310 41918 21362 41970
rect 21870 41918 21922 41970
rect 22206 41918 22258 41970
rect 23550 41918 23602 41970
rect 23998 41918 24050 41970
rect 24670 41918 24722 41970
rect 28030 41918 28082 41970
rect 6974 41806 7026 41858
rect 7534 41806 7586 41858
rect 9886 41806 9938 41858
rect 13022 41806 13074 41858
rect 15150 41806 15202 41858
rect 15822 41806 15874 41858
rect 25230 41806 25282 41858
rect 27358 41806 27410 41858
rect 2718 41694 2770 41746
rect 16270 41694 16322 41746
rect 21646 41694 21698 41746
rect 22206 41694 22258 41746
rect 22878 41694 22930 41746
rect 23326 41694 23378 41746
rect 4616 41526 4668 41578
rect 4720 41526 4772 41578
rect 4824 41526 4876 41578
rect 11420 41526 11472 41578
rect 11524 41526 11576 41578
rect 11628 41526 11680 41578
rect 18224 41526 18276 41578
rect 18328 41526 18380 41578
rect 18432 41526 18484 41578
rect 25028 41526 25080 41578
rect 25132 41526 25184 41578
rect 25236 41526 25288 41578
rect 2718 41358 2770 41410
rect 3054 41358 3106 41410
rect 3278 41358 3330 41410
rect 3950 41358 4002 41410
rect 22430 41358 22482 41410
rect 22766 41358 22818 41410
rect 26350 41358 26402 41410
rect 3950 41246 4002 41298
rect 4846 41246 4898 41298
rect 10558 41246 10610 41298
rect 11790 41246 11842 41298
rect 14590 41246 14642 41298
rect 15598 41246 15650 41298
rect 17726 41246 17778 41298
rect 19518 41246 19570 41298
rect 20414 41246 20466 41298
rect 21422 41246 21474 41298
rect 22766 41246 22818 41298
rect 23998 41246 24050 41298
rect 24670 41246 24722 41298
rect 25118 41246 25170 41298
rect 27358 41246 27410 41298
rect 28030 41246 28082 41298
rect 5854 41134 5906 41186
rect 6862 41134 6914 41186
rect 7646 41134 7698 41186
rect 13582 41134 13634 41186
rect 14030 41134 14082 41186
rect 14814 41134 14866 41186
rect 18846 41134 18898 41186
rect 19406 41134 19458 41186
rect 19966 41134 20018 41186
rect 26350 41134 26402 41186
rect 26686 41134 26738 41186
rect 6302 41022 6354 41074
rect 8430 41022 8482 41074
rect 12238 41022 12290 41074
rect 13470 41022 13522 41074
rect 13806 41022 13858 41074
rect 18286 41022 18338 41074
rect 18622 41022 18674 41074
rect 26910 41022 26962 41074
rect 2046 40910 2098 40962
rect 2382 40910 2434 40962
rect 2830 40910 2882 40962
rect 3502 40910 3554 40962
rect 4398 40910 4450 40962
rect 6190 40910 6242 40962
rect 7310 40910 7362 40962
rect 11342 40910 11394 40962
rect 12798 40910 12850 40962
rect 18510 40910 18562 40962
rect 19630 40910 19682 40962
rect 21870 40910 21922 40962
rect 22318 40910 22370 40962
rect 23550 40910 23602 40962
rect 25790 40910 25842 40962
rect 26798 40910 26850 40962
rect 8018 40742 8070 40794
rect 8122 40742 8174 40794
rect 8226 40742 8278 40794
rect 14822 40742 14874 40794
rect 14926 40742 14978 40794
rect 15030 40742 15082 40794
rect 21626 40742 21678 40794
rect 21730 40742 21782 40794
rect 21834 40742 21886 40794
rect 28430 40742 28482 40794
rect 28534 40742 28586 40794
rect 28638 40742 28690 40794
rect 2718 40574 2770 40626
rect 8430 40574 8482 40626
rect 10334 40574 10386 40626
rect 10782 40574 10834 40626
rect 11566 40574 11618 40626
rect 13246 40574 13298 40626
rect 13582 40574 13634 40626
rect 14030 40574 14082 40626
rect 15150 40574 15202 40626
rect 15598 40574 15650 40626
rect 16046 40574 16098 40626
rect 16718 40574 16770 40626
rect 21086 40574 21138 40626
rect 21534 40574 21586 40626
rect 22430 40574 22482 40626
rect 22878 40574 22930 40626
rect 23326 40574 23378 40626
rect 23886 40574 23938 40626
rect 25342 40574 25394 40626
rect 27470 40574 27522 40626
rect 28142 40574 28194 40626
rect 2046 40462 2098 40514
rect 3166 40462 3218 40514
rect 8206 40462 8258 40514
rect 11118 40462 11170 40514
rect 18510 40462 18562 40514
rect 21982 40462 22034 40514
rect 24110 40462 24162 40514
rect 26350 40462 26402 40514
rect 1710 40350 1762 40402
rect 2494 40350 2546 40402
rect 2942 40350 2994 40402
rect 3614 40350 3666 40402
rect 4286 40350 4338 40402
rect 8430 40350 8482 40402
rect 8990 40350 9042 40402
rect 9886 40350 9938 40402
rect 11342 40350 11394 40402
rect 11790 40350 11842 40402
rect 12574 40350 12626 40402
rect 17726 40350 17778 40402
rect 24334 40350 24386 40402
rect 24670 40350 24722 40402
rect 25790 40350 25842 40402
rect 26798 40350 26850 40402
rect 5070 40238 5122 40290
rect 7198 40238 7250 40290
rect 7870 40238 7922 40290
rect 9550 40238 9602 40290
rect 9662 40238 9714 40290
rect 12238 40238 12290 40290
rect 12350 40238 12402 40290
rect 14478 40238 14530 40290
rect 20638 40238 20690 40290
rect 24222 40238 24274 40290
rect 2606 40126 2658 40178
rect 3726 40126 3778 40178
rect 8766 40126 8818 40178
rect 11678 40126 11730 40178
rect 4616 39958 4668 40010
rect 4720 39958 4772 40010
rect 4824 39958 4876 40010
rect 11420 39958 11472 40010
rect 11524 39958 11576 40010
rect 11628 39958 11680 40010
rect 18224 39958 18276 40010
rect 18328 39958 18380 40010
rect 18432 39958 18484 40010
rect 25028 39958 25080 40010
rect 25132 39958 25184 40010
rect 25236 39958 25288 40010
rect 5966 39790 6018 39842
rect 7310 39790 7362 39842
rect 7870 39790 7922 39842
rect 8766 39790 8818 39842
rect 9662 39790 9714 39842
rect 13582 39790 13634 39842
rect 14478 39790 14530 39842
rect 17838 39790 17890 39842
rect 18734 39790 18786 39842
rect 19406 39790 19458 39842
rect 19630 39790 19682 39842
rect 26798 39790 26850 39842
rect 27358 39790 27410 39842
rect 27694 39790 27746 39842
rect 2494 39678 2546 39730
rect 4622 39678 4674 39730
rect 5070 39678 5122 39730
rect 7198 39678 7250 39730
rect 8094 39678 8146 39730
rect 8542 39678 8594 39730
rect 8990 39678 9042 39730
rect 10782 39678 10834 39730
rect 12910 39678 12962 39730
rect 16046 39678 16098 39730
rect 16382 39678 16434 39730
rect 19406 39678 19458 39730
rect 20414 39678 20466 39730
rect 22654 39678 22706 39730
rect 22990 39678 23042 39730
rect 28142 39678 28194 39730
rect 1822 39566 1874 39618
rect 5630 39566 5682 39618
rect 6190 39566 6242 39618
rect 6414 39566 6466 39618
rect 9998 39566 10050 39618
rect 14142 39566 14194 39618
rect 15150 39566 15202 39618
rect 25902 39566 25954 39618
rect 26238 39566 26290 39618
rect 26462 39566 26514 39618
rect 26910 39566 26962 39618
rect 14590 39454 14642 39506
rect 14926 39454 14978 39506
rect 15486 39454 15538 39506
rect 25118 39454 25170 39506
rect 5630 39342 5682 39394
rect 7758 39342 7810 39394
rect 9550 39342 9602 39394
rect 13582 39342 13634 39394
rect 15150 39342 15202 39394
rect 16942 39342 16994 39394
rect 17838 39342 17890 39394
rect 18174 39342 18226 39394
rect 18622 39342 18674 39394
rect 19854 39342 19906 39394
rect 20750 39342 20802 39394
rect 21422 39342 21474 39394
rect 21870 39342 21922 39394
rect 27022 39342 27074 39394
rect 27470 39342 27522 39394
rect 8018 39174 8070 39226
rect 8122 39174 8174 39226
rect 8226 39174 8278 39226
rect 14822 39174 14874 39226
rect 14926 39174 14978 39226
rect 15030 39174 15082 39226
rect 21626 39174 21678 39226
rect 21730 39174 21782 39226
rect 21834 39174 21886 39226
rect 28430 39174 28482 39226
rect 28534 39174 28586 39226
rect 28638 39174 28690 39226
rect 2270 39006 2322 39058
rect 3390 39006 3442 39058
rect 3950 39006 4002 39058
rect 4398 39006 4450 39058
rect 5518 39006 5570 39058
rect 10110 39006 10162 39058
rect 10894 39006 10946 39058
rect 11342 39006 11394 39058
rect 12798 39006 12850 39058
rect 19630 39006 19682 39058
rect 19966 39006 20018 39058
rect 23998 39006 24050 39058
rect 3502 38894 3554 38946
rect 5070 38894 5122 38946
rect 14702 38894 14754 38946
rect 18062 38894 18114 38946
rect 18846 38894 18898 38946
rect 19854 38894 19906 38946
rect 24110 38894 24162 38946
rect 24334 38894 24386 38946
rect 27358 38894 27410 38946
rect 1822 38782 1874 38834
rect 12350 38782 12402 38834
rect 14030 38782 14082 38834
rect 18510 38782 18562 38834
rect 18734 38782 18786 38834
rect 19406 38782 19458 38834
rect 19742 38782 19794 38834
rect 20638 38782 20690 38834
rect 23662 38782 23714 38834
rect 28030 38782 28082 38834
rect 11678 38670 11730 38722
rect 16830 38670 16882 38722
rect 17502 38670 17554 38722
rect 19070 38670 19122 38722
rect 21310 38670 21362 38722
rect 23438 38670 23490 38722
rect 25230 38670 25282 38722
rect 4616 38390 4668 38442
rect 4720 38390 4772 38442
rect 4824 38390 4876 38442
rect 11420 38390 11472 38442
rect 11524 38390 11576 38442
rect 11628 38390 11680 38442
rect 18224 38390 18276 38442
rect 18328 38390 18380 38442
rect 18432 38390 18484 38442
rect 25028 38390 25080 38442
rect 25132 38390 25184 38442
rect 25236 38390 25288 38442
rect 2382 38222 2434 38274
rect 11790 38222 11842 38274
rect 12126 38222 12178 38274
rect 13694 38222 13746 38274
rect 14030 38222 14082 38274
rect 21982 38222 22034 38274
rect 23550 38222 23602 38274
rect 24110 38222 24162 38274
rect 26462 38222 26514 38274
rect 27246 38222 27298 38274
rect 9102 38110 9154 38162
rect 11790 38110 11842 38162
rect 13582 38110 13634 38162
rect 16494 38110 16546 38162
rect 20190 38110 20242 38162
rect 20750 38110 20802 38162
rect 21534 38110 21586 38162
rect 24110 38110 24162 38162
rect 25230 38110 25282 38162
rect 25678 38110 25730 38162
rect 27022 38110 27074 38162
rect 27470 38110 27522 38162
rect 2382 37998 2434 38050
rect 3390 37998 3442 38050
rect 6190 37998 6242 38050
rect 10110 37998 10162 38050
rect 10558 37998 10610 38050
rect 10782 37998 10834 38050
rect 15934 37998 15986 38050
rect 21758 37998 21810 38050
rect 22094 37998 22146 38050
rect 22766 37998 22818 38050
rect 23102 37998 23154 38050
rect 23662 37998 23714 38050
rect 2718 37886 2770 37938
rect 2942 37886 2994 37938
rect 6974 37886 7026 37938
rect 21422 37886 21474 37938
rect 2494 37774 2546 37826
rect 3838 37774 3890 37826
rect 5854 37774 5906 37826
rect 10334 37774 10386 37826
rect 10446 37774 10498 37826
rect 11230 37774 11282 37826
rect 12238 37774 12290 37826
rect 12910 37774 12962 37826
rect 14142 37774 14194 37826
rect 22654 37774 22706 37826
rect 22878 37774 22930 37826
rect 22990 37774 23042 37826
rect 24782 37774 24834 37826
rect 26126 37774 26178 37826
rect 26574 37774 26626 37826
rect 28142 37774 28194 37826
rect 8018 37606 8070 37658
rect 8122 37606 8174 37658
rect 8226 37606 8278 37658
rect 14822 37606 14874 37658
rect 14926 37606 14978 37658
rect 15030 37606 15082 37658
rect 21626 37606 21678 37658
rect 21730 37606 21782 37658
rect 21834 37606 21886 37658
rect 28430 37606 28482 37658
rect 28534 37606 28586 37658
rect 28638 37606 28690 37658
rect 6414 37438 6466 37490
rect 6862 37438 6914 37490
rect 7310 37438 7362 37490
rect 8206 37438 8258 37490
rect 8430 37438 8482 37490
rect 9662 37438 9714 37490
rect 11454 37438 11506 37490
rect 13582 37438 13634 37490
rect 13918 37438 13970 37490
rect 15262 37438 15314 37490
rect 16046 37438 16098 37490
rect 16830 37438 16882 37490
rect 17502 37438 17554 37490
rect 17614 37438 17666 37490
rect 18398 37438 18450 37490
rect 18846 37438 18898 37490
rect 19070 37438 19122 37490
rect 19854 37438 19906 37490
rect 20862 37438 20914 37490
rect 22318 37438 22370 37490
rect 22990 37438 23042 37490
rect 23438 37438 23490 37490
rect 25230 37438 25282 37490
rect 25678 37438 25730 37490
rect 27358 37438 27410 37490
rect 2494 37326 2546 37378
rect 7534 37326 7586 37378
rect 7758 37326 7810 37378
rect 10110 37326 10162 37378
rect 11006 37326 11058 37378
rect 11230 37326 11282 37378
rect 11790 37326 11842 37378
rect 20414 37326 20466 37378
rect 23998 37326 24050 37378
rect 24334 37326 24386 37378
rect 1822 37214 1874 37266
rect 7086 37214 7138 37266
rect 8318 37214 8370 37266
rect 8766 37214 8818 37266
rect 9998 37214 10050 37266
rect 10334 37214 10386 37266
rect 10558 37214 10610 37266
rect 11454 37214 11506 37266
rect 12126 37214 12178 37266
rect 12574 37214 12626 37266
rect 12798 37214 12850 37266
rect 14254 37214 14306 37266
rect 14478 37214 14530 37266
rect 14590 37214 14642 37266
rect 15038 37214 15090 37266
rect 17390 37214 17442 37266
rect 17950 37214 18002 37266
rect 18958 37214 19010 37266
rect 19182 37214 19234 37266
rect 19406 37214 19458 37266
rect 22542 37214 22594 37266
rect 24558 37214 24610 37266
rect 25342 37214 25394 37266
rect 25454 37214 25506 37266
rect 26910 37214 26962 37266
rect 4622 37102 4674 37154
rect 5070 37102 5122 37154
rect 5966 37102 6018 37154
rect 12686 37102 12738 37154
rect 15598 37102 15650 37154
rect 21310 37102 21362 37154
rect 21758 37102 21810 37154
rect 21982 37102 22034 37154
rect 24110 37102 24162 37154
rect 5854 36990 5906 37042
rect 21310 36990 21362 37042
rect 26238 37102 26290 37154
rect 26798 37102 26850 37154
rect 27918 37102 27970 37154
rect 22206 36990 22258 37042
rect 26574 36990 26626 37042
rect 4616 36822 4668 36874
rect 4720 36822 4772 36874
rect 4824 36822 4876 36874
rect 11420 36822 11472 36874
rect 11524 36822 11576 36874
rect 11628 36822 11680 36874
rect 18224 36822 18276 36874
rect 18328 36822 18380 36874
rect 18432 36822 18484 36874
rect 25028 36822 25080 36874
rect 25132 36822 25184 36874
rect 25236 36822 25288 36874
rect 3166 36654 3218 36706
rect 6862 36654 6914 36706
rect 14366 36654 14418 36706
rect 18622 36654 18674 36706
rect 2494 36542 2546 36594
rect 3278 36542 3330 36594
rect 3950 36542 4002 36594
rect 5070 36542 5122 36594
rect 8654 36542 8706 36594
rect 9326 36542 9378 36594
rect 9998 36542 10050 36594
rect 12126 36542 12178 36594
rect 14590 36542 14642 36594
rect 18398 36542 18450 36594
rect 1710 36430 1762 36482
rect 4734 36430 4786 36482
rect 5630 36430 5682 36482
rect 5966 36430 6018 36482
rect 6078 36430 6130 36482
rect 6750 36430 6802 36482
rect 8206 36430 8258 36482
rect 8430 36430 8482 36482
rect 8878 36430 8930 36482
rect 12910 36430 12962 36482
rect 13694 36430 13746 36482
rect 13918 36430 13970 36482
rect 14030 36430 14082 36482
rect 14702 36430 14754 36482
rect 15150 36430 15202 36482
rect 15262 36430 15314 36482
rect 15486 36430 15538 36482
rect 15710 36430 15762 36482
rect 16494 36430 16546 36482
rect 4958 36318 5010 36370
rect 6414 36318 6466 36370
rect 13470 36318 13522 36370
rect 16046 36318 16098 36370
rect 16606 36318 16658 36370
rect 17614 36318 17666 36370
rect 2046 36206 2098 36258
rect 4398 36206 4450 36258
rect 5630 36206 5682 36258
rect 8654 36206 8706 36258
rect 15374 36206 15426 36258
rect 16270 36206 16322 36258
rect 16382 36206 16434 36258
rect 26798 36654 26850 36706
rect 19966 36542 20018 36594
rect 22430 36542 22482 36594
rect 22766 36542 22818 36594
rect 24110 36542 24162 36594
rect 26238 36542 26290 36594
rect 27806 36542 27858 36594
rect 18958 36430 19010 36482
rect 21310 36430 21362 36482
rect 23438 36430 23490 36482
rect 26574 36430 26626 36482
rect 27022 36430 27074 36482
rect 27358 36430 27410 36482
rect 19406 36318 19458 36370
rect 21422 36318 21474 36370
rect 21646 36318 21698 36370
rect 21870 36318 21922 36370
rect 17166 36206 17218 36258
rect 18734 36206 18786 36258
rect 19070 36206 19122 36258
rect 19182 36206 19234 36258
rect 20414 36206 20466 36258
rect 27246 36206 27298 36258
rect 8018 36038 8070 36090
rect 8122 36038 8174 36090
rect 8226 36038 8278 36090
rect 14822 36038 14874 36090
rect 14926 36038 14978 36090
rect 15030 36038 15082 36090
rect 21626 36038 21678 36090
rect 21730 36038 21782 36090
rect 21834 36038 21886 36090
rect 28430 36038 28482 36090
rect 28534 36038 28586 36090
rect 28638 36038 28690 36090
rect 3726 35870 3778 35922
rect 7422 35870 7474 35922
rect 8542 35870 8594 35922
rect 8990 35870 9042 35922
rect 10110 35870 10162 35922
rect 12462 35870 12514 35922
rect 16718 35870 16770 35922
rect 4846 35758 4898 35810
rect 9662 35758 9714 35810
rect 22990 35758 23042 35810
rect 27358 35758 27410 35810
rect 4062 35646 4114 35698
rect 12126 35646 12178 35698
rect 12238 35646 12290 35698
rect 12574 35646 12626 35698
rect 13358 35646 13410 35698
rect 17390 35646 17442 35698
rect 23774 35646 23826 35698
rect 28030 35646 28082 35698
rect 1822 35534 1874 35586
rect 6974 35534 7026 35586
rect 10782 35534 10834 35586
rect 11678 35534 11730 35586
rect 12350 35534 12402 35586
rect 14142 35534 14194 35586
rect 16270 35534 16322 35586
rect 18174 35534 18226 35586
rect 20302 35534 20354 35586
rect 20862 35534 20914 35586
rect 24222 35534 24274 35586
rect 24670 35534 24722 35586
rect 25230 35534 25282 35586
rect 4616 35254 4668 35306
rect 4720 35254 4772 35306
rect 4824 35254 4876 35306
rect 11420 35254 11472 35306
rect 11524 35254 11576 35306
rect 11628 35254 11680 35306
rect 18224 35254 18276 35306
rect 18328 35254 18380 35306
rect 18432 35254 18484 35306
rect 25028 35254 25080 35306
rect 25132 35254 25184 35306
rect 25236 35254 25288 35306
rect 11678 35086 11730 35138
rect 13582 35086 13634 35138
rect 13918 35086 13970 35138
rect 14478 35086 14530 35138
rect 16382 35086 16434 35138
rect 18622 35086 18674 35138
rect 18958 35086 19010 35138
rect 19182 35086 19234 35138
rect 24782 35086 24834 35138
rect 25118 35086 25170 35138
rect 25902 35086 25954 35138
rect 26574 35086 26626 35138
rect 2942 34974 2994 35026
rect 4846 34974 4898 35026
rect 8654 34974 8706 35026
rect 12910 34974 12962 35026
rect 13582 34974 13634 35026
rect 14814 34974 14866 35026
rect 18062 34974 18114 35026
rect 21534 34974 21586 35026
rect 21982 34974 22034 35026
rect 24670 34974 24722 35026
rect 26238 34974 26290 35026
rect 26574 34974 26626 35026
rect 27134 34974 27186 35026
rect 2830 34862 2882 34914
rect 3502 34862 3554 34914
rect 8094 34862 8146 34914
rect 8318 34862 8370 34914
rect 10110 34862 10162 34914
rect 10670 34862 10722 34914
rect 11342 34862 11394 34914
rect 14142 34862 14194 34914
rect 14702 34862 14754 34914
rect 14926 34862 14978 34914
rect 15934 34862 15986 34914
rect 17950 34862 18002 34914
rect 18174 34862 18226 34914
rect 18510 34862 18562 34914
rect 19630 34862 19682 34914
rect 20190 34862 20242 34914
rect 22542 34862 22594 34914
rect 1710 34750 1762 34802
rect 3390 34750 3442 34802
rect 7758 34750 7810 34802
rect 8654 34750 8706 34802
rect 9550 34750 9602 34802
rect 9774 34750 9826 34802
rect 10334 34750 10386 34802
rect 10782 34750 10834 34802
rect 11006 34750 11058 34802
rect 15710 34750 15762 34802
rect 15822 34750 15874 34802
rect 17614 34750 17666 34802
rect 19742 34750 19794 34802
rect 20078 34750 20130 34802
rect 20638 34750 20690 34802
rect 2046 34638 2098 34690
rect 8542 34638 8594 34690
rect 10110 34638 10162 34690
rect 12462 34638 12514 34690
rect 17054 34638 17106 34690
rect 18958 34638 19010 34690
rect 21870 34638 21922 34690
rect 22094 34638 22146 34690
rect 22878 34638 22930 34690
rect 23326 34638 23378 34690
rect 23886 34638 23938 34690
rect 24222 34638 24274 34690
rect 25118 34638 25170 34690
rect 25678 34638 25730 34690
rect 27694 34638 27746 34690
rect 28142 34638 28194 34690
rect 8018 34470 8070 34522
rect 8122 34470 8174 34522
rect 8226 34470 8278 34522
rect 14822 34470 14874 34522
rect 14926 34470 14978 34522
rect 15030 34470 15082 34522
rect 21626 34470 21678 34522
rect 21730 34470 21782 34522
rect 21834 34470 21886 34522
rect 28430 34470 28482 34522
rect 28534 34470 28586 34522
rect 28638 34470 28690 34522
rect 6414 34302 6466 34354
rect 7198 34302 7250 34354
rect 8990 34302 9042 34354
rect 12126 34302 12178 34354
rect 13918 34302 13970 34354
rect 15822 34302 15874 34354
rect 18622 34302 18674 34354
rect 19070 34302 19122 34354
rect 19966 34302 20018 34354
rect 20190 34302 20242 34354
rect 20750 34302 20802 34354
rect 21198 34302 21250 34354
rect 21758 34302 21810 34354
rect 22766 34302 22818 34354
rect 23326 34302 23378 34354
rect 25342 34302 25394 34354
rect 26686 34302 26738 34354
rect 27806 34302 27858 34354
rect 5742 34190 5794 34242
rect 27134 34190 27186 34242
rect 27358 34190 27410 34242
rect 1822 34078 1874 34130
rect 5182 34078 5234 34130
rect 5966 34078 6018 34130
rect 7870 34078 7922 34130
rect 8094 34078 8146 34130
rect 8318 34078 8370 34130
rect 8430 34078 8482 34130
rect 9550 34078 9602 34130
rect 9774 34078 9826 34130
rect 9998 34078 10050 34130
rect 10110 34078 10162 34130
rect 10558 34078 10610 34130
rect 10782 34078 10834 34130
rect 11118 34078 11170 34130
rect 19630 34078 19682 34130
rect 19854 34078 19906 34130
rect 20078 34078 20130 34130
rect 25902 34078 25954 34130
rect 26126 34078 26178 34130
rect 26462 34078 26514 34130
rect 2494 33966 2546 34018
rect 4622 33966 4674 34018
rect 5854 33966 5906 34018
rect 6526 33966 6578 34018
rect 7534 33966 7586 34018
rect 8206 33966 8258 34018
rect 9886 33966 9938 34018
rect 10670 33966 10722 34018
rect 11566 33966 11618 34018
rect 12462 33966 12514 34018
rect 15374 33966 15426 34018
rect 18062 33966 18114 34018
rect 22094 33966 22146 34018
rect 23662 33966 23714 34018
rect 24222 33966 24274 34018
rect 24670 33966 24722 34018
rect 5406 33854 5458 33906
rect 23998 33854 24050 33906
rect 24670 33854 24722 33906
rect 26462 33854 26514 33906
rect 27022 33854 27074 33906
rect 4616 33686 4668 33738
rect 4720 33686 4772 33738
rect 4824 33686 4876 33738
rect 11420 33686 11472 33738
rect 11524 33686 11576 33738
rect 11628 33686 11680 33738
rect 18224 33686 18276 33738
rect 18328 33686 18380 33738
rect 18432 33686 18484 33738
rect 25028 33686 25080 33738
rect 25132 33686 25184 33738
rect 25236 33686 25288 33738
rect 3726 33518 3778 33570
rect 8990 33518 9042 33570
rect 9550 33518 9602 33570
rect 9774 33518 9826 33570
rect 10110 33518 10162 33570
rect 21422 33518 21474 33570
rect 2606 33406 2658 33458
rect 3502 33406 3554 33458
rect 6414 33406 6466 33458
rect 8542 33406 8594 33458
rect 9102 33406 9154 33458
rect 9550 33406 9602 33458
rect 10110 33406 10162 33458
rect 12798 33406 12850 33458
rect 14926 33406 14978 33458
rect 18062 33406 18114 33458
rect 24894 33406 24946 33458
rect 25230 33406 25282 33458
rect 27358 33406 27410 33458
rect 2382 33294 2434 33346
rect 2830 33294 2882 33346
rect 3390 33294 3442 33346
rect 5742 33294 5794 33346
rect 10446 33294 10498 33346
rect 11118 33294 11170 33346
rect 12014 33294 12066 33346
rect 12350 33294 12402 33346
rect 15150 33294 15202 33346
rect 20078 33294 20130 33346
rect 20190 33294 20242 33346
rect 21310 33294 21362 33346
rect 22430 33294 22482 33346
rect 22654 33294 22706 33346
rect 23998 33294 24050 33346
rect 28030 33294 28082 33346
rect 3054 33182 3106 33234
rect 10558 33182 10610 33234
rect 10670 33182 10722 33234
rect 11678 33182 11730 33234
rect 14814 33182 14866 33234
rect 15598 33182 15650 33234
rect 19070 33182 19122 33234
rect 20526 33182 20578 33234
rect 22878 33182 22930 33234
rect 2606 33070 2658 33122
rect 4398 33070 4450 33122
rect 4846 33070 4898 33122
rect 11342 33070 11394 33122
rect 11902 33070 11954 33122
rect 12126 33070 12178 33122
rect 13582 33070 13634 33122
rect 18510 33070 18562 33122
rect 19518 33070 19570 33122
rect 19966 33070 20018 33122
rect 20302 33070 20354 33122
rect 21422 33070 21474 33122
rect 22318 33070 22370 33122
rect 22542 33070 22594 33122
rect 23438 33070 23490 33122
rect 23550 33070 23602 33122
rect 23662 33070 23714 33122
rect 24446 33070 24498 33122
rect 8018 32902 8070 32954
rect 8122 32902 8174 32954
rect 8226 32902 8278 32954
rect 14822 32902 14874 32954
rect 14926 32902 14978 32954
rect 15030 32902 15082 32954
rect 21626 32902 21678 32954
rect 21730 32902 21782 32954
rect 21834 32902 21886 32954
rect 28430 32902 28482 32954
rect 28534 32902 28586 32954
rect 28638 32902 28690 32954
rect 2606 32734 2658 32786
rect 3054 32734 3106 32786
rect 3502 32734 3554 32786
rect 10446 32734 10498 32786
rect 11006 32734 11058 32786
rect 11454 32734 11506 32786
rect 12574 32734 12626 32786
rect 18734 32734 18786 32786
rect 20190 32734 20242 32786
rect 25678 32734 25730 32786
rect 27134 32734 27186 32786
rect 17390 32622 17442 32674
rect 12910 32510 12962 32562
rect 17726 32510 17778 32562
rect 17838 32510 17890 32562
rect 18398 32510 18450 32562
rect 18622 32510 18674 32562
rect 18846 32510 18898 32562
rect 19070 32510 19122 32562
rect 19518 32510 19570 32562
rect 19966 32510 20018 32562
rect 20078 32510 20130 32562
rect 20302 32510 20354 32562
rect 20526 32510 20578 32562
rect 21870 32510 21922 32562
rect 26014 32510 26066 32562
rect 26350 32510 26402 32562
rect 1822 32398 1874 32450
rect 3950 32398 4002 32450
rect 8766 32398 8818 32450
rect 12126 32398 12178 32450
rect 13694 32398 13746 32450
rect 15822 32398 15874 32450
rect 16270 32398 16322 32450
rect 16830 32398 16882 32450
rect 17502 32398 17554 32450
rect 20974 32398 21026 32450
rect 21422 32398 21474 32450
rect 22542 32398 22594 32450
rect 24670 32398 24722 32450
rect 27918 32398 27970 32450
rect 3166 32286 3218 32338
rect 3502 32286 3554 32338
rect 3950 32286 4002 32338
rect 26350 32286 26402 32338
rect 26686 32286 26738 32338
rect 4616 32118 4668 32170
rect 4720 32118 4772 32170
rect 4824 32118 4876 32170
rect 11420 32118 11472 32170
rect 11524 32118 11576 32170
rect 11628 32118 11680 32170
rect 18224 32118 18276 32170
rect 18328 32118 18380 32170
rect 18432 32118 18484 32170
rect 25028 32118 25080 32170
rect 25132 32118 25184 32170
rect 25236 32118 25288 32170
rect 2494 31950 2546 32002
rect 11902 31950 11954 32002
rect 12798 31950 12850 32002
rect 19182 31950 19234 32002
rect 3390 31838 3442 31890
rect 9102 31838 9154 31890
rect 9998 31838 10050 31890
rect 12462 31838 12514 31890
rect 23102 31838 23154 31890
rect 24222 31838 24274 31890
rect 25230 31838 25282 31890
rect 2830 31726 2882 31778
rect 4062 31726 4114 31778
rect 4734 31726 4786 31778
rect 5854 31726 5906 31778
rect 6302 31726 6354 31778
rect 9774 31726 9826 31778
rect 10222 31726 10274 31778
rect 11566 31726 11618 31778
rect 12014 31726 12066 31778
rect 17278 31726 17330 31778
rect 19406 31726 19458 31778
rect 20190 31726 20242 31778
rect 20750 31726 20802 31778
rect 21310 31726 21362 31778
rect 22990 31726 23042 31778
rect 23550 31726 23602 31778
rect 28030 31726 28082 31778
rect 1710 31614 1762 31666
rect 2046 31614 2098 31666
rect 5070 31614 5122 31666
rect 6974 31614 7026 31666
rect 9550 31614 9602 31666
rect 11342 31614 11394 31666
rect 12574 31614 12626 31666
rect 16718 31614 16770 31666
rect 19518 31614 19570 31666
rect 21534 31614 21586 31666
rect 22206 31614 22258 31666
rect 22542 31614 22594 31666
rect 23326 31614 23378 31666
rect 24670 31614 24722 31666
rect 27358 31614 27410 31666
rect 2606 31502 2658 31554
rect 3278 31502 3330 31554
rect 4174 31502 4226 31554
rect 9998 31502 10050 31554
rect 11006 31502 11058 31554
rect 11454 31502 11506 31554
rect 8018 31334 8070 31386
rect 8122 31334 8174 31386
rect 8226 31334 8278 31386
rect 14822 31334 14874 31386
rect 14926 31334 14978 31386
rect 15030 31334 15082 31386
rect 21626 31334 21678 31386
rect 21730 31334 21782 31386
rect 21834 31334 21886 31386
rect 28430 31334 28482 31386
rect 28534 31334 28586 31386
rect 28638 31334 28690 31386
rect 5070 31166 5122 31218
rect 5742 31166 5794 31218
rect 6302 31166 6354 31218
rect 7086 31166 7138 31218
rect 9886 31166 9938 31218
rect 10222 31166 10274 31218
rect 14142 31166 14194 31218
rect 15934 31166 15986 31218
rect 16046 31166 16098 31218
rect 16494 31166 16546 31218
rect 16942 31166 16994 31218
rect 17950 31166 18002 31218
rect 19070 31166 19122 31218
rect 19518 31166 19570 31218
rect 21646 31166 21698 31218
rect 24110 31166 24162 31218
rect 26686 31166 26738 31218
rect 7198 31054 7250 31106
rect 8206 31054 8258 31106
rect 11342 31054 11394 31106
rect 15486 31054 15538 31106
rect 18174 31054 18226 31106
rect 18734 31054 18786 31106
rect 18846 31054 18898 31106
rect 19854 31054 19906 31106
rect 22542 31054 22594 31106
rect 24334 31054 24386 31106
rect 26126 31054 26178 31106
rect 1822 30942 1874 30994
rect 6974 30942 7026 30994
rect 7534 30942 7586 30994
rect 8430 30942 8482 30994
rect 10670 30942 10722 30994
rect 14030 30942 14082 30994
rect 14254 30942 14306 30994
rect 14590 30942 14642 30994
rect 15710 30942 15762 30994
rect 17614 30942 17666 30994
rect 17838 30942 17890 30994
rect 18062 30942 18114 30994
rect 21534 30942 21586 30994
rect 21982 30942 22034 30994
rect 24670 30942 24722 30994
rect 25902 30942 25954 30994
rect 26350 30942 26402 30994
rect 26462 30942 26514 30994
rect 2494 30830 2546 30882
rect 4622 30830 4674 30882
rect 6638 30830 6690 30882
rect 8094 30830 8146 30882
rect 8878 30830 8930 30882
rect 13470 30830 13522 30882
rect 24222 30830 24274 30882
rect 25342 30830 25394 30882
rect 27134 30830 27186 30882
rect 27582 30830 27634 30882
rect 28142 30830 28194 30882
rect 7534 30718 7586 30770
rect 14590 30718 14642 30770
rect 27246 30718 27298 30770
rect 28142 30718 28194 30770
rect 4616 30550 4668 30602
rect 4720 30550 4772 30602
rect 4824 30550 4876 30602
rect 11420 30550 11472 30602
rect 11524 30550 11576 30602
rect 11628 30550 11680 30602
rect 18224 30550 18276 30602
rect 18328 30550 18380 30602
rect 18432 30550 18484 30602
rect 25028 30550 25080 30602
rect 25132 30550 25184 30602
rect 25236 30550 25288 30602
rect 2606 30382 2658 30434
rect 3502 30382 3554 30434
rect 4062 30382 4114 30434
rect 4734 30382 4786 30434
rect 5070 30382 5122 30434
rect 5854 30382 5906 30434
rect 18846 30382 18898 30434
rect 19070 30382 19122 30434
rect 20638 30382 20690 30434
rect 6862 30270 6914 30322
rect 7646 30270 7698 30322
rect 8318 30270 8370 30322
rect 8430 30270 8482 30322
rect 9774 30270 9826 30322
rect 10894 30270 10946 30322
rect 11454 30270 11506 30322
rect 12574 30270 12626 30322
rect 14814 30270 14866 30322
rect 18398 30270 18450 30322
rect 21422 30270 21474 30322
rect 2046 30158 2098 30210
rect 2270 30158 2322 30210
rect 2830 30158 2882 30210
rect 5070 30158 5122 30210
rect 5630 30158 5682 30210
rect 6414 30158 6466 30210
rect 7198 30158 7250 30210
rect 7422 30158 7474 30210
rect 7870 30158 7922 30210
rect 9550 30158 9602 30210
rect 9886 30158 9938 30210
rect 10334 30158 10386 30210
rect 10558 30158 10610 30210
rect 12014 30158 12066 30210
rect 15598 30158 15650 30210
rect 16270 30158 16322 30210
rect 18846 30158 18898 30210
rect 19854 30158 19906 30210
rect 20750 30158 20802 30210
rect 23998 30158 24050 30210
rect 3054 30046 3106 30098
rect 6190 30046 6242 30098
rect 9326 30046 9378 30098
rect 10894 30046 10946 30098
rect 15150 30046 15202 30098
rect 27918 30046 27970 30098
rect 2606 29934 2658 29986
rect 3614 29934 3666 29986
rect 3950 29934 4002 29986
rect 4398 29934 4450 29986
rect 5630 29934 5682 29986
rect 7310 29934 7362 29986
rect 8542 29934 8594 29986
rect 9774 29934 9826 29986
rect 10782 29934 10834 29986
rect 12910 29934 12962 29986
rect 13806 29934 13858 29986
rect 14142 29934 14194 29986
rect 14590 29934 14642 29986
rect 14702 29934 14754 29986
rect 14926 29934 14978 29986
rect 19294 29934 19346 29986
rect 20190 29934 20242 29986
rect 20638 29934 20690 29986
rect 21870 29934 21922 29986
rect 22542 29934 22594 29986
rect 8018 29766 8070 29818
rect 8122 29766 8174 29818
rect 8226 29766 8278 29818
rect 14822 29766 14874 29818
rect 14926 29766 14978 29818
rect 15030 29766 15082 29818
rect 21626 29766 21678 29818
rect 21730 29766 21782 29818
rect 21834 29766 21886 29818
rect 28430 29766 28482 29818
rect 28534 29766 28586 29818
rect 28638 29766 28690 29818
rect 10558 29598 10610 29650
rect 11902 29598 11954 29650
rect 12350 29598 12402 29650
rect 16158 29598 16210 29650
rect 17726 29598 17778 29650
rect 17838 29598 17890 29650
rect 2046 29486 2098 29538
rect 3614 29486 3666 29538
rect 6862 29486 6914 29538
rect 10334 29486 10386 29538
rect 11230 29486 11282 29538
rect 20190 29486 20242 29538
rect 20414 29486 20466 29538
rect 21086 29486 21138 29538
rect 1710 29374 1762 29426
rect 2830 29374 2882 29426
rect 6078 29374 6130 29426
rect 10446 29374 10498 29426
rect 10894 29374 10946 29426
rect 12798 29374 12850 29426
rect 17390 29374 17442 29426
rect 17950 29374 18002 29426
rect 18846 29374 18898 29426
rect 19854 29374 19906 29426
rect 24670 29374 24722 29426
rect 28142 29374 28194 29426
rect 2494 29262 2546 29314
rect 5742 29262 5794 29314
rect 8990 29262 9042 29314
rect 9662 29262 9714 29314
rect 13582 29262 13634 29314
rect 15710 29262 15762 29314
rect 16606 29262 16658 29314
rect 19294 29262 19346 29314
rect 21422 29262 21474 29314
rect 21758 29262 21810 29314
rect 23886 29262 23938 29314
rect 25230 29262 25282 29314
rect 27358 29262 27410 29314
rect 18510 29150 18562 29202
rect 18846 29150 18898 29202
rect 19070 29150 19122 29202
rect 19630 29150 19682 29202
rect 4616 28982 4668 29034
rect 4720 28982 4772 29034
rect 4824 28982 4876 29034
rect 11420 28982 11472 29034
rect 11524 28982 11576 29034
rect 11628 28982 11680 29034
rect 18224 28982 18276 29034
rect 18328 28982 18380 29034
rect 18432 28982 18484 29034
rect 25028 28982 25080 29034
rect 25132 28982 25184 29034
rect 25236 28982 25288 29034
rect 2046 28814 2098 28866
rect 2270 28814 2322 28866
rect 3838 28814 3890 28866
rect 5966 28814 6018 28866
rect 6414 28814 6466 28866
rect 20414 28814 20466 28866
rect 2046 28702 2098 28754
rect 2718 28702 2770 28754
rect 3502 28702 3554 28754
rect 4286 28702 4338 28754
rect 5182 28702 5234 28754
rect 5966 28702 6018 28754
rect 6414 28702 6466 28754
rect 6862 28702 6914 28754
rect 7310 28702 7362 28754
rect 12462 28702 12514 28754
rect 12910 28702 12962 28754
rect 13806 28702 13858 28754
rect 14814 28702 14866 28754
rect 15710 28702 15762 28754
rect 19742 28702 19794 28754
rect 21870 28702 21922 28754
rect 24670 28702 24722 28754
rect 27134 28702 27186 28754
rect 27470 28702 27522 28754
rect 2382 28590 2434 28642
rect 2942 28590 2994 28642
rect 4174 28590 4226 28642
rect 11230 28590 11282 28642
rect 14030 28590 14082 28642
rect 14142 28590 14194 28642
rect 14254 28590 14306 28642
rect 14926 28590 14978 28642
rect 15150 28590 15202 28642
rect 16046 28590 16098 28642
rect 16942 28590 16994 28642
rect 20302 28590 20354 28642
rect 23662 28590 23714 28642
rect 24222 28590 24274 28642
rect 24446 28590 24498 28642
rect 24782 28590 24834 28642
rect 25006 28590 25058 28642
rect 25230 28590 25282 28642
rect 25454 28590 25506 28642
rect 25678 28590 25730 28642
rect 26462 28590 26514 28642
rect 3166 28478 3218 28530
rect 3614 28478 3666 28530
rect 13694 28478 13746 28530
rect 17614 28478 17666 28530
rect 20750 28478 20802 28530
rect 26126 28478 26178 28530
rect 26350 28478 26402 28530
rect 2382 28366 2434 28418
rect 11790 28366 11842 28418
rect 20526 28366 20578 28418
rect 26574 28366 26626 28418
rect 28142 28366 28194 28418
rect 8018 28198 8070 28250
rect 8122 28198 8174 28250
rect 8226 28198 8278 28250
rect 14822 28198 14874 28250
rect 14926 28198 14978 28250
rect 15030 28198 15082 28250
rect 21626 28198 21678 28250
rect 21730 28198 21782 28250
rect 21834 28198 21886 28250
rect 28430 28198 28482 28250
rect 28534 28198 28586 28250
rect 28638 28198 28690 28250
rect 5070 28030 5122 28082
rect 6638 28030 6690 28082
rect 11454 28030 11506 28082
rect 11566 28030 11618 28082
rect 14254 28030 14306 28082
rect 15710 28030 15762 28082
rect 17726 28030 17778 28082
rect 23998 28030 24050 28082
rect 24670 28030 24722 28082
rect 25678 28030 25730 28082
rect 26686 28030 26738 28082
rect 2494 27918 2546 27970
rect 10222 27918 10274 27970
rect 10446 27918 10498 27970
rect 10782 27918 10834 27970
rect 11006 27918 11058 27970
rect 17838 27918 17890 27970
rect 25902 27918 25954 27970
rect 26126 27918 26178 27970
rect 27134 27918 27186 27970
rect 27358 27918 27410 27970
rect 27806 27918 27858 27970
rect 1822 27806 1874 27858
rect 8990 27806 9042 27858
rect 11342 27806 11394 27858
rect 12014 27806 12066 27858
rect 14926 27806 14978 27858
rect 17614 27806 17666 27858
rect 18174 27806 18226 27858
rect 19630 27806 19682 27858
rect 22878 27806 22930 27858
rect 23102 27806 23154 27858
rect 23326 27806 23378 27858
rect 23550 27806 23602 27858
rect 26462 27806 26514 27858
rect 4622 27694 4674 27746
rect 9662 27694 9714 27746
rect 10558 27694 10610 27746
rect 12350 27694 12402 27746
rect 12798 27694 12850 27746
rect 15262 27694 15314 27746
rect 16158 27694 16210 27746
rect 16942 27694 16994 27746
rect 18846 27694 18898 27746
rect 19294 27694 19346 27746
rect 20414 27694 20466 27746
rect 22542 27694 22594 27746
rect 22990 27694 23042 27746
rect 14926 27582 14978 27634
rect 18174 27582 18226 27634
rect 26350 27582 26402 27634
rect 27022 27582 27074 27634
rect 4616 27414 4668 27466
rect 4720 27414 4772 27466
rect 4824 27414 4876 27466
rect 11420 27414 11472 27466
rect 11524 27414 11576 27466
rect 11628 27414 11680 27466
rect 18224 27414 18276 27466
rect 18328 27414 18380 27466
rect 18432 27414 18484 27466
rect 25028 27414 25080 27466
rect 25132 27414 25184 27466
rect 25236 27414 25288 27466
rect 8542 27246 8594 27298
rect 17950 27246 18002 27298
rect 18510 27246 18562 27298
rect 2494 27134 2546 27186
rect 3838 27134 3890 27186
rect 4286 27134 4338 27186
rect 5070 27134 5122 27186
rect 5630 27134 5682 27186
rect 5966 27134 6018 27186
rect 6414 27134 6466 27186
rect 6862 27134 6914 27186
rect 7758 27134 7810 27186
rect 10334 27134 10386 27186
rect 12462 27134 12514 27186
rect 12910 27134 12962 27186
rect 16382 27134 16434 27186
rect 16830 27134 16882 27186
rect 19070 27134 19122 27186
rect 20302 27134 20354 27186
rect 22318 27134 22370 27186
rect 23998 27134 24050 27186
rect 24670 27246 24722 27298
rect 24446 27134 24498 27186
rect 25230 27134 25282 27186
rect 27358 27134 27410 27186
rect 2942 27022 2994 27074
rect 6750 27022 6802 27074
rect 8318 27022 8370 27074
rect 8878 27022 8930 27074
rect 9662 27022 9714 27074
rect 13582 27022 13634 27074
rect 18622 27022 18674 27074
rect 1710 26910 1762 26962
rect 5854 26910 5906 26962
rect 8094 26966 8146 27018
rect 20414 27022 20466 27074
rect 23662 27022 23714 27074
rect 28142 27022 28194 27074
rect 14254 26910 14306 26962
rect 18286 26910 18338 26962
rect 20190 26910 20242 26962
rect 20750 26910 20802 26962
rect 2046 26798 2098 26850
rect 3390 26798 3442 26850
rect 6302 26798 6354 26850
rect 8206 26798 8258 26850
rect 19854 26798 19906 26850
rect 24894 26798 24946 26850
rect 8018 26630 8070 26682
rect 8122 26630 8174 26682
rect 8226 26630 8278 26682
rect 14822 26630 14874 26682
rect 14926 26630 14978 26682
rect 15030 26630 15082 26682
rect 21626 26630 21678 26682
rect 21730 26630 21782 26682
rect 21834 26630 21886 26682
rect 28430 26630 28482 26682
rect 28534 26630 28586 26682
rect 28638 26630 28690 26682
rect 2830 26462 2882 26514
rect 9662 26462 9714 26514
rect 12574 26462 12626 26514
rect 13470 26462 13522 26514
rect 14254 26462 14306 26514
rect 15262 26462 15314 26514
rect 15710 26462 15762 26514
rect 16382 26462 16434 26514
rect 20190 26462 20242 26514
rect 21310 26462 21362 26514
rect 21422 26462 21474 26514
rect 21534 26462 21586 26514
rect 23886 26462 23938 26514
rect 24334 26462 24386 26514
rect 25230 26462 25282 26514
rect 26238 26462 26290 26514
rect 26910 26462 26962 26514
rect 27358 26462 27410 26514
rect 3390 26350 3442 26402
rect 6078 26350 6130 26402
rect 13358 26350 13410 26402
rect 14030 26350 14082 26402
rect 17390 26350 17442 26402
rect 19294 26350 19346 26402
rect 19742 26350 19794 26402
rect 4958 26238 5010 26290
rect 9886 26238 9938 26290
rect 10782 26238 10834 26290
rect 12798 26238 12850 26290
rect 13134 26238 13186 26290
rect 14366 26238 14418 26290
rect 14814 26238 14866 26290
rect 17614 26238 17666 26290
rect 18174 26238 18226 26290
rect 18510 26238 18562 26290
rect 21982 26238 22034 26290
rect 22654 26238 22706 26290
rect 25454 26238 25506 26290
rect 25902 26238 25954 26290
rect 10334 26126 10386 26178
rect 12126 26126 12178 26178
rect 16830 26126 16882 26178
rect 17502 26126 17554 26178
rect 20974 26126 21026 26178
rect 22318 26126 22370 26178
rect 22766 26126 22818 26178
rect 23438 26126 23490 26178
rect 25342 26126 25394 26178
rect 28142 26126 28194 26178
rect 9550 26014 9602 26066
rect 14590 26014 14642 26066
rect 15150 26014 15202 26066
rect 15822 26014 15874 26066
rect 17838 26014 17890 26066
rect 18510 26014 18562 26066
rect 18846 26014 18898 26066
rect 22990 26014 23042 26066
rect 4616 25846 4668 25898
rect 4720 25846 4772 25898
rect 4824 25846 4876 25898
rect 11420 25846 11472 25898
rect 11524 25846 11576 25898
rect 11628 25846 11680 25898
rect 18224 25846 18276 25898
rect 18328 25846 18380 25898
rect 18432 25846 18484 25898
rect 25028 25846 25080 25898
rect 25132 25846 25184 25898
rect 25236 25846 25288 25898
rect 2494 25678 2546 25730
rect 5966 25678 6018 25730
rect 2270 25566 2322 25618
rect 5070 25566 5122 25618
rect 7870 25566 7922 25618
rect 9998 25566 10050 25618
rect 12910 25566 12962 25618
rect 13806 25566 13858 25618
rect 16718 25566 16770 25618
rect 18846 25566 18898 25618
rect 20190 25566 20242 25618
rect 20750 25566 20802 25618
rect 21646 25566 21698 25618
rect 24894 25566 24946 25618
rect 3502 25454 3554 25506
rect 4062 25454 4114 25506
rect 5742 25454 5794 25506
rect 6190 25454 6242 25506
rect 6414 25454 6466 25506
rect 7198 25454 7250 25506
rect 14142 25454 14194 25506
rect 16046 25454 16098 25506
rect 19294 25454 19346 25506
rect 24558 25454 24610 25506
rect 27806 25454 27858 25506
rect 2718 25342 2770 25394
rect 4622 25342 4674 25394
rect 14478 25342 14530 25394
rect 23774 25342 23826 25394
rect 27022 25342 27074 25394
rect 2606 25230 2658 25282
rect 5630 25230 5682 25282
rect 10446 25230 10498 25282
rect 14366 25230 14418 25282
rect 14926 25230 14978 25282
rect 15374 25230 15426 25282
rect 19742 25230 19794 25282
rect 8018 25062 8070 25114
rect 8122 25062 8174 25114
rect 8226 25062 8278 25114
rect 14822 25062 14874 25114
rect 14926 25062 14978 25114
rect 15030 25062 15082 25114
rect 21626 25062 21678 25114
rect 21730 25062 21782 25114
rect 21834 25062 21886 25114
rect 28430 25062 28482 25114
rect 28534 25062 28586 25114
rect 28638 25062 28690 25114
rect 2382 24894 2434 24946
rect 7758 24894 7810 24946
rect 8990 24894 9042 24946
rect 14254 24894 14306 24946
rect 15150 24894 15202 24946
rect 15710 24894 15762 24946
rect 16942 24894 16994 24946
rect 18734 24894 18786 24946
rect 20190 24894 20242 24946
rect 20974 24894 21026 24946
rect 21198 24894 21250 24946
rect 22990 24894 23042 24946
rect 25678 24894 25730 24946
rect 3614 24782 3666 24834
rect 5182 24782 5234 24834
rect 16270 24782 16322 24834
rect 19630 24782 19682 24834
rect 20078 24782 20130 24834
rect 20414 24782 20466 24834
rect 20862 24782 20914 24834
rect 25454 24782 25506 24834
rect 2046 24670 2098 24722
rect 2382 24670 2434 24722
rect 2942 24670 2994 24722
rect 3166 24670 3218 24722
rect 3502 24670 3554 24722
rect 4062 24670 4114 24722
rect 4510 24670 4562 24722
rect 9662 24670 9714 24722
rect 13358 24670 13410 24722
rect 16158 24670 16210 24722
rect 16606 24670 16658 24722
rect 19854 24670 19906 24722
rect 20638 24670 20690 24722
rect 21422 24670 21474 24722
rect 21646 24670 21698 24722
rect 22206 24670 22258 24722
rect 22542 24670 22594 24722
rect 22878 24670 22930 24722
rect 25342 24670 25394 24722
rect 25902 24670 25954 24722
rect 7310 24558 7362 24610
rect 10334 24558 10386 24610
rect 12462 24558 12514 24610
rect 12910 24558 12962 24610
rect 14702 24558 14754 24610
rect 15934 24558 15986 24610
rect 17614 24558 17666 24610
rect 17950 24558 18002 24610
rect 18398 24558 18450 24610
rect 19294 24558 19346 24610
rect 21534 24558 21586 24610
rect 23438 24558 23490 24610
rect 24222 24558 24274 24610
rect 24670 24558 24722 24610
rect 26238 24558 26290 24610
rect 26910 24558 26962 24610
rect 27358 24558 27410 24610
rect 28142 24558 28194 24610
rect 2606 24446 2658 24498
rect 14254 24446 14306 24498
rect 14926 24446 14978 24498
rect 19070 24446 19122 24498
rect 22766 24446 22818 24498
rect 23102 24446 23154 24498
rect 23438 24446 23490 24498
rect 4616 24278 4668 24330
rect 4720 24278 4772 24330
rect 4824 24278 4876 24330
rect 11420 24278 11472 24330
rect 11524 24278 11576 24330
rect 11628 24278 11680 24330
rect 18224 24278 18276 24330
rect 18328 24278 18380 24330
rect 18432 24278 18484 24330
rect 25028 24278 25080 24330
rect 25132 24278 25184 24330
rect 25236 24278 25288 24330
rect 15822 24110 15874 24162
rect 16606 24110 16658 24162
rect 16942 24110 16994 24162
rect 18510 24110 18562 24162
rect 22094 24110 22146 24162
rect 22878 24110 22930 24162
rect 2494 23998 2546 24050
rect 4622 23998 4674 24050
rect 5742 23998 5794 24050
rect 8990 24024 9042 24076
rect 9774 23998 9826 24050
rect 12798 23998 12850 24050
rect 13470 23998 13522 24050
rect 14030 23998 14082 24050
rect 19294 23998 19346 24050
rect 20190 23998 20242 24050
rect 20638 23998 20690 24050
rect 21422 23998 21474 24050
rect 24558 23998 24610 24050
rect 25342 23998 25394 24050
rect 27246 23998 27298 24050
rect 27694 23998 27746 24050
rect 1822 23886 1874 23938
rect 6078 23886 6130 23938
rect 10110 23886 10162 23938
rect 10446 23886 10498 23938
rect 11230 23886 11282 23938
rect 11566 23886 11618 23938
rect 11790 23886 11842 23938
rect 12350 23886 12402 23938
rect 13694 23886 13746 23938
rect 14478 23886 14530 23938
rect 14926 23886 14978 23938
rect 16718 23886 16770 23938
rect 19854 23886 19906 23938
rect 26238 23886 26290 23938
rect 26350 23886 26402 23938
rect 6862 23774 6914 23826
rect 10670 23774 10722 23826
rect 11678 23774 11730 23826
rect 12014 23774 12066 23826
rect 12686 23774 12738 23826
rect 15150 23774 15202 23826
rect 15710 23774 15762 23826
rect 16270 23774 16322 23826
rect 17502 23774 17554 23826
rect 17950 23774 18002 23826
rect 18398 23774 18450 23826
rect 26574 23774 26626 23826
rect 26798 23774 26850 23826
rect 5070 23662 5122 23714
rect 10334 23662 10386 23714
rect 12910 23662 12962 23714
rect 14702 23662 14754 23714
rect 15822 23662 15874 23714
rect 16494 23662 16546 23714
rect 17054 23662 17106 23714
rect 17278 23662 17330 23714
rect 18174 23662 18226 23714
rect 18846 23662 18898 23714
rect 19294 23662 19346 23714
rect 19518 23662 19570 23714
rect 21870 23662 21922 23714
rect 22318 23662 22370 23714
rect 22766 23662 22818 23714
rect 23214 23662 23266 23714
rect 23998 23662 24050 23714
rect 25006 23662 25058 23714
rect 26686 23662 26738 23714
rect 28142 23662 28194 23714
rect 8018 23494 8070 23546
rect 8122 23494 8174 23546
rect 8226 23494 8278 23546
rect 14822 23494 14874 23546
rect 14926 23494 14978 23546
rect 15030 23494 15082 23546
rect 21626 23494 21678 23546
rect 21730 23494 21782 23546
rect 21834 23494 21886 23546
rect 28430 23494 28482 23546
rect 28534 23494 28586 23546
rect 28638 23494 28690 23546
rect 2046 23326 2098 23378
rect 3166 23326 3218 23378
rect 4622 23326 4674 23378
rect 6974 23326 7026 23378
rect 10894 23326 10946 23378
rect 12686 23326 12738 23378
rect 12798 23326 12850 23378
rect 13246 23326 13298 23378
rect 17614 23326 17666 23378
rect 20078 23326 20130 23378
rect 23214 23326 23266 23378
rect 23662 23326 23714 23378
rect 3838 23214 3890 23266
rect 6638 23214 6690 23266
rect 7534 23214 7586 23266
rect 8654 23214 8706 23266
rect 8878 23214 8930 23266
rect 14254 23214 14306 23266
rect 22430 23214 22482 23266
rect 22654 23214 22706 23266
rect 23774 23214 23826 23266
rect 1710 23102 1762 23154
rect 3390 23102 3442 23154
rect 4510 23102 4562 23154
rect 7198 23102 7250 23154
rect 7758 23102 7810 23154
rect 8542 23102 8594 23154
rect 12238 23102 12290 23154
rect 12462 23102 12514 23154
rect 13582 23102 13634 23154
rect 20526 23102 20578 23154
rect 20750 23102 20802 23154
rect 22990 23102 23042 23154
rect 23998 23102 24050 23154
rect 24222 23102 24274 23154
rect 27358 23102 27410 23154
rect 28030 23102 28082 23154
rect 2718 22990 2770 23042
rect 5518 22990 5570 23042
rect 6190 22990 6242 23042
rect 8318 22990 8370 23042
rect 8990 22990 9042 23042
rect 11902 22990 11954 23042
rect 16382 22990 16434 23042
rect 16830 22990 16882 23042
rect 17950 22990 18002 23042
rect 18622 22990 18674 23042
rect 19070 22990 19122 23042
rect 19518 22990 19570 23042
rect 21198 22990 21250 23042
rect 21870 22990 21922 23042
rect 23886 22990 23938 23042
rect 24670 22990 24722 23042
rect 25230 22990 25282 23042
rect 3054 22878 3106 22930
rect 3726 22878 3778 22930
rect 7310 22878 7362 22930
rect 8206 22878 8258 22930
rect 18622 22878 18674 22930
rect 18958 22878 19010 22930
rect 20414 22878 20466 22930
rect 21870 22878 21922 22930
rect 22206 22878 22258 22930
rect 22990 22878 23042 22930
rect 4616 22710 4668 22762
rect 4720 22710 4772 22762
rect 4824 22710 4876 22762
rect 11420 22710 11472 22762
rect 11524 22710 11576 22762
rect 11628 22710 11680 22762
rect 18224 22710 18276 22762
rect 18328 22710 18380 22762
rect 18432 22710 18484 22762
rect 25028 22710 25080 22762
rect 25132 22710 25184 22762
rect 25236 22710 25288 22762
rect 20190 22542 20242 22594
rect 4622 22430 4674 22482
rect 8878 22430 8930 22482
rect 10222 22430 10274 22482
rect 11006 22430 11058 22482
rect 13022 22430 13074 22482
rect 13694 22430 13746 22482
rect 15710 22430 15762 22482
rect 16606 22430 16658 22482
rect 18622 22430 18674 22482
rect 21870 22430 21922 22482
rect 22318 22430 22370 22482
rect 24558 22430 24610 22482
rect 25006 22430 25058 22482
rect 26910 22430 26962 22482
rect 1822 22318 1874 22370
rect 15822 22318 15874 22370
rect 17054 22318 17106 22370
rect 19070 22318 19122 22370
rect 19854 22318 19906 22370
rect 20302 22318 20354 22370
rect 23214 22318 23266 22370
rect 23662 22318 23714 22370
rect 25230 22318 25282 22370
rect 26014 22318 26066 22370
rect 2494 22206 2546 22258
rect 10446 22206 10498 22258
rect 16046 22206 16098 22258
rect 19630 22206 19682 22258
rect 23998 22206 24050 22258
rect 24894 22206 24946 22258
rect 5070 22094 5122 22146
rect 7982 22094 8034 22146
rect 10334 22094 10386 22146
rect 15598 22094 15650 22146
rect 17502 22094 17554 22146
rect 18174 22094 18226 22146
rect 19742 22094 19794 22146
rect 21422 22094 21474 22146
rect 22878 22094 22930 22146
rect 22990 22094 23042 22146
rect 8018 21926 8070 21978
rect 8122 21926 8174 21978
rect 8226 21926 8278 21978
rect 14822 21926 14874 21978
rect 14926 21926 14978 21978
rect 15030 21926 15082 21978
rect 21626 21926 21678 21978
rect 21730 21926 21782 21978
rect 21834 21926 21886 21978
rect 28430 21926 28482 21978
rect 28534 21926 28586 21978
rect 28638 21926 28690 21978
rect 2718 21758 2770 21810
rect 3950 21758 4002 21810
rect 4398 21758 4450 21810
rect 12910 21758 12962 21810
rect 13358 21758 13410 21810
rect 17950 21758 18002 21810
rect 24334 21758 24386 21810
rect 2046 21646 2098 21698
rect 3278 21646 3330 21698
rect 8430 21646 8482 21698
rect 8654 21646 8706 21698
rect 14478 21646 14530 21698
rect 19742 21646 19794 21698
rect 24222 21646 24274 21698
rect 1822 21534 1874 21586
rect 2718 21534 2770 21586
rect 3054 21534 3106 21586
rect 3502 21534 3554 21586
rect 5070 21534 5122 21586
rect 9662 21534 9714 21586
rect 17614 21534 17666 21586
rect 18958 21534 19010 21586
rect 22766 21534 22818 21586
rect 26014 21534 26066 21586
rect 5854 21422 5906 21474
rect 7982 21422 8034 21474
rect 10334 21422 10386 21474
rect 12462 21422 12514 21474
rect 14254 21422 14306 21474
rect 14366 21422 14418 21474
rect 15038 21422 15090 21474
rect 15486 21422 15538 21474
rect 18398 21422 18450 21474
rect 21870 21422 21922 21474
rect 23438 21422 23490 21474
rect 27022 21422 27074 21474
rect 8318 21310 8370 21362
rect 24446 21310 24498 21362
rect 4616 21142 4668 21194
rect 4720 21142 4772 21194
rect 4824 21142 4876 21194
rect 11420 21142 11472 21194
rect 11524 21142 11576 21194
rect 11628 21142 11680 21194
rect 18224 21142 18276 21194
rect 18328 21142 18380 21194
rect 18432 21142 18484 21194
rect 25028 21142 25080 21194
rect 25132 21142 25184 21194
rect 25236 21142 25288 21194
rect 3054 20974 3106 21026
rect 1822 20862 1874 20914
rect 2382 20862 2434 20914
rect 2718 20750 2770 20802
rect 3502 20750 3554 20802
rect 3614 20750 3666 20802
rect 4286 20974 4338 21026
rect 4846 20974 4898 21026
rect 5854 20974 5906 21026
rect 6414 20974 6466 21026
rect 6862 20974 6914 21026
rect 9998 20974 10050 21026
rect 11006 20974 11058 21026
rect 11678 20974 11730 21026
rect 12014 20974 12066 21026
rect 12238 20974 12290 21026
rect 12462 20974 12514 21026
rect 14030 20974 14082 21026
rect 19518 20974 19570 21026
rect 20078 20974 20130 21026
rect 26350 20974 26402 21026
rect 27134 20974 27186 21026
rect 27470 20974 27522 21026
rect 4846 20862 4898 20914
rect 8206 20862 8258 20914
rect 9102 20862 9154 20914
rect 12462 20862 12514 20914
rect 12910 20862 12962 20914
rect 14926 20862 14978 20914
rect 18622 20862 18674 20914
rect 23326 20862 23378 20914
rect 25454 20862 25506 20914
rect 6638 20750 6690 20802
rect 8654 20750 8706 20802
rect 9774 20750 9826 20802
rect 10222 20750 10274 20802
rect 10782 20750 10834 20802
rect 11342 20750 11394 20802
rect 14254 20750 14306 20802
rect 15822 20750 15874 20802
rect 18958 20750 19010 20802
rect 19182 20750 19234 20802
rect 19518 20750 19570 20802
rect 20078 20750 20130 20802
rect 22654 20750 22706 20802
rect 26126 20750 26178 20802
rect 26350 20750 26402 20802
rect 27134 20750 27186 20802
rect 6190 20638 6242 20690
rect 7086 20638 7138 20690
rect 7310 20638 7362 20690
rect 7758 20638 7810 20690
rect 9438 20638 9490 20690
rect 10558 20638 10610 20690
rect 11790 20638 11842 20690
rect 13470 20638 13522 20690
rect 13694 20638 13746 20690
rect 16494 20638 16546 20690
rect 20414 20638 20466 20690
rect 25790 20638 25842 20690
rect 2942 20526 2994 20578
rect 3390 20526 3442 20578
rect 3950 20526 4002 20578
rect 4398 20526 4450 20578
rect 5742 20526 5794 20578
rect 6526 20526 6578 20578
rect 10222 20526 10274 20578
rect 10670 20526 10722 20578
rect 13582 20526 13634 20578
rect 15374 20526 15426 20578
rect 19070 20526 19122 20578
rect 21422 20526 21474 20578
rect 22094 20526 22146 20578
rect 25902 20526 25954 20578
rect 27918 20526 27970 20578
rect 8018 20358 8070 20410
rect 8122 20358 8174 20410
rect 8226 20358 8278 20410
rect 14822 20358 14874 20410
rect 14926 20358 14978 20410
rect 15030 20358 15082 20410
rect 21626 20358 21678 20410
rect 21730 20358 21782 20410
rect 21834 20358 21886 20410
rect 28430 20358 28482 20410
rect 28534 20358 28586 20410
rect 28638 20358 28690 20410
rect 2494 20190 2546 20242
rect 7198 20190 7250 20242
rect 10446 20190 10498 20242
rect 11454 20190 11506 20242
rect 11678 20190 11730 20242
rect 3054 20078 3106 20130
rect 3278 20078 3330 20130
rect 5406 20078 5458 20130
rect 8878 20078 8930 20130
rect 9998 20078 10050 20130
rect 2606 19966 2658 20018
rect 2830 19966 2882 20018
rect 3950 19966 4002 20018
rect 4958 19854 5010 19906
rect 8318 19854 8370 19906
rect 4510 19742 4562 19794
rect 16494 20190 16546 20242
rect 23102 20190 23154 20242
rect 11902 20078 11954 20130
rect 13022 20078 13074 20130
rect 15710 20078 15762 20130
rect 16046 20078 16098 20130
rect 23662 20078 23714 20130
rect 24670 20078 24722 20130
rect 26014 20078 26066 20130
rect 12350 19966 12402 20018
rect 16270 19966 16322 20018
rect 16606 19966 16658 20018
rect 17614 19966 17666 20018
rect 25342 19966 25394 20018
rect 15150 19854 15202 19906
rect 19406 19854 19458 19906
rect 24110 19854 24162 19906
rect 28142 19854 28194 19906
rect 11902 19742 11954 19794
rect 16606 19742 16658 19794
rect 4616 19574 4668 19626
rect 4720 19574 4772 19626
rect 4824 19574 4876 19626
rect 11420 19574 11472 19626
rect 11524 19574 11576 19626
rect 11628 19574 11680 19626
rect 18224 19574 18276 19626
rect 18328 19574 18380 19626
rect 18432 19574 18484 19626
rect 25028 19574 25080 19626
rect 25132 19574 25184 19626
rect 25236 19574 25288 19626
rect 18174 19406 18226 19458
rect 2494 19294 2546 19346
rect 4622 19294 4674 19346
rect 8654 19294 8706 19346
rect 9774 19294 9826 19346
rect 11902 19294 11954 19346
rect 12462 19294 12514 19346
rect 12910 19294 12962 19346
rect 15374 19294 15426 19346
rect 17054 19294 17106 19346
rect 18286 19294 18338 19346
rect 20526 19294 20578 19346
rect 22654 19294 22706 19346
rect 23102 19294 23154 19346
rect 27022 19294 27074 19346
rect 28030 19294 28082 19346
rect 1822 19182 1874 19234
rect 6078 19182 6130 19234
rect 6414 19182 6466 19234
rect 6638 19182 6690 19234
rect 7758 19182 7810 19234
rect 8206 19182 8258 19234
rect 8990 19182 9042 19234
rect 13358 19182 13410 19234
rect 13806 19182 13858 19234
rect 13918 19182 13970 19234
rect 14590 19182 14642 19234
rect 16046 19182 16098 19234
rect 16494 19182 16546 19234
rect 18510 19182 18562 19234
rect 19518 19182 19570 19234
rect 19742 19182 19794 19234
rect 20078 19182 20130 19234
rect 21646 19182 21698 19234
rect 21870 19182 21922 19234
rect 22318 19182 22370 19234
rect 25902 19182 25954 19234
rect 6974 19070 7026 19122
rect 15598 19070 15650 19122
rect 21758 19070 21810 19122
rect 25230 19070 25282 19122
rect 5070 18958 5122 19010
rect 6526 18958 6578 19010
rect 7534 18958 7586 19010
rect 7646 18958 7698 19010
rect 13582 18958 13634 19010
rect 14702 18958 14754 19010
rect 17502 18958 17554 19010
rect 18958 18958 19010 19010
rect 19630 18958 19682 19010
rect 26462 18958 26514 19010
rect 27358 18958 27410 19010
rect 8018 18790 8070 18842
rect 8122 18790 8174 18842
rect 8226 18790 8278 18842
rect 14822 18790 14874 18842
rect 14926 18790 14978 18842
rect 15030 18790 15082 18842
rect 21626 18790 21678 18842
rect 21730 18790 21782 18842
rect 21834 18790 21886 18842
rect 28430 18790 28482 18842
rect 28534 18790 28586 18842
rect 28638 18790 28690 18842
rect 3278 18622 3330 18674
rect 8990 18622 9042 18674
rect 25342 18622 25394 18674
rect 26126 18622 26178 18674
rect 26350 18622 26402 18674
rect 2046 18510 2098 18562
rect 5966 18510 6018 18562
rect 1710 18398 1762 18450
rect 3726 18398 3778 18450
rect 5182 18398 5234 18450
rect 8542 18398 8594 18450
rect 11566 18398 11618 18450
rect 18510 18398 18562 18450
rect 19182 18398 19234 18450
rect 23998 18398 24050 18450
rect 24670 18398 24722 18450
rect 25230 18398 25282 18450
rect 25454 18398 25506 18450
rect 25678 18398 25730 18450
rect 26238 18398 26290 18450
rect 26798 18398 26850 18450
rect 28030 18398 28082 18450
rect 2494 18286 2546 18338
rect 8094 18286 8146 18338
rect 11230 18286 11282 18338
rect 13582 18286 13634 18338
rect 17502 18286 17554 18338
rect 17950 18286 18002 18338
rect 21310 18286 21362 18338
rect 22206 18286 22258 18338
rect 27134 18286 27186 18338
rect 27582 18286 27634 18338
rect 27134 18174 27186 18226
rect 27806 18174 27858 18226
rect 4616 18006 4668 18058
rect 4720 18006 4772 18058
rect 4824 18006 4876 18058
rect 11420 18006 11472 18058
rect 11524 18006 11576 18058
rect 11628 18006 11680 18058
rect 18224 18006 18276 18058
rect 18328 18006 18380 18058
rect 18432 18006 18484 18058
rect 25028 18006 25080 18058
rect 25132 18006 25184 18058
rect 25236 18006 25288 18058
rect 2718 17838 2770 17890
rect 12686 17838 12738 17890
rect 12910 17838 12962 17890
rect 3502 17726 3554 17778
rect 8542 17726 8594 17778
rect 8990 17726 9042 17778
rect 10110 17726 10162 17778
rect 12910 17726 12962 17778
rect 13918 17726 13970 17778
rect 15262 17726 15314 17778
rect 16942 17726 16994 17778
rect 20750 17726 20802 17778
rect 21310 17726 21362 17778
rect 25230 17726 25282 17778
rect 27582 17726 27634 17778
rect 4174 17614 4226 17666
rect 5742 17614 5794 17666
rect 10446 17614 10498 17666
rect 10782 17614 10834 17666
rect 11006 17614 11058 17666
rect 11566 17614 11618 17666
rect 11678 17614 11730 17666
rect 12014 17614 12066 17666
rect 14030 17614 14082 17666
rect 14926 17614 14978 17666
rect 15374 17614 15426 17666
rect 15934 17614 15986 17666
rect 16494 17614 16546 17666
rect 17054 17614 17106 17666
rect 17838 17614 17890 17666
rect 24110 17614 24162 17666
rect 26574 17614 26626 17666
rect 2942 17502 2994 17554
rect 6414 17502 6466 17554
rect 13806 17502 13858 17554
rect 14702 17502 14754 17554
rect 16270 17502 16322 17554
rect 18622 17502 18674 17554
rect 23438 17502 23490 17554
rect 2830 17390 2882 17442
rect 3390 17390 3442 17442
rect 4734 17390 4786 17442
rect 9438 17390 9490 17442
rect 10558 17390 10610 17442
rect 11454 17390 11506 17442
rect 12462 17390 12514 17442
rect 14254 17390 14306 17442
rect 15150 17390 15202 17442
rect 16046 17390 16098 17442
rect 16830 17390 16882 17442
rect 17278 17390 17330 17442
rect 28030 17390 28082 17442
rect 8018 17222 8070 17274
rect 8122 17222 8174 17274
rect 8226 17222 8278 17274
rect 14822 17222 14874 17274
rect 14926 17222 14978 17274
rect 15030 17222 15082 17274
rect 21626 17222 21678 17274
rect 21730 17222 21782 17274
rect 21834 17222 21886 17274
rect 28430 17222 28482 17274
rect 28534 17222 28586 17274
rect 28638 17222 28690 17274
rect 5070 17054 5122 17106
rect 6526 17054 6578 17106
rect 7646 17054 7698 17106
rect 7870 17054 7922 17106
rect 8990 17054 9042 17106
rect 9662 17054 9714 17106
rect 10334 17054 10386 17106
rect 11230 17054 11282 17106
rect 11678 17054 11730 17106
rect 15934 17054 15986 17106
rect 16718 17054 16770 17106
rect 18062 17054 18114 17106
rect 18510 17054 18562 17106
rect 18958 17054 19010 17106
rect 20302 17054 20354 17106
rect 20750 17054 20802 17106
rect 21310 17054 21362 17106
rect 23102 17054 23154 17106
rect 23550 17054 23602 17106
rect 24334 17054 24386 17106
rect 24670 17054 24722 17106
rect 6974 16942 7026 16994
rect 7758 16942 7810 16994
rect 12798 16942 12850 16994
rect 16270 16942 16322 16994
rect 18846 16942 18898 16994
rect 19182 16942 19234 16994
rect 19406 16942 19458 16994
rect 21198 16942 21250 16994
rect 22654 16942 22706 16994
rect 26350 16942 26402 16994
rect 1822 16830 1874 16882
rect 6078 16830 6130 16882
rect 6302 16830 6354 16882
rect 6750 16830 6802 16882
rect 8318 16830 8370 16882
rect 10782 16830 10834 16882
rect 12126 16830 12178 16882
rect 15374 16830 15426 16882
rect 17614 16830 17666 16882
rect 21534 16830 21586 16882
rect 21646 16830 21698 16882
rect 22206 16830 22258 16882
rect 27582 16830 27634 16882
rect 2494 16718 2546 16770
rect 4622 16718 4674 16770
rect 5294 16718 5346 16770
rect 5630 16718 5682 16770
rect 14926 16718 14978 16770
rect 19854 16718 19906 16770
rect 6078 16606 6130 16658
rect 15262 16606 15314 16658
rect 16494 16606 16546 16658
rect 17278 16606 17330 16658
rect 17838 16606 17890 16658
rect 22206 16606 22258 16658
rect 23214 16606 23266 16658
rect 4616 16438 4668 16490
rect 4720 16438 4772 16490
rect 4824 16438 4876 16490
rect 11420 16438 11472 16490
rect 11524 16438 11576 16490
rect 11628 16438 11680 16490
rect 18224 16438 18276 16490
rect 18328 16438 18380 16490
rect 18432 16438 18484 16490
rect 25028 16438 25080 16490
rect 25132 16438 25184 16490
rect 25236 16438 25288 16490
rect 2830 16270 2882 16322
rect 13582 16270 13634 16322
rect 14142 16270 14194 16322
rect 8878 16158 8930 16210
rect 14142 16158 14194 16210
rect 14590 16158 14642 16210
rect 15822 16158 15874 16210
rect 17950 16158 18002 16210
rect 18398 16158 18450 16210
rect 20750 16158 20802 16210
rect 24110 16158 24162 16210
rect 27022 16158 27074 16210
rect 27582 16158 27634 16210
rect 28142 16158 28194 16210
rect 1822 16046 1874 16098
rect 2606 16046 2658 16098
rect 3054 16046 3106 16098
rect 8206 16046 8258 16098
rect 12574 16046 12626 16098
rect 15150 16046 15202 16098
rect 20302 16046 20354 16098
rect 21310 16046 21362 16098
rect 3278 15934 3330 15986
rect 12798 15934 12850 15986
rect 2046 15822 2098 15874
rect 2494 15822 2546 15874
rect 3726 15822 3778 15874
rect 4174 15822 4226 15874
rect 12350 15822 12402 15874
rect 12462 15822 12514 15874
rect 13694 15822 13746 15874
rect 8018 15654 8070 15706
rect 8122 15654 8174 15706
rect 8226 15654 8278 15706
rect 14822 15654 14874 15706
rect 14926 15654 14978 15706
rect 15030 15654 15082 15706
rect 21626 15654 21678 15706
rect 21730 15654 21782 15706
rect 21834 15654 21886 15706
rect 28430 15654 28482 15706
rect 28534 15654 28586 15706
rect 28638 15654 28690 15706
rect 1822 15486 1874 15538
rect 3054 15486 3106 15538
rect 3502 15486 3554 15538
rect 6078 15486 6130 15538
rect 6526 15486 6578 15538
rect 7758 15486 7810 15538
rect 8990 15486 9042 15538
rect 13022 15486 13074 15538
rect 13358 15486 13410 15538
rect 13582 15486 13634 15538
rect 13806 15486 13858 15538
rect 15374 15486 15426 15538
rect 15598 15486 15650 15538
rect 16158 15486 16210 15538
rect 18958 15486 19010 15538
rect 20638 15486 20690 15538
rect 21758 15486 21810 15538
rect 22206 15486 22258 15538
rect 24222 15486 24274 15538
rect 24334 15486 24386 15538
rect 7422 15374 7474 15426
rect 10334 15374 10386 15426
rect 14254 15374 14306 15426
rect 19742 15374 19794 15426
rect 23774 15374 23826 15426
rect 6862 15262 6914 15314
rect 7982 15262 8034 15314
rect 8318 15262 8370 15314
rect 9662 15262 9714 15314
rect 14478 15262 14530 15314
rect 14814 15262 14866 15314
rect 15150 15262 15202 15314
rect 15262 15262 15314 15314
rect 16606 15262 16658 15314
rect 18734 15262 18786 15314
rect 19294 15262 19346 15314
rect 20190 15262 20242 15314
rect 21982 15262 22034 15314
rect 22654 15262 22706 15314
rect 23214 15262 23266 15314
rect 23326 15262 23378 15314
rect 23550 15262 23602 15314
rect 24110 15262 24162 15314
rect 24670 15262 24722 15314
rect 25790 15262 25842 15314
rect 3950 15150 4002 15202
rect 4398 15150 4450 15202
rect 5630 15150 5682 15202
rect 7870 15150 7922 15202
rect 12462 15150 12514 15202
rect 13470 15150 13522 15202
rect 14366 15150 14418 15202
rect 18846 15150 18898 15202
rect 21198 15150 21250 15202
rect 22094 15150 22146 15202
rect 26350 15150 26402 15202
rect 3166 15038 3218 15090
rect 3950 15038 4002 15090
rect 4616 14870 4668 14922
rect 4720 14870 4772 14922
rect 4824 14870 4876 14922
rect 11420 14870 11472 14922
rect 11524 14870 11576 14922
rect 11628 14870 11680 14922
rect 18224 14870 18276 14922
rect 18328 14870 18380 14922
rect 18432 14870 18484 14922
rect 25028 14870 25080 14922
rect 25132 14870 25184 14922
rect 25236 14870 25288 14922
rect 2046 14590 2098 14642
rect 9438 14590 9490 14642
rect 12686 14590 12738 14642
rect 14366 14590 14418 14642
rect 16494 14590 16546 14642
rect 19854 14590 19906 14642
rect 20750 14590 20802 14642
rect 22430 14590 22482 14642
rect 23550 14590 23602 14642
rect 25678 14590 25730 14642
rect 27022 14590 27074 14642
rect 27806 14590 27858 14642
rect 28142 14590 28194 14642
rect 2270 14478 2322 14530
rect 2606 14478 2658 14530
rect 3614 14478 3666 14530
rect 5070 14478 5122 14530
rect 5518 14478 5570 14530
rect 6190 14478 6242 14530
rect 6638 14478 6690 14530
rect 9886 14478 9938 14530
rect 13694 14478 13746 14530
rect 17054 14478 17106 14530
rect 21198 14478 21250 14530
rect 21534 14478 21586 14530
rect 21870 14478 21922 14530
rect 22766 14478 22818 14530
rect 2830 14366 2882 14418
rect 3054 14366 3106 14418
rect 4622 14366 4674 14418
rect 5966 14366 6018 14418
rect 7310 14366 7362 14418
rect 10558 14366 10610 14418
rect 17726 14366 17778 14418
rect 2606 14254 2658 14306
rect 4174 14254 4226 14306
rect 5742 14254 5794 14306
rect 20302 14254 20354 14306
rect 21422 14254 21474 14306
rect 26126 14254 26178 14306
rect 26574 14254 26626 14306
rect 8018 14086 8070 14138
rect 8122 14086 8174 14138
rect 8226 14086 8278 14138
rect 14822 14086 14874 14138
rect 14926 14086 14978 14138
rect 15030 14086 15082 14138
rect 21626 14086 21678 14138
rect 21730 14086 21782 14138
rect 21834 14086 21886 14138
rect 28430 14086 28482 14138
rect 28534 14086 28586 14138
rect 28638 14086 28690 14138
rect 2270 13918 2322 13970
rect 3278 13918 3330 13970
rect 8542 13918 8594 13970
rect 9662 13918 9714 13970
rect 10670 13918 10722 13970
rect 11566 13918 11618 13970
rect 15262 13918 15314 13970
rect 15710 13918 15762 13970
rect 18174 13918 18226 13970
rect 25454 13918 25506 13970
rect 26686 13918 26738 13970
rect 27134 13918 27186 13970
rect 2718 13806 2770 13858
rect 5294 13806 5346 13858
rect 8766 13806 8818 13858
rect 8990 13806 9042 13858
rect 11118 13806 11170 13858
rect 18622 13806 18674 13858
rect 19070 13806 19122 13858
rect 20974 13806 21026 13858
rect 4510 13694 4562 13746
rect 8094 13694 8146 13746
rect 8318 13694 8370 13746
rect 9550 13694 9602 13746
rect 9774 13694 9826 13746
rect 10110 13694 10162 13746
rect 10446 13694 10498 13746
rect 10782 13694 10834 13746
rect 12014 13694 12066 13746
rect 17950 13694 18002 13746
rect 18398 13694 18450 13746
rect 20190 13694 20242 13746
rect 23550 13694 23602 13746
rect 2494 13582 2546 13634
rect 2830 13582 2882 13634
rect 3390 13582 3442 13634
rect 4174 13582 4226 13634
rect 7422 13582 7474 13634
rect 12686 13582 12738 13634
rect 14814 13582 14866 13634
rect 17726 13582 17778 13634
rect 23102 13582 23154 13634
rect 24222 13582 24274 13634
rect 24670 13582 24722 13634
rect 25790 13582 25842 13634
rect 26238 13582 26290 13634
rect 4616 13302 4668 13354
rect 4720 13302 4772 13354
rect 4824 13302 4876 13354
rect 11420 13302 11472 13354
rect 11524 13302 11576 13354
rect 11628 13302 11680 13354
rect 18224 13302 18276 13354
rect 18328 13302 18380 13354
rect 18432 13302 18484 13354
rect 25028 13302 25080 13354
rect 25132 13302 25184 13354
rect 25236 13302 25288 13354
rect 12014 13134 12066 13186
rect 12686 13134 12738 13186
rect 13022 13134 13074 13186
rect 14366 13134 14418 13186
rect 15038 13134 15090 13186
rect 26462 13134 26514 13186
rect 27022 13134 27074 13186
rect 2494 13022 2546 13074
rect 4622 13022 4674 13074
rect 5070 13022 5122 13074
rect 8094 13022 8146 13074
rect 10894 13022 10946 13074
rect 11342 13022 11394 13074
rect 12238 13022 12290 13074
rect 12686 13022 12738 13074
rect 14590 13022 14642 13074
rect 14926 13022 14978 13074
rect 17054 13022 17106 13074
rect 22094 13022 22146 13074
rect 24446 13022 24498 13074
rect 26238 13022 26290 13074
rect 27022 13022 27074 13074
rect 1822 12910 1874 12962
rect 5518 12910 5570 12962
rect 6974 12910 7026 12962
rect 7198 12910 7250 12962
rect 13470 12910 13522 12962
rect 13694 12910 13746 12962
rect 14142 12910 14194 12962
rect 17614 12910 17666 12962
rect 18958 12910 19010 12962
rect 19742 12910 19794 12962
rect 22766 12910 22818 12962
rect 23438 12910 23490 12962
rect 26574 12910 26626 12962
rect 5966 12798 6018 12850
rect 6190 12798 6242 12850
rect 7086 12798 7138 12850
rect 10110 12798 10162 12850
rect 17390 12798 17442 12850
rect 17950 12798 18002 12850
rect 18398 12798 18450 12850
rect 5742 12686 5794 12738
rect 6638 12686 6690 12738
rect 7422 12686 7474 12738
rect 8542 12686 8594 12738
rect 9326 12686 9378 12738
rect 9662 12686 9714 12738
rect 9774 12686 9826 12738
rect 9886 12686 9938 12738
rect 11790 12686 11842 12738
rect 13806 12686 13858 12738
rect 17502 12686 17554 12738
rect 18286 12686 18338 12738
rect 18510 12686 18562 12738
rect 19294 12686 19346 12738
rect 20190 12686 20242 12738
rect 8018 12518 8070 12570
rect 8122 12518 8174 12570
rect 8226 12518 8278 12570
rect 14822 12518 14874 12570
rect 14926 12518 14978 12570
rect 15030 12518 15082 12570
rect 21626 12518 21678 12570
rect 21730 12518 21782 12570
rect 21834 12518 21886 12570
rect 28430 12518 28482 12570
rect 28534 12518 28586 12570
rect 28638 12518 28690 12570
rect 4062 12350 4114 12402
rect 8206 12350 8258 12402
rect 11454 12350 11506 12402
rect 12014 12350 12066 12402
rect 13246 12350 13298 12402
rect 16382 12350 16434 12402
rect 17726 12350 17778 12402
rect 18174 12350 18226 12402
rect 18958 12350 19010 12402
rect 20974 12350 21026 12402
rect 21758 12350 21810 12402
rect 22990 12350 23042 12402
rect 23550 12350 23602 12402
rect 24110 12350 24162 12402
rect 2046 12238 2098 12290
rect 2382 12238 2434 12290
rect 2606 12238 2658 12290
rect 3390 12238 3442 12290
rect 5182 12238 5234 12290
rect 10558 12238 10610 12290
rect 11006 12238 11058 12290
rect 18734 12238 18786 12290
rect 19854 12238 19906 12290
rect 22206 12238 22258 12290
rect 22542 12238 22594 12290
rect 1710 12126 1762 12178
rect 3054 12126 3106 12178
rect 4510 12126 4562 12178
rect 8990 12126 9042 12178
rect 9662 12126 9714 12178
rect 9774 12126 9826 12178
rect 10222 12126 10274 12178
rect 18622 12126 18674 12178
rect 19518 12126 19570 12178
rect 22094 12126 22146 12178
rect 25230 12126 25282 12178
rect 2606 12014 2658 12066
rect 7310 12014 7362 12066
rect 8542 12014 8594 12066
rect 9998 12014 10050 12066
rect 14366 12014 14418 12066
rect 15262 12014 15314 12066
rect 16830 12014 16882 12066
rect 20526 12014 20578 12066
rect 22430 12014 22482 12066
rect 24670 12014 24722 12066
rect 27134 12014 27186 12066
rect 20414 11902 20466 11954
rect 20862 11902 20914 11954
rect 22766 11902 22818 11954
rect 23438 11902 23490 11954
rect 4616 11734 4668 11786
rect 4720 11734 4772 11786
rect 4824 11734 4876 11786
rect 11420 11734 11472 11786
rect 11524 11734 11576 11786
rect 11628 11734 11680 11786
rect 18224 11734 18276 11786
rect 18328 11734 18380 11786
rect 18432 11734 18484 11786
rect 25028 11734 25080 11786
rect 25132 11734 25184 11786
rect 25236 11734 25288 11786
rect 2606 11566 2658 11618
rect 3950 11566 4002 11618
rect 7198 11454 7250 11506
rect 7646 11454 7698 11506
rect 7870 11454 7922 11506
rect 9998 11454 10050 11506
rect 15822 11454 15874 11506
rect 17054 11454 17106 11506
rect 19182 11454 19234 11506
rect 21310 11454 21362 11506
rect 23438 11454 23490 11506
rect 25790 11454 25842 11506
rect 2270 11342 2322 11394
rect 3054 11342 3106 11394
rect 3390 11342 3442 11394
rect 10670 11342 10722 11394
rect 14478 11342 14530 11394
rect 15934 11342 15986 11394
rect 16382 11342 16434 11394
rect 19630 11342 19682 11394
rect 20078 11342 20130 11394
rect 20190 11342 20242 11394
rect 20750 11342 20802 11394
rect 24110 11342 24162 11394
rect 24670 11342 24722 11394
rect 2830 11230 2882 11282
rect 4286 11230 4338 11282
rect 4958 11230 5010 11282
rect 5070 11230 5122 11282
rect 6302 11230 6354 11282
rect 6526 11230 6578 11282
rect 11230 11230 11282 11282
rect 12910 11230 12962 11282
rect 13582 11230 13634 11282
rect 13918 11230 13970 11282
rect 14142 11230 14194 11282
rect 14702 11230 14754 11282
rect 15822 11230 15874 11282
rect 2046 11118 2098 11170
rect 2606 11118 2658 11170
rect 4398 11118 4450 11170
rect 4510 11118 4562 11170
rect 5966 11118 6018 11170
rect 6414 11118 6466 11170
rect 12014 11118 12066 11170
rect 12462 11118 12514 11170
rect 13806 11118 13858 11170
rect 19854 11118 19906 11170
rect 8018 10950 8070 11002
rect 8122 10950 8174 11002
rect 8226 10950 8278 11002
rect 14822 10950 14874 11002
rect 14926 10950 14978 11002
rect 15030 10950 15082 11002
rect 21626 10950 21678 11002
rect 21730 10950 21782 11002
rect 21834 10950 21886 11002
rect 28430 10950 28482 11002
rect 28534 10950 28586 11002
rect 28638 10950 28690 11002
rect 8654 10782 8706 10834
rect 9886 10782 9938 10834
rect 11678 10782 11730 10834
rect 11902 10782 11954 10834
rect 12126 10782 12178 10834
rect 12798 10782 12850 10834
rect 13582 10782 13634 10834
rect 14590 10782 14642 10834
rect 14702 10782 14754 10834
rect 14926 10782 14978 10834
rect 16382 10782 16434 10834
rect 17950 10782 18002 10834
rect 18622 10782 18674 10834
rect 19630 10782 19682 10834
rect 20302 10782 20354 10834
rect 22318 10782 22370 10834
rect 22430 10782 22482 10834
rect 24110 10782 24162 10834
rect 2270 10670 2322 10722
rect 7758 10670 7810 10722
rect 14030 10670 14082 10722
rect 15710 10670 15762 10722
rect 15934 10670 15986 10722
rect 17614 10670 17666 10722
rect 20862 10670 20914 10722
rect 21646 10670 21698 10722
rect 22654 10670 22706 10722
rect 23214 10670 23266 10722
rect 23662 10670 23714 10722
rect 7310 10558 7362 10610
rect 8094 10558 8146 10610
rect 10222 10558 10274 10610
rect 10446 10558 10498 10610
rect 10782 10558 10834 10610
rect 11118 10558 11170 10610
rect 11790 10558 11842 10610
rect 13806 10558 13858 10610
rect 14478 10558 14530 10610
rect 15262 10558 15314 10610
rect 16270 10558 16322 10610
rect 16494 10558 16546 10610
rect 16830 10558 16882 10610
rect 17390 10558 17442 10610
rect 18510 10558 18562 10610
rect 19966 10558 20018 10610
rect 20302 10558 20354 10610
rect 21198 10558 21250 10610
rect 21310 10558 21362 10610
rect 21422 10558 21474 10610
rect 22206 10558 22258 10610
rect 25566 10558 25618 10610
rect 10670 10446 10722 10498
rect 13358 10446 13410 10498
rect 13694 10446 13746 10498
rect 15486 10446 15538 10498
rect 24558 10446 24610 10498
rect 26350 10446 26402 10498
rect 7646 10334 7698 10386
rect 4616 10166 4668 10218
rect 4720 10166 4772 10218
rect 4824 10166 4876 10218
rect 11420 10166 11472 10218
rect 11524 10166 11576 10218
rect 11628 10166 11680 10218
rect 18224 10166 18276 10218
rect 18328 10166 18380 10218
rect 18432 10166 18484 10218
rect 25028 10166 25080 10218
rect 25132 10166 25184 10218
rect 25236 10166 25288 10218
rect 2494 9886 2546 9938
rect 4622 9886 4674 9938
rect 8766 9886 8818 9938
rect 10446 9886 10498 9938
rect 12574 9886 12626 9938
rect 14254 9886 14306 9938
rect 16382 9886 16434 9938
rect 18622 9886 18674 9938
rect 20750 9912 20802 9964
rect 21534 9886 21586 9938
rect 21982 9886 22034 9938
rect 22990 9886 23042 9938
rect 1822 9774 1874 9826
rect 5966 9774 6018 9826
rect 9774 9774 9826 9826
rect 13470 9774 13522 9826
rect 16718 9774 16770 9826
rect 17054 9774 17106 9826
rect 17838 9774 17890 9826
rect 24894 9774 24946 9826
rect 25566 9774 25618 9826
rect 26014 9774 26066 9826
rect 6638 9662 6690 9714
rect 17390 9662 17442 9714
rect 5070 9550 5122 9602
rect 9214 9550 9266 9602
rect 17054 9550 17106 9602
rect 8018 9382 8070 9434
rect 8122 9382 8174 9434
rect 8226 9382 8278 9434
rect 14822 9382 14874 9434
rect 14926 9382 14978 9434
rect 15030 9382 15082 9434
rect 21626 9382 21678 9434
rect 21730 9382 21782 9434
rect 21834 9382 21886 9434
rect 28430 9382 28482 9434
rect 28534 9382 28586 9434
rect 28638 9382 28690 9434
rect 6526 9214 6578 9266
rect 7534 9214 7586 9266
rect 7870 9214 7922 9266
rect 8878 9214 8930 9266
rect 12462 9214 12514 9266
rect 12798 9214 12850 9266
rect 15038 9214 15090 9266
rect 17614 9214 17666 9266
rect 18062 9214 18114 9266
rect 18174 9214 18226 9266
rect 19070 9214 19122 9266
rect 19518 9214 19570 9266
rect 19966 9214 20018 9266
rect 24222 9214 24274 9266
rect 2382 9102 2434 9154
rect 3166 9102 3218 9154
rect 4510 9102 4562 9154
rect 6302 9102 6354 9154
rect 13134 9102 13186 9154
rect 13694 9102 13746 9154
rect 14142 9102 14194 9154
rect 16830 9102 16882 9154
rect 17950 9102 18002 9154
rect 4398 8990 4450 9042
rect 6078 8990 6130 9042
rect 6526 8990 6578 9042
rect 6638 8990 6690 9042
rect 7758 8990 7810 9042
rect 13358 8990 13410 9042
rect 15486 8990 15538 9042
rect 18622 8990 18674 9042
rect 23438 8990 23490 9042
rect 2158 8878 2210 8930
rect 5518 8878 5570 8930
rect 13246 8878 13298 8930
rect 14702 8878 14754 8930
rect 16158 8878 16210 8930
rect 20974 8878 21026 8930
rect 4616 8598 4668 8650
rect 4720 8598 4772 8650
rect 4824 8598 4876 8650
rect 11420 8598 11472 8650
rect 11524 8598 11576 8650
rect 11628 8598 11680 8650
rect 18224 8598 18276 8650
rect 18328 8598 18380 8650
rect 18432 8598 18484 8650
rect 25028 8598 25080 8650
rect 25132 8598 25184 8650
rect 25236 8598 25288 8650
rect 6862 8430 6914 8482
rect 16942 8430 16994 8482
rect 17166 8430 17218 8482
rect 1822 8318 1874 8370
rect 5070 8318 5122 8370
rect 7534 8318 7586 8370
rect 14254 8318 14306 8370
rect 16382 8318 16434 8370
rect 16942 8318 16994 8370
rect 17390 8318 17442 8370
rect 17838 8318 17890 8370
rect 18174 8318 18226 8370
rect 18846 8318 18898 8370
rect 21422 8318 21474 8370
rect 22654 8318 22706 8370
rect 2270 8206 2322 8258
rect 6638 8206 6690 8258
rect 6862 8206 6914 8258
rect 13582 8206 13634 8258
rect 19294 8206 19346 8258
rect 20078 8206 20130 8258
rect 20638 8206 20690 8258
rect 22094 8206 22146 8258
rect 22318 8206 22370 8258
rect 24558 8206 24610 8258
rect 24782 8206 24834 8258
rect 2942 8094 2994 8146
rect 6302 8094 6354 8146
rect 7422 8094 7474 8146
rect 8094 8094 8146 8146
rect 8206 8094 8258 8146
rect 19742 8094 19794 8146
rect 20302 8094 20354 8146
rect 20750 8094 20802 8146
rect 23998 8094 24050 8146
rect 6078 7982 6130 8034
rect 6750 7982 6802 8034
rect 7646 7982 7698 8034
rect 8654 7982 8706 8034
rect 24446 7982 24498 8034
rect 8018 7814 8070 7866
rect 8122 7814 8174 7866
rect 8226 7814 8278 7866
rect 14822 7814 14874 7866
rect 14926 7814 14978 7866
rect 15030 7814 15082 7866
rect 21626 7814 21678 7866
rect 21730 7814 21782 7866
rect 21834 7814 21886 7866
rect 28430 7814 28482 7866
rect 28534 7814 28586 7866
rect 28638 7814 28690 7866
rect 2046 7646 2098 7698
rect 2830 7646 2882 7698
rect 3726 7646 3778 7698
rect 5070 7646 5122 7698
rect 9662 7646 9714 7698
rect 13582 7646 13634 7698
rect 20638 7646 20690 7698
rect 22766 7646 22818 7698
rect 23214 7646 23266 7698
rect 5518 7534 5570 7586
rect 6862 7534 6914 7586
rect 14702 7534 14754 7586
rect 19854 7534 19906 7586
rect 1710 7422 1762 7474
rect 3278 7422 3330 7474
rect 4734 7422 4786 7474
rect 5182 7422 5234 7474
rect 6190 7422 6242 7474
rect 13918 7422 13970 7474
rect 20526 7422 20578 7474
rect 21198 7422 21250 7474
rect 22430 7422 22482 7474
rect 23662 7422 23714 7474
rect 23774 7422 23826 7474
rect 23886 7422 23938 7474
rect 8990 7310 9042 7362
rect 16830 7310 16882 7362
rect 19070 7310 19122 7362
rect 4958 7198 5010 7250
rect 4616 7030 4668 7082
rect 4720 7030 4772 7082
rect 4824 7030 4876 7082
rect 11420 7030 11472 7082
rect 11524 7030 11576 7082
rect 11628 7030 11680 7082
rect 18224 7030 18276 7082
rect 18328 7030 18380 7082
rect 18432 7030 18484 7082
rect 25028 7030 25080 7082
rect 25132 7030 25184 7082
rect 25236 7030 25288 7082
rect 5854 6862 5906 6914
rect 6302 6862 6354 6914
rect 6638 6862 6690 6914
rect 22430 6862 22482 6914
rect 2494 6750 2546 6802
rect 3390 6750 3442 6802
rect 5854 6750 5906 6802
rect 6638 6750 6690 6802
rect 18958 6750 19010 6802
rect 19518 6750 19570 6802
rect 24670 6750 24722 6802
rect 4734 6638 4786 6690
rect 4846 6638 4898 6690
rect 6190 6638 6242 6690
rect 16158 6638 16210 6690
rect 16830 6638 16882 6690
rect 20078 6638 20130 6690
rect 21646 6638 21698 6690
rect 22094 6638 22146 6690
rect 24446 6638 24498 6690
rect 4398 6526 4450 6578
rect 20526 6526 20578 6578
rect 21310 6526 21362 6578
rect 22542 6526 22594 6578
rect 23886 6526 23938 6578
rect 3838 6414 3890 6466
rect 24894 6414 24946 6466
rect 8018 6246 8070 6298
rect 8122 6246 8174 6298
rect 8226 6246 8278 6298
rect 14822 6246 14874 6298
rect 14926 6246 14978 6298
rect 15030 6246 15082 6298
rect 21626 6246 21678 6298
rect 21730 6246 21782 6298
rect 21834 6246 21886 6298
rect 28430 6246 28482 6298
rect 28534 6246 28586 6298
rect 28638 6246 28690 6298
rect 5182 6078 5234 6130
rect 5854 6078 5906 6130
rect 18734 6078 18786 6130
rect 21422 6078 21474 6130
rect 25454 6078 25506 6130
rect 20078 5966 20130 6018
rect 21870 5966 21922 6018
rect 22542 5966 22594 6018
rect 24222 5966 24274 6018
rect 26014 5966 26066 6018
rect 19854 5854 19906 5906
rect 21758 5854 21810 5906
rect 22990 5854 23042 5906
rect 23102 5854 23154 5906
rect 23438 5854 23490 5906
rect 23662 5854 23714 5906
rect 23886 5854 23938 5906
rect 25902 5854 25954 5906
rect 24110 5742 24162 5794
rect 25566 5742 25618 5794
rect 4616 5462 4668 5514
rect 4720 5462 4772 5514
rect 4824 5462 4876 5514
rect 11420 5462 11472 5514
rect 11524 5462 11576 5514
rect 11628 5462 11680 5514
rect 18224 5462 18276 5514
rect 18328 5462 18380 5514
rect 18432 5462 18484 5514
rect 25028 5462 25080 5514
rect 25132 5462 25184 5514
rect 25236 5462 25288 5514
rect 22542 5182 22594 5234
rect 1710 5070 1762 5122
rect 2494 5070 2546 5122
rect 18734 5070 18786 5122
rect 20638 5070 20690 5122
rect 21534 5070 21586 5122
rect 22990 5070 23042 5122
rect 25454 5070 25506 5122
rect 26910 5070 26962 5122
rect 27358 5070 27410 5122
rect 27806 5070 27858 5122
rect 2046 4958 2098 5010
rect 19742 4958 19794 5010
rect 20414 4958 20466 5010
rect 23214 4958 23266 5010
rect 23886 4958 23938 5010
rect 19070 4846 19122 4898
rect 19854 4846 19906 4898
rect 20078 4846 20130 4898
rect 20526 4846 20578 4898
rect 21310 4846 21362 4898
rect 26014 4846 26066 4898
rect 26462 4846 26514 4898
rect 8018 4678 8070 4730
rect 8122 4678 8174 4730
rect 8226 4678 8278 4730
rect 14822 4678 14874 4730
rect 14926 4678 14978 4730
rect 15030 4678 15082 4730
rect 21626 4678 21678 4730
rect 21730 4678 21782 4730
rect 21834 4678 21886 4730
rect 28430 4678 28482 4730
rect 28534 4678 28586 4730
rect 28638 4678 28690 4730
rect 19630 4510 19682 4562
rect 22430 4510 22482 4562
rect 11790 4398 11842 4450
rect 18510 4398 18562 4450
rect 18846 4398 18898 4450
rect 19182 4398 19234 4450
rect 20638 4398 20690 4450
rect 22990 4398 23042 4450
rect 25230 4398 25282 4450
rect 11230 4286 11282 4338
rect 11566 4286 11618 4338
rect 19406 4286 19458 4338
rect 21534 4286 21586 4338
rect 23438 4286 23490 4338
rect 24222 4286 24274 4338
rect 25342 4286 25394 4338
rect 25790 4286 25842 4338
rect 10782 4174 10834 4226
rect 11678 4174 11730 4226
rect 12238 4174 12290 4226
rect 17838 4174 17890 4226
rect 18286 4174 18338 4226
rect 21870 4174 21922 4226
rect 23214 4174 23266 4226
rect 24110 4174 24162 4226
rect 24670 4174 24722 4226
rect 26462 4174 26514 4226
rect 26910 4174 26962 4226
rect 27358 4174 27410 4226
rect 27806 4174 27858 4226
rect 19742 4062 19794 4114
rect 24558 4062 24610 4114
rect 27022 4062 27074 4114
rect 27806 4062 27858 4114
rect 4616 3894 4668 3946
rect 4720 3894 4772 3946
rect 4824 3894 4876 3946
rect 11420 3894 11472 3946
rect 11524 3894 11576 3946
rect 11628 3894 11680 3946
rect 18224 3894 18276 3946
rect 18328 3894 18380 3946
rect 18432 3894 18484 3946
rect 25028 3894 25080 3946
rect 25132 3894 25184 3946
rect 25236 3894 25288 3946
rect 20078 3726 20130 3778
rect 22206 3726 22258 3778
rect 11006 3614 11058 3666
rect 13022 3614 13074 3666
rect 21422 3614 21474 3666
rect 21982 3614 22034 3666
rect 27918 3614 27970 3666
rect 7646 3502 7698 3554
rect 9662 3502 9714 3554
rect 11790 3502 11842 3554
rect 15150 3502 15202 3554
rect 17278 3502 17330 3554
rect 19294 3502 19346 3554
rect 20078 3502 20130 3554
rect 20302 3502 20354 3554
rect 22318 3502 22370 3554
rect 22654 3502 22706 3554
rect 23662 3502 23714 3554
rect 24110 3502 24162 3554
rect 24558 3502 24610 3554
rect 26126 3502 26178 3554
rect 5182 3390 5234 3442
rect 5630 3390 5682 3442
rect 5742 3390 5794 3442
rect 7758 3390 7810 3442
rect 10222 3390 10274 3442
rect 12126 3390 12178 3442
rect 12350 3390 12402 3442
rect 16270 3390 16322 3442
rect 17726 3390 17778 3442
rect 19630 3390 19682 3442
rect 23326 3390 23378 3442
rect 25678 3390 25730 3442
rect 27134 3390 27186 3442
rect 27470 3390 27522 3442
rect 4622 3278 4674 3330
rect 5966 3278 6018 3330
rect 6302 3278 6354 3330
rect 6862 3278 6914 3330
rect 7422 3278 7474 3330
rect 13582 3278 13634 3330
rect 18846 3278 18898 3330
rect 21310 3278 21362 3330
rect 8018 3110 8070 3162
rect 8122 3110 8174 3162
rect 8226 3110 8278 3162
rect 14822 3110 14874 3162
rect 14926 3110 14978 3162
rect 15030 3110 15082 3162
rect 21626 3110 21678 3162
rect 21730 3110 21782 3162
rect 21834 3110 21886 3162
rect 28430 3110 28482 3162
rect 28534 3110 28586 3162
rect 28638 3110 28690 3162
rect 6190 2942 6242 2994
rect 9102 2942 9154 2994
rect 12014 2942 12066 2994
rect 12574 2942 12626 2994
rect 17502 2942 17554 2994
rect 24334 2942 24386 2994
rect 25342 2942 25394 2994
rect 9998 2830 10050 2882
rect 17950 2830 18002 2882
rect 19518 2830 19570 2882
rect 20750 2830 20802 2882
rect 21646 2830 21698 2882
rect 25454 2830 25506 2882
rect 26126 2830 26178 2882
rect 26686 2830 26738 2882
rect 27358 2830 27410 2882
rect 2942 2718 2994 2770
rect 6190 2718 6242 2770
rect 6302 2718 6354 2770
rect 9662 2718 9714 2770
rect 10558 2718 10610 2770
rect 11678 2718 11730 2770
rect 12686 2718 12738 2770
rect 17390 2718 17442 2770
rect 18398 2718 18450 2770
rect 18958 2718 19010 2770
rect 21198 2718 21250 2770
rect 22990 2718 23042 2770
rect 24110 2718 24162 2770
rect 24334 2718 24386 2770
rect 25342 2718 25394 2770
rect 27022 2718 27074 2770
rect 27582 2718 27634 2770
rect 4062 2606 4114 2658
rect 5966 2606 6018 2658
rect 7758 2606 7810 2658
rect 8206 2606 8258 2658
rect 8654 2606 8706 2658
rect 11118 2606 11170 2658
rect 11454 2606 11506 2658
rect 13694 2606 13746 2658
rect 14142 2606 14194 2658
rect 14814 2606 14866 2658
rect 15486 2606 15538 2658
rect 16270 2606 16322 2658
rect 16718 2606 16770 2658
rect 18622 2606 18674 2658
rect 20862 2606 20914 2658
rect 23774 2606 23826 2658
rect 28142 2606 28194 2658
rect 10446 2494 10498 2546
rect 10782 2494 10834 2546
rect 11006 2494 11058 2546
rect 12574 2494 12626 2546
rect 12910 2494 12962 2546
rect 13134 2494 13186 2546
rect 4616 2326 4668 2378
rect 4720 2326 4772 2378
rect 4824 2326 4876 2378
rect 11420 2326 11472 2378
rect 11524 2326 11576 2378
rect 11628 2326 11680 2378
rect 18224 2326 18276 2378
rect 18328 2326 18380 2378
rect 18432 2326 18484 2378
rect 25028 2326 25080 2378
rect 25132 2326 25184 2378
rect 25236 2326 25288 2378
rect 18958 2046 19010 2098
rect 20750 2046 20802 2098
rect 20974 2046 21026 2098
rect 21870 2046 21922 2098
rect 22878 2046 22930 2098
rect 24670 2046 24722 2098
rect 25454 2046 25506 2098
rect 26462 2046 26514 2098
rect 1934 1934 1986 1986
rect 2718 1934 2770 1986
rect 4062 1934 4114 1986
rect 4734 1934 4786 1986
rect 6078 1934 6130 1986
rect 6526 1934 6578 1986
rect 7198 1934 7250 1986
rect 7870 1934 7922 1986
rect 8542 1934 8594 1986
rect 9662 1934 9714 1986
rect 10334 1934 10386 1986
rect 11230 1934 11282 1986
rect 11678 1934 11730 1986
rect 12350 1934 12402 1986
rect 13470 1934 13522 1986
rect 13918 1934 13970 1986
rect 14702 1934 14754 1986
rect 17614 1934 17666 1986
rect 18622 1934 18674 1986
rect 19854 1934 19906 1986
rect 20190 1934 20242 1986
rect 21086 1934 21138 1986
rect 22430 1934 22482 1986
rect 23214 1934 23266 1986
rect 23998 1934 24050 1986
rect 25006 1934 25058 1986
rect 25902 1934 25954 1986
rect 26910 1934 26962 1986
rect 27582 1934 27634 1986
rect 2942 1822 2994 1874
rect 3278 1822 3330 1874
rect 3614 1822 3666 1874
rect 4286 1822 4338 1874
rect 4958 1822 5010 1874
rect 5742 1822 5794 1874
rect 6750 1822 6802 1874
rect 7422 1822 7474 1874
rect 8094 1822 8146 1874
rect 8766 1822 8818 1874
rect 9886 1822 9938 1874
rect 10558 1822 10610 1874
rect 11902 1822 11954 1874
rect 12574 1822 12626 1874
rect 13694 1822 13746 1874
rect 14366 1822 14418 1874
rect 15038 1822 15090 1874
rect 15374 1822 15426 1874
rect 15710 1822 15762 1874
rect 16046 1822 16098 1874
rect 16942 1822 16994 1874
rect 17278 1822 17330 1874
rect 17950 1822 18002 1874
rect 18510 1822 18562 1874
rect 19294 1822 19346 1874
rect 19630 1822 19682 1874
rect 20078 1822 20130 1874
rect 23662 1822 23714 1874
rect 27358 1822 27410 1874
rect 2382 1710 2434 1762
rect 10894 1710 10946 1762
rect 8018 1542 8070 1594
rect 8122 1542 8174 1594
rect 8226 1542 8278 1594
rect 14822 1542 14874 1594
rect 14926 1542 14978 1594
rect 15030 1542 15082 1594
rect 21626 1542 21678 1594
rect 21730 1542 21782 1594
rect 21834 1542 21886 1594
rect 28430 1542 28482 1594
rect 28534 1542 28586 1594
rect 28638 1542 28690 1594
<< metal2 >>
rect 1344 119600 1456 120000
rect 3136 119600 3248 120000
rect 4928 119600 5040 120000
rect 6720 119600 6832 120000
rect 8512 119600 8624 120000
rect 10304 119600 10416 120000
rect 12096 119600 12208 120000
rect 13888 119600 14000 120000
rect 15680 119600 15792 120000
rect 17472 119600 17584 120000
rect 19264 119600 19376 120000
rect 21056 119600 21168 120000
rect 22848 119600 22960 120000
rect 23660 119644 24388 119700
rect 1372 118692 1428 119600
rect 1372 118636 1764 118692
rect 1708 117906 1764 118636
rect 1708 117854 1710 117906
rect 1762 117854 1764 117906
rect 1708 117842 1764 117854
rect 3164 117908 3220 119600
rect 4956 118804 5012 119600
rect 4956 118748 5572 118804
rect 4614 118412 4878 118422
rect 4670 118356 4718 118412
rect 4774 118356 4822 118412
rect 4614 118346 4878 118356
rect 3388 117908 3444 117918
rect 3164 117906 3444 117908
rect 3164 117854 3390 117906
rect 3442 117854 3444 117906
rect 3164 117852 3444 117854
rect 3388 117842 3444 117852
rect 5516 117906 5572 118748
rect 5516 117854 5518 117906
rect 5570 117854 5572 117906
rect 5516 117842 5572 117854
rect 6748 117908 6804 119600
rect 8540 118802 8596 119600
rect 8540 118750 8542 118802
rect 8594 118750 8596 118802
rect 8540 118738 8596 118750
rect 9324 118802 9380 118814
rect 9324 118750 9326 118802
rect 9378 118750 9380 118802
rect 6972 117908 7028 117918
rect 6748 117906 7028 117908
rect 6748 117854 6974 117906
rect 7026 117854 7028 117906
rect 6748 117852 7028 117854
rect 6972 117842 7028 117852
rect 9324 117906 9380 118750
rect 9324 117854 9326 117906
rect 9378 117854 9380 117906
rect 9324 117842 9380 117854
rect 10332 117908 10388 119600
rect 11418 118412 11682 118422
rect 11474 118356 11522 118412
rect 11578 118356 11626 118412
rect 11418 118346 11682 118356
rect 10556 117908 10612 117918
rect 10332 117906 10612 117908
rect 10332 117854 10558 117906
rect 10610 117854 10612 117906
rect 10332 117852 10612 117854
rect 12124 117908 12180 119600
rect 13916 118804 13972 119600
rect 13356 118748 13972 118804
rect 12348 117908 12404 117918
rect 12124 117906 12404 117908
rect 12124 117854 12350 117906
rect 12402 117854 12404 117906
rect 12124 117852 12404 117854
rect 10556 117842 10612 117852
rect 12348 117842 12404 117852
rect 13356 117906 13412 118748
rect 13356 117854 13358 117906
rect 13410 117854 13412 117906
rect 13356 117842 13412 117854
rect 13804 118018 13860 118030
rect 13804 117966 13806 118018
rect 13858 117966 13860 118018
rect 8016 117628 8280 117638
rect 8072 117572 8120 117628
rect 8176 117572 8224 117628
rect 8016 117562 8280 117572
rect 13804 117236 13860 117966
rect 14700 118018 14756 118030
rect 14700 117966 14702 118018
rect 14754 117966 14756 118018
rect 13804 117234 13972 117236
rect 13804 117182 13806 117234
rect 13858 117182 13972 117234
rect 13804 117180 13972 117182
rect 13804 117170 13860 117180
rect 4614 116844 4878 116854
rect 4670 116788 4718 116844
rect 4774 116788 4822 116844
rect 4614 116778 4878 116788
rect 11418 116844 11682 116854
rect 11474 116788 11522 116844
rect 11578 116788 11626 116844
rect 11418 116778 11682 116788
rect 10780 116450 10836 116462
rect 10780 116398 10782 116450
rect 10834 116398 10836 116450
rect 8016 116060 8280 116070
rect 8072 116004 8120 116060
rect 8176 116004 8224 116060
rect 8016 115994 8280 116004
rect 1708 115778 1764 115790
rect 1708 115726 1710 115778
rect 1762 115726 1764 115778
rect 1708 114996 1764 115726
rect 10780 115668 10836 116398
rect 11452 116450 11508 116462
rect 11452 116398 11454 116450
rect 11506 116398 11508 116450
rect 10780 115602 10836 115612
rect 11228 115668 11284 115678
rect 11452 115668 11508 116398
rect 13916 116450 13972 117180
rect 13916 116398 13918 116450
rect 13970 116398 13972 116450
rect 13020 116228 13076 116238
rect 13580 116228 13636 116238
rect 12684 116226 13748 116228
rect 12684 116174 13022 116226
rect 13074 116174 13582 116226
rect 13634 116174 13748 116226
rect 12684 116172 13748 116174
rect 12684 115890 12740 116172
rect 13020 116162 13076 116172
rect 13580 116162 13636 116172
rect 12684 115838 12686 115890
rect 12738 115838 12740 115890
rect 12684 115826 12740 115838
rect 11228 115666 11508 115668
rect 11228 115614 11230 115666
rect 11282 115614 11508 115666
rect 11228 115612 11508 115614
rect 12236 115668 12292 115678
rect 10108 115442 10164 115454
rect 10108 115390 10110 115442
rect 10162 115390 10164 115442
rect 4614 115276 4878 115286
rect 4670 115220 4718 115276
rect 4774 115220 4822 115276
rect 4614 115210 4878 115220
rect 1708 114930 1764 114940
rect 8016 114492 8280 114502
rect 8072 114436 8120 114492
rect 8176 114436 8224 114492
rect 8016 114426 8280 114436
rect 10108 114212 10164 115390
rect 11228 114268 11284 115612
rect 12236 115574 12292 115612
rect 13356 115668 13412 115678
rect 13468 115668 13524 115678
rect 13412 115666 13524 115668
rect 13412 115614 13470 115666
rect 13522 115614 13524 115666
rect 13412 115612 13524 115614
rect 11418 115276 11682 115286
rect 11474 115220 11522 115276
rect 11578 115220 11626 115276
rect 11418 115210 11682 115220
rect 13356 114268 13412 115612
rect 13468 115602 13524 115612
rect 10108 113874 10164 114156
rect 11116 114212 11284 114268
rect 13020 114212 13636 114268
rect 11116 114146 11172 114156
rect 10108 113822 10110 113874
rect 10162 113822 10164 113874
rect 4614 113708 4878 113718
rect 4670 113652 4718 113708
rect 4774 113652 4822 113708
rect 4614 113642 4878 113652
rect 7980 113314 8036 113326
rect 7980 113262 7982 113314
rect 8034 113262 8036 113314
rect 7980 113204 8036 113262
rect 7980 113138 8036 113148
rect 8876 113314 8932 113326
rect 8876 113262 8878 113314
rect 8930 113262 8932 113314
rect 8016 112924 8280 112934
rect 8072 112868 8120 112924
rect 8176 112868 8224 112924
rect 8016 112858 8280 112868
rect 8428 112644 8484 112654
rect 8428 112532 8484 112588
rect 8876 112644 8932 113262
rect 8876 112578 8932 112588
rect 9212 113204 9268 113214
rect 8316 112476 8484 112532
rect 3948 112308 4004 112318
rect 1708 109620 1764 109630
rect 1708 105586 1764 109564
rect 3948 106484 4004 112252
rect 4614 112140 4878 112150
rect 4670 112084 4718 112140
rect 4774 112084 4822 112140
rect 4614 112074 4878 112084
rect 8316 111746 8372 112476
rect 9212 111748 9268 113148
rect 10108 113092 10164 113822
rect 10556 114100 10612 114110
rect 10556 113314 10612 114044
rect 10556 113262 10558 113314
rect 10610 113262 10612 113314
rect 10556 113204 10612 113262
rect 10556 113138 10612 113148
rect 11228 114098 11284 114110
rect 11228 114046 11230 114098
rect 11282 114046 11284 114098
rect 11228 113314 11284 114046
rect 12124 114100 12180 114110
rect 12124 114006 12180 114044
rect 12684 114100 12740 114110
rect 11418 113708 11682 113718
rect 11474 113652 11522 113708
rect 11578 113652 11626 113708
rect 11418 113642 11682 113652
rect 11228 113262 11230 113314
rect 11282 113262 11284 113314
rect 10220 113092 10276 113102
rect 10108 113090 10276 113092
rect 10108 113038 10222 113090
rect 10274 113038 10276 113090
rect 10108 113036 10276 113038
rect 9548 111748 9604 111758
rect 8316 111694 8318 111746
rect 8370 111694 8372 111746
rect 8316 111682 8372 111694
rect 8876 111746 9604 111748
rect 8876 111694 9214 111746
rect 9266 111694 9550 111746
rect 9602 111694 9604 111746
rect 8876 111692 9604 111694
rect 6860 111522 6916 111534
rect 6860 111470 6862 111522
rect 6914 111470 6916 111522
rect 6860 110964 6916 111470
rect 8016 111356 8280 111366
rect 8072 111300 8120 111356
rect 8176 111300 8224 111356
rect 8016 111290 8280 111300
rect 6860 110898 6916 110908
rect 4614 110572 4878 110582
rect 4670 110516 4718 110572
rect 4774 110516 4822 110572
rect 4614 110506 4878 110516
rect 8876 110178 8932 111692
rect 9212 111682 9268 111692
rect 9548 110962 9604 111692
rect 9548 110910 9550 110962
rect 9602 110910 9604 110962
rect 9548 110898 9604 110910
rect 9548 110740 9604 110750
rect 8876 110126 8878 110178
rect 8930 110126 8932 110178
rect 8876 110114 8932 110126
rect 8988 110180 9044 110190
rect 8016 109788 8280 109798
rect 8072 109732 8120 109788
rect 8176 109732 8224 109788
rect 8016 109722 8280 109732
rect 4614 109004 4878 109014
rect 4670 108948 4718 109004
rect 4774 108948 4822 109004
rect 4614 108938 4878 108948
rect 8988 108722 9044 110124
rect 9548 109228 9604 110684
rect 10220 110740 10276 113036
rect 10220 110674 10276 110684
rect 10332 112644 10388 112654
rect 10332 111746 10388 112588
rect 11228 112644 11284 113262
rect 11228 112578 11284 112588
rect 12124 113092 12180 113102
rect 11452 112532 11508 112542
rect 11452 112438 11508 112476
rect 12124 112530 12180 113036
rect 12124 112478 12126 112530
rect 12178 112478 12180 112530
rect 11418 112140 11682 112150
rect 11474 112084 11522 112140
rect 11578 112084 11626 112140
rect 11418 112074 11682 112084
rect 10332 111694 10334 111746
rect 10386 111694 10388 111746
rect 10332 110962 10388 111694
rect 10332 110910 10334 110962
rect 10386 110910 10388 110962
rect 9660 110180 9716 110190
rect 9660 110086 9716 110124
rect 10332 110180 10388 110910
rect 11676 111972 11732 111982
rect 12124 111972 12180 112478
rect 11676 111970 12180 111972
rect 11676 111918 11678 111970
rect 11730 111918 12180 111970
rect 11676 111916 12180 111918
rect 11004 110740 11060 110750
rect 11004 110402 11060 110684
rect 11676 110740 11732 111916
rect 12348 111524 12404 111534
rect 12348 111522 12516 111524
rect 12348 111470 12350 111522
rect 12402 111470 12516 111522
rect 12348 111468 12516 111470
rect 12348 111458 12404 111468
rect 12124 110964 12180 110974
rect 12012 110962 12180 110964
rect 12012 110910 12126 110962
rect 12178 110910 12180 110962
rect 12012 110908 12180 110910
rect 11676 110674 11732 110684
rect 11788 110852 11844 110862
rect 11418 110572 11682 110582
rect 11474 110516 11522 110572
rect 11578 110516 11626 110572
rect 11418 110506 11682 110516
rect 11004 110350 11006 110402
rect 11058 110350 11060 110402
rect 11004 110338 11060 110350
rect 11452 110292 11508 110302
rect 11452 110198 11508 110236
rect 10332 110114 10388 110124
rect 10780 110180 10836 110190
rect 10780 109394 10836 110124
rect 11676 110180 11732 110190
rect 11676 110086 11732 110124
rect 10780 109342 10782 109394
rect 10834 109342 10836 109394
rect 10780 109330 10836 109342
rect 11676 109396 11732 109406
rect 11788 109396 11844 110796
rect 12012 110402 12068 110908
rect 12124 110898 12180 110908
rect 12012 110350 12014 110402
rect 12066 110350 12068 110402
rect 12012 110338 12068 110350
rect 12460 110292 12516 111468
rect 12684 111074 12740 114044
rect 12796 113092 12852 113102
rect 12796 112998 12852 113036
rect 12684 111022 12686 111074
rect 12738 111022 12740 111074
rect 12684 110852 12740 111022
rect 12684 110786 12740 110796
rect 13020 112532 13076 114212
rect 13580 114098 13636 114212
rect 13580 114046 13582 114098
rect 13634 114046 13636 114098
rect 13580 114034 13636 114046
rect 13356 113092 13412 113102
rect 13692 113092 13748 116172
rect 13916 115668 13972 116398
rect 14700 117234 14756 117966
rect 14820 117628 15084 117638
rect 14876 117572 14924 117628
rect 14980 117572 15028 117628
rect 14820 117562 15084 117572
rect 14700 117182 14702 117234
rect 14754 117182 14756 117234
rect 14700 116452 14756 117182
rect 15708 117012 15764 119600
rect 16044 117794 16100 117806
rect 16044 117742 16046 117794
rect 16098 117742 16100 117794
rect 16044 117124 16100 117742
rect 16380 117794 16436 117806
rect 16380 117742 16382 117794
rect 16434 117742 16436 117794
rect 16380 117124 16436 117742
rect 17388 117234 17444 117246
rect 17388 117182 17390 117234
rect 17442 117182 17444 117234
rect 16828 117124 16884 117134
rect 16044 117122 16884 117124
rect 16044 117070 16046 117122
rect 16098 117070 16382 117122
rect 16434 117070 16830 117122
rect 16882 117070 16884 117122
rect 16044 117068 16884 117070
rect 16044 117058 16100 117068
rect 15484 116956 15764 117012
rect 14924 116452 14980 116462
rect 15148 116452 15204 116462
rect 14700 116450 15148 116452
rect 14700 116398 14926 116450
rect 14978 116398 15148 116450
rect 14700 116396 15148 116398
rect 13916 115602 13972 115612
rect 14476 115668 14532 115678
rect 14700 115668 14756 116396
rect 14924 116386 14980 116396
rect 15148 116386 15204 116396
rect 14820 116060 15084 116070
rect 14876 116004 14924 116060
rect 14980 116004 15028 116060
rect 14820 115994 15084 116004
rect 14476 115666 14756 115668
rect 14476 115614 14478 115666
rect 14530 115614 14756 115666
rect 14476 115612 14756 115614
rect 14476 115602 14532 115612
rect 14820 114492 15084 114502
rect 14876 114436 14924 114492
rect 14980 114436 15028 114492
rect 14820 114426 15084 114436
rect 15484 114268 15540 116956
rect 16268 116564 16324 116574
rect 16380 116564 16436 117068
rect 16268 116562 16436 116564
rect 16268 116510 16270 116562
rect 16322 116510 16436 116562
rect 16268 116508 16436 116510
rect 16828 116564 16884 117068
rect 16268 116452 16324 116508
rect 16828 116498 16884 116508
rect 16156 115892 16212 115902
rect 16268 115892 16324 116396
rect 16716 116452 16772 116462
rect 16716 116358 16772 116396
rect 17388 116452 17444 117182
rect 17500 117012 17556 119600
rect 18222 118412 18486 118422
rect 18278 118356 18326 118412
rect 18382 118356 18430 118412
rect 18222 118346 18486 118356
rect 17836 117794 17892 117806
rect 17836 117742 17838 117794
rect 17890 117742 17892 117794
rect 17500 116956 17668 117012
rect 16156 115890 16324 115892
rect 16156 115838 16158 115890
rect 16210 115838 16324 115890
rect 16156 115836 16324 115838
rect 16156 115826 16212 115836
rect 17388 115668 17444 116396
rect 17500 115668 17556 115678
rect 17388 115666 17556 115668
rect 17388 115614 17502 115666
rect 17554 115614 17556 115666
rect 17388 115612 17556 115614
rect 15596 115442 15652 115454
rect 15596 115390 15598 115442
rect 15650 115390 15652 115442
rect 15596 114996 15652 115390
rect 15708 114996 15764 115006
rect 15596 114994 15764 114996
rect 15596 114942 15710 114994
rect 15762 114942 15764 114994
rect 15596 114940 15764 114942
rect 15260 114212 15540 114268
rect 14588 114100 14644 114110
rect 14588 114098 14756 114100
rect 14588 114046 14590 114098
rect 14642 114046 14756 114098
rect 14588 114044 14756 114046
rect 14588 114034 14644 114044
rect 13804 113092 13860 113102
rect 13412 113090 13860 113092
rect 13412 113038 13806 113090
rect 13858 113038 13860 113090
rect 13412 113036 13860 113038
rect 13356 113026 13412 113036
rect 12348 109954 12404 109966
rect 12348 109902 12350 109954
rect 12402 109902 12404 109954
rect 11676 109394 11844 109396
rect 11676 109342 11678 109394
rect 11730 109342 11844 109394
rect 11676 109340 11844 109342
rect 12124 109506 12180 109518
rect 12124 109454 12126 109506
rect 12178 109454 12180 109506
rect 11676 109330 11732 109340
rect 9548 109172 9716 109228
rect 8988 108670 8990 108722
rect 9042 108670 9044 108722
rect 8988 108658 9044 108670
rect 9660 109170 9716 109172
rect 9660 109118 9662 109170
rect 9714 109118 9716 109170
rect 9660 108834 9716 109118
rect 11418 109004 11682 109014
rect 11474 108948 11522 109004
rect 11578 108948 11626 109004
rect 11418 108938 11682 108948
rect 9660 108782 9662 108834
rect 9714 108782 9716 108834
rect 9212 108500 9268 108510
rect 9268 108444 9380 108500
rect 9212 108406 9268 108444
rect 8016 108220 8280 108230
rect 8072 108164 8120 108220
rect 8176 108164 8224 108220
rect 8016 108154 8280 108164
rect 7532 107716 7588 107726
rect 7420 107660 7532 107716
rect 4614 107436 4878 107446
rect 4670 107380 4718 107436
rect 4774 107380 4822 107436
rect 4614 107370 4878 107380
rect 3948 106418 4004 106428
rect 4284 106932 4340 106942
rect 3164 106370 3220 106382
rect 3164 106318 3166 106370
rect 3218 106318 3220 106370
rect 3164 106148 3220 106318
rect 3164 106082 3220 106092
rect 3276 106146 3332 106158
rect 3276 106094 3278 106146
rect 3330 106094 3332 106146
rect 3276 105700 3332 106094
rect 3836 106148 3892 106158
rect 3836 106054 3892 106092
rect 3388 106036 3444 106046
rect 3388 106034 3780 106036
rect 3388 105982 3390 106034
rect 3442 105982 3780 106034
rect 3388 105980 3780 105982
rect 3388 105970 3444 105980
rect 3724 105924 3780 105980
rect 3724 105868 4004 105924
rect 3276 105644 3892 105700
rect 1708 105534 1710 105586
rect 1762 105534 1764 105586
rect 1708 104916 1764 105534
rect 3836 105586 3892 105644
rect 3836 105534 3838 105586
rect 3890 105534 3892 105586
rect 3836 105522 3892 105534
rect 1708 104850 1764 104860
rect 3836 104916 3892 104926
rect 3836 104822 3892 104860
rect 3948 104914 4004 105868
rect 3948 104862 3950 104914
rect 4002 104862 4004 104914
rect 3948 104850 4004 104862
rect 4060 105700 4116 105710
rect 4060 104914 4116 105644
rect 4284 105252 4340 106876
rect 5628 106484 5684 106494
rect 4732 106146 4788 106158
rect 4732 106094 4734 106146
rect 4786 106094 4788 106146
rect 4732 106036 4788 106094
rect 4956 106148 5012 106158
rect 4844 106036 4900 106046
rect 4732 105980 4844 106036
rect 4844 105970 4900 105980
rect 4614 105868 4878 105878
rect 4670 105812 4718 105868
rect 4774 105812 4822 105868
rect 4614 105802 4878 105812
rect 4508 105476 4564 105486
rect 4284 105186 4340 105196
rect 4396 105420 4508 105476
rect 4060 104862 4062 104914
rect 4114 104862 4116 104914
rect 4060 104850 4116 104862
rect 4284 104804 4340 104814
rect 4284 104710 4340 104748
rect 3724 104692 3780 104702
rect 3388 104636 3724 104692
rect 2828 104580 2884 104590
rect 3276 104580 3332 104590
rect 2828 104578 2996 104580
rect 2828 104526 2830 104578
rect 2882 104526 2996 104578
rect 2828 104524 2996 104526
rect 2828 104514 2884 104524
rect 2940 104466 2996 104524
rect 3276 104486 3332 104524
rect 2940 104414 2942 104466
rect 2994 104414 2996 104466
rect 1708 104020 1764 104030
rect 1708 103348 1764 103964
rect 1708 103282 1764 103292
rect 2604 103124 2660 103134
rect 2604 103030 2660 103068
rect 2156 103010 2212 103022
rect 2156 102958 2158 103010
rect 2210 102958 2212 103010
rect 1708 101668 1764 101678
rect 1708 101442 1764 101612
rect 1708 101390 1710 101442
rect 1762 101390 1764 101442
rect 1708 101378 1764 101390
rect 2156 100546 2212 102958
rect 2940 103010 2996 104414
rect 3388 104466 3444 104636
rect 3724 104598 3780 104636
rect 3388 104414 3390 104466
rect 3442 104414 3444 104466
rect 3388 104402 3444 104414
rect 4396 104580 4452 105420
rect 4508 105382 4564 105420
rect 4396 103908 4452 104524
rect 4732 104580 4788 104590
rect 4956 104580 5012 106092
rect 5292 106146 5348 106158
rect 5292 106094 5294 106146
rect 5346 106094 5348 106146
rect 5292 105476 5348 106094
rect 5628 105588 5684 106428
rect 6076 106258 6132 106270
rect 6076 106206 6078 106258
rect 6130 106206 6132 106258
rect 5740 106148 5796 106158
rect 6076 106148 6132 106206
rect 5796 106092 6132 106148
rect 6300 106146 6356 106158
rect 6300 106094 6302 106146
rect 6354 106094 6356 106146
rect 5740 106054 5796 106092
rect 6300 105588 6356 106094
rect 7308 106146 7364 106158
rect 7308 106094 7310 106146
rect 7362 106094 7364 106146
rect 6412 106036 6468 106046
rect 6412 106034 6692 106036
rect 6412 105982 6414 106034
rect 6466 105982 6692 106034
rect 6412 105980 6692 105982
rect 6412 105970 6468 105980
rect 5628 105586 6244 105588
rect 5628 105534 5630 105586
rect 5682 105534 6244 105586
rect 5628 105532 6244 105534
rect 5628 105522 5684 105532
rect 5292 105410 5348 105420
rect 5180 105250 5236 105262
rect 5180 105198 5182 105250
rect 5234 105198 5236 105250
rect 5180 104692 5236 105198
rect 5180 104598 5236 104636
rect 5852 105252 5908 105262
rect 4732 104578 5012 104580
rect 4732 104526 4734 104578
rect 4786 104526 5012 104578
rect 4732 104524 5012 104526
rect 4732 104514 4788 104524
rect 4614 104300 4878 104310
rect 4670 104244 4718 104300
rect 4774 104244 4822 104300
rect 4614 104234 4878 104244
rect 4844 104020 4900 104030
rect 4508 103908 4564 103918
rect 4396 103906 4564 103908
rect 4396 103854 4510 103906
rect 4562 103854 4564 103906
rect 4396 103852 4564 103854
rect 3836 103794 3892 103806
rect 3836 103742 3838 103794
rect 3890 103742 3892 103794
rect 2940 102958 2942 103010
rect 2994 102958 2996 103010
rect 2940 102508 2996 102958
rect 2716 102452 2996 102508
rect 3276 103684 3332 103694
rect 3276 103122 3332 103628
rect 3500 103236 3556 103246
rect 3500 103142 3556 103180
rect 3724 103236 3780 103246
rect 3836 103236 3892 103742
rect 4284 103348 4340 103358
rect 4284 103254 4340 103292
rect 3724 103234 3892 103236
rect 3724 103182 3726 103234
rect 3778 103182 3892 103234
rect 3724 103180 3892 103182
rect 4060 103236 4116 103246
rect 3724 103170 3780 103180
rect 4060 103142 4116 103180
rect 3276 103070 3278 103122
rect 3330 103070 3332 103122
rect 2716 102228 2772 102452
rect 2604 102116 2660 102126
rect 2716 102116 2772 102172
rect 2604 102114 2772 102116
rect 2604 102062 2606 102114
rect 2658 102062 2772 102114
rect 2604 102060 2772 102062
rect 2604 102050 2660 102060
rect 2604 100660 2660 100670
rect 2604 100566 2660 100604
rect 2156 100494 2158 100546
rect 2210 100494 2212 100546
rect 2156 99874 2212 100494
rect 2156 99822 2158 99874
rect 2210 99822 2212 99874
rect 2156 99762 2212 99822
rect 2156 99710 2158 99762
rect 2210 99710 2212 99762
rect 2156 99698 2212 99710
rect 2604 99874 2660 99886
rect 2604 99822 2606 99874
rect 2658 99822 2660 99874
rect 1708 99314 1764 99326
rect 1708 99262 1710 99314
rect 1762 99262 1764 99314
rect 1708 98868 1764 99262
rect 1708 98802 1764 98812
rect 2380 98420 2436 98430
rect 2380 98306 2436 98364
rect 2380 98254 2382 98306
rect 2434 98254 2436 98306
rect 2380 98196 2436 98254
rect 2156 98140 2436 98196
rect 1932 96852 1988 96862
rect 2156 96852 2212 98140
rect 2604 97748 2660 99822
rect 2716 98420 2772 102060
rect 3052 102114 3108 102126
rect 3052 102062 3054 102114
rect 3106 102062 3108 102114
rect 3052 101556 3108 102062
rect 3052 101490 3108 101500
rect 3276 100772 3332 103070
rect 3948 103124 4004 103134
rect 4396 103124 4452 103134
rect 3948 103030 4004 103068
rect 4284 103122 4452 103124
rect 4284 103070 4398 103122
rect 4450 103070 4452 103122
rect 4284 103068 4452 103070
rect 3612 103012 3668 103022
rect 3388 102340 3444 102350
rect 3388 102246 3444 102284
rect 3500 102114 3556 102126
rect 3500 102062 3502 102114
rect 3554 102062 3556 102114
rect 3500 101668 3556 102062
rect 3500 101602 3556 101612
rect 3612 101444 3668 102956
rect 4172 102562 4228 102574
rect 4172 102510 4174 102562
rect 4226 102510 4228 102562
rect 2940 100770 3332 100772
rect 2940 100718 3278 100770
rect 3330 100718 3332 100770
rect 2940 100716 3332 100718
rect 2940 99986 2996 100716
rect 3276 100706 3332 100716
rect 3388 101388 3668 101444
rect 3724 102114 3780 102126
rect 3724 102062 3726 102114
rect 3778 102062 3780 102114
rect 3052 100546 3108 100558
rect 3052 100494 3054 100546
rect 3106 100494 3108 100546
rect 3052 100324 3108 100494
rect 3052 100268 3332 100324
rect 3164 99988 3220 99998
rect 2940 99934 2942 99986
rect 2994 99934 2996 99986
rect 2828 99876 2884 99886
rect 2940 99876 2996 99934
rect 2828 99874 2996 99876
rect 2828 99822 2830 99874
rect 2882 99822 2996 99874
rect 2828 99820 2996 99822
rect 2828 99810 2884 99820
rect 2828 98756 2884 98766
rect 2828 98642 2884 98700
rect 2828 98590 2830 98642
rect 2882 98590 2884 98642
rect 2828 98578 2884 98590
rect 2716 98354 2772 98364
rect 2604 97682 2660 97692
rect 2828 97410 2884 97422
rect 2828 97358 2830 97410
rect 2882 97358 2884 97410
rect 2828 97076 2884 97358
rect 2940 97076 2996 99820
rect 3052 99986 3220 99988
rect 3052 99934 3166 99986
rect 3218 99934 3220 99986
rect 3052 99932 3220 99934
rect 3052 98642 3108 99932
rect 3164 99922 3220 99932
rect 3276 99764 3332 100268
rect 3388 100100 3444 101388
rect 3724 101332 3780 102062
rect 3500 101276 3780 101332
rect 3836 101442 3892 101454
rect 3836 101390 3838 101442
rect 3890 101390 3892 101442
rect 3500 100770 3556 101276
rect 3724 100884 3780 100894
rect 3836 100884 3892 101390
rect 3724 100882 3892 100884
rect 3724 100830 3726 100882
rect 3778 100830 3892 100882
rect 3724 100828 3892 100830
rect 3724 100818 3780 100828
rect 3500 100718 3502 100770
rect 3554 100718 3556 100770
rect 3500 100706 3556 100718
rect 3948 100770 4004 100782
rect 3948 100718 3950 100770
rect 4002 100718 4004 100770
rect 3948 100548 4004 100718
rect 3948 100482 4004 100492
rect 4172 100212 4228 102510
rect 4284 102340 4340 103068
rect 4396 103058 4452 103068
rect 4508 102900 4564 103852
rect 4844 103124 4900 103964
rect 4956 103684 5012 104524
rect 5628 104578 5684 104590
rect 5628 104526 5630 104578
rect 5682 104526 5684 104578
rect 4956 103348 5012 103628
rect 4956 103282 5012 103292
rect 5068 104132 5124 104142
rect 5068 103682 5124 104076
rect 5068 103630 5070 103682
rect 5122 103630 5124 103682
rect 4844 103058 4900 103068
rect 4396 102844 4564 102900
rect 5068 102898 5124 103630
rect 5292 103908 5348 103918
rect 5292 103346 5348 103852
rect 5292 103294 5294 103346
rect 5346 103294 5348 103346
rect 5292 103282 5348 103294
rect 5628 103012 5684 104526
rect 5852 104468 5908 105196
rect 5852 104018 5908 104412
rect 5852 103966 5854 104018
rect 5906 103966 5908 104018
rect 5852 103954 5908 103966
rect 6076 104578 6132 104590
rect 6076 104526 6078 104578
rect 6130 104526 6132 104578
rect 6076 103236 6132 104526
rect 6188 104468 6244 105532
rect 6300 105522 6356 105532
rect 6636 104916 6692 105980
rect 7308 106034 7364 106094
rect 7308 105982 7310 106034
rect 7362 105982 7364 106034
rect 7308 105970 7364 105982
rect 6748 104916 6804 104926
rect 6636 104914 6804 104916
rect 6636 104862 6750 104914
rect 6802 104862 6804 104914
rect 6636 104860 6804 104862
rect 6748 104850 6804 104860
rect 6860 104916 6916 104926
rect 6524 104692 6580 104702
rect 6524 104598 6580 104636
rect 6636 104690 6692 104702
rect 6636 104638 6638 104690
rect 6690 104638 6692 104690
rect 6636 104468 6692 104638
rect 6188 104412 6692 104468
rect 6860 104690 6916 104860
rect 7308 104804 7364 104814
rect 7196 104802 7364 104804
rect 7196 104750 7310 104802
rect 7362 104750 7364 104802
rect 7196 104748 7364 104750
rect 6860 104638 6862 104690
rect 6914 104638 6916 104690
rect 6860 104356 6916 104638
rect 7084 104690 7140 104702
rect 7084 104638 7086 104690
rect 7138 104638 7140 104690
rect 7084 104580 7140 104638
rect 7084 104514 7140 104524
rect 6524 104300 6916 104356
rect 6412 103236 6468 103246
rect 5964 103180 6412 103236
rect 5628 103010 5796 103012
rect 5628 102958 5630 103010
rect 5682 102958 5796 103010
rect 5628 102956 5796 102958
rect 5628 102946 5684 102956
rect 5068 102846 5070 102898
rect 5122 102846 5124 102898
rect 4396 102564 4452 102844
rect 4614 102732 4878 102742
rect 4670 102676 4718 102732
rect 4774 102676 4822 102732
rect 4614 102666 4878 102676
rect 4396 102508 4676 102564
rect 4284 102274 4340 102284
rect 4284 102116 4340 102126
rect 4284 102022 4340 102060
rect 4396 101556 4452 101566
rect 4508 101556 4564 101566
rect 4620 101556 4676 102508
rect 5068 102562 5124 102846
rect 5068 102510 5070 102562
rect 5122 102510 5124 102562
rect 5068 102498 5124 102510
rect 4452 101554 4676 101556
rect 4452 101502 4510 101554
rect 4562 101502 4676 101554
rect 4452 101500 4676 101502
rect 4732 102116 4788 102126
rect 4396 100548 4452 101500
rect 4508 101490 4564 101500
rect 4732 101332 4788 102060
rect 5068 102114 5124 102126
rect 5068 102062 5070 102114
rect 5122 102062 5124 102114
rect 5068 101556 5124 102062
rect 5740 101556 5796 102956
rect 5964 102450 6020 103180
rect 6412 103170 6468 103180
rect 6076 103010 6132 103022
rect 6076 102958 6078 103010
rect 6130 102958 6132 103010
rect 6076 102898 6132 102958
rect 6076 102846 6078 102898
rect 6130 102846 6132 102898
rect 6076 102834 6132 102846
rect 6524 103010 6580 104300
rect 7084 103796 7140 103806
rect 6972 103348 7028 103358
rect 6972 103254 7028 103292
rect 7084 103346 7140 103740
rect 7084 103294 7086 103346
rect 7138 103294 7140 103346
rect 7084 103282 7140 103294
rect 7196 103234 7252 104748
rect 7308 104738 7364 104748
rect 7196 103182 7198 103234
rect 7250 103182 7252 103234
rect 7196 103170 7252 103182
rect 6524 102958 6526 103010
rect 6578 102958 6580 103010
rect 6524 102564 6580 102958
rect 6860 102900 6916 102910
rect 6524 102498 6580 102508
rect 6748 102844 6860 102900
rect 7420 102900 7476 107660
rect 7532 107650 7588 107660
rect 8988 107714 9044 107726
rect 8988 107662 8990 107714
rect 9042 107662 9044 107714
rect 8540 107266 8596 107278
rect 8540 107214 8542 107266
rect 8594 107214 8596 107266
rect 7532 106820 7588 106830
rect 8092 106820 8148 106830
rect 7532 106818 8148 106820
rect 7532 106766 7534 106818
rect 7586 106766 8094 106818
rect 8146 106766 8148 106818
rect 7532 106764 8148 106766
rect 7532 105812 7588 106764
rect 8092 106754 8148 106764
rect 8540 106818 8596 107214
rect 8988 107266 9044 107662
rect 8988 107214 8990 107266
rect 9042 107214 9044 107266
rect 8988 107202 9044 107214
rect 8540 106766 8542 106818
rect 8594 106766 8596 106818
rect 8016 106652 8280 106662
rect 8072 106596 8120 106652
rect 8176 106596 8224 106652
rect 8016 106586 8280 106596
rect 8540 106372 8596 106766
rect 9100 106820 9156 106830
rect 9100 106818 9268 106820
rect 9100 106766 9102 106818
rect 9154 106766 9268 106818
rect 9100 106764 9268 106766
rect 9100 106754 9156 106764
rect 9100 106372 9156 106382
rect 8540 106316 8820 106372
rect 8092 106260 8148 106270
rect 8092 106166 8148 106204
rect 7644 106148 7700 106158
rect 7644 106054 7700 106092
rect 8540 106148 8596 106158
rect 8316 106034 8372 106046
rect 8316 105982 8318 106034
rect 8370 105982 8372 106034
rect 8316 105924 8372 105982
rect 8540 106034 8596 106092
rect 8540 105982 8542 106034
rect 8594 105982 8596 106034
rect 8540 105970 8596 105982
rect 8316 105868 8484 105924
rect 8428 105812 8596 105868
rect 7532 105140 7588 105756
rect 7756 105588 7812 105598
rect 7756 105494 7812 105532
rect 8540 105474 8596 105812
rect 8540 105422 8542 105474
rect 8594 105422 8596 105474
rect 7532 105074 7588 105084
rect 8016 105084 8280 105094
rect 8072 105028 8120 105084
rect 8176 105028 8224 105084
rect 8016 105018 8280 105028
rect 7980 104916 8036 104926
rect 7532 104914 8036 104916
rect 7532 104862 7982 104914
rect 8034 104862 8036 104914
rect 7532 104860 8036 104862
rect 7532 104802 7588 104860
rect 7980 104850 8036 104860
rect 8092 104916 8148 104926
rect 8092 104822 8148 104860
rect 8316 104916 8372 104926
rect 7532 104750 7534 104802
rect 7586 104750 7588 104802
rect 7532 104738 7588 104750
rect 8316 104802 8372 104860
rect 8316 104750 8318 104802
rect 8370 104750 8372 104802
rect 8316 104738 8372 104750
rect 7644 104692 7700 104702
rect 7868 104692 7924 104702
rect 7644 104598 7700 104636
rect 7756 104690 7924 104692
rect 7756 104638 7870 104690
rect 7922 104638 7924 104690
rect 7756 104636 7924 104638
rect 7532 104468 7588 104478
rect 7756 104468 7812 104636
rect 7868 104626 7924 104636
rect 7588 104412 7812 104468
rect 7868 104468 7924 104478
rect 7532 104402 7588 104412
rect 7644 103684 7700 103694
rect 7644 103122 7700 103628
rect 7868 103346 7924 104412
rect 8540 104356 8596 105422
rect 8540 104290 8596 104300
rect 8652 104690 8708 104702
rect 8652 104638 8654 104690
rect 8706 104638 8708 104690
rect 8316 104244 8372 104254
rect 7980 103796 8036 103806
rect 7980 103702 8036 103740
rect 8316 103684 8372 104188
rect 8652 104244 8708 104638
rect 8652 104178 8708 104188
rect 8764 104132 8820 106316
rect 9100 106278 9156 106316
rect 9100 106036 9156 106046
rect 9212 106036 9268 106764
rect 9100 106034 9268 106036
rect 9100 105982 9102 106034
rect 9154 105982 9268 106034
rect 9100 105980 9268 105982
rect 9100 105970 9156 105980
rect 8876 105364 8932 105374
rect 8876 105270 8932 105308
rect 8988 105252 9044 105262
rect 8988 105250 9156 105252
rect 8988 105198 8990 105250
rect 9042 105198 9156 105250
rect 8988 105196 9156 105198
rect 8988 105186 9044 105196
rect 8988 104802 9044 104814
rect 8988 104750 8990 104802
rect 9042 104750 9044 104802
rect 8988 104692 9044 104750
rect 8988 104626 9044 104636
rect 8988 104132 9044 104142
rect 8764 104076 8988 104132
rect 8652 103908 8708 103918
rect 8540 103906 8708 103908
rect 8540 103854 8654 103906
rect 8706 103854 8708 103906
rect 8540 103852 8708 103854
rect 8540 103796 8596 103852
rect 8652 103842 8708 103852
rect 8876 103908 8932 103918
rect 8316 103628 8484 103684
rect 8016 103516 8280 103526
rect 8072 103460 8120 103516
rect 8176 103460 8224 103516
rect 8016 103450 8280 103460
rect 7868 103294 7870 103346
rect 7922 103294 7924 103346
rect 7868 103282 7924 103294
rect 8204 103348 8260 103358
rect 7756 103236 7812 103246
rect 7756 103142 7812 103180
rect 7644 103070 7646 103122
rect 7698 103070 7700 103122
rect 7644 103058 7700 103070
rect 8092 103122 8148 103134
rect 8092 103070 8094 103122
rect 8146 103070 8148 103122
rect 8092 102900 8148 103070
rect 7420 102844 8148 102900
rect 5964 102398 5966 102450
rect 6018 102398 6020 102450
rect 5964 102386 6020 102398
rect 6524 102114 6580 102126
rect 6524 102062 6526 102114
rect 6578 102062 6580 102114
rect 5852 101556 5908 101566
rect 6524 101556 6580 102062
rect 5740 101500 5852 101556
rect 5068 101490 5124 101500
rect 5180 101444 5236 101454
rect 5236 101388 5460 101444
rect 5180 101350 5236 101388
rect 4732 101276 5012 101332
rect 4614 101164 4878 101174
rect 4670 101108 4718 101164
rect 4774 101108 4822 101164
rect 4614 101098 4878 101108
rect 4956 100996 5012 101276
rect 4844 100940 5012 100996
rect 4844 100660 4900 100940
rect 4844 100566 4900 100604
rect 4508 100548 4564 100558
rect 4396 100546 4564 100548
rect 4396 100494 4510 100546
rect 4562 100494 4564 100546
rect 4396 100492 4564 100494
rect 4284 100212 4340 100222
rect 4172 100156 4284 100212
rect 4284 100118 4340 100156
rect 3500 100100 3556 100110
rect 3388 100098 3556 100100
rect 3388 100046 3502 100098
rect 3554 100046 3556 100098
rect 3388 100044 3556 100046
rect 3500 100034 3556 100044
rect 4508 99988 4564 100492
rect 4956 100546 5012 100558
rect 4956 100494 4958 100546
rect 5010 100494 5012 100546
rect 4956 100436 5012 100494
rect 4956 100370 5012 100380
rect 5180 100546 5236 100558
rect 5180 100494 5182 100546
rect 5234 100494 5236 100546
rect 5180 100100 5236 100494
rect 5292 100100 5348 100110
rect 5180 100098 5348 100100
rect 5180 100046 5294 100098
rect 5346 100046 5348 100098
rect 5180 100044 5348 100046
rect 5292 100034 5348 100044
rect 4620 99988 4676 99998
rect 4508 99986 5012 99988
rect 4508 99934 4622 99986
rect 4674 99934 5012 99986
rect 4508 99932 5012 99934
rect 4620 99922 4676 99932
rect 3164 99708 3332 99764
rect 3388 99874 3444 99886
rect 3388 99822 3390 99874
rect 3442 99822 3444 99874
rect 3164 98756 3220 99708
rect 3388 99540 3444 99822
rect 4614 99596 4878 99606
rect 4670 99540 4718 99596
rect 4774 99540 4822 99596
rect 3388 99484 3892 99540
rect 4614 99530 4878 99540
rect 3836 99314 3892 99484
rect 3836 99262 3838 99314
rect 3890 99262 3892 99314
rect 3836 99250 3892 99262
rect 4620 99202 4676 99214
rect 4620 99150 4622 99202
rect 4674 99150 4676 99202
rect 3164 98690 3220 98700
rect 3276 98868 3332 98878
rect 3052 98590 3054 98642
rect 3106 98590 3108 98642
rect 3052 98578 3108 98590
rect 3276 98642 3332 98812
rect 3276 98590 3278 98642
rect 3330 98590 3332 98642
rect 3276 98578 3332 98590
rect 4396 98644 4452 98654
rect 4396 98550 4452 98588
rect 4060 98532 4116 98542
rect 4060 98438 4116 98476
rect 3388 98420 3444 98430
rect 3388 98326 3444 98364
rect 4620 98308 4676 99150
rect 4956 99092 5012 99932
rect 5404 99876 5460 101388
rect 5628 101442 5684 101454
rect 5628 101390 5630 101442
rect 5682 101390 5684 101442
rect 5628 100772 5684 101390
rect 5628 100706 5684 100716
rect 5740 100770 5796 100782
rect 5740 100718 5742 100770
rect 5794 100718 5796 100770
rect 5292 99820 5460 99876
rect 5740 100660 5796 100718
rect 5180 99428 5236 99438
rect 5180 99314 5236 99372
rect 5180 99262 5182 99314
rect 5234 99262 5236 99314
rect 5180 99250 5236 99262
rect 4956 99036 5124 99092
rect 4844 98308 4900 98318
rect 4956 98308 5012 98318
rect 4620 98306 4956 98308
rect 4620 98254 4846 98306
rect 4898 98254 4956 98306
rect 4620 98252 4956 98254
rect 4844 98242 4900 98252
rect 4614 98028 4878 98038
rect 4670 97972 4718 98028
rect 4774 97972 4822 98028
rect 4614 97962 4878 97972
rect 4620 97860 4676 97870
rect 3276 97748 3332 97758
rect 3276 97654 3332 97692
rect 4620 97746 4676 97804
rect 4620 97694 4622 97746
rect 4674 97694 4676 97746
rect 3836 97636 3892 97646
rect 3836 97542 3892 97580
rect 4620 97468 4676 97694
rect 4172 97410 4228 97422
rect 4172 97358 4174 97410
rect 4226 97358 4228 97410
rect 2716 97020 3108 97076
rect 1932 96850 2212 96852
rect 1932 96798 1934 96850
rect 1986 96798 2158 96850
rect 2210 96798 2212 96850
rect 1932 96796 2212 96798
rect 1932 96786 1988 96796
rect 1708 96180 1764 96190
rect 1708 96086 1764 96124
rect 2156 94276 2212 96796
rect 2268 96962 2324 96974
rect 2268 96910 2270 96962
rect 2322 96910 2324 96962
rect 2268 96180 2324 96910
rect 2716 96962 2772 97020
rect 2716 96910 2718 96962
rect 2770 96910 2772 96962
rect 2716 96898 2772 96910
rect 2492 96850 2548 96862
rect 2492 96798 2494 96850
rect 2546 96798 2548 96850
rect 2492 96740 2548 96798
rect 2940 96850 2996 96862
rect 2940 96798 2942 96850
rect 2994 96798 2996 96850
rect 2940 96740 2996 96798
rect 2492 96684 2996 96740
rect 3052 96628 3108 97020
rect 3276 96850 3332 96862
rect 3276 96798 3278 96850
rect 3330 96798 3332 96850
rect 3164 96740 3220 96750
rect 3164 96646 3220 96684
rect 2268 96114 2324 96124
rect 2940 96572 3108 96628
rect 2380 95508 2436 95518
rect 2380 95414 2436 95452
rect 2828 95396 2884 95406
rect 2828 95302 2884 95340
rect 2492 94276 2548 94286
rect 2156 94274 2548 94276
rect 2156 94222 2494 94274
rect 2546 94222 2548 94274
rect 2156 94220 2548 94222
rect 2492 94052 2548 94220
rect 2492 93986 2548 93996
rect 2492 93828 2548 93838
rect 2940 93828 2996 96572
rect 3276 95732 3332 96798
rect 3836 96740 3892 96750
rect 3276 95666 3332 95676
rect 3388 96628 3444 96638
rect 3276 95508 3332 95518
rect 3388 95508 3444 96572
rect 3836 96178 3892 96684
rect 4172 96740 4228 97358
rect 4172 96646 4228 96684
rect 4396 97412 4676 97468
rect 4956 97748 5012 98252
rect 3836 96126 3838 96178
rect 3890 96126 3892 96178
rect 3836 96114 3892 96126
rect 3276 95506 3444 95508
rect 3276 95454 3278 95506
rect 3330 95454 3444 95506
rect 3276 95452 3444 95454
rect 3276 95442 3332 95452
rect 3724 95172 3780 95182
rect 3724 95078 3780 95116
rect 4060 95170 4116 95182
rect 4060 95118 4062 95170
rect 4114 95118 4116 95170
rect 3948 95060 4004 95070
rect 3052 94612 3108 94622
rect 3388 94612 3444 94622
rect 3052 94518 3108 94556
rect 3164 94610 3444 94612
rect 3164 94558 3390 94610
rect 3442 94558 3444 94610
rect 3164 94556 3444 94558
rect 2492 93826 2996 93828
rect 2492 93774 2494 93826
rect 2546 93774 2942 93826
rect 2994 93774 2996 93826
rect 2492 93772 2996 93774
rect 2492 93762 2548 93772
rect 1708 93492 1764 93502
rect 1708 93042 1764 93436
rect 1708 92990 1710 93042
rect 1762 92990 1764 93042
rect 1708 92978 1764 92990
rect 2940 92372 2996 93772
rect 3164 93826 3220 94556
rect 3388 94546 3444 94556
rect 3724 94612 3780 94622
rect 3724 94498 3780 94556
rect 3724 94446 3726 94498
rect 3778 94446 3780 94498
rect 3724 94434 3780 94446
rect 3948 94498 4004 95004
rect 3948 94446 3950 94498
rect 4002 94446 4004 94498
rect 3948 94434 4004 94446
rect 3388 94276 3444 94286
rect 3276 94274 3444 94276
rect 3276 94222 3390 94274
rect 3442 94222 3444 94274
rect 3276 94220 3444 94222
rect 3276 94052 3332 94220
rect 3388 94210 3444 94220
rect 3500 94274 3556 94286
rect 3500 94222 3502 94274
rect 3554 94222 3556 94274
rect 3276 93986 3332 93996
rect 3164 93774 3166 93826
rect 3218 93774 3220 93826
rect 3164 93762 3220 93774
rect 3052 93604 3108 93614
rect 3052 93510 3108 93548
rect 3500 93492 3556 94222
rect 4060 94276 4116 95118
rect 4396 95058 4452 97412
rect 4614 96460 4878 96470
rect 4670 96404 4718 96460
rect 4774 96404 4822 96460
rect 4614 96394 4878 96404
rect 4620 96068 4676 96078
rect 4956 96068 5012 97692
rect 5068 97524 5124 99036
rect 5180 98420 5236 98430
rect 5180 98326 5236 98364
rect 5068 97458 5124 97468
rect 4620 96066 5012 96068
rect 4620 96014 4622 96066
rect 4674 96014 5012 96066
rect 4620 96012 5012 96014
rect 4620 96002 4676 96012
rect 4956 95620 5012 96012
rect 5068 95844 5124 95854
rect 5068 95842 5236 95844
rect 5068 95790 5070 95842
rect 5122 95790 5236 95842
rect 5068 95788 5236 95790
rect 5068 95778 5124 95788
rect 4956 95564 5124 95620
rect 4508 95172 4564 95182
rect 4508 95078 4564 95116
rect 4956 95170 5012 95182
rect 4956 95118 4958 95170
rect 5010 95118 5012 95170
rect 4396 95006 4398 95058
rect 4450 95006 4452 95058
rect 4396 94994 4452 95006
rect 4956 95058 5012 95118
rect 4956 95006 4958 95058
rect 5010 95006 5012 95058
rect 4956 94994 5012 95006
rect 4614 94892 4878 94902
rect 4670 94836 4718 94892
rect 4774 94836 4822 94892
rect 4614 94826 4878 94836
rect 4844 94724 4900 94734
rect 4620 94668 4844 94724
rect 4620 94610 4676 94668
rect 4620 94558 4622 94610
rect 4674 94558 4676 94610
rect 4620 94546 4676 94558
rect 4060 93938 4116 94220
rect 4060 93886 4062 93938
rect 4114 93886 4116 93938
rect 4060 93874 4116 93886
rect 4844 93716 4900 94668
rect 5068 94610 5124 95564
rect 5180 95172 5236 95788
rect 5180 94836 5236 95116
rect 5180 94770 5236 94780
rect 5068 94558 5070 94610
rect 5122 94558 5124 94610
rect 5068 94546 5124 94558
rect 4844 93714 5012 93716
rect 4844 93662 4846 93714
rect 4898 93662 5012 93714
rect 4844 93660 5012 93662
rect 4844 93650 4900 93660
rect 3500 93426 3556 93436
rect 3836 93604 3892 93614
rect 3836 93042 3892 93548
rect 4508 93604 4564 93614
rect 4508 93510 4564 93548
rect 4614 93324 4878 93334
rect 4670 93268 4718 93324
rect 4774 93268 4822 93324
rect 4614 93258 4878 93268
rect 3836 92990 3838 93042
rect 3890 92990 3892 93042
rect 3836 92978 3892 92990
rect 4620 92932 4676 92942
rect 4956 92932 5012 93660
rect 5292 93604 5348 99820
rect 5740 99204 5796 100604
rect 5852 99988 5908 101500
rect 6076 101500 6580 101556
rect 5964 100660 6020 100670
rect 6076 100660 6132 101500
rect 6636 101444 6692 101454
rect 6300 101442 6692 101444
rect 6300 101390 6638 101442
rect 6690 101390 6692 101442
rect 6300 101388 6692 101390
rect 6300 100882 6356 101388
rect 6636 101378 6692 101388
rect 6300 100830 6302 100882
rect 6354 100830 6356 100882
rect 6300 100818 6356 100830
rect 6524 100772 6580 100782
rect 6020 100604 6132 100660
rect 6412 100660 6468 100670
rect 5964 100594 6020 100604
rect 6412 100566 6468 100604
rect 6188 100546 6244 100558
rect 6188 100494 6190 100546
rect 6242 100494 6244 100546
rect 6188 100324 6244 100494
rect 6244 100268 6356 100324
rect 6188 100258 6244 100268
rect 5852 99932 6020 99988
rect 5740 99138 5796 99148
rect 5852 99202 5908 99214
rect 5852 99150 5854 99202
rect 5906 99150 5908 99202
rect 5852 98532 5908 99150
rect 5404 98306 5460 98318
rect 5404 98254 5406 98306
rect 5458 98254 5460 98306
rect 5404 95844 5460 98254
rect 5516 98194 5572 98206
rect 5516 98142 5518 98194
rect 5570 98142 5572 98194
rect 5516 96180 5572 98142
rect 5852 98084 5908 98476
rect 5964 98418 6020 99932
rect 5964 98366 5966 98418
rect 6018 98366 6020 98418
rect 5964 98308 6020 98366
rect 5964 98242 6020 98252
rect 6076 99202 6132 99214
rect 6300 99204 6356 100268
rect 6524 99988 6580 100716
rect 6076 99150 6078 99202
rect 6130 99150 6132 99202
rect 6076 98084 6132 99150
rect 5852 98028 6132 98084
rect 6188 99202 6356 99204
rect 6188 99150 6302 99202
rect 6354 99150 6356 99202
rect 6188 99148 6356 99150
rect 6188 98644 6244 99148
rect 6300 99138 6356 99148
rect 6412 99932 6580 99988
rect 5516 96114 5572 96124
rect 5628 97636 5684 97646
rect 5404 95778 5460 95788
rect 5628 95396 5684 97580
rect 5740 97634 5796 97646
rect 5740 97582 5742 97634
rect 5794 97582 5796 97634
rect 5740 96740 5796 97582
rect 5852 97636 5908 97646
rect 5852 97542 5908 97580
rect 5964 97468 6020 98028
rect 6076 97636 6132 97674
rect 6076 97570 6132 97580
rect 6188 97634 6244 98588
rect 6188 97582 6190 97634
rect 6242 97582 6244 97634
rect 5964 97412 6132 97468
rect 5740 96404 5796 96684
rect 5964 96404 6020 96414
rect 5740 96348 5964 96404
rect 5180 93044 5236 93054
rect 5180 92950 5236 92988
rect 4620 92930 5012 92932
rect 4620 92878 4622 92930
rect 4674 92878 5012 92930
rect 4620 92876 5012 92878
rect 2940 92306 2996 92316
rect 4284 92372 4340 92382
rect 2492 92260 2548 92270
rect 2492 92166 2548 92204
rect 3276 92260 3332 92270
rect 3276 92166 3332 92204
rect 3052 92148 3108 92158
rect 2940 92146 3108 92148
rect 2940 92094 3054 92146
rect 3106 92094 3108 92146
rect 2940 92092 3108 92094
rect 1820 92036 1876 92046
rect 1820 91362 1876 91980
rect 2828 92036 2884 92046
rect 2828 91942 2884 91980
rect 2940 91588 2996 92092
rect 3052 92082 3108 92092
rect 3388 92146 3444 92158
rect 3388 92094 3390 92146
rect 3442 92094 3444 92146
rect 2492 91532 2996 91588
rect 3388 91588 3444 92094
rect 2492 91474 2548 91532
rect 3388 91522 3444 91532
rect 2492 91422 2494 91474
rect 2546 91422 2548 91474
rect 2492 91410 2548 91422
rect 1820 91310 1822 91362
rect 1874 91310 1876 91362
rect 1820 91298 1876 91310
rect 1708 90580 1764 90590
rect 1708 88898 1764 90524
rect 1708 88846 1710 88898
rect 1762 88846 1764 88898
rect 1708 88834 1764 88846
rect 2492 88900 2548 88910
rect 1708 88116 1764 88126
rect 1708 87668 1764 88060
rect 2492 88114 2548 88844
rect 3836 88900 3892 88910
rect 3836 88806 3892 88844
rect 2492 88062 2494 88114
rect 2546 88062 2548 88114
rect 2492 88050 2548 88062
rect 2828 88114 2884 88126
rect 2828 88062 2830 88114
rect 2882 88062 2884 88114
rect 2044 88002 2100 88014
rect 2044 87950 2046 88002
rect 2098 87950 2100 88002
rect 1820 87668 1876 87678
rect 1708 87666 1876 87668
rect 1708 87614 1822 87666
rect 1874 87614 1876 87666
rect 1708 87612 1876 87614
rect 1820 87602 1876 87612
rect 2044 87556 2100 87950
rect 2828 88004 2884 88062
rect 2828 87938 2884 87948
rect 3388 88004 3444 88014
rect 3388 87910 3444 87948
rect 2044 87490 2100 87500
rect 3052 87444 3108 87454
rect 2044 85988 2100 85998
rect 2044 85894 2100 85932
rect 1708 85874 1764 85886
rect 1708 85822 1710 85874
rect 1762 85822 1764 85874
rect 1708 85428 1764 85822
rect 3052 85874 3108 87388
rect 3836 86546 3892 86558
rect 3836 86494 3838 86546
rect 3890 86494 3892 86546
rect 3500 86436 3556 86446
rect 3836 86436 3892 86494
rect 4172 86436 4228 86446
rect 3500 86434 3780 86436
rect 3500 86382 3502 86434
rect 3554 86382 3780 86434
rect 3500 86380 3780 86382
rect 3836 86434 4228 86436
rect 3836 86382 4174 86434
rect 4226 86382 4228 86434
rect 3836 86380 4228 86382
rect 3500 86370 3556 86380
rect 3724 85986 3780 86380
rect 4172 86370 4228 86380
rect 3724 85934 3726 85986
rect 3778 85934 3780 85986
rect 3724 85922 3780 85934
rect 3052 85822 3054 85874
rect 3106 85822 3108 85874
rect 3052 85810 3108 85822
rect 1708 85362 1764 85372
rect 2492 85762 2548 85774
rect 2492 85710 2494 85762
rect 2546 85710 2548 85762
rect 2492 85428 2548 85710
rect 4284 85708 4340 92316
rect 4620 92036 4676 92876
rect 4620 91970 4676 91980
rect 4614 91756 4878 91766
rect 4670 91700 4718 91756
rect 4774 91700 4822 91756
rect 4614 91690 4878 91700
rect 4620 91474 4676 91486
rect 4620 91422 4622 91474
rect 4674 91422 4676 91474
rect 4620 90804 4676 91422
rect 4732 90804 4788 90814
rect 4620 90802 4788 90804
rect 4620 90750 4734 90802
rect 4786 90750 4788 90802
rect 4620 90748 4788 90750
rect 4732 90738 4788 90748
rect 4508 90692 4564 90702
rect 4508 90598 4564 90636
rect 4614 90188 4878 90198
rect 4670 90132 4718 90188
rect 4774 90132 4822 90188
rect 4614 90122 4878 90132
rect 4844 89908 4900 89918
rect 4956 89908 5012 92876
rect 5068 92146 5124 92158
rect 5068 92094 5070 92146
rect 5122 92094 5124 92146
rect 5068 91140 5124 92094
rect 5068 91046 5124 91084
rect 5292 90804 5348 93548
rect 5404 95284 5460 95294
rect 5404 95170 5460 95228
rect 5404 95118 5406 95170
rect 5458 95118 5460 95170
rect 5404 95058 5460 95118
rect 5404 95006 5406 95058
rect 5458 95006 5460 95058
rect 5404 92260 5460 95006
rect 5628 95284 5684 95340
rect 5964 95394 6020 96348
rect 6076 95956 6132 97412
rect 6076 95862 6132 95900
rect 5964 95342 5966 95394
rect 6018 95342 6020 95394
rect 5964 95330 6020 95342
rect 6076 95508 6132 95518
rect 5852 95284 5908 95294
rect 5628 95282 5908 95284
rect 5628 95230 5854 95282
rect 5906 95230 5908 95282
rect 5628 95228 5908 95230
rect 5628 94108 5684 95228
rect 5852 94948 5908 95228
rect 6076 95284 6132 95452
rect 6188 95284 6244 97582
rect 6300 97748 6356 97758
rect 6300 96962 6356 97692
rect 6300 96910 6302 96962
rect 6354 96910 6356 96962
rect 6300 96898 6356 96910
rect 6412 95732 6468 99932
rect 6748 99876 6804 102844
rect 6860 102834 6916 102844
rect 7644 102340 7700 102350
rect 8204 102340 8260 103292
rect 8316 103236 8372 103246
rect 8316 103122 8372 103180
rect 8316 103070 8318 103122
rect 8370 103070 8372 103122
rect 8316 102788 8372 103070
rect 8316 102722 8372 102732
rect 8316 102564 8372 102574
rect 8428 102564 8484 103628
rect 8316 102562 8484 102564
rect 8316 102510 8318 102562
rect 8370 102510 8484 102562
rect 8316 102508 8484 102510
rect 8316 102498 8372 102508
rect 7644 102338 8260 102340
rect 7644 102286 7646 102338
rect 7698 102286 8260 102338
rect 7644 102284 8260 102286
rect 6860 102116 6916 102126
rect 7308 102116 7364 102126
rect 6860 101556 6916 102060
rect 6860 101490 6916 101500
rect 7196 102114 7364 102116
rect 7196 102062 7310 102114
rect 7362 102062 7364 102114
rect 7196 102060 7364 102062
rect 6524 99820 6804 99876
rect 7084 99876 7140 99886
rect 6524 99090 6580 99820
rect 6636 99204 6692 99214
rect 6636 99110 6692 99148
rect 6748 99202 6804 99214
rect 6748 99150 6750 99202
rect 6802 99150 6804 99202
rect 6524 99038 6526 99090
rect 6578 99038 6580 99090
rect 6524 99026 6580 99038
rect 6748 98756 6804 99150
rect 6860 99092 6916 99102
rect 6860 98978 6916 99036
rect 7084 99090 7140 99820
rect 7084 99038 7086 99090
rect 7138 99038 7140 99090
rect 7084 99026 7140 99038
rect 6860 98926 6862 98978
rect 6914 98926 6916 98978
rect 6860 98868 6916 98926
rect 7196 98868 7252 102060
rect 7308 102050 7364 102060
rect 7644 101108 7700 102284
rect 7756 102114 7812 102126
rect 7756 102062 7758 102114
rect 7810 102062 7812 102114
rect 7756 101332 7812 102062
rect 8540 102116 8596 103740
rect 8876 103572 8932 103852
rect 8876 103236 8932 103516
rect 8988 103346 9044 104076
rect 8988 103294 8990 103346
rect 9042 103294 9044 103346
rect 8988 103282 9044 103294
rect 8764 103180 8932 103236
rect 8764 103122 8820 103180
rect 8764 103070 8766 103122
rect 8818 103070 8820 103122
rect 8764 103058 8820 103070
rect 8988 103124 9044 103134
rect 8876 103012 8932 103022
rect 8988 103012 9044 103068
rect 8876 103010 9044 103012
rect 8876 102958 8878 103010
rect 8930 102958 9044 103010
rect 8876 102956 9044 102958
rect 8876 102946 8932 102956
rect 8988 102788 9044 102798
rect 8988 102564 9044 102732
rect 8652 102508 9044 102564
rect 8652 102450 8708 102508
rect 8652 102398 8654 102450
rect 8706 102398 8708 102450
rect 8652 102386 8708 102398
rect 8764 102340 8820 102350
rect 8652 102116 8708 102126
rect 8540 102060 8652 102116
rect 8652 102050 8708 102060
rect 8016 101948 8280 101958
rect 8072 101892 8120 101948
rect 8176 101892 8224 101948
rect 8016 101882 8280 101892
rect 8540 101892 8596 101902
rect 7756 101266 7812 101276
rect 7308 101052 7700 101108
rect 7308 100770 7364 101052
rect 7420 100884 7476 100922
rect 7420 100818 7476 100828
rect 7308 100718 7310 100770
rect 7362 100718 7364 100770
rect 7308 100436 7364 100718
rect 7420 100660 7476 100670
rect 7420 100548 7476 100604
rect 7756 100658 7812 100670
rect 7756 100606 7758 100658
rect 7810 100606 7812 100658
rect 7420 100546 7588 100548
rect 7420 100494 7422 100546
rect 7474 100494 7588 100546
rect 7420 100492 7588 100494
rect 7420 100482 7476 100492
rect 7308 99876 7364 100380
rect 7532 99988 7588 100492
rect 7756 100324 7812 100606
rect 8016 100380 8280 100390
rect 8072 100324 8120 100380
rect 8176 100324 8224 100380
rect 8016 100314 8280 100324
rect 7756 100258 7812 100268
rect 7532 99922 7588 99932
rect 8540 100098 8596 101836
rect 8764 101442 8820 102284
rect 8764 101390 8766 101442
rect 8818 101390 8820 101442
rect 8764 100884 8820 101390
rect 8876 102338 8932 102350
rect 8876 102286 8878 102338
rect 8930 102286 8932 102338
rect 8876 100996 8932 102286
rect 8876 100930 8932 100940
rect 8988 102228 9044 102238
rect 8764 100818 8820 100828
rect 8988 100660 9044 102172
rect 9100 100772 9156 105196
rect 9212 104132 9268 105980
rect 9212 104066 9268 104076
rect 9324 104020 9380 108444
rect 9660 107602 9716 108782
rect 10780 108610 10836 108622
rect 10780 108558 10782 108610
rect 10834 108558 10836 108610
rect 9660 107550 9662 107602
rect 9714 107550 9716 107602
rect 9436 107266 9492 107278
rect 9436 107214 9438 107266
rect 9490 107214 9492 107266
rect 9436 107154 9492 107214
rect 9436 107102 9438 107154
rect 9490 107102 9492 107154
rect 9436 107090 9492 107102
rect 9660 106820 9716 107550
rect 9660 106754 9716 106764
rect 9772 107828 9828 107838
rect 9772 106370 9828 107772
rect 10780 107826 10836 108558
rect 10780 107774 10782 107826
rect 10834 107774 10836 107826
rect 9884 107604 9940 107614
rect 9884 107266 9940 107548
rect 9884 107214 9886 107266
rect 9938 107214 9940 107266
rect 9884 107154 9940 107214
rect 9884 107102 9886 107154
rect 9938 107102 9940 107154
rect 9884 107090 9940 107102
rect 9996 107044 10052 107054
rect 9884 106484 9940 106494
rect 9996 106484 10052 106988
rect 10780 107044 10836 107774
rect 11676 108612 11732 108622
rect 12124 108612 12180 109454
rect 12348 109394 12404 109902
rect 12348 109342 12350 109394
rect 12402 109342 12404 109394
rect 12348 109330 12404 109342
rect 12460 109284 12516 110236
rect 11676 108610 12180 108612
rect 11676 108558 11678 108610
rect 11730 108558 12180 108610
rect 11676 108556 12180 108558
rect 12348 109172 12516 109228
rect 12684 110178 12740 110190
rect 12684 110126 12686 110178
rect 12738 110126 12740 110178
rect 11676 107828 11732 108556
rect 11676 107826 11844 107828
rect 11676 107774 11678 107826
rect 11730 107774 11844 107826
rect 11676 107772 11844 107774
rect 11676 107762 11732 107772
rect 11418 107436 11682 107446
rect 11474 107380 11522 107436
rect 11578 107380 11626 107436
rect 11418 107370 11682 107380
rect 9884 106482 10052 106484
rect 9884 106430 9886 106482
rect 9938 106430 10052 106482
rect 9884 106428 10052 106430
rect 10108 106820 10164 106830
rect 9884 106418 9940 106428
rect 10108 106372 10164 106764
rect 9772 106318 9774 106370
rect 9826 106318 9828 106370
rect 9772 105924 9828 106318
rect 9548 105868 9828 105924
rect 9996 106316 10164 106372
rect 9996 106260 10052 106316
rect 9324 103964 9492 104020
rect 9324 103794 9380 103806
rect 9324 103742 9326 103794
rect 9378 103742 9380 103794
rect 9212 103682 9268 103694
rect 9212 103630 9214 103682
rect 9266 103630 9268 103682
rect 9212 102900 9268 103630
rect 9212 102834 9268 102844
rect 9212 102676 9268 102686
rect 9212 102338 9268 102620
rect 9212 102286 9214 102338
rect 9266 102286 9268 102338
rect 9212 101892 9268 102286
rect 9324 102340 9380 103742
rect 9436 103124 9492 103964
rect 9548 103796 9604 105868
rect 9660 105700 9716 105710
rect 9996 105700 10052 106204
rect 9660 105698 10052 105700
rect 9660 105646 9662 105698
rect 9714 105646 10052 105698
rect 9660 105644 10052 105646
rect 9660 104690 9716 105644
rect 10780 105474 10836 106988
rect 11452 107044 11508 107054
rect 11452 106950 11508 106988
rect 11788 107044 11844 107772
rect 12124 107826 12180 107838
rect 12124 107774 12126 107826
rect 12178 107774 12180 107826
rect 12124 107604 12180 107774
rect 12348 107826 12404 109172
rect 12572 108612 12628 108622
rect 12684 108612 12740 110126
rect 12908 110178 12964 110190
rect 12908 110126 12910 110178
rect 12962 110126 12964 110178
rect 12796 110068 12852 110078
rect 12796 108834 12852 110012
rect 12908 109284 12964 110126
rect 12908 109218 12964 109228
rect 13020 109282 13076 112476
rect 13468 112306 13524 113036
rect 13804 113026 13860 113036
rect 13468 112254 13470 112306
rect 13522 112254 13524 112306
rect 13468 112242 13524 112254
rect 13916 112530 13972 112542
rect 13916 112478 13918 112530
rect 13970 112478 13972 112530
rect 13916 111746 13972 112478
rect 13916 111694 13918 111746
rect 13970 111694 13972 111746
rect 13692 111522 13748 111534
rect 13692 111470 13694 111522
rect 13746 111470 13748 111522
rect 13132 110852 13188 110862
rect 13580 110852 13636 110862
rect 13692 110852 13748 111470
rect 13132 110850 13748 110852
rect 13132 110798 13134 110850
rect 13186 110798 13582 110850
rect 13634 110798 13748 110850
rect 13132 110796 13748 110798
rect 13916 110962 13972 111694
rect 13916 110910 13918 110962
rect 13970 110910 13972 110962
rect 13132 110786 13188 110796
rect 13020 109230 13022 109282
rect 13074 109230 13076 109282
rect 13020 109218 13076 109230
rect 13468 110066 13524 110796
rect 13580 110786 13636 110796
rect 13468 110014 13470 110066
rect 13522 110014 13524 110066
rect 13468 109284 13524 110014
rect 13916 110178 13972 110910
rect 14700 112532 14756 114044
rect 14820 112924 15084 112934
rect 14876 112868 14924 112924
rect 14980 112868 15028 112924
rect 14820 112858 15084 112868
rect 14700 111746 14756 112476
rect 14700 111694 14702 111746
rect 14754 111694 14756 111746
rect 14700 110962 14756 111694
rect 14820 111356 15084 111366
rect 14876 111300 14924 111356
rect 14980 111300 15028 111356
rect 14820 111290 15084 111300
rect 14700 110910 14702 110962
rect 14754 110910 14756 110962
rect 14476 110740 14532 110750
rect 13916 110126 13918 110178
rect 13970 110126 13972 110178
rect 13916 110068 13972 110126
rect 13916 110002 13972 110012
rect 14252 110180 14308 110190
rect 13580 109954 13636 109966
rect 13580 109902 13582 109954
rect 13634 109902 13636 109954
rect 13580 109394 13636 109902
rect 14252 109506 14308 110124
rect 14252 109454 14254 109506
rect 14306 109454 14308 109506
rect 13580 109342 13582 109394
rect 13634 109342 13636 109394
rect 13580 109330 13636 109342
rect 14028 109396 14084 109406
rect 13468 109218 13524 109228
rect 12796 108782 12798 108834
rect 12850 108782 12852 108834
rect 12796 108770 12852 108782
rect 14028 108722 14084 109340
rect 14252 108834 14308 109454
rect 14252 108782 14254 108834
rect 14306 108782 14308 108834
rect 14252 108770 14308 108782
rect 14476 110180 14532 110684
rect 14700 110180 14756 110910
rect 14476 110178 14756 110180
rect 14476 110126 14702 110178
rect 14754 110126 14756 110178
rect 14476 110124 14756 110126
rect 14028 108670 14030 108722
rect 14082 108670 14084 108722
rect 12796 108612 12852 108622
rect 12684 108610 12852 108612
rect 12684 108558 12798 108610
rect 12850 108558 12852 108610
rect 12684 108556 12852 108558
rect 12572 108518 12628 108556
rect 12796 107940 12852 108556
rect 13692 108610 13748 108622
rect 13692 108558 13694 108610
rect 13746 108558 13748 108610
rect 13692 108500 13748 108558
rect 13692 108434 13748 108444
rect 13132 107940 13188 107950
rect 12796 107938 13188 107940
rect 12796 107886 13134 107938
rect 13186 107886 13188 107938
rect 12796 107884 13188 107886
rect 13132 107874 13188 107884
rect 12348 107774 12350 107826
rect 12402 107774 12404 107826
rect 12236 107716 12292 107726
rect 12236 107622 12292 107660
rect 12124 107538 12180 107548
rect 10780 105422 10782 105474
rect 10834 105422 10836 105474
rect 10780 105410 10836 105422
rect 11228 106146 11284 106158
rect 11228 106094 11230 106146
rect 11282 106094 11284 106146
rect 10444 105364 10500 105374
rect 10444 104802 10500 105308
rect 10444 104750 10446 104802
rect 10498 104750 10500 104802
rect 10444 104738 10500 104750
rect 9660 104638 9662 104690
rect 9714 104638 9716 104690
rect 9660 104626 9716 104638
rect 11228 104690 11284 106094
rect 11418 105868 11682 105878
rect 11474 105812 11522 105868
rect 11578 105812 11626 105868
rect 11418 105802 11682 105812
rect 11788 105700 11844 106988
rect 11676 105644 11844 105700
rect 12348 106372 12404 107774
rect 12684 107826 12740 107838
rect 12684 107774 12686 107826
rect 12738 107774 12740 107826
rect 12460 107044 12516 107054
rect 12460 106950 12516 106988
rect 12348 105700 12404 106316
rect 12684 105924 12740 107774
rect 13580 107828 13636 107838
rect 13580 107734 13636 107772
rect 14028 107714 14084 108670
rect 14476 108050 14532 110124
rect 14700 110114 14756 110124
rect 14820 109788 15084 109798
rect 14876 109732 14924 109788
rect 14980 109732 15028 109788
rect 14820 109722 15084 109732
rect 15036 109284 15092 109294
rect 15036 108722 15092 109228
rect 15036 108670 15038 108722
rect 15090 108670 15092 108722
rect 15036 108658 15092 108670
rect 14924 108612 14980 108622
rect 14924 108518 14980 108556
rect 14820 108220 15084 108230
rect 14876 108164 14924 108220
rect 14980 108164 15028 108220
rect 14820 108154 15084 108164
rect 14476 107998 14478 108050
rect 14530 107998 14532 108050
rect 14476 107986 14532 107998
rect 14924 108052 14980 108062
rect 14028 107662 14030 107714
rect 14082 107662 14084 107714
rect 14028 107156 14084 107662
rect 14924 107266 14980 107996
rect 14924 107214 14926 107266
rect 14978 107214 14980 107266
rect 14924 107202 14980 107214
rect 14252 107156 14308 107166
rect 14028 107154 14308 107156
rect 14028 107102 14254 107154
rect 14306 107102 14308 107154
rect 14028 107100 14308 107102
rect 13580 107044 13636 107054
rect 13580 106950 13636 106988
rect 13468 106932 13524 106942
rect 13468 106838 13524 106876
rect 13020 106818 13076 106830
rect 13020 106766 13022 106818
rect 13074 106766 13076 106818
rect 13020 105868 13076 106766
rect 12684 105858 12740 105868
rect 12908 105812 13076 105868
rect 13580 105924 13636 105934
rect 12684 105700 12740 105710
rect 12348 105644 12684 105700
rect 11676 105474 11732 105644
rect 11676 105422 11678 105474
rect 11730 105422 11732 105474
rect 11676 105410 11732 105422
rect 12684 105474 12740 105644
rect 12684 105422 12686 105474
rect 12738 105422 12740 105474
rect 12684 105410 12740 105422
rect 12796 105588 12852 105598
rect 12460 105250 12516 105262
rect 12460 105198 12462 105250
rect 12514 105198 12516 105250
rect 11228 104638 11230 104690
rect 11282 104638 11284 104690
rect 11228 104626 11284 104638
rect 11788 104692 11844 104702
rect 11788 104598 11844 104636
rect 11228 104468 11284 104478
rect 10108 104132 10164 104142
rect 9884 103908 9940 103918
rect 9884 103814 9940 103852
rect 9548 103730 9604 103740
rect 9660 103794 9716 103806
rect 9660 103742 9662 103794
rect 9714 103742 9716 103794
rect 9548 103348 9604 103358
rect 9548 103254 9604 103292
rect 9660 103124 9716 103742
rect 10108 103796 10164 104076
rect 11228 104018 11284 104412
rect 12460 104468 12516 105198
rect 12796 105250 12852 105532
rect 12796 105198 12798 105250
rect 12850 105198 12852 105250
rect 12460 104402 12516 104412
rect 12684 104916 12740 104926
rect 11418 104300 11682 104310
rect 11474 104244 11522 104300
rect 11578 104244 11626 104300
rect 11418 104234 11682 104244
rect 11228 103966 11230 104018
rect 11282 103966 11284 104018
rect 11228 103954 11284 103966
rect 12012 104076 12292 104132
rect 9436 103068 9604 103124
rect 9436 102898 9492 102910
rect 9436 102846 9438 102898
rect 9490 102846 9492 102898
rect 9436 102788 9492 102846
rect 9436 102722 9492 102732
rect 9324 102284 9492 102340
rect 9212 101826 9268 101836
rect 9324 100884 9380 100894
rect 9212 100772 9268 100782
rect 9100 100716 9212 100772
rect 9212 100706 9268 100716
rect 9324 100770 9380 100828
rect 9324 100718 9326 100770
rect 9378 100718 9380 100770
rect 9324 100706 9380 100718
rect 8540 100046 8542 100098
rect 8594 100046 8596 100098
rect 7420 99876 7476 99886
rect 8204 99876 8260 99886
rect 7308 99874 7476 99876
rect 7308 99822 7422 99874
rect 7474 99822 7476 99874
rect 7308 99820 7476 99822
rect 7420 99764 7476 99820
rect 7868 99874 8260 99876
rect 7868 99822 8206 99874
rect 8258 99822 8260 99874
rect 7868 99820 8260 99822
rect 7420 99708 7588 99764
rect 7420 99202 7476 99214
rect 7420 99150 7422 99202
rect 7474 99150 7476 99202
rect 7420 99092 7476 99150
rect 7420 99026 7476 99036
rect 6860 98812 7140 98868
rect 7196 98812 7364 98868
rect 6636 98700 6804 98756
rect 6636 98530 6692 98700
rect 6636 98478 6638 98530
rect 6690 98478 6692 98530
rect 6636 98466 6692 98478
rect 7084 97860 7140 98812
rect 6860 97748 6916 97758
rect 6748 97636 6804 97674
rect 6748 97570 6804 97580
rect 6860 97634 6916 97692
rect 6860 97582 6862 97634
rect 6914 97582 6916 97634
rect 6860 97570 6916 97582
rect 6636 97524 6692 97534
rect 7084 97524 7140 97804
rect 7196 97524 7252 97534
rect 7084 97522 7252 97524
rect 7084 97470 7198 97522
rect 7250 97470 7252 97522
rect 7084 97468 7252 97470
rect 6636 97412 6916 97468
rect 7196 97458 7252 97468
rect 6860 96852 6916 97412
rect 6972 97412 7028 97422
rect 6972 97410 7140 97412
rect 6972 97358 6974 97410
rect 7026 97358 7140 97410
rect 6972 97356 7140 97358
rect 6972 97346 7028 97356
rect 6972 96852 7028 96862
rect 6748 96850 7028 96852
rect 6748 96798 6974 96850
rect 7026 96798 7028 96850
rect 6748 96796 7028 96798
rect 6636 96180 6692 96190
rect 6636 96086 6692 96124
rect 6412 95676 6692 95732
rect 6524 95508 6580 95518
rect 6076 95282 6244 95284
rect 6076 95230 6078 95282
rect 6130 95230 6244 95282
rect 6076 95228 6244 95230
rect 6076 95218 6132 95228
rect 5852 94882 5908 94892
rect 5740 94612 5796 94622
rect 5740 94518 5796 94556
rect 6076 94274 6132 94286
rect 6076 94222 6078 94274
rect 6130 94222 6132 94274
rect 5628 94052 5796 94108
rect 5516 93604 5572 93614
rect 5516 93510 5572 93548
rect 5404 92194 5460 92204
rect 5740 91812 5796 94052
rect 6076 93940 6132 94222
rect 6188 94164 6244 95228
rect 6412 95452 6524 95508
rect 6188 94098 6244 94108
rect 6300 95172 6356 95182
rect 6076 93874 6132 93884
rect 6188 93604 6244 93614
rect 6076 93380 6132 93390
rect 6076 92930 6132 93324
rect 6188 93042 6244 93548
rect 6188 92990 6190 93042
rect 6242 92990 6244 93042
rect 6188 92978 6244 92990
rect 6076 92878 6078 92930
rect 6130 92878 6132 92930
rect 5292 90690 5348 90748
rect 5292 90638 5294 90690
rect 5346 90638 5348 90690
rect 5292 90626 5348 90638
rect 5628 91756 5796 91812
rect 5852 92706 5908 92718
rect 5852 92654 5854 92706
rect 5906 92654 5908 92706
rect 5852 92260 5908 92654
rect 4844 89906 5012 89908
rect 4844 89854 4846 89906
rect 4898 89854 5012 89906
rect 4844 89852 5012 89854
rect 4844 89842 4900 89852
rect 4620 89012 4676 89022
rect 4956 89012 5012 89852
rect 5628 89124 5684 91756
rect 5740 91588 5796 91598
rect 5740 91494 5796 91532
rect 5740 90692 5796 90702
rect 5852 90692 5908 92204
rect 6076 91476 6132 92878
rect 6300 92930 6356 95116
rect 6412 94722 6468 95452
rect 6524 95414 6580 95452
rect 6636 95284 6692 95676
rect 6412 94670 6414 94722
rect 6466 94670 6468 94722
rect 6412 94658 6468 94670
rect 6524 95228 6692 95284
rect 6412 93940 6468 93950
rect 6412 93492 6468 93884
rect 6412 93426 6468 93436
rect 6524 93044 6580 95228
rect 6636 94836 6692 94846
rect 6636 94610 6692 94780
rect 6636 94558 6638 94610
rect 6690 94558 6692 94610
rect 6636 94546 6692 94558
rect 6748 94724 6804 96796
rect 6972 96786 7028 96796
rect 7084 95620 7140 97356
rect 6860 95564 7140 95620
rect 7196 96068 7252 96078
rect 6860 95508 6916 95564
rect 6860 95394 6916 95452
rect 6860 95342 6862 95394
rect 6914 95342 6916 95394
rect 6860 95330 6916 95342
rect 7196 95282 7252 96012
rect 7196 95230 7198 95282
rect 7250 95230 7252 95282
rect 6972 95172 7028 95182
rect 6972 95078 7028 95116
rect 6300 92878 6302 92930
rect 6354 92878 6356 92930
rect 6300 92866 6356 92878
rect 6412 92988 6524 93044
rect 6076 91382 6132 91420
rect 5796 90636 5908 90692
rect 5740 90598 5796 90636
rect 6412 90580 6468 92988
rect 6524 92978 6580 92988
rect 6636 94164 6692 94174
rect 5852 90578 6468 90580
rect 5852 90526 6414 90578
rect 6466 90526 6468 90578
rect 5852 90524 6468 90526
rect 5852 89906 5908 90524
rect 5852 89854 5854 89906
rect 5906 89854 5908 89906
rect 5852 89842 5908 89854
rect 5404 89068 6244 89124
rect 5068 89012 5124 89022
rect 4620 89010 5124 89012
rect 4620 88958 4622 89010
rect 4674 88958 5070 89010
rect 5122 88958 5124 89010
rect 4620 88956 5124 88958
rect 4620 88946 4676 88956
rect 4614 88620 4878 88630
rect 4670 88564 4718 88620
rect 4774 88564 4822 88620
rect 4614 88554 4878 88564
rect 5068 88340 5124 88956
rect 4732 87556 4788 87566
rect 4396 87554 4788 87556
rect 4396 87502 4734 87554
rect 4786 87502 4788 87554
rect 4396 87500 4788 87502
rect 4396 86884 4452 87500
rect 4732 87490 4788 87500
rect 5068 87444 5124 88284
rect 5068 87378 5124 87388
rect 5292 87556 5348 87566
rect 4508 87332 4564 87342
rect 4508 87330 5012 87332
rect 4508 87278 4510 87330
rect 4562 87278 5012 87330
rect 4508 87276 5012 87278
rect 4508 87266 4564 87276
rect 4614 87052 4878 87062
rect 4670 86996 4718 87052
rect 4774 86996 4822 87052
rect 4614 86986 4878 86996
rect 4508 86884 4564 86894
rect 4396 86882 4564 86884
rect 4396 86830 4510 86882
rect 4562 86830 4564 86882
rect 4396 86828 4564 86830
rect 4508 86818 4564 86828
rect 4732 86772 4788 86782
rect 4956 86772 5012 87276
rect 4732 86770 5012 86772
rect 4732 86718 4734 86770
rect 4786 86718 5012 86770
rect 4732 86716 5012 86718
rect 4732 86706 4788 86716
rect 2492 85362 2548 85372
rect 3948 85652 4340 85708
rect 3948 85202 4004 85652
rect 4614 85484 4878 85494
rect 4670 85428 4718 85484
rect 4774 85428 4822 85484
rect 4614 85418 4878 85428
rect 3948 85150 3950 85202
rect 4002 85150 4004 85202
rect 3052 85092 3108 85102
rect 2940 85036 3052 85092
rect 2492 84194 2548 84206
rect 2492 84142 2494 84194
rect 2546 84142 2548 84194
rect 1708 83412 1764 83422
rect 1708 82740 1764 83356
rect 2492 83412 2548 84142
rect 2492 83346 2548 83356
rect 1708 82674 1764 82684
rect 2044 83298 2100 83310
rect 2044 83246 2046 83298
rect 2098 83246 2100 83298
rect 2044 82740 2100 83246
rect 2828 83298 2884 83310
rect 2828 83246 2830 83298
rect 2882 83246 2884 83298
rect 2828 82964 2884 83246
rect 2044 82674 2100 82684
rect 2268 82908 2884 82964
rect 2268 82738 2324 82908
rect 2268 82686 2270 82738
rect 2322 82686 2324 82738
rect 1820 82292 1876 82302
rect 1820 81954 1876 82236
rect 1820 81902 1822 81954
rect 1874 81902 1876 81954
rect 1820 81890 1876 81902
rect 2268 81956 2324 82686
rect 2604 82738 2660 82750
rect 2604 82686 2606 82738
rect 2658 82686 2660 82738
rect 2380 82626 2436 82638
rect 2380 82574 2382 82626
rect 2434 82574 2436 82626
rect 2380 82068 2436 82574
rect 2492 82068 2548 82078
rect 2380 82066 2548 82068
rect 2380 82014 2494 82066
rect 2546 82014 2548 82066
rect 2380 82012 2548 82014
rect 2492 82002 2548 82012
rect 2268 81890 2324 81900
rect 2604 81284 2660 82686
rect 2828 82516 2884 82526
rect 2828 82422 2884 82460
rect 2604 81218 2660 81228
rect 2828 80500 2884 80510
rect 2940 80500 2996 85036
rect 3052 84998 3108 85036
rect 3276 83412 3332 83422
rect 3052 83356 3276 83412
rect 3052 82738 3108 83356
rect 3276 83318 3332 83356
rect 3836 83298 3892 83310
rect 3836 83246 3838 83298
rect 3890 83246 3892 83298
rect 3052 82686 3054 82738
rect 3106 82686 3108 82738
rect 3052 82674 3108 82686
rect 3276 82740 3332 82750
rect 3388 82740 3444 82750
rect 3332 82738 3444 82740
rect 3332 82686 3390 82738
rect 3442 82686 3444 82738
rect 3332 82684 3444 82686
rect 3052 82180 3108 82190
rect 3052 81170 3108 82124
rect 3052 81118 3054 81170
rect 3106 81118 3108 81170
rect 3052 81106 3108 81118
rect 2828 80498 2996 80500
rect 2828 80446 2830 80498
rect 2882 80446 2996 80498
rect 2828 80444 2996 80446
rect 2828 80434 2884 80444
rect 2940 80388 2996 80444
rect 3052 80388 3108 80398
rect 2940 80386 3220 80388
rect 2940 80334 3054 80386
rect 3106 80334 3220 80386
rect 2940 80332 3220 80334
rect 3052 80322 3108 80332
rect 1708 80162 1764 80174
rect 1708 80110 1710 80162
rect 1762 80110 1764 80162
rect 1708 80052 1764 80110
rect 2044 80164 2100 80174
rect 2044 80070 2100 80108
rect 1708 79986 1764 79996
rect 2492 80052 2548 80062
rect 2492 79826 2548 79996
rect 2492 79774 2494 79826
rect 2546 79774 2548 79826
rect 2492 79762 2548 79774
rect 3164 78988 3220 80332
rect 3276 79602 3332 82684
rect 3388 82674 3444 82684
rect 3388 82516 3444 82526
rect 3388 82422 3444 82460
rect 3724 82516 3780 82526
rect 3836 82516 3892 83246
rect 3724 82514 3892 82516
rect 3724 82462 3726 82514
rect 3778 82462 3892 82514
rect 3724 82460 3892 82462
rect 3724 81956 3780 82460
rect 3724 81890 3780 81900
rect 3276 79550 3278 79602
rect 3330 79550 3332 79602
rect 3276 79538 3332 79550
rect 3612 79380 3668 79390
rect 3612 79378 3892 79380
rect 3612 79326 3614 79378
rect 3666 79326 3892 79378
rect 3612 79324 3892 79326
rect 3612 79314 3668 79324
rect 3164 78932 3444 78988
rect 1820 78818 1876 78830
rect 1820 78766 1822 78818
rect 1874 78766 1876 78818
rect 1708 78034 1764 78046
rect 1708 77982 1710 78034
rect 1762 77982 1764 78034
rect 1708 77364 1764 77982
rect 1708 77298 1764 77308
rect 1820 76580 1876 78766
rect 2492 78706 2548 78718
rect 2492 78654 2494 78706
rect 2546 78654 2548 78706
rect 2380 78260 2436 78270
rect 2492 78260 2548 78654
rect 3164 78596 3220 78606
rect 2380 78258 2548 78260
rect 2380 78206 2382 78258
rect 2434 78206 2548 78258
rect 2380 78204 2548 78206
rect 2828 78260 2884 78270
rect 2380 78194 2436 78204
rect 2044 78146 2100 78158
rect 2044 78094 2046 78146
rect 2098 78094 2100 78146
rect 1708 76524 1876 76580
rect 1932 77364 1988 77374
rect 1708 75684 1764 76524
rect 1820 76356 1876 76366
rect 1932 76356 1988 77308
rect 2044 77140 2100 78094
rect 2604 78036 2660 78046
rect 2828 78036 2884 78204
rect 3164 78146 3220 78540
rect 3164 78094 3166 78146
rect 3218 78094 3220 78146
rect 2604 78034 2884 78036
rect 2604 77982 2606 78034
rect 2658 77982 2884 78034
rect 2604 77980 2884 77982
rect 2604 77970 2660 77980
rect 2716 77810 2772 77822
rect 2716 77758 2718 77810
rect 2770 77758 2772 77810
rect 2716 77362 2772 77758
rect 2828 77700 2884 77980
rect 2940 78036 2996 78046
rect 2940 77942 2996 77980
rect 2828 77644 3108 77700
rect 2716 77310 2718 77362
rect 2770 77310 2772 77362
rect 2716 77298 2772 77310
rect 2044 77074 2100 77084
rect 2492 77138 2548 77150
rect 2492 77086 2494 77138
rect 2546 77086 2548 77138
rect 2156 77028 2212 77038
rect 2492 77028 2548 77086
rect 2716 77140 2772 77150
rect 2716 77046 2772 77084
rect 2156 77026 2548 77028
rect 2156 76974 2158 77026
rect 2210 76974 2548 77026
rect 2156 76972 2548 76974
rect 2156 76962 2212 76972
rect 1820 76354 1988 76356
rect 1820 76302 1822 76354
rect 1874 76302 1988 76354
rect 1820 76300 1988 76302
rect 2268 76354 2324 76972
rect 2828 76578 2884 76590
rect 2828 76526 2830 76578
rect 2882 76526 2884 76578
rect 2268 76302 2270 76354
rect 2322 76302 2324 76354
rect 1820 76290 1876 76300
rect 2268 76244 2324 76302
rect 2716 76354 2772 76366
rect 2716 76302 2718 76354
rect 2770 76302 2772 76354
rect 2604 76244 2660 76254
rect 2268 76242 2660 76244
rect 2268 76190 2606 76242
rect 2658 76190 2660 76242
rect 2268 76188 2660 76190
rect 1708 75682 1988 75684
rect 1708 75630 1710 75682
rect 1762 75630 1988 75682
rect 1708 75628 1988 75630
rect 1708 75618 1764 75628
rect 1708 74898 1764 74910
rect 1708 74846 1710 74898
rect 1762 74846 1764 74898
rect 1708 74676 1764 74846
rect 1708 74610 1764 74620
rect 1820 73890 1876 73902
rect 1820 73838 1822 73890
rect 1874 73838 1876 73890
rect 1708 73332 1764 73342
rect 1820 73332 1876 73838
rect 1708 73330 1876 73332
rect 1708 73278 1710 73330
rect 1762 73278 1876 73330
rect 1708 73276 1876 73278
rect 1708 71988 1764 73276
rect 1820 72548 1876 72558
rect 1932 72548 1988 75628
rect 2492 75570 2548 75582
rect 2492 75518 2494 75570
rect 2546 75518 2548 75570
rect 2380 75124 2436 75134
rect 2492 75124 2548 75518
rect 2380 75122 2548 75124
rect 2380 75070 2382 75122
rect 2434 75070 2548 75122
rect 2380 75068 2548 75070
rect 2380 75058 2436 75068
rect 2044 75010 2100 75022
rect 2044 74958 2046 75010
rect 2098 74958 2100 75010
rect 2044 74900 2100 74958
rect 2044 74834 2100 74844
rect 2492 74898 2548 74910
rect 2492 74846 2494 74898
rect 2546 74846 2548 74898
rect 2268 74676 2324 74686
rect 2268 74226 2324 74620
rect 2268 74174 2270 74226
rect 2322 74174 2324 74226
rect 2268 74162 2324 74174
rect 2492 74228 2548 74846
rect 2492 74162 2548 74172
rect 2604 73892 2660 76188
rect 2716 74898 2772 76302
rect 2716 74846 2718 74898
rect 2770 74846 2772 74898
rect 2716 74834 2772 74846
rect 2828 74900 2884 76526
rect 2940 75684 2996 75694
rect 2940 75010 2996 75628
rect 2940 74958 2942 75010
rect 2994 74958 2996 75010
rect 2940 74946 2996 74958
rect 2828 74834 2884 74844
rect 2940 74228 2996 74238
rect 3052 74228 3108 77644
rect 3164 75010 3220 78094
rect 3388 76580 3444 78932
rect 3500 78036 3556 78046
rect 3500 77942 3556 77980
rect 3724 78034 3780 78046
rect 3724 77982 3726 78034
rect 3778 77982 3780 78034
rect 3612 77924 3668 77934
rect 3724 77924 3780 77982
rect 3612 77922 3780 77924
rect 3612 77870 3614 77922
rect 3666 77870 3780 77922
rect 3612 77868 3780 77870
rect 3500 77252 3556 77262
rect 3500 77158 3556 77196
rect 3500 76580 3556 76590
rect 3388 76524 3500 76580
rect 3500 76514 3556 76524
rect 3612 76244 3668 77868
rect 3724 76580 3780 76590
rect 3724 76466 3780 76524
rect 3724 76414 3726 76466
rect 3778 76414 3780 76466
rect 3724 76402 3780 76414
rect 3612 76188 3780 76244
rect 3164 74958 3166 75010
rect 3218 74958 3220 75010
rect 3164 74340 3220 74958
rect 3612 74900 3668 74910
rect 3612 74806 3668 74844
rect 3220 74284 3332 74340
rect 3164 74274 3220 74284
rect 2996 74172 3108 74228
rect 2940 74162 2996 74172
rect 2940 73892 2996 73902
rect 2604 73890 2996 73892
rect 2604 73838 2942 73890
rect 2994 73838 2996 73890
rect 2604 73836 2996 73838
rect 2940 73556 2996 73836
rect 2940 73490 2996 73500
rect 2044 73444 2100 73454
rect 2044 73350 2100 73388
rect 2716 73444 2772 73454
rect 1876 72492 1988 72548
rect 2380 73332 2436 73342
rect 2380 73106 2436 73276
rect 2716 73332 2772 73388
rect 3164 73332 3220 73342
rect 2716 73330 3220 73332
rect 2716 73278 2718 73330
rect 2770 73278 3166 73330
rect 3218 73278 3220 73330
rect 2716 73276 3220 73278
rect 2716 73266 2772 73276
rect 3164 73266 3220 73276
rect 2380 73054 2382 73106
rect 2434 73054 2436 73106
rect 1820 72454 1876 72492
rect 1708 71922 1764 71932
rect 2268 71876 2324 71886
rect 2268 71782 2324 71820
rect 1820 70978 1876 70990
rect 1820 70926 1822 70978
rect 1874 70926 1876 70978
rect 1820 70532 1876 70926
rect 1708 69410 1764 69422
rect 1708 69358 1710 69410
rect 1762 69358 1764 69410
rect 1708 67284 1764 69358
rect 1820 69300 1876 70476
rect 1932 70756 1988 70766
rect 1932 69972 1988 70700
rect 2044 70754 2100 70766
rect 2044 70702 2046 70754
rect 2098 70702 2100 70754
rect 2044 70420 2100 70702
rect 2380 70756 2436 73054
rect 2716 73106 2772 73118
rect 2716 73054 2718 73106
rect 2770 73054 2772 73106
rect 2492 72434 2548 72446
rect 2492 72382 2494 72434
rect 2546 72382 2548 72434
rect 2492 71986 2548 72382
rect 2492 71934 2494 71986
rect 2546 71934 2548 71986
rect 2492 71922 2548 71934
rect 2604 71764 2660 71774
rect 2604 71670 2660 71708
rect 2716 71762 2772 73054
rect 2716 71710 2718 71762
rect 2770 71710 2772 71762
rect 2716 71698 2772 71710
rect 3052 72212 3108 72222
rect 3052 71762 3108 72156
rect 3052 71710 3054 71762
rect 3106 71710 3108 71762
rect 3052 71698 3108 71710
rect 3276 71876 3332 74284
rect 3612 74228 3668 74238
rect 3612 74114 3668 74172
rect 3612 74062 3614 74114
rect 3666 74062 3668 74114
rect 3500 73218 3556 73230
rect 3500 73166 3502 73218
rect 3554 73166 3556 73218
rect 3500 72436 3556 73166
rect 3500 72370 3556 72380
rect 2604 70756 2660 70766
rect 2380 70700 2604 70756
rect 2604 70662 2660 70700
rect 3052 70754 3108 70766
rect 3276 70756 3332 71820
rect 3612 72212 3668 74062
rect 3388 71764 3444 71774
rect 3388 71670 3444 71708
rect 3500 71650 3556 71662
rect 3500 71598 3502 71650
rect 3554 71598 3556 71650
rect 3500 71204 3556 71598
rect 3052 70702 3054 70754
rect 3106 70702 3108 70754
rect 3052 70532 3108 70702
rect 3052 70466 3108 70476
rect 3164 70700 3276 70756
rect 2268 70420 2324 70430
rect 2044 70418 2548 70420
rect 2044 70366 2270 70418
rect 2322 70366 2548 70418
rect 2044 70364 2548 70366
rect 2268 70354 2324 70364
rect 2492 70196 2548 70364
rect 2716 70196 2772 70206
rect 2492 70194 2772 70196
rect 2492 70142 2718 70194
rect 2770 70142 2772 70194
rect 2492 70140 2772 70142
rect 2716 70130 2772 70140
rect 3052 70084 3108 70094
rect 3052 69990 3108 70028
rect 2044 69972 2100 69982
rect 1932 69970 2324 69972
rect 1932 69918 2046 69970
rect 2098 69918 2324 69970
rect 1932 69916 2324 69918
rect 2044 69906 2100 69916
rect 1820 69234 1876 69244
rect 1596 67228 1764 67284
rect 1820 67618 1876 67630
rect 1820 67566 1822 67618
rect 1874 67566 1876 67618
rect 1596 67060 1652 67228
rect 1596 66388 1652 67004
rect 1708 67060 1764 67070
rect 1820 67060 1876 67566
rect 2044 67172 2100 67182
rect 2044 67078 2100 67116
rect 1708 67058 1876 67060
rect 1708 67006 1710 67058
rect 1762 67006 1876 67058
rect 1708 67004 1876 67006
rect 1708 66612 1764 67004
rect 2268 66836 2324 69916
rect 2380 69970 2436 69982
rect 2380 69918 2382 69970
rect 2434 69918 2436 69970
rect 2380 68404 2436 69918
rect 2492 69300 2548 69310
rect 2492 69298 2660 69300
rect 2492 69246 2494 69298
rect 2546 69246 2660 69298
rect 2492 69244 2660 69246
rect 2492 69234 2548 69244
rect 2604 68850 2660 69244
rect 2604 68798 2606 68850
rect 2658 68798 2660 68850
rect 2604 68786 2660 68798
rect 3052 68740 3108 68750
rect 3164 68740 3220 70700
rect 3276 70690 3332 70700
rect 3388 71202 3556 71204
rect 3388 71150 3502 71202
rect 3554 71150 3556 71202
rect 3388 71148 3556 71150
rect 3388 69076 3444 71148
rect 3500 71138 3556 71148
rect 3388 69010 3444 69020
rect 3500 70980 3556 70990
rect 3612 70980 3668 72156
rect 3500 70978 3668 70980
rect 3500 70926 3502 70978
rect 3554 70926 3668 70978
rect 3500 70924 3668 70926
rect 3500 68852 3556 70924
rect 3724 70588 3780 76188
rect 3836 71092 3892 79324
rect 3948 72324 4004 85150
rect 4956 85092 5012 86716
rect 5292 85708 5348 87500
rect 5404 87444 5460 89068
rect 6076 88900 6132 88910
rect 5628 88450 5684 88462
rect 5628 88398 5630 88450
rect 5682 88398 5684 88450
rect 5404 87442 5572 87444
rect 5404 87390 5406 87442
rect 5458 87390 5572 87442
rect 5404 87388 5572 87390
rect 5404 87378 5460 87388
rect 5516 85764 5572 87388
rect 5628 87442 5684 88398
rect 5740 88340 5796 88350
rect 6076 88340 6132 88844
rect 5796 88284 6132 88340
rect 5740 88246 5796 88284
rect 5628 87390 5630 87442
rect 5682 87390 5684 87442
rect 5628 87378 5684 87390
rect 6076 87442 6132 88284
rect 6188 88338 6244 89068
rect 6412 89012 6468 90524
rect 6524 91362 6580 91374
rect 6524 91310 6526 91362
rect 6578 91310 6580 91362
rect 6524 90804 6580 91310
rect 6524 89236 6580 90748
rect 6524 89170 6580 89180
rect 6468 88956 6580 89012
rect 6412 88946 6468 88956
rect 6188 88286 6190 88338
rect 6242 88286 6244 88338
rect 6188 88274 6244 88286
rect 6076 87390 6078 87442
rect 6130 87390 6132 87442
rect 6076 86770 6132 87390
rect 6076 86718 6078 86770
rect 6130 86718 6132 86770
rect 5852 85764 5908 85774
rect 5516 85708 5852 85764
rect 4956 84532 5012 85036
rect 4956 84466 5012 84476
rect 5068 85652 5348 85708
rect 5852 85670 5908 85708
rect 4614 83916 4878 83926
rect 4670 83860 4718 83916
rect 4774 83860 4822 83916
rect 4614 83850 4878 83860
rect 4172 83412 4228 83422
rect 4060 83300 4116 83310
rect 4060 82738 4116 83244
rect 4060 82686 4062 82738
rect 4114 82686 4116 82738
rect 4060 82516 4116 82686
rect 4060 82450 4116 82460
rect 4172 83298 4228 83356
rect 4172 83246 4174 83298
rect 4226 83246 4228 83298
rect 4060 80500 4116 80510
rect 4172 80500 4228 83246
rect 4620 83300 4676 83310
rect 4620 83206 4676 83244
rect 5068 83298 5124 85652
rect 6076 84868 6132 86718
rect 6524 86772 6580 88956
rect 6636 88450 6692 94108
rect 6748 92258 6804 94668
rect 6748 92206 6750 92258
rect 6802 92206 6804 92258
rect 6748 92194 6804 92206
rect 6860 94836 6916 94846
rect 6636 88398 6638 88450
rect 6690 88398 6692 88450
rect 6636 88338 6692 88398
rect 6636 88286 6638 88338
rect 6690 88286 6692 88338
rect 6636 88274 6692 88286
rect 6748 91140 6804 91150
rect 6748 87444 6804 91084
rect 6860 89460 6916 94780
rect 7196 94836 7252 95230
rect 7196 94770 7252 94780
rect 7084 94388 7140 94398
rect 7084 94274 7140 94332
rect 7084 94222 7086 94274
rect 7138 94222 7140 94274
rect 7084 94164 7140 94222
rect 7308 94276 7364 98812
rect 7532 98084 7588 99708
rect 7644 99204 7700 99214
rect 7644 99110 7700 99148
rect 7532 98018 7588 98028
rect 7868 97634 7924 99820
rect 8204 99810 8260 99820
rect 8540 99428 8596 100046
rect 8540 99362 8596 99372
rect 8764 100604 9044 100660
rect 8764 100210 8820 100604
rect 8764 100158 8766 100210
rect 8818 100158 8820 100210
rect 8764 98980 8820 100158
rect 8988 100212 9044 100222
rect 8764 98914 8820 98924
rect 8876 99874 8932 99886
rect 8876 99822 8878 99874
rect 8930 99822 8932 99874
rect 8016 98812 8280 98822
rect 8072 98756 8120 98812
rect 8176 98756 8224 98812
rect 8016 98746 8280 98756
rect 8764 98420 8820 98430
rect 8764 98306 8820 98364
rect 8764 98254 8766 98306
rect 8818 98254 8820 98306
rect 8764 98242 8820 98254
rect 7868 97582 7870 97634
rect 7922 97582 7924 97634
rect 7868 97468 7924 97582
rect 8876 97468 8932 99822
rect 7308 94210 7364 94220
rect 7420 97412 7924 97468
rect 8540 97412 8932 97468
rect 7084 94098 7140 94108
rect 6972 92932 7028 92942
rect 6972 92838 7028 92876
rect 7308 91476 7364 91486
rect 7308 91362 7364 91420
rect 7308 91310 7310 91362
rect 7362 91310 7364 91362
rect 7308 91298 7364 91310
rect 6972 91138 7028 91150
rect 6972 91086 6974 91138
rect 7026 91086 7028 91138
rect 6972 90578 7028 91086
rect 7196 91138 7252 91150
rect 7196 91086 7198 91138
rect 7250 91086 7252 91138
rect 7196 90804 7252 91086
rect 7420 91140 7476 97412
rect 7532 97300 7588 97310
rect 7532 97074 7588 97244
rect 8016 97244 8280 97254
rect 8072 97188 8120 97244
rect 8176 97188 8224 97244
rect 8016 97178 8280 97188
rect 7532 97022 7534 97074
rect 7586 97022 7588 97074
rect 7532 97010 7588 97022
rect 8540 96850 8596 97412
rect 8988 97300 9044 100156
rect 9436 98532 9492 102284
rect 9548 102338 9604 103068
rect 9660 102788 9716 103068
rect 9772 103122 9828 103134
rect 9772 103070 9774 103122
rect 9826 103070 9828 103122
rect 9772 102900 9828 103070
rect 9996 103122 10052 103134
rect 9996 103070 9998 103122
rect 10050 103070 10052 103122
rect 9884 102900 9940 102910
rect 9772 102844 9884 102900
rect 9884 102834 9940 102844
rect 9660 102722 9716 102732
rect 9548 102286 9550 102338
rect 9602 102286 9604 102338
rect 9548 101668 9604 102286
rect 9660 102228 9716 102238
rect 9660 102134 9716 102172
rect 9772 102114 9828 102126
rect 9772 102062 9774 102114
rect 9826 102062 9828 102114
rect 9772 101892 9828 102062
rect 9884 102116 9940 102126
rect 9996 102116 10052 103070
rect 10108 102676 10164 103740
rect 10668 103906 10724 103918
rect 10892 103908 10948 103918
rect 10668 103854 10670 103906
rect 10722 103854 10724 103906
rect 10668 103796 10724 103854
rect 10668 103730 10724 103740
rect 10780 103906 10948 103908
rect 10780 103854 10894 103906
rect 10946 103854 10948 103906
rect 10780 103852 10948 103854
rect 10220 103682 10276 103694
rect 10220 103630 10222 103682
rect 10274 103630 10276 103682
rect 10220 103348 10276 103630
rect 10780 103348 10836 103852
rect 10892 103842 10948 103852
rect 11116 103796 11172 103806
rect 11116 103702 11172 103740
rect 11340 103684 11396 103694
rect 10220 103282 10276 103292
rect 10556 103292 10836 103348
rect 11228 103682 11396 103684
rect 11228 103630 11342 103682
rect 11394 103630 11396 103682
rect 11228 103628 11396 103630
rect 10108 102610 10164 102620
rect 10220 103122 10276 103134
rect 10220 103070 10222 103122
rect 10274 103070 10276 103122
rect 10220 102564 10276 103070
rect 10220 102498 10276 102508
rect 10332 102788 10388 102798
rect 10108 102340 10164 102350
rect 10108 102246 10164 102284
rect 9940 102060 10052 102116
rect 9884 102050 9940 102060
rect 10332 102004 10388 102732
rect 9996 101948 10388 102004
rect 9996 101892 10052 101948
rect 9772 101836 10052 101892
rect 9548 101602 9604 101612
rect 9884 101668 9940 101678
rect 9884 101574 9940 101612
rect 9772 101332 9828 101342
rect 9772 100884 9828 101276
rect 9548 100658 9604 100670
rect 9548 100606 9550 100658
rect 9602 100606 9604 100658
rect 9548 100436 9604 100606
rect 9548 100370 9604 100380
rect 9436 98466 9492 98476
rect 9548 98420 9604 98430
rect 9548 98326 9604 98364
rect 9772 98418 9828 100828
rect 9884 100212 9940 100222
rect 9996 100212 10052 101836
rect 10220 101554 10276 101566
rect 10220 101502 10222 101554
rect 10274 101502 10276 101554
rect 10220 101444 10276 101502
rect 10220 101378 10276 101388
rect 10444 100770 10500 100782
rect 10444 100718 10446 100770
rect 10498 100718 10500 100770
rect 10444 100660 10500 100718
rect 10444 100594 10500 100604
rect 10108 100436 10164 100446
rect 10164 100380 10276 100436
rect 10108 100370 10164 100380
rect 9940 100156 10052 100212
rect 9884 100146 9940 100156
rect 10108 99988 10164 99998
rect 10108 99894 10164 99932
rect 9884 99092 9940 99102
rect 9884 98530 9940 99036
rect 9884 98478 9886 98530
rect 9938 98478 9940 98530
rect 9884 98466 9940 98478
rect 9772 98366 9774 98418
rect 9826 98366 9828 98418
rect 9772 97636 9828 98366
rect 10108 98420 10164 98430
rect 10220 98420 10276 100380
rect 10556 99092 10612 103292
rect 10668 103124 10724 103162
rect 10668 103058 10724 103068
rect 10892 103124 10948 103134
rect 11116 103124 11172 103134
rect 10892 103122 11060 103124
rect 10892 103070 10894 103122
rect 10946 103070 11060 103122
rect 10892 103068 11060 103070
rect 10892 103058 10948 103068
rect 10780 103012 10836 103022
rect 10780 102918 10836 102956
rect 10668 102900 10724 102910
rect 10668 101442 10724 102844
rect 10668 101390 10670 101442
rect 10722 101390 10724 101442
rect 10668 100882 10724 101390
rect 10668 100830 10670 100882
rect 10722 100830 10724 100882
rect 10668 100436 10724 100830
rect 10668 100370 10724 100380
rect 10780 100996 10836 101006
rect 10780 99874 10836 100940
rect 10780 99822 10782 99874
rect 10834 99822 10836 99874
rect 10780 99810 10836 99822
rect 11004 99316 11060 103068
rect 11116 102900 11172 103068
rect 11116 102450 11172 102844
rect 11228 103012 11284 103628
rect 11340 103618 11396 103628
rect 11788 103460 11844 103470
rect 11788 103122 11844 103404
rect 11788 103070 11790 103122
rect 11842 103070 11844 103122
rect 11788 103058 11844 103070
rect 11228 102788 11284 102956
rect 11228 102722 11284 102732
rect 11418 102732 11682 102742
rect 11474 102676 11522 102732
rect 11578 102676 11626 102732
rect 11418 102666 11682 102676
rect 11116 102398 11118 102450
rect 11170 102398 11172 102450
rect 11116 102386 11172 102398
rect 11116 101554 11172 101566
rect 11116 101502 11118 101554
rect 11170 101502 11172 101554
rect 11116 100996 11172 101502
rect 12012 101332 12068 104076
rect 12124 103906 12180 103918
rect 12124 103854 12126 103906
rect 12178 103854 12180 103906
rect 12124 103122 12180 103854
rect 12236 103906 12292 104076
rect 12236 103854 12238 103906
rect 12290 103854 12292 103906
rect 12236 103842 12292 103854
rect 12348 104018 12404 104030
rect 12348 103966 12350 104018
rect 12402 103966 12404 104018
rect 12124 103070 12126 103122
rect 12178 103070 12180 103122
rect 12124 102340 12180 103070
rect 12236 103012 12292 103022
rect 12348 103012 12404 103966
rect 12572 103236 12628 103246
rect 12572 103122 12628 103180
rect 12572 103070 12574 103122
rect 12626 103070 12628 103122
rect 12572 103058 12628 103070
rect 12236 103010 12404 103012
rect 12236 102958 12238 103010
rect 12290 102958 12404 103010
rect 12236 102956 12404 102958
rect 12236 102564 12292 102956
rect 12684 102898 12740 104860
rect 12796 104804 12852 105198
rect 12796 104738 12852 104748
rect 12908 105250 12964 105812
rect 13468 105252 13524 105262
rect 12908 105198 12910 105250
rect 12962 105198 12964 105250
rect 12908 104132 12964 105198
rect 12908 104066 12964 104076
rect 13132 105250 13524 105252
rect 13132 105198 13470 105250
rect 13522 105198 13524 105250
rect 13132 105196 13524 105198
rect 13020 103682 13076 103694
rect 13020 103630 13022 103682
rect 13074 103630 13076 103682
rect 13020 103236 13076 103630
rect 13020 103170 13076 103180
rect 13132 103122 13188 105196
rect 13468 105186 13524 105196
rect 13580 104018 13636 105868
rect 13804 105474 13860 105486
rect 13804 105422 13806 105474
rect 13858 105422 13860 105474
rect 13804 104468 13860 105422
rect 13804 104402 13860 104412
rect 14028 105474 14084 105486
rect 14028 105422 14030 105474
rect 14082 105422 14084 105474
rect 14028 104132 14084 105422
rect 13580 103966 13582 104018
rect 13634 103966 13636 104018
rect 13580 103954 13636 103966
rect 13804 104076 14084 104132
rect 14252 104692 14308 107100
rect 14588 107042 14644 107054
rect 14588 106990 14590 107042
rect 14642 106990 14644 107042
rect 14588 106932 14644 106990
rect 14588 105924 14644 106876
rect 14820 106652 15084 106662
rect 14876 106596 14924 106652
rect 14980 106596 15028 106652
rect 14820 106586 15084 106596
rect 14588 105858 14644 105868
rect 13132 103070 13134 103122
rect 13186 103070 13188 103122
rect 13132 103058 13188 103070
rect 13804 103794 13860 104076
rect 13804 103742 13806 103794
rect 13858 103742 13860 103794
rect 13804 103012 13860 103742
rect 13804 102946 13860 102956
rect 13916 103906 13972 103918
rect 13916 103854 13918 103906
rect 13970 103854 13972 103906
rect 12684 102846 12686 102898
rect 12738 102846 12740 102898
rect 12684 102834 12740 102846
rect 12236 102562 12516 102564
rect 12236 102510 12238 102562
rect 12290 102510 12516 102562
rect 12236 102508 12516 102510
rect 12236 102498 12292 102508
rect 12124 102274 12180 102284
rect 12348 102338 12404 102350
rect 12348 102286 12350 102338
rect 12402 102286 12404 102338
rect 12236 102114 12292 102126
rect 12236 102062 12238 102114
rect 12290 102062 12292 102114
rect 12236 101554 12292 102062
rect 12236 101502 12238 101554
rect 12290 101502 12292 101554
rect 12236 101490 12292 101502
rect 12012 101266 12068 101276
rect 11418 101164 11682 101174
rect 11474 101108 11522 101164
rect 11578 101108 11626 101164
rect 11418 101098 11682 101108
rect 11116 100930 11172 100940
rect 12236 100996 12292 101006
rect 11004 99250 11060 99260
rect 11116 100098 11172 100110
rect 11116 100046 11118 100098
rect 11170 100046 11172 100098
rect 10556 99026 10612 99036
rect 10892 98644 10948 98654
rect 11116 98644 11172 100046
rect 11788 99986 11844 99998
rect 11788 99934 11790 99986
rect 11842 99934 11844 99986
rect 11418 99596 11682 99606
rect 11474 99540 11522 99596
rect 11578 99540 11626 99596
rect 11418 99530 11682 99540
rect 11788 99316 11844 99934
rect 10444 98642 11172 98644
rect 10444 98590 10894 98642
rect 10946 98590 11172 98642
rect 10444 98588 11172 98590
rect 11228 99314 11844 99316
rect 11228 99262 11790 99314
rect 11842 99262 11844 99314
rect 11228 99260 11844 99262
rect 10108 98418 10276 98420
rect 10108 98366 10110 98418
rect 10162 98366 10276 98418
rect 10108 98364 10276 98366
rect 10332 98420 10388 98430
rect 10444 98420 10500 98588
rect 10892 98578 10948 98588
rect 10332 98418 10500 98420
rect 10332 98366 10334 98418
rect 10386 98366 10500 98418
rect 10332 98364 10500 98366
rect 10780 98418 10836 98430
rect 10780 98366 10782 98418
rect 10834 98366 10836 98418
rect 9996 97636 10052 97646
rect 9772 97580 9996 97636
rect 9996 97570 10052 97580
rect 10108 97468 10164 98364
rect 10332 98354 10388 98364
rect 8988 97234 9044 97244
rect 9996 97412 10164 97468
rect 10332 98084 10388 98094
rect 9996 97188 10052 97412
rect 9996 97122 10052 97132
rect 10108 97300 10164 97310
rect 8876 97076 8932 97086
rect 8876 96982 8932 97020
rect 8540 96798 8542 96850
rect 8594 96798 8596 96850
rect 8540 96786 8596 96798
rect 8764 96852 8820 96862
rect 9100 96852 9156 96862
rect 8764 96758 8820 96796
rect 8876 96850 9156 96852
rect 8876 96798 9102 96850
rect 9154 96798 9156 96850
rect 8876 96796 9156 96798
rect 8092 96738 8148 96750
rect 8092 96686 8094 96738
rect 8146 96686 8148 96738
rect 7868 96626 7924 96638
rect 7868 96574 7870 96626
rect 7922 96574 7924 96626
rect 7756 95844 7812 95854
rect 7644 95172 7700 95182
rect 7532 95116 7644 95172
rect 7532 94948 7588 95116
rect 7644 95078 7700 95116
rect 7532 94882 7588 94892
rect 7644 94836 7700 94846
rect 7532 94276 7588 94286
rect 7532 94182 7588 94220
rect 7644 93602 7700 94780
rect 7644 93550 7646 93602
rect 7698 93550 7700 93602
rect 7644 93538 7700 93550
rect 7756 92930 7812 95788
rect 7868 95508 7924 96574
rect 8092 95844 8148 96686
rect 8092 95788 8484 95844
rect 8428 95732 8484 95788
rect 8016 95676 8280 95686
rect 8072 95620 8120 95676
rect 8176 95620 8224 95676
rect 8428 95666 8484 95676
rect 8016 95610 8280 95620
rect 8540 95620 8596 95630
rect 7868 95442 7924 95452
rect 8540 95282 8596 95564
rect 8540 95230 8542 95282
rect 8594 95230 8596 95282
rect 8092 95170 8148 95182
rect 8092 95118 8094 95170
rect 8146 95118 8148 95170
rect 8092 94724 8148 95118
rect 8092 94658 8148 94668
rect 8540 94276 8596 95230
rect 8016 94108 8280 94118
rect 8072 94052 8120 94108
rect 8176 94052 8224 94108
rect 8016 94042 8280 94052
rect 7756 92878 7758 92930
rect 7810 92878 7812 92930
rect 7756 92866 7812 92878
rect 8316 93940 8372 93950
rect 8316 92932 8372 93884
rect 8428 93714 8484 93726
rect 8428 93662 8430 93714
rect 8482 93662 8484 93714
rect 8428 93156 8484 93662
rect 8540 93716 8596 94220
rect 8876 94164 8932 96796
rect 9100 96786 9156 96796
rect 10108 96740 10164 97244
rect 10332 96964 10388 98028
rect 10220 96740 10276 96750
rect 10108 96738 10276 96740
rect 10108 96686 10222 96738
rect 10274 96686 10276 96738
rect 10108 96684 10276 96686
rect 10220 96628 10276 96684
rect 10220 96562 10276 96572
rect 10220 95508 10276 95518
rect 9660 95394 9716 95406
rect 9660 95342 9662 95394
rect 9714 95342 9716 95394
rect 9548 95284 9604 95294
rect 9212 95282 9604 95284
rect 9212 95230 9550 95282
rect 9602 95230 9604 95282
rect 9212 95228 9604 95230
rect 8988 95172 9044 95182
rect 9212 95172 9268 95228
rect 9548 95218 9604 95228
rect 9660 95284 9716 95342
rect 10220 95394 10276 95452
rect 10220 95342 10222 95394
rect 10274 95342 10276 95394
rect 10220 95330 10276 95342
rect 9660 95218 9716 95228
rect 10332 95282 10388 96908
rect 10332 95230 10334 95282
rect 10386 95230 10388 95282
rect 10332 95218 10388 95230
rect 10444 97972 10500 97982
rect 10444 97522 10500 97916
rect 10444 97470 10446 97522
rect 10498 97470 10500 97522
rect 8988 95170 9268 95172
rect 8988 95118 8990 95170
rect 9042 95118 9268 95170
rect 8988 95116 9268 95118
rect 8988 95106 9044 95116
rect 9660 95058 9716 95070
rect 9660 95006 9662 95058
rect 9714 95006 9716 95058
rect 9660 94612 9716 95006
rect 9772 94612 9828 94622
rect 9660 94610 9828 94612
rect 9660 94558 9774 94610
rect 9826 94558 9828 94610
rect 9660 94556 9828 94558
rect 9772 94546 9828 94556
rect 10444 94498 10500 97470
rect 10780 97468 10836 98366
rect 10780 97412 11060 97468
rect 10556 97188 10612 97198
rect 10556 95282 10612 97132
rect 10892 96850 10948 96862
rect 10892 96798 10894 96850
rect 10946 96798 10948 96850
rect 10780 96180 10836 96190
rect 10556 95230 10558 95282
rect 10610 95230 10612 95282
rect 10556 95218 10612 95230
rect 10668 95732 10724 95742
rect 10444 94446 10446 94498
rect 10498 94446 10500 94498
rect 8876 94108 9380 94164
rect 8764 93996 9044 94052
rect 8652 93940 8708 93950
rect 8764 93940 8820 93996
rect 8652 93938 8820 93940
rect 8652 93886 8654 93938
rect 8706 93886 8820 93938
rect 8652 93884 8820 93886
rect 8988 93940 9044 93996
rect 8988 93884 9268 93940
rect 8652 93874 8708 93884
rect 8652 93716 8708 93726
rect 8540 93714 8708 93716
rect 8540 93662 8654 93714
rect 8706 93662 8708 93714
rect 8540 93660 8708 93662
rect 8652 93650 8708 93660
rect 8764 93716 8820 93726
rect 8428 93100 8596 93156
rect 8428 92932 8484 92942
rect 8372 92930 8484 92932
rect 8372 92878 8430 92930
rect 8482 92878 8484 92930
rect 8372 92876 8484 92878
rect 8316 92838 8372 92876
rect 7532 92706 7588 92718
rect 8092 92708 8148 92718
rect 7532 92654 7534 92706
rect 7586 92654 7588 92706
rect 7532 92260 7588 92654
rect 7868 92706 8148 92708
rect 7868 92654 8094 92706
rect 8146 92654 8148 92706
rect 7868 92652 8148 92654
rect 7868 92484 7924 92652
rect 8092 92642 8148 92652
rect 7532 92194 7588 92204
rect 7644 92428 7924 92484
rect 8016 92540 8280 92550
rect 8072 92484 8120 92540
rect 8176 92484 8224 92540
rect 8016 92474 8280 92484
rect 7420 91074 7476 91084
rect 7196 90738 7252 90748
rect 7532 90692 7588 90702
rect 6972 90526 6974 90578
rect 7026 90526 7028 90578
rect 6972 90514 7028 90526
rect 7084 90580 7140 90590
rect 7420 90580 7476 90590
rect 7084 90578 7476 90580
rect 7084 90526 7086 90578
rect 7138 90526 7422 90578
rect 7474 90526 7476 90578
rect 7084 90524 7476 90526
rect 7084 90514 7140 90524
rect 7420 90514 7476 90524
rect 6860 89404 7140 89460
rect 6860 89236 6916 89246
rect 6860 89010 6916 89180
rect 6860 88958 6862 89010
rect 6914 88958 6916 89010
rect 6860 88946 6916 88958
rect 7084 88786 7140 89404
rect 7196 89012 7252 89022
rect 7196 88918 7252 88956
rect 7084 88734 7086 88786
rect 7138 88734 7140 88786
rect 6860 88450 6916 88462
rect 6860 88398 6862 88450
rect 6914 88398 6916 88450
rect 6860 87554 6916 88398
rect 7084 88340 7140 88734
rect 7532 88788 7588 90636
rect 7644 89012 7700 92428
rect 7980 91364 8036 91374
rect 8428 91364 8484 92876
rect 7980 91362 8484 91364
rect 7980 91310 7982 91362
rect 8034 91310 8484 91362
rect 7980 91308 8484 91310
rect 7980 91298 8036 91308
rect 8016 90972 8280 90982
rect 8072 90916 8120 90972
rect 8176 90916 8224 90972
rect 8016 90906 8280 90916
rect 8428 90804 8484 90814
rect 8540 90804 8596 93100
rect 8484 90748 8596 90804
rect 8652 91250 8708 91262
rect 8652 91198 8654 91250
rect 8706 91198 8708 91250
rect 8652 90802 8708 91198
rect 8652 90750 8654 90802
rect 8706 90750 8708 90802
rect 8428 90690 8484 90748
rect 8652 90738 8708 90750
rect 8428 90638 8430 90690
rect 8482 90638 8484 90690
rect 8428 90626 8484 90638
rect 8764 90692 8820 93660
rect 8988 93714 9044 93726
rect 8988 93662 8990 93714
rect 9042 93662 9044 93714
rect 8988 92372 9044 93662
rect 9212 93042 9268 93884
rect 9212 92990 9214 93042
rect 9266 92990 9268 93042
rect 9212 92978 9268 92990
rect 8988 92306 9044 92316
rect 8764 90598 8820 90636
rect 7756 90580 7812 90590
rect 8876 90580 8932 90590
rect 7756 90578 8036 90580
rect 7756 90526 7758 90578
rect 7810 90526 8036 90578
rect 7756 90524 8036 90526
rect 7756 90514 7812 90524
rect 7980 89906 8036 90524
rect 8092 90468 8148 90478
rect 8092 90374 8148 90412
rect 7980 89854 7982 89906
rect 8034 89854 8036 89906
rect 7980 89842 8036 89854
rect 8652 89794 8708 89806
rect 8652 89742 8654 89794
rect 8706 89742 8708 89794
rect 8016 89404 8280 89414
rect 8072 89348 8120 89404
rect 8176 89348 8224 89404
rect 8016 89338 8280 89348
rect 7644 88946 7700 88956
rect 7756 89236 7812 89246
rect 8652 89236 8708 89742
rect 7756 89010 7812 89180
rect 7756 88958 7758 89010
rect 7810 88958 7812 89010
rect 7756 88946 7812 88958
rect 8092 89180 8708 89236
rect 8092 88900 8148 89180
rect 8876 89124 8932 90524
rect 8988 90580 9044 90590
rect 9212 90580 9268 90590
rect 8988 90578 9212 90580
rect 8988 90526 8990 90578
rect 9042 90526 9212 90578
rect 8988 90524 9212 90526
rect 9324 90580 9380 94108
rect 9996 93940 10052 93950
rect 9884 93826 9940 93838
rect 9884 93774 9886 93826
rect 9938 93774 9940 93826
rect 9548 93714 9604 93726
rect 9548 93662 9550 93714
rect 9602 93662 9604 93714
rect 9548 93492 9604 93662
rect 9548 93426 9604 93436
rect 9884 93492 9940 93774
rect 9884 93044 9940 93436
rect 9884 92978 9940 92988
rect 9772 92260 9828 92270
rect 9772 92166 9828 92204
rect 9660 90804 9716 90814
rect 9660 90690 9716 90748
rect 9660 90638 9662 90690
rect 9714 90638 9716 90690
rect 9660 90626 9716 90638
rect 9772 90580 9828 90590
rect 9324 90524 9492 90580
rect 8988 90514 9044 90524
rect 9212 90514 9268 90524
rect 8652 89068 8932 89124
rect 8652 89010 8708 89068
rect 8652 88958 8654 89010
rect 8706 88958 8708 89010
rect 8652 88946 8708 88958
rect 8092 88806 8148 88844
rect 9100 88898 9156 88910
rect 9100 88846 9102 88898
rect 9154 88846 9156 88898
rect 7532 88732 7700 88788
rect 7196 88340 7252 88350
rect 7084 88338 7252 88340
rect 7084 88286 7198 88338
rect 7250 88286 7252 88338
rect 7084 88284 7252 88286
rect 7196 88274 7252 88284
rect 6860 87502 6862 87554
rect 6914 87502 6916 87554
rect 6860 87490 6916 87502
rect 6748 87378 6804 87388
rect 6524 86678 6580 86716
rect 7084 86882 7140 86894
rect 7084 86830 7086 86882
rect 7138 86830 7140 86882
rect 7084 86770 7140 86830
rect 7084 86718 7086 86770
rect 7138 86718 7140 86770
rect 7084 86706 7140 86718
rect 7532 86660 7588 86670
rect 7308 86100 7364 86110
rect 7308 86006 7364 86044
rect 7084 85988 7140 85998
rect 6972 85764 7028 85774
rect 6972 85670 7028 85708
rect 6524 85090 6580 85102
rect 6524 85038 6526 85090
rect 6578 85038 6580 85090
rect 6524 84868 6580 85038
rect 6076 84866 6580 84868
rect 6076 84814 6078 84866
rect 6130 84814 6580 84866
rect 6076 84812 6580 84814
rect 6076 84802 6132 84812
rect 5740 84532 5796 84542
rect 5740 84438 5796 84476
rect 5404 84194 5460 84206
rect 5404 84142 5406 84194
rect 5458 84142 5460 84194
rect 5404 83860 5460 84142
rect 5404 83804 6356 83860
rect 5740 83522 5796 83534
rect 5740 83470 5742 83522
rect 5794 83470 5796 83522
rect 5740 83412 5796 83470
rect 5740 83346 5796 83356
rect 5964 83522 6020 83534
rect 5964 83470 5966 83522
rect 6018 83470 6020 83522
rect 5068 83246 5070 83298
rect 5122 83246 5124 83298
rect 4844 82852 4900 82862
rect 4844 82758 4900 82796
rect 5068 82404 5124 83246
rect 5628 83298 5684 83310
rect 5628 83246 5630 83298
rect 5682 83246 5684 83298
rect 5628 82852 5684 83246
rect 5628 82786 5684 82796
rect 4614 82348 4878 82358
rect 5068 82348 5796 82404
rect 4670 82292 4718 82348
rect 4774 82292 4822 82348
rect 4614 82282 4878 82292
rect 4620 82068 4676 82078
rect 4956 82068 5012 82078
rect 4620 82066 5012 82068
rect 4620 82014 4622 82066
rect 4674 82014 4958 82066
rect 5010 82014 5012 82066
rect 4620 82012 5012 82014
rect 4620 82002 4676 82012
rect 4956 82002 5012 82012
rect 5740 81956 5796 82348
rect 5964 82178 6020 83470
rect 6188 83412 6244 83422
rect 6300 83412 6356 83804
rect 6412 83412 6468 83422
rect 6300 83410 6468 83412
rect 6300 83358 6414 83410
rect 6466 83358 6468 83410
rect 6300 83356 6468 83358
rect 6188 83318 6244 83356
rect 5964 82126 5966 82178
rect 6018 82126 6020 82178
rect 5964 82114 6020 82126
rect 5964 81956 6020 81966
rect 5740 81954 6020 81956
rect 5740 81902 5966 81954
rect 6018 81902 6020 81954
rect 5740 81900 6020 81902
rect 4844 81844 4900 81854
rect 4844 81058 4900 81788
rect 5628 81844 5684 81854
rect 5068 81732 5124 81742
rect 5068 81638 5124 81676
rect 4844 81006 4846 81058
rect 4898 81006 4900 81058
rect 4844 80948 4900 81006
rect 5628 81060 5684 81788
rect 5740 81060 5796 81070
rect 5628 81058 5796 81060
rect 5628 81006 5742 81058
rect 5794 81006 5796 81058
rect 5628 81004 5796 81006
rect 5180 80948 5236 80958
rect 4844 80892 5180 80948
rect 4614 80780 4878 80790
rect 4670 80724 4718 80780
rect 4774 80724 4822 80780
rect 4614 80714 4878 80724
rect 4060 80498 4228 80500
rect 4060 80446 4062 80498
rect 4114 80446 4228 80498
rect 4060 80444 4228 80446
rect 4060 79490 4116 80444
rect 5068 80162 5124 80174
rect 5068 80110 5070 80162
rect 5122 80110 5124 80162
rect 5068 80052 5124 80110
rect 5068 79986 5124 79996
rect 4508 79604 4564 79614
rect 4060 79438 4062 79490
rect 4114 79438 4116 79490
rect 4060 78708 4116 79438
rect 4396 79602 4564 79604
rect 4396 79550 4510 79602
rect 4562 79550 4564 79602
rect 4396 79548 4564 79550
rect 4396 78932 4452 79548
rect 4508 79538 4564 79548
rect 4614 79212 4878 79222
rect 4670 79156 4718 79212
rect 4774 79156 4822 79212
rect 4614 79146 4878 79156
rect 4508 78932 4564 78942
rect 4396 78876 4508 78932
rect 4508 78866 4564 78876
rect 4620 78930 4676 78942
rect 4620 78878 4622 78930
rect 4674 78878 4676 78930
rect 4060 78260 4116 78652
rect 4060 78194 4116 78204
rect 4060 77924 4116 77934
rect 4620 77924 4676 78878
rect 4844 78932 4900 78942
rect 4844 78260 4900 78876
rect 5068 78596 5124 78606
rect 5180 78596 5236 80892
rect 5740 80274 5796 81004
rect 5740 80222 5742 80274
rect 5794 80222 5796 80274
rect 5740 80052 5796 80222
rect 5740 79986 5796 79996
rect 5852 80162 5908 80174
rect 5852 80110 5854 80162
rect 5906 80110 5908 80162
rect 5124 78540 5236 78596
rect 5292 79490 5348 79502
rect 5292 79438 5294 79490
rect 5346 79438 5348 79490
rect 5292 78596 5348 79438
rect 5852 79042 5908 80110
rect 5852 78990 5854 79042
rect 5906 78990 5908 79042
rect 5852 78978 5908 78990
rect 5852 78818 5908 78830
rect 5852 78766 5854 78818
rect 5906 78766 5908 78818
rect 5852 78708 5908 78766
rect 5852 78642 5908 78652
rect 5628 78596 5684 78606
rect 5292 78594 5684 78596
rect 5292 78542 5630 78594
rect 5682 78542 5684 78594
rect 5292 78540 5684 78542
rect 5068 78502 5124 78540
rect 5628 78530 5684 78540
rect 5292 78260 5348 78270
rect 4844 78258 5684 78260
rect 4844 78206 4846 78258
rect 4898 78206 5294 78258
rect 5346 78206 5684 78258
rect 4844 78204 5684 78206
rect 4844 78194 4900 78204
rect 5292 78194 5348 78204
rect 4060 77922 4676 77924
rect 4060 77870 4062 77922
rect 4114 77870 4676 77922
rect 4060 77868 4676 77870
rect 4060 77810 4116 77868
rect 4060 77758 4062 77810
rect 4114 77758 4116 77810
rect 4060 77746 4116 77758
rect 4614 77644 4878 77654
rect 4670 77588 4718 77644
rect 4774 77588 4822 77644
rect 4614 77578 4878 77588
rect 5628 77250 5684 78204
rect 5964 78148 6020 81900
rect 6188 81060 6244 81070
rect 6412 81060 6468 83356
rect 6524 83300 6580 84812
rect 7084 83748 7140 85932
rect 7196 85650 7252 85662
rect 7196 85598 7198 85650
rect 7250 85598 7252 85650
rect 7196 85202 7252 85598
rect 7196 85150 7198 85202
rect 7250 85150 7252 85202
rect 7196 85138 7252 85150
rect 7420 83748 7476 83758
rect 7084 83746 7476 83748
rect 7084 83694 7422 83746
rect 7474 83694 7476 83746
rect 7084 83692 7476 83694
rect 6524 81954 6580 83244
rect 6748 83412 6804 83422
rect 6748 83298 6804 83356
rect 6860 83412 6916 83422
rect 6860 83410 7028 83412
rect 6860 83358 6862 83410
rect 6914 83358 7028 83410
rect 6860 83356 7028 83358
rect 6860 83346 6916 83356
rect 6748 83246 6750 83298
rect 6802 83246 6804 83298
rect 6748 82516 6804 83246
rect 6972 82626 7028 83356
rect 7308 83300 7364 83310
rect 6972 82574 6974 82626
rect 7026 82574 7028 82626
rect 6972 82562 7028 82574
rect 7084 83298 7364 83300
rect 7084 83246 7310 83298
rect 7362 83246 7364 83298
rect 7084 83244 7364 83246
rect 6748 82450 6804 82460
rect 6524 81902 6526 81954
rect 6578 81902 6580 81954
rect 6524 81844 6580 81902
rect 7084 81844 7140 83244
rect 7308 83234 7364 83244
rect 7420 82962 7476 83692
rect 7420 82910 7422 82962
rect 7474 82910 7476 82962
rect 7420 82898 7476 82910
rect 7420 82626 7476 82638
rect 7420 82574 7422 82626
rect 7474 82574 7476 82626
rect 6524 81788 7140 81844
rect 7196 81842 7252 81854
rect 7196 81790 7198 81842
rect 7250 81790 7252 81842
rect 6636 81060 6692 81070
rect 6412 81058 6692 81060
rect 6412 81006 6638 81058
rect 6690 81006 6692 81058
rect 6412 81004 6692 81006
rect 6188 80966 6244 81004
rect 6636 80948 6692 81004
rect 6636 80882 6692 80892
rect 6748 80500 6804 81788
rect 7196 81394 7252 81790
rect 7196 81342 7198 81394
rect 7250 81342 7252 81394
rect 7196 81330 7252 81342
rect 6972 81170 7028 81182
rect 6972 81118 6974 81170
rect 7026 81118 7028 81170
rect 6972 80948 7028 81118
rect 7308 81172 7364 81182
rect 7308 81078 7364 81116
rect 7420 81170 7476 82574
rect 7420 81118 7422 81170
rect 7474 81118 7476 81170
rect 7420 81106 7476 81118
rect 6972 80882 7028 80892
rect 7084 80500 7140 80510
rect 6748 80498 7140 80500
rect 6748 80446 7086 80498
rect 7138 80446 7140 80498
rect 6748 80444 7140 80446
rect 7084 80434 7140 80444
rect 6076 80386 6132 80398
rect 6076 80334 6078 80386
rect 6130 80334 6132 80386
rect 6076 80164 6132 80334
rect 6076 80098 6132 80108
rect 6524 80162 6580 80174
rect 6524 80110 6526 80162
rect 6578 80110 6580 80162
rect 6524 80052 6580 80110
rect 6524 79986 6580 79996
rect 7532 79716 7588 86604
rect 7644 82740 7700 88732
rect 8204 88786 8260 88798
rect 8204 88734 8206 88786
rect 8258 88734 8260 88786
rect 7756 88450 7812 88462
rect 7756 88398 7758 88450
rect 7810 88398 7812 88450
rect 7756 88340 7812 88398
rect 8092 88340 8148 88350
rect 7756 88338 8148 88340
rect 7756 88286 8094 88338
rect 8146 88286 8148 88338
rect 7756 88284 8148 88286
rect 8092 88274 8148 88284
rect 8204 88226 8260 88734
rect 9100 88452 9156 88846
rect 9436 88788 9492 90524
rect 9772 90486 9828 90524
rect 9884 90578 9940 90590
rect 9884 90526 9886 90578
rect 9938 90526 9940 90578
rect 9884 90468 9940 90526
rect 9884 90402 9940 90412
rect 9436 88722 9492 88732
rect 9548 89908 9604 89918
rect 9100 88386 9156 88396
rect 8204 88174 8206 88226
rect 8258 88174 8260 88226
rect 8204 88162 8260 88174
rect 8540 88228 8596 88238
rect 9100 88228 9156 88238
rect 8540 88226 9156 88228
rect 8540 88174 8542 88226
rect 8594 88174 9102 88226
rect 9154 88174 9156 88226
rect 8540 88172 9156 88174
rect 8540 88162 8596 88172
rect 9100 88162 9156 88172
rect 9548 88228 9604 89852
rect 9996 89906 10052 93884
rect 10444 93940 10500 94446
rect 10668 94500 10724 95676
rect 10780 95282 10836 96124
rect 10780 95230 10782 95282
rect 10834 95230 10836 95282
rect 10780 95218 10836 95230
rect 10668 94434 10724 94444
rect 10780 94724 10836 94734
rect 10444 93874 10500 93884
rect 10332 93828 10388 93838
rect 10332 93734 10388 93772
rect 10780 93826 10836 94668
rect 10780 93774 10782 93826
rect 10834 93774 10836 93826
rect 10780 93762 10836 93774
rect 10332 93044 10388 93054
rect 10220 92372 10276 92382
rect 10220 92278 10276 92316
rect 10332 92370 10388 92988
rect 10556 92372 10612 92382
rect 10332 92318 10334 92370
rect 10386 92318 10388 92370
rect 10332 92306 10388 92318
rect 10444 92370 10612 92372
rect 10444 92318 10558 92370
rect 10610 92318 10612 92370
rect 10444 92316 10612 92318
rect 10444 92260 10500 92316
rect 10556 92306 10612 92316
rect 10892 92372 10948 96798
rect 11004 95956 11060 97412
rect 11228 96066 11284 99260
rect 11788 99250 11844 99260
rect 11900 98980 11956 98990
rect 11788 98532 11844 98542
rect 11788 98438 11844 98476
rect 11418 98028 11682 98038
rect 11474 97972 11522 98028
rect 11578 97972 11626 98028
rect 11418 97962 11682 97972
rect 11900 96962 11956 98924
rect 11900 96910 11902 96962
rect 11954 96910 11956 96962
rect 11900 96898 11956 96910
rect 12012 97188 12068 97198
rect 11788 96850 11844 96862
rect 11788 96798 11790 96850
rect 11842 96798 11844 96850
rect 11418 96460 11682 96470
rect 11474 96404 11522 96460
rect 11578 96404 11626 96460
rect 11418 96394 11682 96404
rect 11228 96014 11230 96066
rect 11282 96014 11284 96066
rect 11228 96002 11284 96014
rect 11788 96068 11844 96798
rect 12012 96738 12068 97132
rect 12012 96686 12014 96738
rect 12066 96686 12068 96738
rect 12012 96292 12068 96686
rect 12012 96226 12068 96236
rect 12124 97076 12180 97086
rect 12124 96180 12180 97020
rect 12236 96852 12292 100940
rect 12348 98308 12404 102286
rect 12348 98242 12404 98252
rect 12460 97076 12516 102508
rect 13580 102452 13636 102462
rect 12572 102340 12628 102350
rect 12572 102246 12628 102284
rect 12796 102338 12852 102350
rect 12796 102286 12798 102338
rect 12850 102286 12852 102338
rect 12796 101332 12852 102286
rect 13468 102340 13524 102350
rect 13468 102226 13524 102284
rect 13468 102174 13470 102226
rect 13522 102174 13524 102226
rect 13468 101444 13524 102174
rect 13580 102226 13636 102396
rect 13804 102340 13860 102350
rect 13916 102340 13972 103854
rect 14140 103682 14196 103694
rect 14140 103630 14142 103682
rect 14194 103630 14196 103682
rect 13804 102338 13972 102340
rect 13804 102286 13806 102338
rect 13858 102286 13972 102338
rect 13804 102284 13972 102286
rect 14028 103122 14084 103134
rect 14028 103070 14030 103122
rect 14082 103070 14084 103122
rect 13804 102274 13860 102284
rect 13580 102174 13582 102226
rect 13634 102174 13636 102226
rect 13580 102162 13636 102174
rect 13468 101388 13636 101444
rect 12796 101266 12852 101276
rect 12908 100996 12964 101006
rect 12572 100884 12628 100894
rect 12572 100790 12628 100828
rect 12908 100770 12964 100940
rect 12908 100718 12910 100770
rect 12962 100718 12964 100770
rect 12908 100706 12964 100718
rect 13468 100772 13524 100782
rect 13468 100678 13524 100716
rect 13580 100548 13636 101388
rect 14028 100996 14084 103070
rect 14140 102340 14196 103630
rect 14252 103572 14308 104636
rect 14588 105474 14644 105486
rect 14588 105422 14590 105474
rect 14642 105422 14644 105474
rect 14252 103010 14308 103516
rect 14252 102958 14254 103010
rect 14306 102958 14308 103010
rect 14252 102946 14308 102958
rect 14364 103682 14420 103694
rect 14364 103630 14366 103682
rect 14418 103630 14420 103682
rect 14140 102274 14196 102284
rect 14252 102338 14308 102350
rect 14252 102286 14254 102338
rect 14306 102286 14308 102338
rect 14028 100930 14084 100940
rect 14252 101442 14308 102286
rect 14252 101390 14254 101442
rect 14306 101390 14308 101442
rect 13468 100492 13636 100548
rect 12460 97010 12516 97020
rect 12572 99428 12628 99438
rect 12348 96852 12404 96862
rect 12236 96850 12404 96852
rect 12236 96798 12350 96850
rect 12402 96798 12404 96850
rect 12236 96796 12404 96798
rect 12348 96404 12404 96796
rect 12348 96338 12404 96348
rect 12572 96852 12628 99372
rect 13468 97076 13524 100492
rect 13580 99876 13636 99886
rect 13580 99782 13636 99820
rect 14252 99202 14308 101390
rect 14252 99150 14254 99202
rect 14306 99150 14308 99202
rect 14252 99138 14308 99150
rect 14140 97524 14196 97562
rect 14140 97458 14196 97468
rect 13804 97412 13860 97422
rect 13804 97410 13972 97412
rect 13804 97358 13806 97410
rect 13858 97358 13972 97410
rect 13804 97356 13972 97358
rect 13804 97346 13860 97356
rect 13468 96962 13524 97020
rect 13804 97074 13860 97086
rect 13804 97022 13806 97074
rect 13858 97022 13860 97074
rect 13468 96910 13470 96962
rect 13522 96910 13524 96962
rect 13468 96898 13524 96910
rect 13692 96964 13748 96974
rect 13692 96870 13748 96908
rect 12124 96086 12180 96124
rect 11788 96002 11844 96012
rect 12012 96066 12068 96078
rect 12012 96014 12014 96066
rect 12066 96014 12068 96066
rect 11004 95890 11060 95900
rect 11900 95956 11956 95966
rect 11340 95732 11396 95742
rect 11116 95508 11172 95518
rect 11004 95282 11060 95294
rect 11004 95230 11006 95282
rect 11058 95230 11060 95282
rect 11004 93156 11060 95230
rect 11116 94498 11172 95452
rect 11228 95396 11284 95406
rect 11228 94610 11284 95340
rect 11340 95172 11396 95676
rect 11340 95106 11396 95116
rect 11788 95060 11844 95070
rect 11788 94966 11844 95004
rect 11418 94892 11682 94902
rect 11474 94836 11522 94892
rect 11578 94836 11626 94892
rect 11418 94826 11682 94836
rect 11228 94558 11230 94610
rect 11282 94558 11284 94610
rect 11228 94546 11284 94558
rect 11676 94612 11732 94622
rect 11116 94446 11118 94498
rect 11170 94446 11172 94498
rect 11116 94434 11172 94446
rect 11340 94500 11396 94510
rect 11340 94406 11396 94444
rect 11676 94498 11732 94556
rect 11676 94446 11678 94498
rect 11730 94446 11732 94498
rect 11676 94434 11732 94446
rect 11228 94388 11284 94398
rect 11116 93940 11172 93950
rect 11116 93846 11172 93884
rect 11004 93090 11060 93100
rect 11228 92820 11284 94332
rect 11418 93324 11682 93334
rect 11474 93268 11522 93324
rect 11578 93268 11626 93324
rect 11418 93258 11682 93268
rect 11564 93156 11620 93166
rect 11564 93062 11620 93100
rect 11340 93044 11396 93054
rect 11340 92950 11396 92988
rect 11676 92820 11732 92830
rect 11228 92818 11732 92820
rect 11228 92766 11678 92818
rect 11730 92766 11732 92818
rect 11228 92764 11732 92766
rect 11676 92754 11732 92764
rect 11900 92708 11956 95900
rect 12012 95284 12068 96014
rect 12124 95956 12180 95966
rect 12124 95862 12180 95900
rect 12012 95282 12292 95284
rect 12012 95230 12014 95282
rect 12066 95230 12292 95282
rect 12012 95228 12292 95230
rect 12012 95218 12068 95228
rect 12236 93940 12292 95228
rect 12348 95282 12404 95294
rect 12348 95230 12350 95282
rect 12402 95230 12404 95282
rect 12348 95172 12404 95230
rect 12348 95106 12404 95116
rect 12460 94612 12516 94622
rect 12572 94612 12628 96796
rect 13132 96738 13188 96750
rect 13132 96686 13134 96738
rect 13186 96686 13188 96738
rect 13132 96516 13188 96686
rect 13132 96450 13188 96460
rect 13356 96628 13412 96638
rect 13356 95844 13412 96572
rect 13356 95778 13412 95788
rect 13692 95842 13748 95854
rect 13692 95790 13694 95842
rect 13746 95790 13748 95842
rect 13244 95508 13300 95518
rect 13692 95508 13748 95790
rect 13244 95414 13300 95452
rect 13468 95452 13748 95508
rect 12460 94610 12628 94612
rect 12460 94558 12462 94610
rect 12514 94558 12628 94610
rect 12460 94556 12628 94558
rect 13468 94836 13524 95452
rect 13580 95284 13636 95294
rect 13580 95190 13636 95228
rect 13692 95172 13748 95182
rect 13692 95078 13748 95116
rect 13692 94836 13748 94846
rect 13468 94780 13692 94836
rect 12460 94546 12516 94556
rect 12796 94498 12852 94510
rect 12796 94446 12798 94498
rect 12850 94446 12852 94498
rect 12348 93940 12404 93950
rect 12236 93938 12404 93940
rect 12236 93886 12350 93938
rect 12402 93886 12404 93938
rect 12236 93884 12404 93886
rect 12124 93714 12180 93726
rect 12124 93662 12126 93714
rect 12178 93662 12180 93714
rect 12124 93492 12180 93662
rect 12124 93426 12180 93436
rect 12236 92930 12292 93884
rect 12348 93874 12404 93884
rect 12796 93938 12852 94446
rect 12796 93886 12798 93938
rect 12850 93886 12852 93938
rect 12796 93874 12852 93886
rect 13468 93828 13524 94780
rect 13692 94770 13748 94780
rect 13692 94500 13748 94510
rect 13804 94500 13860 97022
rect 13916 96292 13972 97356
rect 14028 97410 14084 97422
rect 14028 97358 14030 97410
rect 14082 97358 14084 97410
rect 14028 96964 14084 97358
rect 14252 97410 14308 97422
rect 14252 97358 14254 97410
rect 14306 97358 14308 97410
rect 14252 97300 14308 97358
rect 14252 97234 14308 97244
rect 14140 97188 14196 97198
rect 14140 97076 14196 97132
rect 14364 97188 14420 103630
rect 14588 100772 14644 105422
rect 14820 105084 15084 105094
rect 14876 105028 14924 105084
rect 14980 105028 15028 105084
rect 14820 105018 15084 105028
rect 15260 104580 15316 114212
rect 15708 113988 15764 114940
rect 17276 114996 17332 115006
rect 17276 114882 17332 114940
rect 17276 114830 17278 114882
rect 17330 114830 17332 114882
rect 17276 114818 17332 114830
rect 17500 114884 17556 115612
rect 17500 114098 17556 114828
rect 17500 114046 17502 114098
rect 17554 114046 17556 114098
rect 17500 114034 17556 114046
rect 16268 113988 16324 113998
rect 15708 113986 16324 113988
rect 15708 113934 16270 113986
rect 16322 113934 16324 113986
rect 15708 113932 16324 113934
rect 15708 113874 15764 113932
rect 15708 113822 15710 113874
rect 15762 113822 15764 113874
rect 15708 112532 15764 113822
rect 16268 113428 16324 113932
rect 16380 113428 16436 113438
rect 16268 113426 16436 113428
rect 16268 113374 16382 113426
rect 16434 113374 16436 113426
rect 16268 113372 16436 113374
rect 16380 113362 16436 113372
rect 16604 112532 16660 112542
rect 15764 112476 16100 112532
rect 15708 112466 15764 112476
rect 16044 112306 16100 112476
rect 16604 112438 16660 112476
rect 17388 112532 17444 112542
rect 16044 112254 16046 112306
rect 16098 112254 16100 112306
rect 16044 111970 16100 112254
rect 16044 111918 16046 111970
rect 16098 111918 16100 111970
rect 16044 110738 16100 111918
rect 16716 111746 16772 111758
rect 16716 111694 16718 111746
rect 16770 111694 16772 111746
rect 16716 110964 16772 111694
rect 17388 111748 17444 112476
rect 17388 111654 17444 111692
rect 16716 110898 16772 110908
rect 17500 110964 17556 110974
rect 17500 110870 17556 110908
rect 16044 110686 16046 110738
rect 16098 110686 16100 110738
rect 16044 110404 16100 110686
rect 16604 110850 16660 110862
rect 16604 110798 16606 110850
rect 16658 110798 16660 110850
rect 16604 110404 16660 110798
rect 16044 110402 16660 110404
rect 16044 110350 16046 110402
rect 16098 110350 16660 110402
rect 16044 110348 16660 110350
rect 16044 110338 16100 110348
rect 16604 110290 16660 110348
rect 16604 110238 16606 110290
rect 16658 110238 16660 110290
rect 16604 110226 16660 110238
rect 15372 109396 15428 109406
rect 15372 109302 15428 109340
rect 15820 109396 15876 109406
rect 15820 109302 15876 109340
rect 16716 109396 16772 109406
rect 16716 109302 16772 109340
rect 16156 109284 16212 109294
rect 16156 109190 16212 109228
rect 16940 108836 16996 108874
rect 16940 108770 16996 108780
rect 17388 108724 17444 108734
rect 17164 108722 17444 108724
rect 17164 108670 17390 108722
rect 17442 108670 17444 108722
rect 17164 108668 17444 108670
rect 16940 108610 16996 108622
rect 16940 108558 16942 108610
rect 16994 108558 16996 108610
rect 16044 108500 16100 108510
rect 16044 108406 16100 108444
rect 16604 108498 16660 108510
rect 16604 108446 16606 108498
rect 16658 108446 16660 108498
rect 15708 108386 15764 108398
rect 15708 108334 15710 108386
rect 15762 108334 15764 108386
rect 15708 108052 15764 108334
rect 16604 108276 16660 108446
rect 16940 108388 16996 108558
rect 16940 108322 16996 108332
rect 16604 108210 16660 108220
rect 15708 107996 16772 108052
rect 15484 107044 15540 107054
rect 15708 107044 15764 107996
rect 15484 107042 15764 107044
rect 15484 106990 15486 107042
rect 15538 106990 15764 107042
rect 15484 106988 15764 106990
rect 16044 107826 16100 107838
rect 16044 107774 16046 107826
rect 16098 107774 16100 107826
rect 16044 107044 16100 107774
rect 16268 107828 16324 107838
rect 16156 107044 16212 107054
rect 16044 106988 16156 107044
rect 15484 106978 15540 106988
rect 16156 106950 16212 106988
rect 15260 104514 15316 104524
rect 15484 106258 15540 106270
rect 15484 106206 15486 106258
rect 15538 106206 15540 106258
rect 15484 104578 15540 106206
rect 15932 106258 15988 106270
rect 15932 106206 15934 106258
rect 15986 106206 15988 106258
rect 15820 106034 15876 106046
rect 15820 105982 15822 106034
rect 15874 105982 15876 106034
rect 15484 104526 15486 104578
rect 15538 104526 15540 104578
rect 15036 104356 15092 104366
rect 14700 104132 14756 104142
rect 14700 104038 14756 104076
rect 15036 103906 15092 104300
rect 15036 103854 15038 103906
rect 15090 103854 15092 103906
rect 15036 103842 15092 103854
rect 15484 103906 15540 104526
rect 15484 103854 15486 103906
rect 15538 103854 15540 103906
rect 15484 103842 15540 103854
rect 15708 105924 15764 105934
rect 14812 103684 14868 103722
rect 14812 103618 14868 103628
rect 14820 103516 15084 103526
rect 14876 103460 14924 103516
rect 14980 103460 15028 103516
rect 14820 103450 15084 103460
rect 14924 103124 14980 103134
rect 14924 103030 14980 103068
rect 14820 101948 15084 101958
rect 14876 101892 14924 101948
rect 14980 101892 15028 101948
rect 14820 101882 15084 101892
rect 14588 100706 14644 100716
rect 15484 100660 15540 100670
rect 15540 100604 15652 100660
rect 15484 100566 15540 100604
rect 14820 100380 15084 100390
rect 14876 100324 14924 100380
rect 14980 100324 15028 100380
rect 14820 100314 15084 100324
rect 15484 99316 15540 99326
rect 15484 99222 15540 99260
rect 15148 99092 15204 99102
rect 14820 98812 15084 98822
rect 14876 98756 14924 98812
rect 14980 98756 15028 98812
rect 14820 98746 15084 98756
rect 15148 97858 15204 99036
rect 15148 97806 15150 97858
rect 15202 97806 15204 97858
rect 15148 97794 15204 97806
rect 15484 99092 15540 99102
rect 15036 97748 15092 97758
rect 14700 97636 14756 97646
rect 14700 97542 14756 97580
rect 15036 97634 15092 97692
rect 15036 97582 15038 97634
rect 15090 97582 15092 97634
rect 15036 97570 15092 97582
rect 14364 97122 14420 97132
rect 14588 97524 14644 97534
rect 14140 97020 14308 97076
rect 14028 96870 14084 96908
rect 14252 96852 14308 97020
rect 14364 96852 14420 96862
rect 14252 96850 14420 96852
rect 14252 96798 14366 96850
rect 14418 96798 14420 96850
rect 14252 96796 14420 96798
rect 14364 96786 14420 96796
rect 13916 96226 13972 96236
rect 14028 96404 14084 96414
rect 14252 96404 14308 96414
rect 14028 96066 14084 96348
rect 14028 96014 14030 96066
rect 14082 96014 14084 96066
rect 14028 96002 14084 96014
rect 14140 96348 14252 96404
rect 14140 95844 14196 96348
rect 14252 96338 14308 96348
rect 14364 95844 14420 95854
rect 13916 95788 14196 95844
rect 14252 95788 14364 95844
rect 13916 95394 13972 95788
rect 13916 95342 13918 95394
rect 13970 95342 13972 95394
rect 13916 95330 13972 95342
rect 13692 94498 13860 94500
rect 13692 94446 13694 94498
rect 13746 94446 13860 94498
rect 13692 94444 13860 94446
rect 14028 95282 14084 95294
rect 14028 95230 14030 95282
rect 14082 95230 14084 95282
rect 13692 94434 13748 94444
rect 13916 94388 13972 94398
rect 13916 94294 13972 94332
rect 14028 94274 14084 95230
rect 14028 94222 14030 94274
rect 14082 94222 14084 94274
rect 14028 94210 14084 94222
rect 14140 95284 14196 95294
rect 14140 94722 14196 95228
rect 14140 94670 14142 94722
rect 14194 94670 14196 94722
rect 13916 94164 13972 94174
rect 13916 93940 13972 94108
rect 13468 93762 13524 93772
rect 13580 93938 13972 93940
rect 13580 93886 13918 93938
rect 13970 93886 13972 93938
rect 13580 93884 13972 93886
rect 12460 93716 12516 93726
rect 12460 93622 12516 93660
rect 13132 93716 13188 93726
rect 13132 93622 13188 93660
rect 12236 92878 12238 92930
rect 12290 92878 12292 92930
rect 12236 92866 12292 92878
rect 13356 93602 13412 93614
rect 13356 93550 13358 93602
rect 13410 93550 13412 93602
rect 13356 93492 13412 93550
rect 13356 92820 13412 93436
rect 13356 92754 13412 92764
rect 12684 92708 12740 92718
rect 11900 92614 11956 92652
rect 12572 92706 12740 92708
rect 12572 92654 12686 92706
rect 12738 92654 12740 92706
rect 12572 92652 12740 92654
rect 10892 92306 10948 92316
rect 12348 92372 12404 92382
rect 10108 92146 10164 92158
rect 10108 92094 10110 92146
rect 10162 92094 10164 92146
rect 10108 90804 10164 92094
rect 10108 90738 10164 90748
rect 9996 89854 9998 89906
rect 10050 89854 10052 89906
rect 9996 88228 10052 89854
rect 10332 90580 10388 90590
rect 10444 90580 10500 92204
rect 11004 92146 11060 92158
rect 11004 92094 11006 92146
rect 11058 92094 11060 92146
rect 10780 91474 10836 91486
rect 10780 91422 10782 91474
rect 10834 91422 10836 91474
rect 10556 90804 10612 90814
rect 10556 90690 10612 90748
rect 10556 90638 10558 90690
rect 10610 90638 10612 90690
rect 10556 90626 10612 90638
rect 10332 90578 10444 90580
rect 10332 90526 10334 90578
rect 10386 90526 10444 90578
rect 10332 90524 10444 90526
rect 10332 89908 10388 90524
rect 10444 90486 10500 90524
rect 10332 89842 10388 89852
rect 10668 90466 10724 90478
rect 10668 90414 10670 90466
rect 10722 90414 10724 90466
rect 10108 89012 10164 89022
rect 10108 88918 10164 88956
rect 10668 88340 10724 90414
rect 10780 89794 10836 91422
rect 10892 90692 10948 90702
rect 10892 90598 10948 90636
rect 10780 89742 10782 89794
rect 10834 89742 10836 89794
rect 10780 89730 10836 89742
rect 11004 88900 11060 92094
rect 11418 91756 11682 91766
rect 11474 91700 11522 91756
rect 11578 91700 11626 91756
rect 11418 91690 11682 91700
rect 11452 91140 11508 91150
rect 11340 91138 11508 91140
rect 11340 91086 11454 91138
rect 11506 91086 11508 91138
rect 11340 91084 11508 91086
rect 11116 90578 11172 90590
rect 11116 90526 11118 90578
rect 11170 90526 11172 90578
rect 11116 90356 11172 90526
rect 11228 90580 11284 90590
rect 11340 90580 11396 91084
rect 11452 91074 11508 91084
rect 12012 91138 12068 91150
rect 12012 91086 12014 91138
rect 12066 91086 12068 91138
rect 11452 90804 11508 90814
rect 11452 90710 11508 90748
rect 11900 90690 11956 90702
rect 11900 90638 11902 90690
rect 11954 90638 11956 90690
rect 11284 90524 11396 90580
rect 11676 90580 11732 90590
rect 11900 90580 11956 90638
rect 11676 90578 11844 90580
rect 11676 90526 11678 90578
rect 11730 90526 11844 90578
rect 11676 90524 11844 90526
rect 11228 90514 11284 90524
rect 11676 90514 11732 90524
rect 11564 90466 11620 90478
rect 11564 90414 11566 90466
rect 11618 90414 11620 90466
rect 11564 90356 11620 90414
rect 11116 90300 11620 90356
rect 11418 90188 11682 90198
rect 11474 90132 11522 90188
rect 11578 90132 11626 90188
rect 11418 90122 11682 90132
rect 11788 89796 11844 90524
rect 11900 90514 11956 90524
rect 12012 90692 12068 91086
rect 12012 90468 12068 90636
rect 12012 89908 12068 90412
rect 12348 90466 12404 92316
rect 12348 90414 12350 90466
rect 12402 90414 12404 90466
rect 12348 90402 12404 90414
rect 12460 89908 12516 89918
rect 12012 89906 12516 89908
rect 12012 89854 12462 89906
rect 12514 89854 12516 89906
rect 12012 89852 12516 89854
rect 11788 89730 11844 89740
rect 11116 88900 11172 88910
rect 11004 88844 11116 88900
rect 11116 88834 11172 88844
rect 11418 88620 11682 88630
rect 11474 88564 11522 88620
rect 11578 88564 11626 88620
rect 11418 88554 11682 88564
rect 10780 88340 10836 88350
rect 10668 88338 10836 88340
rect 10668 88286 10782 88338
rect 10834 88286 10836 88338
rect 10668 88284 10836 88286
rect 10780 88274 10836 88284
rect 10108 88228 10164 88238
rect 9548 88226 9716 88228
rect 9548 88174 9550 88226
rect 9602 88174 9716 88226
rect 9548 88172 9716 88174
rect 9996 88226 10164 88228
rect 9996 88174 10110 88226
rect 10162 88174 10164 88226
rect 9996 88172 10164 88174
rect 9548 88162 9604 88172
rect 7756 88116 7812 88126
rect 7756 88022 7812 88060
rect 7980 88114 8036 88126
rect 7980 88062 7982 88114
rect 8034 88062 8036 88114
rect 7980 88004 8036 88062
rect 9212 88116 9268 88126
rect 9212 88022 9268 88060
rect 7980 87938 8036 87948
rect 8876 88004 8932 88014
rect 8988 88004 9044 88014
rect 8932 88002 9044 88004
rect 8932 87950 8990 88002
rect 9042 87950 9044 88002
rect 8932 87948 9044 87950
rect 8016 87836 8280 87846
rect 8072 87780 8120 87836
rect 8176 87780 8224 87836
rect 8016 87770 8280 87780
rect 7868 87332 7924 87342
rect 7868 86882 7924 87276
rect 8876 87108 8932 87948
rect 8988 87938 9044 87948
rect 9548 87444 9604 87454
rect 8988 87442 9604 87444
rect 8988 87390 9550 87442
rect 9602 87390 9604 87442
rect 8988 87388 9604 87390
rect 8988 87330 9044 87388
rect 9548 87378 9604 87388
rect 8988 87278 8990 87330
rect 9042 87278 9044 87330
rect 8988 87266 9044 87278
rect 9660 87332 9716 88172
rect 10108 88162 10164 88172
rect 12348 88116 12404 88126
rect 9660 87266 9716 87276
rect 10108 87332 10164 87342
rect 8876 87052 9156 87108
rect 7868 86830 7870 86882
rect 7922 86830 7924 86882
rect 7868 86770 7924 86830
rect 7868 86718 7870 86770
rect 7922 86718 7924 86770
rect 7868 86706 7924 86718
rect 8428 86772 8484 86782
rect 8988 86772 9044 86782
rect 8428 86770 8932 86772
rect 8428 86718 8430 86770
rect 8482 86718 8932 86770
rect 8428 86716 8932 86718
rect 8428 86706 8484 86716
rect 8652 86546 8708 86558
rect 8652 86494 8654 86546
rect 8706 86494 8708 86546
rect 8652 86436 8708 86494
rect 8428 86380 8652 86436
rect 8016 86268 8280 86278
rect 8072 86212 8120 86268
rect 8176 86212 8224 86268
rect 8016 86202 8280 86212
rect 8428 86100 8484 86380
rect 8652 86370 8708 86380
rect 8764 86434 8820 86446
rect 8764 86382 8766 86434
rect 8818 86382 8820 86434
rect 8092 86044 8484 86100
rect 8092 85986 8148 86044
rect 8092 85934 8094 85986
rect 8146 85934 8148 85986
rect 8092 85922 8148 85934
rect 8652 85988 8708 85998
rect 8652 85894 8708 85932
rect 7756 85876 7812 85886
rect 7756 85782 7812 85820
rect 8316 85874 8372 85886
rect 8316 85822 8318 85874
rect 8370 85822 8372 85874
rect 8204 85762 8260 85774
rect 8204 85710 8206 85762
rect 8258 85710 8260 85762
rect 8204 85708 8260 85710
rect 7868 85652 8260 85708
rect 8316 85764 8372 85822
rect 8316 85698 8372 85708
rect 7868 85650 7924 85652
rect 7868 85598 7870 85650
rect 7922 85598 7924 85650
rect 7868 85586 7924 85598
rect 8016 84700 8280 84710
rect 8072 84644 8120 84700
rect 8176 84644 8224 84700
rect 8016 84634 8280 84644
rect 8764 84084 8820 86382
rect 8876 85652 8932 86716
rect 8988 86658 9044 86716
rect 8988 86606 8990 86658
rect 9042 86606 9044 86658
rect 8988 86594 9044 86606
rect 8988 86436 9044 86446
rect 9100 86436 9156 87052
rect 10108 86772 10164 87276
rect 11418 87052 11682 87062
rect 11474 86996 11522 87052
rect 11578 86996 11626 87052
rect 11418 86986 11682 86996
rect 10108 86658 10164 86716
rect 10108 86606 10110 86658
rect 10162 86606 10164 86658
rect 10108 86594 10164 86606
rect 11228 86772 11284 86782
rect 9212 86548 9268 86558
rect 9212 86454 9268 86492
rect 10892 86548 10948 86558
rect 10892 86454 10948 86492
rect 11228 86546 11284 86716
rect 12236 86660 12292 86670
rect 12236 86566 12292 86604
rect 11228 86494 11230 86546
rect 11282 86494 11284 86546
rect 9044 86380 9156 86436
rect 9548 86436 9604 86446
rect 8988 86370 9044 86380
rect 9548 86342 9604 86380
rect 9660 86434 9716 86446
rect 9660 86382 9662 86434
rect 9714 86382 9716 86434
rect 9660 85988 9716 86382
rect 9660 85922 9716 85932
rect 9772 86434 9828 86446
rect 9772 86382 9774 86434
rect 9826 86382 9828 86434
rect 9772 86100 9828 86382
rect 9772 85708 9828 86044
rect 10780 86436 10836 86446
rect 10780 85986 10836 86380
rect 10780 85934 10782 85986
rect 10834 85934 10836 85986
rect 10780 85922 10836 85934
rect 11004 86434 11060 86446
rect 11004 86382 11006 86434
rect 11058 86382 11060 86434
rect 11004 85876 11060 86382
rect 11004 85810 11060 85820
rect 11228 85708 11284 86494
rect 9772 85652 10276 85708
rect 8876 84532 8932 85596
rect 9324 85202 9380 85214
rect 9324 85150 9326 85202
rect 9378 85150 9380 85202
rect 9324 85092 9380 85150
rect 9660 85092 9716 85102
rect 9324 85090 9716 85092
rect 9324 85038 9662 85090
rect 9714 85038 9716 85090
rect 9324 85036 9716 85038
rect 9660 85026 9716 85036
rect 8988 84532 9044 84542
rect 8876 84476 8988 84532
rect 8988 84438 9044 84476
rect 10220 84420 10276 85652
rect 10892 85652 11284 85708
rect 12012 86434 12068 86446
rect 12012 86382 12014 86434
rect 12066 86382 12068 86434
rect 12012 85652 12068 86382
rect 10220 84326 10276 84364
rect 10332 84532 10388 84542
rect 9884 84308 9940 84318
rect 9772 84196 9828 84206
rect 9884 84196 9940 84252
rect 9772 84194 9940 84196
rect 9772 84142 9774 84194
rect 9826 84142 9940 84194
rect 9772 84140 9940 84142
rect 9772 84130 9828 84140
rect 8764 84018 8820 84028
rect 7756 83746 7812 83758
rect 7756 83694 7758 83746
rect 7810 83694 7812 83746
rect 7756 83300 7812 83694
rect 9548 83524 9604 83534
rect 9884 83524 9940 84140
rect 9548 83522 9940 83524
rect 9548 83470 9550 83522
rect 9602 83470 9940 83522
rect 9548 83468 9940 83470
rect 9548 83458 9604 83468
rect 7756 83298 7924 83300
rect 7756 83246 7758 83298
rect 7810 83246 7924 83298
rect 7756 83244 7924 83246
rect 7756 83234 7812 83244
rect 7644 82684 7812 82740
rect 7644 82514 7700 82526
rect 7644 82462 7646 82514
rect 7698 82462 7700 82514
rect 7644 81844 7700 82462
rect 7756 81956 7812 82684
rect 7756 81890 7812 81900
rect 7644 81778 7700 81788
rect 7756 81170 7812 81182
rect 7756 81118 7758 81170
rect 7810 81118 7812 81170
rect 7756 81060 7812 81118
rect 7756 79828 7812 81004
rect 7868 80500 7924 83244
rect 8016 83132 8280 83142
rect 8072 83076 8120 83132
rect 8176 83076 8224 83132
rect 8016 83066 8280 83076
rect 9884 82962 9940 83468
rect 9884 82910 9886 82962
rect 9938 82910 9940 82962
rect 9884 82898 9940 82910
rect 10108 84084 10164 84094
rect 8092 82626 8148 82638
rect 8092 82574 8094 82626
rect 8146 82574 8148 82626
rect 8092 81844 8148 82574
rect 9324 82124 9716 82180
rect 9324 82066 9380 82124
rect 9324 82014 9326 82066
rect 9378 82014 9380 82066
rect 9324 82002 9380 82014
rect 9660 82066 9716 82124
rect 9660 82014 9662 82066
rect 9714 82014 9716 82066
rect 9660 82002 9716 82014
rect 8092 81778 8148 81788
rect 9548 81956 9604 81966
rect 8016 81564 8280 81574
rect 8072 81508 8120 81564
rect 8176 81508 8224 81564
rect 8016 81498 8280 81508
rect 7868 80434 7924 80444
rect 9436 81396 9492 81406
rect 9436 80386 9492 81340
rect 9436 80334 9438 80386
rect 9490 80334 9492 80386
rect 9436 80322 9492 80334
rect 8016 79996 8280 80006
rect 8072 79940 8120 79996
rect 8176 79940 8224 79996
rect 8016 79930 8280 79940
rect 7756 79772 8036 79828
rect 7308 79660 7588 79716
rect 6188 78820 6244 78830
rect 6188 78726 6244 78764
rect 6412 78706 6468 78718
rect 6412 78654 6414 78706
rect 6466 78654 6468 78706
rect 6412 78596 6468 78654
rect 6412 78258 6468 78540
rect 6860 78596 6916 78606
rect 6860 78502 6916 78540
rect 6412 78206 6414 78258
rect 6466 78206 6468 78258
rect 6412 78194 6468 78206
rect 5964 78082 6020 78092
rect 5628 77198 5630 77250
rect 5682 77198 5684 77250
rect 4060 77026 4116 77038
rect 4060 76974 4062 77026
rect 4114 76974 4116 77026
rect 4060 76468 4116 76974
rect 4732 77026 4788 77038
rect 4732 76974 4734 77026
rect 4786 76974 4788 77026
rect 4060 76402 4116 76412
rect 4620 76692 4676 76702
rect 4620 76356 4676 76636
rect 4396 76354 4676 76356
rect 4396 76302 4622 76354
rect 4674 76302 4676 76354
rect 4396 76300 4676 76302
rect 4396 75572 4452 76300
rect 4620 76290 4676 76300
rect 4732 76244 4788 76974
rect 5068 77026 5124 77038
rect 5068 76974 5070 77026
rect 5122 76974 5124 77026
rect 5068 76692 5124 76974
rect 5068 76636 5460 76692
rect 5068 76580 5124 76636
rect 5068 76514 5124 76524
rect 5292 76468 5348 76478
rect 5292 76374 5348 76412
rect 4732 76188 5012 76244
rect 4614 76076 4878 76086
rect 4670 76020 4718 76076
rect 4774 76020 4822 76076
rect 4614 76010 4878 76020
rect 4956 75908 5012 76188
rect 4620 75852 5124 75908
rect 4620 75794 4676 75852
rect 4620 75742 4622 75794
rect 4674 75742 4676 75794
rect 4620 75730 4676 75742
rect 4956 75684 5012 75694
rect 4956 75590 5012 75628
rect 5068 75682 5124 75852
rect 5068 75630 5070 75682
rect 5122 75630 5124 75682
rect 4396 75516 4900 75572
rect 4172 74788 4228 74798
rect 4172 74694 4228 74732
rect 4060 74340 4116 74350
rect 4060 73890 4116 74284
rect 4396 73948 4452 75516
rect 4844 75122 4900 75516
rect 4844 75070 4846 75122
rect 4898 75070 4900 75122
rect 4844 75058 4900 75070
rect 4614 74508 4878 74518
rect 4670 74452 4718 74508
rect 4774 74452 4822 74508
rect 4614 74442 4878 74452
rect 5068 73948 5124 75630
rect 5292 74788 5348 74798
rect 5292 74694 5348 74732
rect 5404 73948 5460 76636
rect 5516 76356 5572 76366
rect 5516 75012 5572 76300
rect 5628 75684 5684 77198
rect 6076 77922 6132 77934
rect 6076 77870 6078 77922
rect 6130 77870 6132 77922
rect 6076 76580 6132 77870
rect 6972 77924 7028 77934
rect 7308 77924 7364 79660
rect 7756 79604 7812 79614
rect 7420 79602 7812 79604
rect 7420 79550 7758 79602
rect 7810 79550 7812 79602
rect 7420 79548 7812 79550
rect 7420 79490 7476 79548
rect 7756 79538 7812 79548
rect 7420 79438 7422 79490
rect 7474 79438 7476 79490
rect 7420 79426 7476 79438
rect 7868 79378 7924 79390
rect 7868 79326 7870 79378
rect 7922 79326 7924 79378
rect 7868 78820 7924 79326
rect 7868 78754 7924 78764
rect 7868 78596 7924 78606
rect 7980 78596 8036 79772
rect 8316 79490 8372 79502
rect 9100 79492 9156 79502
rect 8316 79438 8318 79490
rect 8370 79438 8372 79490
rect 8316 78932 8372 79438
rect 8316 78866 8372 78876
rect 8988 79490 9156 79492
rect 8988 79438 9102 79490
rect 9154 79438 9156 79490
rect 8988 79436 9156 79438
rect 8428 78820 8484 78830
rect 8988 78820 9044 79436
rect 9100 79426 9156 79436
rect 8428 78818 9044 78820
rect 8428 78766 8430 78818
rect 8482 78766 9044 78818
rect 8428 78764 9044 78766
rect 8428 78754 8484 78764
rect 7924 78540 8036 78596
rect 7868 78502 7924 78540
rect 8764 78484 8820 78494
rect 8016 78428 8280 78438
rect 8072 78372 8120 78428
rect 8176 78372 8224 78428
rect 8016 78362 8280 78372
rect 7868 78036 7924 78046
rect 7868 77942 7924 77980
rect 8204 78034 8260 78046
rect 8204 77982 8206 78034
rect 8258 77982 8260 78034
rect 6972 77922 7364 77924
rect 6972 77870 6974 77922
rect 7026 77870 7364 77922
rect 6972 77868 7364 77870
rect 7420 77922 7476 77934
rect 7420 77870 7422 77922
rect 7474 77870 7476 77922
rect 6972 77700 7028 77868
rect 6972 77634 7028 77644
rect 7420 77810 7476 77870
rect 7420 77758 7422 77810
rect 7474 77758 7476 77810
rect 6412 77138 6468 77150
rect 6412 77086 6414 77138
rect 6466 77086 6468 77138
rect 6412 76692 6468 77086
rect 6636 76692 6692 76702
rect 7420 76692 7476 77758
rect 7980 77812 8036 77822
rect 8204 77812 8260 77982
rect 7980 77810 8260 77812
rect 7980 77758 7982 77810
rect 8034 77758 8260 77810
rect 7980 77756 8260 77758
rect 8540 78034 8596 78046
rect 8540 77982 8542 78034
rect 8594 77982 8596 78034
rect 7980 77746 8036 77756
rect 8540 77700 8596 77982
rect 8764 78034 8820 78428
rect 8764 77982 8766 78034
rect 8818 77982 8820 78034
rect 8764 77970 8820 77982
rect 8540 77634 8596 77644
rect 8764 77810 8820 77822
rect 8764 77758 8766 77810
rect 8818 77758 8820 77810
rect 8540 77364 8596 77374
rect 8428 77362 8596 77364
rect 8428 77310 8542 77362
rect 8594 77310 8596 77362
rect 8428 77308 8596 77310
rect 8016 76860 8280 76870
rect 8072 76804 8120 76860
rect 8176 76804 8224 76860
rect 8016 76794 8280 76804
rect 6412 76690 6692 76692
rect 6412 76638 6638 76690
rect 6690 76638 6692 76690
rect 6412 76636 6692 76638
rect 6636 76626 6692 76636
rect 7196 76636 7476 76692
rect 7084 76580 7140 76590
rect 6132 76524 6244 76580
rect 6076 76514 6132 76524
rect 5740 76356 5796 76366
rect 5740 76262 5796 76300
rect 5628 75682 5796 75684
rect 5628 75630 5630 75682
rect 5682 75630 5796 75682
rect 5628 75628 5796 75630
rect 5628 75618 5684 75628
rect 5628 75012 5684 75022
rect 5516 75010 5684 75012
rect 5516 74958 5630 75010
rect 5682 74958 5684 75010
rect 5516 74956 5684 74958
rect 4396 73892 4676 73948
rect 4060 73838 4062 73890
rect 4114 73838 4116 73890
rect 4060 73826 4116 73838
rect 4172 73218 4228 73230
rect 4620 73220 4676 73892
rect 4844 73892 4900 73902
rect 5068 73892 5348 73948
rect 5404 73892 5572 73948
rect 4844 73332 4900 73836
rect 4956 73332 5012 73342
rect 4844 73330 5012 73332
rect 4844 73278 4958 73330
rect 5010 73278 5012 73330
rect 4844 73276 5012 73278
rect 4172 73166 4174 73218
rect 4226 73166 4228 73218
rect 4172 72548 4228 73166
rect 4396 73218 4676 73220
rect 4396 73166 4622 73218
rect 4674 73166 4676 73218
rect 4396 73164 4676 73166
rect 4396 72772 4452 73164
rect 4620 73154 4676 73164
rect 4614 72940 4878 72950
rect 4670 72884 4718 72940
rect 4774 72884 4822 72940
rect 4614 72874 4878 72884
rect 4396 72716 4564 72772
rect 4396 72548 4452 72558
rect 4172 72492 4396 72548
rect 3948 72268 4340 72324
rect 4172 71876 4228 71886
rect 3948 71652 4004 71662
rect 3948 71202 4004 71596
rect 3948 71150 3950 71202
rect 4002 71150 4004 71202
rect 3948 71138 4004 71150
rect 3836 71026 3892 71036
rect 3948 70756 4004 70766
rect 3948 70662 4004 70700
rect 4172 70756 4228 71820
rect 3724 70532 4116 70588
rect 3500 68786 3556 68796
rect 3052 68738 3220 68740
rect 3052 68686 3054 68738
rect 3106 68686 3220 68738
rect 3052 68684 3220 68686
rect 3052 68674 3108 68684
rect 2492 68628 2548 68666
rect 2492 68562 2548 68572
rect 2828 68628 2884 68638
rect 2828 68534 2884 68572
rect 2492 68404 2548 68414
rect 2380 68402 2548 68404
rect 2380 68350 2494 68402
rect 2546 68350 2548 68402
rect 2380 68348 2548 68350
rect 2492 68338 2548 68348
rect 3164 67956 3220 68684
rect 3388 68628 3444 68638
rect 3388 68534 3444 68572
rect 3500 68514 3556 68526
rect 3500 68462 3502 68514
rect 3554 68462 3556 68514
rect 3500 68404 3556 68462
rect 3500 68338 3556 68348
rect 3948 68514 4004 68526
rect 3948 68462 3950 68514
rect 4002 68462 4004 68514
rect 3948 68404 4004 68462
rect 3948 68310 4004 68348
rect 3276 67956 3332 67966
rect 3164 67954 3332 67956
rect 3164 67902 3278 67954
rect 3330 67902 3332 67954
rect 3164 67900 3332 67902
rect 2716 67172 2772 67182
rect 2716 67060 2772 67116
rect 3052 67060 3108 67070
rect 2716 67058 3108 67060
rect 2716 67006 2718 67058
rect 2770 67006 3054 67058
rect 3106 67006 3108 67058
rect 2716 67004 3108 67006
rect 2716 66994 2772 67004
rect 3052 66994 3108 67004
rect 2380 66836 2436 66846
rect 2268 66780 2380 66836
rect 1708 66546 1764 66556
rect 1596 66332 1764 66388
rect 1708 66276 1764 66332
rect 1708 66274 1876 66276
rect 1708 66222 1710 66274
rect 1762 66222 1876 66274
rect 1708 66220 1876 66222
rect 1708 66210 1764 66220
rect 1708 64596 1764 64606
rect 1708 64502 1764 64540
rect 1820 64148 1876 66220
rect 1708 64092 1876 64148
rect 1932 64596 1988 64606
rect 1708 63138 1764 64092
rect 1820 63924 1876 63934
rect 1932 63924 1988 64540
rect 2268 64596 2324 64606
rect 2380 64596 2436 66780
rect 2716 66834 2772 66846
rect 2716 66782 2718 66834
rect 2770 66782 2772 66834
rect 2492 66162 2548 66174
rect 2492 66110 2494 66162
rect 2546 66110 2548 66162
rect 2492 65716 2548 66110
rect 2604 65716 2660 65726
rect 2492 65714 2660 65716
rect 2492 65662 2606 65714
rect 2658 65662 2660 65714
rect 2492 65660 2660 65662
rect 2604 65650 2660 65660
rect 2492 65492 2548 65502
rect 2492 64820 2548 65436
rect 2604 65492 2660 65502
rect 2716 65492 2772 66782
rect 3164 66834 3220 66846
rect 3164 66782 3166 66834
rect 3218 66782 3220 66834
rect 2828 65828 2884 65838
rect 2828 65602 2884 65772
rect 2828 65550 2830 65602
rect 2882 65550 2884 65602
rect 2828 65538 2884 65550
rect 3052 65604 3108 65614
rect 3052 65510 3108 65548
rect 2604 65490 2772 65492
rect 2604 65438 2606 65490
rect 2658 65438 2772 65490
rect 2604 65436 2772 65438
rect 2604 65426 2660 65436
rect 2492 64764 2660 64820
rect 2324 64540 2436 64596
rect 2044 64484 2100 64494
rect 2044 64390 2100 64428
rect 1876 63868 1988 63924
rect 1820 63830 1876 63868
rect 1708 63086 1710 63138
rect 1762 63086 1764 63138
rect 1708 62188 1764 63086
rect 2268 62188 2324 64540
rect 2492 64148 2548 64158
rect 2380 64146 2548 64148
rect 2380 64094 2494 64146
rect 2546 64094 2548 64146
rect 2380 64092 2548 64094
rect 2380 63252 2436 64092
rect 2492 64082 2548 64092
rect 2604 63924 2660 64764
rect 3052 64596 3108 64606
rect 3052 64502 3108 64540
rect 2828 64484 2884 64494
rect 2828 64390 2884 64428
rect 2940 64482 2996 64494
rect 2940 64430 2942 64482
rect 2994 64430 2996 64482
rect 2716 63924 2772 63934
rect 2604 63868 2716 63924
rect 2492 63252 2548 63262
rect 2380 63250 2548 63252
rect 2380 63198 2494 63250
rect 2546 63198 2548 63250
rect 2380 63196 2548 63198
rect 2492 63186 2548 63196
rect 1708 62132 1876 62188
rect 1708 61458 1764 61470
rect 1708 61406 1710 61458
rect 1762 61406 1764 61458
rect 1708 61236 1764 61406
rect 1708 61170 1764 61180
rect 1820 60002 1876 62132
rect 2156 62132 2324 62188
rect 2492 62242 2548 62254
rect 2492 62190 2494 62242
rect 2546 62190 2548 62242
rect 2044 61460 2100 61470
rect 2044 61366 2100 61404
rect 2044 61012 2100 61022
rect 2156 61012 2212 62132
rect 2044 61010 2212 61012
rect 2044 60958 2046 61010
rect 2098 60958 2212 61010
rect 2044 60956 2212 60958
rect 2044 60946 2100 60956
rect 2156 60676 2212 60956
rect 2380 61348 2436 61358
rect 2380 60786 2436 61292
rect 2492 61236 2548 62190
rect 2716 61348 2772 63868
rect 2828 63924 2884 63934
rect 2940 63924 2996 64430
rect 2828 63922 2996 63924
rect 2828 63870 2830 63922
rect 2882 63870 2996 63922
rect 2828 63868 2996 63870
rect 3052 63922 3108 63934
rect 3052 63870 3054 63922
rect 3106 63870 3108 63922
rect 2828 63858 2884 63868
rect 3052 63812 3108 63870
rect 3052 63746 3108 63756
rect 3164 63028 3220 66782
rect 3276 65604 3332 67900
rect 3836 66948 3892 66958
rect 3836 66854 3892 66892
rect 3500 65828 3556 65838
rect 3388 65716 3444 65726
rect 3500 65716 3556 65772
rect 3388 65714 3556 65716
rect 3388 65662 3390 65714
rect 3442 65662 3556 65714
rect 3388 65660 3556 65662
rect 3388 65650 3444 65660
rect 3276 65538 3332 65548
rect 3500 65380 3556 65390
rect 3836 65380 3892 65390
rect 3500 65378 3836 65380
rect 3500 65326 3502 65378
rect 3554 65326 3836 65378
rect 3500 65324 3836 65326
rect 3500 65314 3556 65324
rect 3724 64930 3780 64942
rect 3724 64878 3726 64930
rect 3778 64878 3780 64930
rect 3724 64482 3780 64878
rect 3724 64430 3726 64482
rect 3778 64430 3780 64482
rect 3164 62962 3220 62972
rect 3276 64148 3332 64158
rect 3276 64034 3332 64092
rect 3276 63982 3278 64034
rect 3330 63982 3332 64034
rect 3276 62804 3332 63982
rect 3724 63924 3780 64430
rect 3724 63858 3780 63868
rect 2828 62748 3332 62804
rect 3500 63812 3556 63822
rect 2828 61684 2884 62748
rect 3500 62578 3556 63756
rect 3500 62526 3502 62578
rect 3554 62526 3556 62578
rect 3500 62514 3556 62526
rect 3724 63252 3780 63262
rect 3612 62468 3668 62478
rect 3724 62468 3780 63196
rect 3612 62466 3780 62468
rect 3612 62414 3614 62466
rect 3666 62414 3780 62466
rect 3612 62412 3780 62414
rect 3612 62402 3668 62412
rect 3500 61796 3556 61806
rect 2828 61682 3108 61684
rect 2828 61630 2830 61682
rect 2882 61630 3108 61682
rect 2828 61628 3108 61630
rect 2828 61618 2884 61628
rect 2716 61282 2772 61292
rect 2492 61170 2548 61180
rect 2604 61012 2660 61022
rect 2380 60734 2382 60786
rect 2434 60734 2436 60786
rect 2212 60620 2324 60676
rect 2156 60610 2212 60620
rect 1820 59950 1822 60002
rect 1874 59950 1876 60002
rect 1708 59218 1764 59230
rect 1708 59166 1710 59218
rect 1762 59166 1764 59218
rect 1708 58548 1764 59166
rect 1708 58482 1764 58492
rect 1820 57876 1876 59950
rect 2044 59330 2100 59342
rect 2044 59278 2046 59330
rect 2098 59278 2100 59330
rect 2044 58436 2100 59278
rect 2044 58370 2100 58380
rect 2268 58212 2324 60620
rect 2380 58660 2436 60734
rect 2492 61010 2660 61012
rect 2492 60958 2606 61010
rect 2658 60958 2660 61010
rect 2492 60956 2660 60958
rect 2492 60114 2548 60956
rect 2604 60946 2660 60956
rect 3052 60900 3108 61628
rect 3500 61682 3556 61740
rect 3500 61630 3502 61682
rect 3554 61630 3556 61682
rect 3500 61618 3556 61630
rect 3276 61570 3332 61582
rect 3276 61518 3278 61570
rect 3330 61518 3332 61570
rect 3276 61460 3332 61518
rect 3052 60898 3220 60900
rect 3052 60846 3054 60898
rect 3106 60846 3220 60898
rect 3052 60844 3220 60846
rect 3052 60834 3108 60844
rect 2828 60788 2884 60798
rect 2828 60786 2996 60788
rect 2828 60734 2830 60786
rect 2882 60734 2996 60786
rect 2828 60732 2996 60734
rect 2828 60722 2884 60732
rect 2604 60564 2660 60574
rect 2604 60470 2660 60508
rect 2492 60062 2494 60114
rect 2546 60062 2548 60114
rect 2492 60050 2548 60062
rect 2940 59444 2996 60732
rect 3164 60116 3220 60844
rect 3276 60788 3332 61404
rect 3724 60900 3780 62412
rect 3836 61012 3892 65324
rect 3948 65378 4004 65390
rect 3948 65326 3950 65378
rect 4002 65326 4004 65378
rect 3948 64930 4004 65326
rect 3948 64878 3950 64930
rect 4002 64878 4004 64930
rect 3948 64866 4004 64878
rect 3948 64484 4004 64494
rect 3948 63922 4004 64428
rect 3948 63870 3950 63922
rect 4002 63870 4004 63922
rect 3948 63858 4004 63870
rect 4060 61124 4116 70532
rect 4172 68404 4228 70700
rect 4172 68338 4228 68348
rect 4284 65268 4340 72268
rect 4396 71762 4452 72492
rect 4508 71876 4564 72716
rect 4508 71810 4564 71820
rect 4620 72658 4676 72670
rect 4620 72606 4622 72658
rect 4674 72606 4676 72658
rect 4396 71710 4398 71762
rect 4450 71710 4452 71762
rect 4396 70084 4452 71710
rect 4508 71652 4564 71662
rect 4620 71652 4676 72606
rect 4956 72548 5012 73276
rect 4956 72482 5012 72492
rect 5068 72436 5124 72446
rect 5068 72342 5124 72380
rect 5068 71764 5124 71774
rect 5068 71762 5236 71764
rect 5068 71710 5070 71762
rect 5122 71710 5236 71762
rect 5068 71708 5236 71710
rect 5068 71698 5124 71708
rect 4564 71596 4676 71652
rect 5180 71652 5236 71708
rect 4508 71586 4564 71596
rect 5180 71586 5236 71596
rect 4614 71372 4878 71382
rect 4670 71316 4718 71372
rect 4774 71316 4822 71372
rect 4614 71306 4878 71316
rect 4620 70866 4676 70878
rect 4620 70814 4622 70866
rect 4674 70814 4676 70866
rect 4508 70756 4564 70766
rect 4620 70756 4676 70814
rect 4564 70700 4676 70756
rect 5180 70754 5236 70766
rect 5180 70702 5182 70754
rect 5234 70702 5236 70754
rect 4508 70690 4564 70700
rect 5068 70644 5124 70654
rect 5068 70308 5124 70588
rect 5180 70532 5236 70702
rect 5180 70466 5236 70476
rect 5068 70252 5236 70308
rect 5068 70084 5124 70094
rect 4396 70082 5124 70084
rect 4396 70030 5070 70082
rect 5122 70030 5124 70082
rect 4396 70028 5124 70030
rect 4614 69804 4878 69814
rect 4670 69748 4718 69804
rect 4774 69748 4822 69804
rect 4614 69738 4878 69748
rect 4620 69524 4676 69534
rect 4508 69522 4676 69524
rect 4508 69470 4622 69522
rect 4674 69470 4676 69522
rect 4508 69468 4676 69470
rect 4396 68516 4452 68526
rect 4396 68422 4452 68460
rect 4508 68402 4564 69468
rect 4620 69458 4676 69468
rect 5068 69188 5124 70028
rect 4956 69186 5124 69188
rect 4956 69134 5070 69186
rect 5122 69134 5124 69186
rect 4956 69132 5124 69134
rect 4844 68628 4900 68638
rect 4956 68628 5012 69132
rect 5068 69122 5124 69132
rect 5180 68964 5236 70252
rect 4844 68626 5012 68628
rect 4844 68574 4846 68626
rect 4898 68574 5012 68626
rect 4844 68572 5012 68574
rect 4844 68562 4900 68572
rect 4508 68350 4510 68402
rect 4562 68350 4564 68402
rect 4508 68338 4564 68350
rect 4614 68236 4878 68246
rect 4670 68180 4718 68236
rect 4774 68180 4822 68236
rect 4614 68170 4878 68180
rect 4956 67956 5012 68572
rect 4732 67060 4788 67070
rect 4956 67060 5012 67900
rect 4788 67004 5012 67060
rect 4732 66966 4788 67004
rect 4614 66668 4878 66678
rect 4670 66612 4718 66668
rect 4774 66612 4822 66668
rect 4614 66602 4878 66612
rect 4620 66386 4676 66398
rect 4620 66334 4622 66386
rect 4674 66334 4676 66386
rect 4396 65604 4452 65614
rect 4396 65510 4452 65548
rect 4620 65380 4676 66334
rect 4620 65314 4676 65324
rect 4844 65380 4900 65390
rect 4956 65380 5012 67004
rect 4844 65378 5012 65380
rect 4844 65326 4846 65378
rect 4898 65326 5012 65378
rect 4844 65324 5012 65326
rect 4844 65314 4900 65324
rect 4284 65202 4340 65212
rect 4614 65100 4878 65110
rect 4670 65044 4718 65100
rect 4774 65044 4822 65100
rect 4614 65034 4878 65044
rect 4284 64820 4340 64830
rect 4172 64708 4228 64718
rect 4172 64148 4228 64652
rect 4172 64082 4228 64092
rect 4172 61348 4228 61358
rect 4172 61254 4228 61292
rect 4060 61068 4228 61124
rect 3836 60956 4116 61012
rect 3724 60844 4004 60900
rect 3388 60788 3444 60798
rect 3276 60786 3444 60788
rect 3276 60734 3390 60786
rect 3442 60734 3444 60786
rect 3276 60732 3444 60734
rect 3388 60722 3444 60732
rect 3724 60676 3780 60686
rect 3724 60582 3780 60620
rect 3388 60564 3444 60574
rect 3388 60470 3444 60508
rect 3836 60564 3892 60574
rect 3164 60060 3444 60116
rect 3276 59892 3332 59902
rect 3164 59444 3220 59454
rect 2940 59442 3220 59444
rect 2940 59390 3166 59442
rect 3218 59390 3220 59442
rect 2940 59388 3220 59390
rect 3164 59378 3220 59388
rect 3276 59330 3332 59836
rect 3276 59278 3278 59330
rect 3330 59278 3332 59330
rect 3276 59266 3332 59278
rect 2380 58594 2436 58604
rect 2492 59106 2548 59118
rect 2492 59054 2494 59106
rect 2546 59054 2548 59106
rect 2492 58548 2548 59054
rect 3388 58828 3444 60060
rect 3724 59106 3780 59118
rect 3724 59054 3726 59106
rect 3778 59054 3780 59106
rect 3724 58828 3780 59054
rect 3388 58772 3780 58828
rect 2940 58660 2996 58670
rect 2940 58566 2996 58604
rect 2492 58482 2548 58492
rect 2828 58548 2884 58558
rect 2828 58434 2884 58492
rect 2828 58382 2830 58434
rect 2882 58382 2884 58434
rect 2828 58370 2884 58382
rect 3164 58322 3220 58334
rect 3164 58270 3166 58322
rect 3218 58270 3220 58322
rect 2604 58212 2660 58222
rect 2268 58118 2324 58156
rect 2492 58210 2660 58212
rect 2492 58158 2606 58210
rect 2658 58158 2660 58210
rect 2492 58156 2660 58158
rect 1820 57650 1876 57820
rect 2492 57762 2548 58156
rect 2604 58146 2660 58156
rect 2492 57710 2494 57762
rect 2546 57710 2548 57762
rect 2492 57698 2548 57710
rect 1820 57598 1822 57650
rect 1874 57598 1876 57650
rect 1820 57586 1876 57598
rect 3164 57092 3220 58270
rect 3388 58324 3444 58334
rect 3612 58324 3668 58772
rect 3724 58660 3780 58670
rect 3724 58566 3780 58604
rect 3836 58436 3892 60508
rect 3388 58322 3668 58324
rect 3388 58270 3390 58322
rect 3442 58270 3668 58322
rect 3388 58268 3668 58270
rect 3388 58258 3444 58268
rect 3612 57316 3668 58268
rect 3612 57250 3668 57260
rect 3724 58380 3892 58436
rect 3164 57026 3220 57036
rect 3500 57092 3556 57102
rect 3500 56998 3556 57036
rect 3612 56756 3668 56766
rect 3612 56662 3668 56700
rect 3500 56644 3556 56654
rect 3388 56420 3444 56430
rect 2044 56196 2100 56206
rect 2044 56194 2436 56196
rect 2044 56142 2046 56194
rect 2098 56142 2436 56194
rect 2044 56140 2436 56142
rect 2044 56130 2100 56140
rect 1708 56082 1764 56094
rect 1708 56030 1710 56082
rect 1762 56030 1764 56082
rect 1708 55860 1764 56030
rect 1708 55794 1764 55804
rect 1820 55298 1876 55310
rect 1820 55246 1822 55298
rect 1874 55246 1876 55298
rect 1820 53732 1876 55246
rect 2156 54516 2212 54526
rect 2156 54422 2212 54460
rect 2380 53732 2436 56140
rect 2492 55970 2548 55982
rect 2492 55918 2494 55970
rect 2546 55918 2548 55970
rect 2492 55860 2548 55918
rect 2492 55794 2548 55804
rect 2492 55186 2548 55198
rect 2492 55134 2494 55186
rect 2546 55134 2548 55186
rect 2492 55076 2548 55134
rect 2492 55020 2996 55076
rect 2940 54738 2996 55020
rect 2940 54686 2942 54738
rect 2994 54686 2996 54738
rect 2940 54674 2996 54686
rect 2604 54628 2660 54638
rect 2828 54628 2884 54638
rect 2604 54626 2828 54628
rect 2604 54574 2606 54626
rect 2658 54574 2828 54626
rect 2604 54572 2828 54574
rect 2604 54562 2660 54572
rect 2828 54534 2884 54572
rect 3052 54628 3108 54638
rect 3052 54626 3332 54628
rect 3052 54574 3054 54626
rect 3106 54574 3332 54626
rect 3052 54572 3332 54574
rect 3052 54562 3108 54572
rect 3276 54516 3332 54572
rect 3276 54450 3332 54460
rect 3388 54514 3444 56364
rect 3500 54628 3556 56588
rect 3612 56196 3668 56206
rect 3612 56102 3668 56140
rect 3724 54740 3780 58380
rect 3836 58212 3892 58222
rect 3836 58118 3892 58156
rect 3836 56196 3892 56206
rect 3948 56196 4004 60844
rect 4060 58548 4116 60956
rect 4172 58772 4228 61068
rect 4172 58706 4228 58716
rect 4060 58492 4228 58548
rect 4060 58324 4116 58334
rect 4060 58230 4116 58268
rect 4060 56756 4116 56766
rect 4060 56662 4116 56700
rect 4172 56308 4228 58492
rect 4284 56532 4340 64764
rect 4620 64596 4676 64606
rect 4620 64502 4676 64540
rect 4508 63924 4564 63934
rect 4508 63830 4564 63868
rect 4614 63532 4878 63542
rect 4670 63476 4718 63532
rect 4774 63476 4822 63532
rect 4614 63466 4878 63476
rect 4620 63252 4676 63262
rect 4956 63252 5012 65324
rect 5068 68908 5236 68964
rect 5068 63476 5124 68908
rect 5180 67732 5236 67742
rect 5180 67638 5236 67676
rect 5180 66164 5236 66174
rect 5180 66070 5236 66108
rect 5068 63410 5124 63420
rect 5180 63924 5236 63934
rect 5068 63252 5124 63262
rect 4956 63250 5124 63252
rect 4956 63198 5070 63250
rect 5122 63198 5124 63250
rect 4956 63196 5124 63198
rect 4620 63158 4676 63196
rect 5068 63186 5124 63196
rect 4956 62916 5012 62926
rect 4614 61964 4878 61974
rect 4670 61908 4718 61964
rect 4774 61908 4822 61964
rect 4614 61898 4878 61908
rect 4620 61684 4676 61694
rect 4620 61590 4676 61628
rect 4396 60786 4452 60798
rect 4396 60734 4398 60786
rect 4450 60734 4452 60786
rect 4396 60564 4452 60734
rect 4396 60498 4452 60508
rect 4614 60396 4878 60406
rect 4670 60340 4718 60396
rect 4774 60340 4822 60396
rect 4614 60330 4878 60340
rect 4620 60114 4676 60126
rect 4620 60062 4622 60114
rect 4674 60062 4676 60114
rect 4620 59892 4676 60062
rect 4620 58996 4676 59836
rect 4620 58930 4676 58940
rect 4614 58828 4878 58838
rect 4670 58772 4718 58828
rect 4774 58772 4822 58828
rect 4614 58762 4878 58772
rect 4620 58548 4676 58558
rect 4620 58454 4676 58492
rect 4620 57538 4676 57550
rect 4620 57486 4622 57538
rect 4674 57486 4676 57538
rect 4620 57428 4676 57486
rect 4396 57372 4676 57428
rect 4396 56756 4452 57372
rect 4614 57260 4878 57270
rect 4670 57204 4718 57260
rect 4774 57204 4822 57260
rect 4614 57194 4878 57204
rect 4396 56690 4452 56700
rect 4620 56868 4676 56878
rect 4284 56466 4340 56476
rect 4172 56252 4340 56308
rect 3948 56140 4116 56196
rect 3836 56102 3892 56140
rect 3948 55970 4004 55982
rect 3948 55918 3950 55970
rect 4002 55918 4004 55970
rect 3724 54674 3780 54684
rect 3836 55636 3892 55646
rect 3500 54562 3556 54572
rect 3388 54462 3390 54514
rect 3442 54462 3444 54514
rect 3276 54292 3332 54302
rect 3276 54198 3332 54236
rect 3388 53844 3444 54462
rect 3836 53956 3892 55580
rect 3948 54292 4004 55918
rect 3948 54226 4004 54236
rect 3276 53842 3444 53844
rect 3276 53790 3390 53842
rect 3442 53790 3444 53842
rect 3276 53788 3444 53790
rect 2492 53732 2548 53742
rect 2380 53730 2548 53732
rect 2380 53678 2494 53730
rect 2546 53678 2548 53730
rect 2380 53676 2548 53678
rect 1708 53620 1764 53630
rect 1708 53526 1764 53564
rect 1820 50594 1876 53676
rect 1820 50542 1822 50594
rect 1874 50542 1876 50594
rect 1708 50484 1764 50494
rect 1708 49810 1764 50428
rect 1708 49758 1710 49810
rect 1762 49758 1764 49810
rect 1708 47572 1764 49758
rect 1820 49700 1876 50542
rect 1820 49364 1876 49644
rect 1820 49298 1876 49308
rect 1932 53620 1988 53630
rect 1932 53172 1988 53564
rect 2044 53508 2100 53518
rect 2044 53506 2436 53508
rect 2044 53454 2046 53506
rect 2098 53454 2436 53506
rect 2044 53452 2436 53454
rect 2044 53442 2100 53452
rect 1820 49140 1876 49150
rect 1932 49140 1988 53116
rect 2380 52948 2436 53452
rect 2492 53170 2548 53676
rect 2828 53620 2884 53630
rect 2828 53618 2996 53620
rect 2828 53566 2830 53618
rect 2882 53566 2996 53618
rect 2828 53564 2996 53566
rect 2828 53554 2884 53564
rect 2940 53508 2996 53564
rect 2492 53118 2494 53170
rect 2546 53118 2548 53170
rect 2492 53106 2548 53118
rect 2828 53172 2884 53182
rect 2380 52892 2548 52948
rect 2156 52836 2212 52846
rect 2156 52742 2212 52780
rect 2492 52162 2548 52892
rect 2492 52110 2494 52162
rect 2546 52110 2548 52162
rect 2268 52052 2324 52062
rect 2268 51958 2324 51996
rect 2492 51602 2548 52110
rect 2492 51550 2494 51602
rect 2546 51550 2548 51602
rect 2492 51538 2548 51550
rect 2604 52834 2660 52846
rect 2604 52782 2606 52834
rect 2658 52782 2660 52834
rect 2604 51380 2660 52782
rect 2268 51324 2660 51380
rect 2716 52724 2772 52734
rect 2044 51266 2100 51278
rect 2044 51214 2046 51266
rect 2098 51214 2100 51266
rect 2044 51156 2100 51214
rect 2044 51090 2100 51100
rect 2156 50148 2212 50158
rect 2044 49924 2100 49934
rect 2044 49830 2100 49868
rect 1820 49138 1988 49140
rect 1820 49086 1822 49138
rect 1874 49086 1988 49138
rect 1820 49084 1988 49086
rect 1820 49074 1876 49084
rect 1708 47506 1764 47516
rect 1820 48916 1876 48926
rect 1820 48242 1876 48860
rect 1820 48190 1822 48242
rect 1874 48190 1876 48242
rect 1708 47348 1764 47358
rect 1708 47254 1764 47292
rect 1820 46900 1876 48190
rect 2156 47460 2212 50092
rect 2044 47236 2100 47246
rect 2044 47142 2100 47180
rect 1708 46674 1764 46686
rect 1708 46622 1710 46674
rect 1762 46622 1764 46674
rect 1708 45108 1764 46622
rect 1820 45890 1876 46844
rect 2044 46788 2100 46798
rect 1820 45838 1822 45890
rect 1874 45838 1876 45890
rect 1820 45826 1876 45838
rect 1932 46786 2100 46788
rect 1932 46734 2046 46786
rect 2098 46734 2100 46786
rect 1932 46732 2100 46734
rect 1708 43764 1764 45052
rect 1932 44884 1988 46732
rect 2044 46722 2100 46732
rect 2156 46564 2212 47404
rect 1932 44818 1988 44828
rect 2044 46508 2212 46564
rect 2044 44994 2100 46508
rect 2268 46004 2324 51324
rect 2156 45948 2324 46004
rect 2380 51154 2436 51166
rect 2380 51102 2382 51154
rect 2434 51102 2436 51154
rect 2156 45556 2212 45948
rect 2380 45780 2436 51102
rect 2716 51156 2772 52668
rect 2828 52276 2884 53116
rect 2828 52182 2884 52220
rect 2716 51062 2772 51100
rect 2492 50484 2548 50494
rect 2492 50390 2548 50428
rect 2940 50148 2996 53452
rect 3276 53170 3332 53788
rect 3388 53778 3444 53788
rect 3724 53900 3892 53956
rect 4060 53956 4116 56140
rect 4172 56084 4228 56094
rect 4172 55990 4228 56028
rect 4284 55860 4340 56252
rect 4620 56082 4676 56812
rect 4956 56308 5012 62860
rect 5180 62132 5236 63868
rect 5292 62188 5348 73892
rect 5516 70196 5572 73892
rect 5628 73668 5684 74956
rect 5740 74226 5796 75628
rect 5964 74898 6020 74910
rect 5964 74846 5966 74898
rect 6018 74846 6020 74898
rect 5964 74788 6020 74846
rect 6076 74900 6132 74910
rect 6076 74806 6132 74844
rect 6188 74898 6244 76524
rect 6524 76466 6580 76478
rect 6524 76414 6526 76466
rect 6578 76414 6580 76466
rect 6300 76354 6356 76366
rect 6300 76302 6302 76354
rect 6354 76302 6356 76354
rect 6300 76244 6356 76302
rect 6524 76356 6580 76414
rect 6524 76290 6580 76300
rect 6860 76468 6916 76478
rect 6300 76178 6356 76188
rect 6860 75908 6916 76412
rect 7084 76466 7140 76524
rect 7084 76414 7086 76466
rect 7138 76414 7140 76466
rect 7084 76402 7140 76414
rect 7084 76242 7140 76254
rect 7084 76190 7086 76242
rect 7138 76190 7140 76242
rect 7084 76132 7140 76190
rect 7196 76132 7252 76636
rect 7980 76468 8036 76478
rect 8428 76468 8484 77308
rect 8540 77298 8596 77308
rect 8764 76692 8820 77758
rect 8764 76626 8820 76636
rect 7980 76466 8484 76468
rect 7980 76414 7982 76466
rect 8034 76414 8484 76466
rect 7980 76412 8484 76414
rect 7980 76402 8036 76412
rect 7756 76354 7812 76366
rect 7756 76302 7758 76354
rect 7810 76302 7812 76354
rect 7644 76244 7700 76254
rect 7196 76076 7364 76132
rect 7084 76066 7140 76076
rect 6860 75842 6916 75852
rect 6412 75570 6468 75582
rect 6412 75518 6414 75570
rect 6466 75518 6468 75570
rect 6412 75122 6468 75518
rect 6412 75070 6414 75122
rect 6466 75070 6468 75122
rect 6412 75058 6468 75070
rect 6972 75460 7028 75470
rect 6972 75122 7028 75404
rect 6972 75070 6974 75122
rect 7026 75070 7028 75122
rect 6972 75058 7028 75070
rect 6188 74846 6190 74898
rect 6242 74846 6244 74898
rect 6188 74834 6244 74846
rect 6860 74900 6916 74910
rect 6860 74806 6916 74844
rect 5964 74340 6020 74732
rect 6748 74676 6804 74686
rect 6748 74674 6916 74676
rect 6748 74622 6750 74674
rect 6802 74622 6916 74674
rect 6748 74620 6916 74622
rect 6748 74610 6804 74620
rect 5964 74274 6020 74284
rect 5740 74174 5742 74226
rect 5794 74174 5796 74226
rect 5740 73892 5796 74174
rect 6524 74004 6580 74014
rect 6580 73948 6692 74004
rect 6524 73938 6580 73948
rect 5740 73826 5796 73836
rect 6636 73892 6692 73948
rect 6748 73892 6804 73902
rect 6636 73890 6804 73892
rect 6636 73838 6750 73890
rect 6802 73838 6804 73890
rect 6636 73836 6804 73838
rect 6636 73668 6692 73836
rect 6748 73826 6804 73836
rect 5628 73612 6692 73668
rect 5628 72436 5684 73612
rect 5740 73220 5796 73230
rect 5740 73218 5908 73220
rect 5740 73166 5742 73218
rect 5794 73166 5908 73218
rect 5740 73164 5908 73166
rect 5740 73154 5796 73164
rect 5852 72658 5908 73164
rect 5852 72606 5854 72658
rect 5906 72606 5908 72658
rect 5852 72594 5908 72606
rect 6188 72660 6244 72670
rect 6188 72566 6244 72604
rect 6076 72546 6132 72558
rect 6076 72494 6078 72546
rect 6130 72494 6132 72546
rect 5740 72436 5796 72446
rect 5628 72434 5796 72436
rect 5628 72382 5742 72434
rect 5794 72382 5796 72434
rect 5628 72380 5796 72382
rect 5628 70866 5684 72380
rect 5740 72370 5796 72380
rect 6076 72436 6132 72494
rect 6076 72370 6132 72380
rect 6300 72546 6356 72558
rect 6300 72494 6302 72546
rect 6354 72494 6356 72546
rect 5740 71652 5796 71662
rect 5740 71090 5796 71596
rect 5740 71038 5742 71090
rect 5794 71038 5796 71090
rect 5740 71026 5796 71038
rect 6076 70980 6132 70990
rect 6076 70886 6132 70924
rect 6188 70980 6244 70990
rect 6300 70980 6356 72494
rect 6188 70978 6356 70980
rect 6188 70926 6190 70978
rect 6242 70926 6356 70978
rect 6188 70924 6356 70926
rect 6636 72436 6692 72446
rect 6860 72436 6916 74620
rect 7196 74004 7252 74042
rect 7196 73938 7252 73948
rect 7196 72772 7252 72782
rect 6972 72660 7028 72670
rect 6972 72566 7028 72604
rect 7196 72546 7252 72716
rect 7196 72494 7198 72546
rect 7250 72494 7252 72546
rect 7196 72482 7252 72494
rect 5628 70814 5630 70866
rect 5682 70814 5684 70866
rect 5628 70644 5684 70814
rect 5628 70578 5684 70588
rect 5852 70866 5908 70878
rect 5852 70814 5854 70866
rect 5906 70814 5908 70866
rect 5516 70130 5572 70140
rect 5852 70532 5908 70814
rect 5964 70756 6020 70766
rect 6188 70756 6244 70924
rect 6020 70700 6244 70756
rect 5964 70690 6020 70700
rect 5852 68964 5908 70476
rect 5852 68908 6244 68964
rect 5516 68516 5572 68526
rect 5516 68514 6132 68516
rect 5516 68462 5518 68514
rect 5570 68462 6132 68514
rect 5516 68460 6132 68462
rect 5516 68450 5572 68460
rect 6076 67954 6132 68460
rect 6076 67902 6078 67954
rect 6130 67902 6132 67954
rect 6076 67890 6132 67902
rect 5964 67730 6020 67742
rect 5964 67678 5966 67730
rect 6018 67678 6020 67730
rect 5964 67620 6020 67678
rect 5964 67554 6020 67564
rect 5404 66946 5460 66958
rect 5404 66894 5406 66946
rect 5458 66894 5460 66946
rect 5404 66500 5460 66894
rect 5404 66444 6020 66500
rect 5964 66386 6020 66444
rect 5964 66334 5966 66386
rect 6018 66334 6020 66386
rect 5964 66322 6020 66334
rect 6076 66274 6132 66286
rect 6076 66222 6078 66274
rect 6130 66222 6132 66274
rect 5852 66162 5908 66174
rect 5852 66110 5854 66162
rect 5906 66110 5908 66162
rect 5852 66052 5908 66110
rect 5852 65986 5908 65996
rect 6076 66164 6132 66222
rect 5740 64820 5796 64830
rect 5740 64706 5796 64764
rect 5740 64654 5742 64706
rect 5794 64654 5796 64706
rect 5740 64642 5796 64654
rect 6076 64484 6132 66108
rect 6076 64418 6132 64428
rect 6188 64036 6244 68908
rect 6300 67732 6356 67742
rect 6300 67638 6356 67676
rect 6524 67730 6580 67742
rect 6524 67678 6526 67730
rect 6578 67678 6580 67730
rect 6412 66948 6468 66958
rect 6412 66274 6468 66892
rect 6412 66222 6414 66274
rect 6466 66222 6468 66274
rect 6412 66210 6468 66222
rect 6524 65716 6580 67678
rect 6524 65650 6580 65660
rect 6636 65492 6692 72380
rect 6748 72434 6916 72436
rect 6748 72382 6862 72434
rect 6914 72382 6916 72434
rect 6748 72380 6916 72382
rect 6748 70868 6804 72380
rect 6860 72370 6916 72380
rect 7308 71876 7364 76076
rect 6972 71820 7364 71876
rect 7532 75124 7588 75134
rect 7644 75124 7700 76188
rect 7756 76132 7812 76302
rect 7756 76066 7812 76076
rect 8016 75292 8280 75302
rect 8072 75236 8120 75292
rect 8176 75236 8224 75292
rect 8016 75226 8280 75236
rect 7532 75122 7700 75124
rect 7532 75070 7534 75122
rect 7586 75070 7700 75122
rect 7532 75068 7700 75070
rect 7980 75124 8036 75134
rect 8428 75124 8484 76412
rect 8540 76356 8596 76366
rect 8540 76262 8596 76300
rect 8540 75794 8596 75806
rect 8540 75742 8542 75794
rect 8594 75742 8596 75794
rect 8540 75460 8596 75742
rect 8876 75684 8932 78764
rect 9100 78706 9156 78718
rect 9100 78654 9102 78706
rect 9154 78654 9156 78706
rect 8988 78260 9044 78270
rect 9100 78260 9156 78654
rect 8988 78258 9156 78260
rect 8988 78206 8990 78258
rect 9042 78206 9156 78258
rect 8988 78204 9156 78206
rect 8988 78194 9044 78204
rect 9324 77026 9380 77038
rect 9324 76974 9326 77026
rect 9378 76974 9380 77026
rect 9324 76468 9380 76974
rect 9548 76916 9604 81900
rect 9772 81730 9828 81742
rect 9772 81678 9774 81730
rect 9826 81678 9828 81730
rect 9772 81172 9828 81678
rect 9772 80276 9828 81116
rect 10108 80498 10164 84028
rect 10220 83410 10276 83422
rect 10220 83358 10222 83410
rect 10274 83358 10276 83410
rect 10220 83076 10276 83358
rect 10220 83010 10276 83020
rect 10332 82964 10388 84476
rect 10668 84308 10724 84318
rect 10668 84214 10724 84252
rect 10332 82870 10388 82908
rect 10780 82964 10836 82974
rect 10780 82870 10836 82908
rect 10220 82178 10276 82190
rect 10220 82126 10222 82178
rect 10274 82126 10276 82178
rect 10220 82066 10276 82126
rect 10220 82014 10222 82066
rect 10274 82014 10276 82066
rect 10220 82002 10276 82014
rect 10668 81730 10724 81742
rect 10668 81678 10670 81730
rect 10722 81678 10724 81730
rect 10668 81620 10724 81678
rect 10668 81554 10724 81564
rect 10780 81732 10836 81742
rect 10220 81396 10276 81406
rect 10220 81302 10276 81340
rect 10108 80446 10110 80498
rect 10162 80446 10164 80498
rect 10108 80434 10164 80446
rect 10556 81170 10612 81182
rect 10556 81118 10558 81170
rect 10610 81118 10612 81170
rect 9772 80220 10164 80276
rect 9996 79604 10052 79614
rect 9884 79044 9940 79054
rect 9884 78036 9940 78988
rect 9884 77942 9940 77980
rect 9660 77252 9716 77262
rect 9660 77158 9716 77196
rect 9548 76850 9604 76860
rect 9772 76468 9828 76478
rect 9324 76412 9772 76468
rect 9772 76374 9828 76412
rect 8988 76354 9044 76366
rect 8988 76302 8990 76354
rect 9042 76302 9044 76354
rect 8988 76244 9044 76302
rect 8988 76178 9044 76188
rect 9772 75796 9828 75806
rect 9772 75702 9828 75740
rect 9100 75684 9156 75694
rect 8876 75682 9268 75684
rect 8876 75630 9102 75682
rect 9154 75630 9268 75682
rect 8876 75628 9268 75630
rect 9100 75618 9156 75628
rect 8540 75394 8596 75404
rect 8652 75572 8708 75582
rect 8540 75124 8596 75134
rect 8428 75122 8596 75124
rect 8428 75070 8542 75122
rect 8594 75070 8596 75122
rect 8428 75068 8596 75070
rect 6860 70980 6916 70990
rect 6860 70886 6916 70924
rect 6748 65828 6804 70812
rect 6972 67844 7028 71820
rect 7196 71650 7252 71662
rect 7196 71598 7198 71650
rect 7250 71598 7252 71650
rect 7084 70980 7140 70990
rect 7196 70980 7252 71598
rect 7532 71538 7588 75068
rect 7980 75030 8036 75068
rect 8540 75058 8596 75068
rect 8428 74898 8484 74910
rect 8428 74846 8430 74898
rect 8482 74846 8484 74898
rect 8016 73724 8280 73734
rect 8072 73668 8120 73724
rect 8176 73668 8224 73724
rect 8016 73658 8280 73668
rect 8428 73556 8484 74846
rect 8652 74228 8708 75516
rect 8764 75124 8820 75134
rect 8764 75030 8820 75068
rect 8988 74898 9044 74910
rect 8988 74846 8990 74898
rect 9042 74846 9044 74898
rect 8876 74674 8932 74686
rect 8876 74622 8878 74674
rect 8930 74622 8932 74674
rect 8652 74226 8820 74228
rect 8652 74174 8654 74226
rect 8706 74174 8820 74226
rect 8652 74172 8820 74174
rect 8652 74162 8708 74172
rect 8764 73892 8820 74172
rect 8764 73826 8820 73836
rect 8876 73668 8932 74622
rect 8988 74340 9044 74846
rect 9100 74340 9156 74350
rect 8988 74338 9156 74340
rect 8988 74286 9102 74338
rect 9154 74286 9156 74338
rect 8988 74284 9156 74286
rect 9100 74226 9156 74284
rect 9100 74174 9102 74226
rect 9154 74174 9156 74226
rect 7868 73218 7924 73230
rect 8316 73220 8372 73230
rect 7868 73166 7870 73218
rect 7922 73166 7924 73218
rect 7868 72772 7924 73166
rect 7868 72706 7924 72716
rect 8204 73218 8372 73220
rect 8204 73166 8318 73218
rect 8370 73166 8372 73218
rect 8204 73164 8372 73166
rect 7980 72660 8036 72670
rect 7980 72566 8036 72604
rect 7644 72548 7700 72558
rect 7644 71986 7700 72492
rect 8092 72548 8148 72558
rect 8204 72548 8260 73164
rect 8316 73154 8372 73164
rect 8428 72996 8484 73500
rect 8148 72492 8260 72548
rect 8316 72940 8484 72996
rect 8652 73612 8932 73668
rect 8988 74004 9044 74014
rect 8316 72546 8372 72940
rect 8316 72494 8318 72546
rect 8370 72494 8372 72546
rect 8092 72482 8148 72492
rect 8316 72482 8372 72494
rect 8428 72770 8484 72782
rect 8428 72718 8430 72770
rect 8482 72718 8484 72770
rect 8016 72156 8280 72166
rect 8072 72100 8120 72156
rect 8176 72100 8224 72156
rect 8016 72090 8280 72100
rect 7644 71934 7646 71986
rect 7698 71934 7700 71986
rect 7644 71922 7700 71934
rect 8428 71988 8484 72718
rect 8540 72772 8596 72782
rect 8540 72546 8596 72716
rect 8540 72494 8542 72546
rect 8594 72494 8596 72546
rect 8540 72482 8596 72494
rect 8540 71988 8596 71998
rect 8428 71986 8596 71988
rect 8428 71934 8542 71986
rect 8594 71934 8596 71986
rect 8428 71932 8596 71934
rect 8540 71922 8596 71932
rect 8428 71764 8484 71774
rect 7532 71486 7534 71538
rect 7586 71486 7588 71538
rect 7084 70978 7252 70980
rect 7084 70926 7086 70978
rect 7138 70926 7252 70978
rect 7084 70924 7252 70926
rect 7308 71202 7364 71214
rect 7308 71150 7310 71202
rect 7362 71150 7364 71202
rect 7084 70420 7140 70924
rect 7084 70354 7140 70364
rect 6972 67788 7252 67844
rect 7084 67620 7140 67630
rect 6860 66052 6916 66062
rect 7084 66052 7140 67564
rect 6916 65996 7140 66052
rect 6860 65958 6916 65996
rect 6748 65772 6916 65828
rect 6524 65436 6692 65492
rect 6412 64596 6468 64606
rect 6300 64594 6468 64596
rect 6300 64542 6414 64594
rect 6466 64542 6468 64594
rect 6300 64540 6468 64542
rect 6300 64146 6356 64540
rect 6412 64530 6468 64540
rect 6300 64094 6302 64146
rect 6354 64094 6356 64146
rect 6300 64082 6356 64094
rect 6412 64148 6468 64158
rect 6188 63970 6244 63980
rect 5740 63922 5796 63934
rect 5740 63870 5742 63922
rect 5794 63870 5796 63922
rect 5740 63700 5796 63870
rect 6076 63924 6132 63934
rect 6076 63830 6132 63868
rect 6300 63922 6356 63934
rect 6300 63870 6302 63922
rect 6354 63870 6356 63922
rect 6300 63700 6356 63870
rect 5740 63644 6356 63700
rect 5740 62188 5796 63644
rect 5292 62132 5460 62188
rect 5068 62076 5180 62132
rect 5068 61682 5124 62076
rect 5180 62066 5236 62076
rect 5068 61630 5070 61682
rect 5122 61630 5124 61682
rect 5068 61618 5124 61630
rect 5292 61796 5348 61806
rect 5180 61124 5236 61134
rect 5068 61068 5180 61124
rect 5068 60898 5124 61068
rect 5180 61058 5236 61068
rect 5068 60846 5070 60898
rect 5122 60846 5124 60898
rect 5068 60834 5124 60846
rect 5068 59778 5124 59790
rect 5068 59726 5070 59778
rect 5122 59726 5124 59778
rect 5068 57876 5124 59726
rect 5068 57782 5124 57820
rect 5180 59444 5236 59454
rect 5068 56980 5124 56990
rect 5180 56980 5236 59388
rect 5068 56978 5236 56980
rect 5068 56926 5070 56978
rect 5122 56926 5236 56978
rect 5068 56924 5236 56926
rect 5068 56914 5124 56924
rect 5180 56532 5236 56924
rect 5292 56756 5348 61740
rect 5404 56980 5460 62132
rect 5404 56914 5460 56924
rect 5516 62132 5796 62188
rect 5852 63476 5908 63486
rect 5852 62244 5908 63420
rect 5292 56690 5348 56700
rect 5516 56756 5572 62132
rect 5852 61572 5908 62188
rect 5628 61516 5908 61572
rect 5964 62132 6020 62142
rect 5964 61570 6020 62076
rect 6188 61684 6244 61694
rect 5964 61518 5966 61570
rect 6018 61518 6020 61570
rect 5628 61458 5684 61516
rect 5964 61506 6020 61518
rect 6076 61572 6132 61582
rect 6076 61478 6132 61516
rect 6188 61570 6244 61628
rect 6188 61518 6190 61570
rect 6242 61518 6244 61570
rect 5628 61406 5630 61458
rect 5682 61406 5684 61458
rect 5628 58828 5684 61406
rect 5740 61346 5796 61358
rect 5740 61294 5742 61346
rect 5794 61294 5796 61346
rect 5740 61124 5796 61294
rect 5740 61058 5796 61068
rect 5740 60564 5796 60574
rect 5740 60228 5796 60508
rect 6188 60340 6244 61518
rect 5740 60002 5796 60172
rect 5740 59950 5742 60002
rect 5794 59950 5796 60002
rect 5740 59938 5796 59950
rect 5852 60284 6244 60340
rect 5740 59444 5796 59454
rect 5852 59444 5908 60284
rect 6412 60228 6468 64092
rect 6524 63364 6580 65436
rect 6636 64820 6692 64830
rect 6636 64148 6692 64764
rect 6636 64092 6804 64148
rect 6636 63922 6692 63934
rect 6636 63870 6638 63922
rect 6690 63870 6692 63922
rect 6636 63812 6692 63870
rect 6636 63746 6692 63756
rect 6636 63364 6692 63374
rect 6524 63308 6636 63364
rect 6636 63298 6692 63308
rect 6748 63138 6804 64092
rect 6748 63086 6750 63138
rect 6802 63086 6804 63138
rect 6748 62580 6804 63086
rect 6748 62514 6804 62524
rect 5796 59388 5908 59444
rect 5964 60172 6468 60228
rect 6524 62356 6580 62366
rect 5740 59350 5796 59388
rect 5628 58772 5796 58828
rect 5628 58436 5684 58446
rect 5628 58342 5684 58380
rect 5516 56690 5572 56700
rect 5628 57316 5684 57326
rect 5628 56866 5684 57260
rect 5740 56980 5796 58772
rect 5852 57988 5908 57998
rect 5964 57988 6020 60172
rect 6524 60116 6580 62300
rect 6636 62244 6692 62282
rect 6860 62188 6916 65772
rect 6972 63924 7028 65996
rect 7196 65828 7252 67788
rect 7084 65772 7252 65828
rect 7084 65268 7140 65772
rect 7308 65716 7364 71150
rect 7420 70868 7476 70878
rect 7532 70868 7588 71486
rect 8092 71650 8148 71662
rect 8092 71598 8094 71650
rect 8146 71598 8148 71650
rect 8092 71538 8148 71598
rect 8092 71486 8094 71538
rect 8146 71486 8148 71538
rect 8092 71474 8148 71486
rect 8092 71202 8148 71214
rect 8092 71150 8094 71202
rect 8146 71150 8148 71202
rect 7980 71092 8036 71102
rect 7476 70812 7588 70868
rect 7420 70802 7476 70812
rect 7532 70754 7588 70812
rect 7532 70702 7534 70754
rect 7586 70702 7588 70754
rect 7532 70690 7588 70702
rect 7868 71036 7980 71092
rect 8092 71092 8148 71150
rect 8428 71202 8484 71708
rect 8652 71652 8708 73612
rect 8988 73556 9044 73948
rect 8764 73554 9044 73556
rect 8764 73502 8990 73554
rect 9042 73502 9044 73554
rect 8764 73500 9044 73502
rect 8764 72546 8820 73500
rect 8988 73490 9044 73500
rect 8764 72494 8766 72546
rect 8818 72494 8820 72546
rect 8764 72482 8820 72494
rect 8876 72548 8932 72558
rect 8876 71986 8932 72492
rect 8988 72548 9044 72558
rect 9100 72548 9156 74174
rect 9212 74004 9268 75628
rect 9772 75460 9828 75470
rect 9772 75122 9828 75404
rect 9772 75070 9774 75122
rect 9826 75070 9828 75122
rect 9772 75058 9828 75070
rect 9996 75124 10052 79548
rect 10108 79602 10164 80220
rect 10108 79550 10110 79602
rect 10162 79550 10164 79602
rect 10108 79538 10164 79550
rect 10332 79602 10388 79614
rect 10332 79550 10334 79602
rect 10386 79550 10388 79602
rect 10332 78932 10388 79550
rect 10556 79490 10612 81118
rect 10780 81170 10836 81676
rect 10780 81118 10782 81170
rect 10834 81118 10836 81170
rect 10780 81106 10836 81118
rect 10556 79438 10558 79490
rect 10610 79438 10612 79490
rect 10556 79380 10612 79438
rect 10556 79314 10612 79324
rect 10668 79378 10724 79390
rect 10668 79326 10670 79378
rect 10722 79326 10724 79378
rect 10332 78866 10388 78876
rect 10332 78708 10388 78718
rect 10108 77252 10164 77262
rect 10108 77158 10164 77196
rect 10108 76468 10164 76478
rect 10108 76374 10164 76412
rect 10220 76354 10276 76366
rect 10220 76302 10222 76354
rect 10274 76302 10276 76354
rect 10220 75796 10276 76302
rect 10220 75730 10276 75740
rect 9548 74898 9604 74910
rect 9548 74846 9550 74898
rect 9602 74846 9604 74898
rect 9324 74004 9380 74014
rect 9212 73948 9324 74004
rect 8988 72546 9156 72548
rect 8988 72494 8990 72546
rect 9042 72494 9156 72546
rect 8988 72492 9156 72494
rect 9324 72660 9380 73948
rect 9548 73890 9604 74846
rect 9996 74226 10052 75068
rect 10220 75012 10276 75022
rect 10332 75012 10388 78652
rect 10668 76692 10724 79326
rect 10780 77140 10836 77150
rect 10780 77046 10836 77084
rect 10556 76636 10724 76692
rect 10444 76580 10500 76590
rect 10444 75572 10500 76524
rect 10444 75506 10500 75516
rect 9996 74174 9998 74226
rect 10050 74174 10052 74226
rect 9996 74116 10052 74174
rect 9548 73838 9550 73890
rect 9602 73838 9604 73890
rect 9548 73556 9604 73838
rect 9772 73892 9828 73902
rect 9772 73780 9828 73836
rect 9772 73724 9940 73780
rect 9660 73556 9716 73566
rect 9604 73554 9716 73556
rect 9604 73502 9662 73554
rect 9714 73502 9716 73554
rect 9604 73500 9716 73502
rect 9548 73490 9604 73500
rect 9660 73490 9716 73500
rect 9324 72546 9380 72604
rect 9324 72494 9326 72546
rect 9378 72494 9380 72546
rect 8988 72482 9044 72492
rect 8876 71934 8878 71986
rect 8930 71934 8932 71986
rect 8876 71922 8932 71934
rect 9100 72324 9156 72334
rect 8764 71764 8820 71774
rect 8764 71670 8820 71708
rect 8988 71762 9044 71774
rect 8988 71710 8990 71762
rect 9042 71710 9044 71762
rect 8428 71150 8430 71202
rect 8482 71150 8484 71202
rect 8428 71138 8484 71150
rect 8540 71596 8708 71652
rect 8988 71652 9044 71710
rect 8316 71092 8372 71102
rect 8092 71090 8372 71092
rect 8092 71038 8318 71090
rect 8370 71038 8372 71090
rect 8092 71036 8372 71038
rect 8540 71092 8596 71596
rect 8988 71586 9044 71596
rect 8876 71092 8932 71102
rect 8540 71036 8820 71092
rect 7868 70194 7924 71036
rect 7980 71026 8036 71036
rect 8316 71026 8372 71036
rect 7980 70756 8036 70794
rect 7980 70690 8036 70700
rect 8540 70644 8596 70654
rect 8016 70588 8280 70598
rect 8072 70532 8120 70588
rect 8176 70532 8224 70588
rect 8016 70522 8280 70532
rect 8428 70588 8540 70644
rect 8428 70420 8484 70588
rect 8540 70578 8596 70588
rect 7868 70142 7870 70194
rect 7922 70142 7924 70194
rect 7868 70130 7924 70142
rect 8316 70364 8484 70420
rect 8316 69634 8372 70364
rect 8316 69582 8318 69634
rect 8370 69582 8372 69634
rect 8316 69570 8372 69582
rect 8204 69412 8260 69422
rect 7644 69410 8260 69412
rect 7644 69358 8206 69410
rect 8258 69358 8260 69410
rect 7644 69356 8260 69358
rect 7644 68516 7700 69356
rect 8204 69346 8260 69356
rect 8764 69410 8820 71036
rect 8876 70998 8932 71036
rect 9100 69524 9156 72268
rect 9324 72100 9380 72494
rect 8764 69358 8766 69410
rect 8818 69358 8820 69410
rect 8764 69346 8820 69358
rect 8876 69468 9156 69524
rect 9212 72044 9380 72100
rect 9212 69524 9268 72044
rect 9548 71764 9604 71774
rect 9436 71762 9604 71764
rect 9436 71710 9550 71762
rect 9602 71710 9604 71762
rect 9436 71708 9604 71710
rect 9436 71652 9492 71708
rect 9548 71698 9604 71708
rect 9772 71762 9828 71774
rect 9772 71710 9774 71762
rect 9826 71710 9828 71762
rect 9436 70754 9492 71596
rect 9660 71652 9716 71662
rect 9660 71558 9716 71596
rect 9548 71540 9604 71550
rect 9548 71090 9604 71484
rect 9548 71038 9550 71090
rect 9602 71038 9604 71090
rect 9548 71026 9604 71038
rect 9436 70702 9438 70754
rect 9490 70702 9492 70754
rect 9436 69860 9492 70702
rect 9660 70754 9716 70766
rect 9660 70702 9662 70754
rect 9714 70702 9716 70754
rect 9548 70308 9604 70318
rect 9548 70214 9604 70252
rect 9436 69794 9492 69804
rect 9212 69468 9604 69524
rect 7420 68514 7700 68516
rect 7420 68462 7646 68514
rect 7698 68462 7700 68514
rect 7420 68460 7700 68462
rect 7420 66724 7476 68460
rect 7644 68450 7700 68460
rect 7868 69186 7924 69198
rect 7868 69134 7870 69186
rect 7922 69134 7924 69186
rect 7756 67956 7812 67966
rect 7868 67956 7924 69134
rect 8428 69188 8484 69198
rect 8016 69020 8280 69030
rect 8072 68964 8120 69020
rect 8176 68964 8224 69020
rect 8016 68954 8280 68964
rect 8428 68850 8484 69132
rect 8428 68798 8430 68850
rect 8482 68798 8484 68850
rect 8428 68786 8484 68798
rect 7812 67900 7924 67956
rect 8316 68514 8372 68526
rect 8316 68462 8318 68514
rect 8370 68462 8372 68514
rect 7756 67862 7812 67900
rect 8316 67620 8372 68462
rect 8876 68068 8932 69468
rect 9212 69412 9268 69468
rect 8988 69356 9268 69412
rect 8988 68850 9044 69356
rect 9324 69300 9380 69310
rect 9324 69206 9380 69244
rect 9212 69188 9268 69198
rect 9212 69094 9268 69132
rect 9436 69188 9492 69198
rect 8988 68798 8990 68850
rect 9042 68798 9044 68850
rect 8988 68786 9044 68798
rect 9436 68068 9492 69132
rect 8652 68012 8932 68068
rect 9212 68012 9492 68068
rect 9548 68626 9604 69468
rect 9548 68574 9550 68626
rect 9602 68574 9604 68626
rect 8316 67564 8484 67620
rect 8016 67452 8280 67462
rect 8072 67396 8120 67452
rect 8176 67396 8224 67452
rect 8016 67386 8280 67396
rect 8092 67284 8148 67294
rect 8428 67284 8484 67564
rect 7532 67282 8484 67284
rect 7532 67230 8094 67282
rect 8146 67230 8484 67282
rect 7532 67228 8484 67230
rect 7532 66946 7588 67228
rect 8092 67218 8148 67228
rect 7532 66894 7534 66946
rect 7586 66894 7588 66946
rect 7532 66882 7588 66894
rect 7868 67058 7924 67070
rect 7868 67006 7870 67058
rect 7922 67006 7924 67058
rect 7868 66836 7924 67006
rect 8428 67058 8484 67070
rect 8428 67006 8430 67058
rect 8482 67006 8484 67058
rect 7980 66948 8036 66958
rect 7980 66854 8036 66892
rect 8428 66946 8484 67006
rect 8428 66894 8430 66946
rect 8482 66894 8484 66946
rect 7868 66770 7924 66780
rect 7420 66668 7588 66724
rect 7196 65660 7364 65716
rect 7420 65716 7476 65726
rect 7196 65492 7252 65660
rect 7196 65426 7252 65436
rect 7308 65490 7364 65502
rect 7308 65438 7310 65490
rect 7362 65438 7364 65490
rect 7084 65212 7252 65268
rect 7196 64708 7252 65212
rect 7084 63924 7140 63934
rect 6972 63868 7084 63924
rect 7084 63810 7140 63868
rect 7084 63758 7086 63810
rect 7138 63758 7140 63810
rect 7084 62356 7140 63758
rect 7084 62290 7140 62300
rect 7196 62188 7252 64652
rect 6636 62178 6692 62188
rect 6748 62132 6916 62188
rect 6972 62132 7252 62188
rect 7308 63924 7364 65438
rect 7420 65490 7476 65660
rect 7532 65714 7588 66668
rect 8316 66388 8372 66398
rect 8316 66274 8372 66332
rect 8316 66222 8318 66274
rect 8370 66222 8372 66274
rect 8316 66210 8372 66222
rect 8016 65884 8280 65894
rect 8072 65828 8120 65884
rect 8176 65828 8224 65884
rect 8016 65818 8280 65828
rect 8428 65716 8484 66894
rect 7532 65662 7534 65714
rect 7586 65662 7588 65714
rect 7532 65650 7588 65662
rect 8316 65660 8484 65716
rect 7420 65438 7422 65490
rect 7474 65438 7476 65490
rect 7420 65426 7476 65438
rect 7644 65492 7700 65502
rect 7644 64146 7700 65436
rect 7980 65490 8036 65502
rect 7980 65438 7982 65490
rect 8034 65438 8036 65490
rect 7980 65380 8036 65438
rect 8316 65380 8372 65660
rect 7980 65378 8372 65380
rect 7980 65326 8318 65378
rect 8370 65326 8372 65378
rect 7980 65324 8372 65326
rect 8316 64596 8372 65324
rect 8428 65492 8484 65502
rect 8428 64820 8484 65436
rect 8540 64820 8596 64830
rect 8428 64818 8596 64820
rect 8428 64766 8542 64818
rect 8594 64766 8596 64818
rect 8428 64764 8596 64766
rect 8540 64754 8596 64764
rect 8316 64540 8484 64596
rect 8016 64316 8280 64326
rect 8072 64260 8120 64316
rect 8176 64260 8224 64316
rect 8016 64250 8280 64260
rect 7644 64094 7646 64146
rect 7698 64094 7700 64146
rect 7644 64082 7700 64094
rect 7420 63924 7476 63934
rect 7308 63868 7420 63924
rect 6748 61458 6804 62132
rect 6860 61572 6916 61582
rect 6860 61478 6916 61516
rect 6748 61406 6750 61458
rect 6802 61406 6804 61458
rect 6748 61348 6804 61406
rect 6972 61348 7028 62132
rect 6748 61282 6804 61292
rect 6860 61292 7028 61348
rect 7084 61570 7140 61582
rect 7084 61518 7086 61570
rect 7138 61518 7140 61570
rect 7084 61460 7140 61518
rect 6300 60060 6580 60116
rect 6748 60452 6804 60462
rect 6188 59108 6244 59118
rect 5908 57932 6020 57988
rect 5852 57922 5908 57932
rect 5964 57874 6020 57932
rect 5964 57822 5966 57874
rect 6018 57822 6020 57874
rect 5964 57810 6020 57822
rect 6076 58546 6132 58558
rect 6076 58494 6078 58546
rect 6130 58494 6132 58546
rect 6076 57764 6132 58494
rect 6076 57698 6132 57708
rect 6188 57540 6244 59052
rect 6300 58828 6356 60060
rect 6412 59890 6468 59902
rect 6412 59838 6414 59890
rect 6466 59838 6468 59890
rect 6412 59444 6468 59838
rect 6636 59444 6692 59454
rect 6412 59442 6692 59444
rect 6412 59390 6638 59442
rect 6690 59390 6692 59442
rect 6412 59388 6692 59390
rect 6636 59378 6692 59388
rect 6524 59220 6580 59230
rect 6524 59126 6580 59164
rect 6748 59218 6804 60396
rect 6748 59166 6750 59218
rect 6802 59166 6804 59218
rect 6748 59108 6804 59166
rect 6860 59220 6916 61292
rect 7084 60676 7140 61404
rect 7196 60676 7252 60686
rect 7084 60674 7252 60676
rect 7084 60622 7198 60674
rect 7250 60622 7252 60674
rect 7084 60620 7252 60622
rect 7196 60610 7252 60620
rect 7308 59444 7364 63868
rect 7420 63830 7476 63868
rect 8092 63924 8148 63934
rect 8428 63924 8484 64540
rect 8092 63922 8484 63924
rect 8092 63870 8094 63922
rect 8146 63870 8430 63922
rect 8482 63870 8484 63922
rect 8092 63868 8484 63870
rect 8092 63858 8148 63868
rect 7532 63812 7588 63822
rect 7532 63718 7588 63756
rect 7532 63028 7588 63038
rect 7532 63026 7924 63028
rect 7532 62974 7534 63026
rect 7586 62974 7924 63026
rect 7532 62972 7924 62974
rect 7532 62962 7588 62972
rect 7868 62578 7924 62972
rect 8428 62916 8484 63868
rect 8428 62850 8484 62860
rect 8016 62748 8280 62758
rect 8072 62692 8120 62748
rect 8176 62692 8224 62748
rect 8016 62682 8280 62692
rect 7868 62526 7870 62578
rect 7922 62526 7924 62578
rect 7868 62514 7924 62526
rect 7980 62580 8036 62590
rect 7756 62356 7812 62366
rect 7756 62262 7812 62300
rect 7420 62242 7476 62254
rect 7420 62190 7422 62242
rect 7474 62190 7476 62242
rect 7420 62188 7476 62190
rect 7420 62132 7812 62188
rect 7756 61460 7812 62132
rect 7980 61682 8036 62524
rect 8428 62580 8484 62590
rect 8316 62468 8372 62478
rect 8316 62374 8372 62412
rect 7980 61630 7982 61682
rect 8034 61630 8036 61682
rect 7980 61618 8036 61630
rect 8092 62354 8148 62366
rect 8092 62302 8094 62354
rect 8146 62302 8148 62354
rect 8092 61460 8148 62302
rect 7756 61404 8148 61460
rect 7532 61348 7588 61358
rect 7532 60788 7588 61292
rect 7532 60562 7588 60732
rect 7532 60510 7534 60562
rect 7586 60510 7588 60562
rect 6860 59154 6916 59164
rect 6972 59388 7364 59444
rect 7420 59444 7476 59454
rect 6748 59042 6804 59052
rect 6300 58772 6580 58828
rect 6300 57876 6356 57886
rect 6300 57762 6356 57820
rect 6300 57710 6302 57762
rect 6354 57710 6356 57762
rect 6300 57698 6356 57710
rect 6076 57484 6244 57540
rect 6412 57538 6468 57550
rect 6412 57486 6414 57538
rect 6466 57486 6468 57538
rect 6076 57204 6132 57484
rect 6412 57316 6468 57486
rect 6076 57138 6132 57148
rect 6188 57260 6468 57316
rect 6188 57090 6244 57260
rect 6188 57038 6190 57090
rect 6242 57038 6244 57090
rect 6188 57026 6244 57038
rect 6412 56980 6468 56990
rect 5740 56924 6020 56980
rect 5628 56814 5630 56866
rect 5682 56814 5684 56866
rect 5628 56644 5684 56814
rect 5852 56756 5908 56766
rect 5852 56662 5908 56700
rect 5628 56578 5684 56588
rect 5740 56642 5796 56654
rect 5740 56590 5742 56642
rect 5794 56590 5796 56642
rect 5180 56466 5236 56476
rect 5740 56308 5796 56590
rect 4956 56252 5236 56308
rect 4620 56030 4622 56082
rect 4674 56030 4676 56082
rect 4620 56018 4676 56030
rect 4956 56084 5012 56094
rect 4284 55794 4340 55804
rect 4614 55692 4878 55702
rect 4670 55636 4718 55692
rect 4774 55636 4822 55692
rect 4614 55626 4878 55636
rect 4956 55524 5012 56028
rect 4620 55468 5012 55524
rect 4620 55410 4676 55468
rect 4620 55358 4622 55410
rect 4674 55358 4676 55410
rect 4620 55346 4676 55358
rect 5068 55074 5124 55086
rect 5068 55022 5070 55074
rect 5122 55022 5124 55074
rect 3276 53118 3278 53170
rect 3330 53118 3332 53170
rect 2940 50082 2996 50092
rect 3052 51156 3108 51166
rect 2828 49922 2884 49934
rect 2828 49870 2830 49922
rect 2882 49870 2884 49922
rect 2604 49812 2660 49822
rect 2828 49812 2884 49870
rect 2660 49756 2884 49812
rect 2492 49698 2548 49710
rect 2492 49646 2494 49698
rect 2546 49646 2548 49698
rect 2492 49588 2548 49646
rect 2492 49522 2548 49532
rect 2604 49138 2660 49756
rect 2604 49086 2606 49138
rect 2658 49086 2660 49138
rect 2604 49074 2660 49086
rect 2492 48132 2548 48142
rect 2492 48038 2548 48076
rect 2492 47572 2548 47582
rect 2492 47478 2548 47516
rect 2828 47460 2884 49756
rect 2940 48804 2996 48814
rect 3052 48804 3108 51100
rect 3164 50484 3220 50494
rect 3164 50034 3220 50428
rect 3164 49982 3166 50034
rect 3218 49982 3220 50034
rect 3164 49970 3220 49982
rect 3276 50036 3332 53118
rect 3724 52388 3780 53900
rect 4060 53890 4116 53900
rect 4396 54628 4452 54638
rect 3836 53732 3892 53742
rect 4396 53732 4452 54572
rect 4956 54402 5012 54414
rect 4956 54350 4958 54402
rect 5010 54350 5012 54402
rect 4614 54124 4878 54134
rect 4670 54068 4718 54124
rect 4774 54068 4822 54124
rect 4614 54058 4878 54068
rect 3836 53638 3892 53676
rect 4284 53730 4452 53732
rect 4284 53678 4398 53730
rect 4450 53678 4452 53730
rect 4284 53676 4452 53678
rect 4172 53620 4228 53630
rect 4172 53526 4228 53564
rect 3836 53284 3892 53294
rect 3836 53170 3892 53228
rect 3836 53118 3838 53170
rect 3890 53118 3892 53170
rect 3836 53106 3892 53118
rect 4284 53170 4340 53676
rect 4396 53666 4452 53676
rect 4508 53956 4564 53966
rect 4284 53118 4286 53170
rect 4338 53118 4340 53170
rect 4060 52948 4116 52958
rect 3724 52322 3780 52332
rect 3948 52946 4116 52948
rect 3948 52894 4062 52946
rect 4114 52894 4116 52946
rect 3948 52892 4116 52894
rect 3388 52276 3444 52286
rect 3388 52182 3444 52220
rect 3724 52164 3780 52174
rect 3948 52164 4004 52892
rect 4060 52882 4116 52892
rect 4284 52276 4340 53118
rect 4508 53170 4564 53900
rect 4732 53956 4788 53966
rect 4620 53844 4676 53854
rect 4620 53730 4676 53788
rect 4732 53842 4788 53900
rect 4732 53790 4734 53842
rect 4786 53790 4788 53842
rect 4732 53778 4788 53790
rect 4620 53678 4622 53730
rect 4674 53678 4676 53730
rect 4620 53666 4676 53678
rect 4956 53620 5012 54350
rect 5068 54290 5124 55022
rect 5068 54238 5070 54290
rect 5122 54238 5124 54290
rect 5068 54226 5124 54238
rect 4956 53554 5012 53564
rect 4732 53506 4788 53518
rect 5180 53508 5236 56252
rect 5292 56252 5796 56308
rect 5292 56194 5348 56252
rect 5292 56142 5294 56194
rect 5346 56142 5348 56194
rect 5292 56130 5348 56142
rect 5516 55860 5572 55870
rect 5292 54740 5348 54750
rect 5292 53844 5348 54684
rect 5292 53778 5348 53788
rect 5404 54628 5460 54638
rect 4732 53454 4734 53506
rect 4786 53454 4788 53506
rect 4508 53118 4510 53170
rect 4562 53118 4564 53170
rect 4508 53106 4564 53118
rect 4620 53172 4676 53182
rect 4732 53172 4788 53454
rect 5068 53452 5236 53508
rect 5068 53284 5124 53452
rect 4620 53170 4788 53172
rect 4620 53118 4622 53170
rect 4674 53118 4788 53170
rect 4620 53116 4788 53118
rect 4620 53106 4676 53116
rect 4620 52948 4676 52958
rect 4620 52834 4676 52892
rect 4620 52782 4622 52834
rect 4674 52782 4676 52834
rect 4620 52770 4676 52782
rect 4732 52724 4788 53116
rect 4732 52658 4788 52668
rect 4956 53228 5124 53284
rect 5180 53284 5236 53294
rect 4614 52556 4878 52566
rect 4670 52500 4718 52556
rect 4774 52500 4822 52556
rect 4614 52490 4878 52500
rect 3780 52108 4004 52164
rect 4172 52162 4228 52174
rect 4172 52110 4174 52162
rect 4226 52110 4228 52162
rect 3724 52070 3780 52108
rect 4060 51490 4116 51502
rect 4060 51438 4062 51490
rect 4114 51438 4116 51490
rect 3612 51380 3668 51418
rect 3612 51314 3668 51324
rect 3948 51266 4004 51278
rect 3948 51214 3950 51266
rect 4002 51214 4004 51266
rect 3836 51156 3892 51166
rect 3836 51062 3892 51100
rect 3276 49924 3332 49980
rect 3276 49868 3444 49924
rect 2940 48802 3108 48804
rect 2940 48750 2942 48802
rect 2994 48750 3108 48802
rect 2940 48748 3108 48750
rect 3164 49812 3220 49822
rect 2940 48356 2996 48748
rect 2940 48290 2996 48300
rect 3052 48132 3108 48142
rect 3052 47570 3108 48076
rect 3164 47684 3220 49756
rect 3388 49810 3444 49868
rect 3388 49758 3390 49810
rect 3442 49758 3444 49810
rect 3388 49746 3444 49758
rect 3388 49588 3444 49598
rect 3948 49588 4004 51214
rect 4060 50820 4116 51438
rect 4060 50754 4116 50764
rect 3388 49586 4004 49588
rect 3388 49534 3390 49586
rect 3442 49534 4004 49586
rect 3388 49532 4004 49534
rect 4172 49698 4228 52110
rect 4284 52162 4340 52220
rect 4284 52110 4286 52162
rect 4338 52110 4340 52162
rect 4284 50260 4340 52110
rect 4732 52388 4788 52398
rect 4732 52162 4788 52332
rect 4732 52110 4734 52162
rect 4786 52110 4788 52162
rect 4732 52098 4788 52110
rect 4508 52052 4564 52062
rect 4396 51940 4452 51950
rect 4396 51846 4452 51884
rect 4508 51940 4564 51996
rect 4956 51940 5012 53228
rect 5068 53060 5124 53070
rect 5068 52946 5124 53004
rect 5068 52894 5070 52946
rect 5122 52894 5124 52946
rect 5068 52882 5124 52894
rect 4508 51938 5012 51940
rect 4508 51886 4510 51938
rect 4562 51886 5012 51938
rect 4508 51884 5012 51886
rect 4508 51874 4564 51884
rect 5180 51716 5236 53228
rect 5292 53172 5348 53182
rect 5404 53172 5460 54572
rect 5292 53170 5460 53172
rect 5292 53118 5294 53170
rect 5346 53118 5460 53170
rect 5292 53116 5460 53118
rect 5516 53170 5572 55804
rect 5964 55412 6020 56924
rect 6188 56866 6244 56878
rect 6188 56814 6190 56866
rect 6242 56814 6244 56866
rect 6188 56532 6244 56814
rect 6188 56466 6244 56476
rect 5740 55356 6020 55412
rect 5740 54738 5796 55356
rect 5740 54686 5742 54738
rect 5794 54686 5796 54738
rect 5740 54674 5796 54686
rect 5628 54290 5684 54302
rect 5628 54238 5630 54290
rect 5682 54238 5684 54290
rect 5628 53732 5684 54238
rect 5628 53638 5684 53676
rect 5852 53844 5908 53854
rect 5516 53118 5518 53170
rect 5570 53118 5572 53170
rect 5292 53106 5348 53116
rect 5516 53106 5572 53118
rect 5628 53172 5684 53182
rect 5628 53170 5796 53172
rect 5628 53118 5630 53170
rect 5682 53118 5796 53170
rect 5628 53116 5796 53118
rect 5628 53106 5684 53116
rect 5740 53060 5796 53116
rect 5740 52994 5796 53004
rect 5628 52836 5684 52846
rect 5628 52834 5796 52836
rect 5628 52782 5630 52834
rect 5682 52782 5796 52834
rect 5628 52780 5796 52782
rect 5628 52770 5684 52780
rect 5740 52724 5796 52780
rect 5740 52658 5796 52668
rect 5852 52500 5908 53788
rect 5964 53060 6020 55356
rect 6076 55074 6132 55086
rect 6076 55022 6078 55074
rect 6130 55022 6132 55074
rect 6076 54628 6132 55022
rect 6076 54562 6132 54572
rect 6188 54404 6244 54414
rect 6188 54310 6244 54348
rect 6300 53844 6356 53854
rect 6412 53844 6468 56924
rect 6356 53788 6468 53844
rect 6300 53778 6356 53788
rect 6300 53620 6356 53630
rect 6300 53284 6356 53564
rect 6076 53060 6132 53070
rect 5964 53058 6132 53060
rect 5964 53006 6078 53058
rect 6130 53006 6132 53058
rect 5964 53004 6132 53006
rect 6076 52994 6132 53004
rect 6300 53058 6356 53228
rect 6412 53618 6468 53630
rect 6412 53566 6414 53618
rect 6466 53566 6468 53618
rect 6412 53170 6468 53566
rect 6412 53118 6414 53170
rect 6466 53118 6468 53170
rect 6412 53106 6468 53118
rect 6300 53006 6302 53058
rect 6354 53006 6356 53058
rect 6300 52994 6356 53006
rect 5740 52444 5908 52500
rect 5068 51660 5236 51716
rect 5628 52052 5684 52062
rect 4732 51604 4788 51614
rect 4732 51510 4788 51548
rect 4614 50988 4878 50998
rect 4670 50932 4718 50988
rect 4774 50932 4822 50988
rect 4614 50922 4878 50932
rect 4620 50820 4676 50830
rect 4620 50706 4676 50764
rect 4620 50654 4622 50706
rect 4674 50654 4676 50706
rect 4620 50642 4676 50654
rect 4284 50204 4452 50260
rect 4172 49646 4174 49698
rect 4226 49646 4228 49698
rect 3388 49522 3444 49532
rect 4172 49476 4228 49646
rect 3724 49420 4228 49476
rect 4284 50036 4340 50046
rect 3612 49028 3668 49038
rect 3612 48934 3668 48972
rect 3612 48804 3668 48814
rect 3164 47618 3220 47628
rect 3500 47684 3556 47694
rect 3500 47590 3556 47628
rect 3052 47518 3054 47570
rect 3106 47518 3108 47570
rect 3052 47506 3108 47518
rect 2940 47460 2996 47470
rect 2828 47458 2996 47460
rect 2828 47406 2942 47458
rect 2994 47406 2996 47458
rect 2828 47404 2996 47406
rect 2604 47348 2660 47358
rect 2604 46340 2660 47292
rect 2716 46564 2772 46574
rect 2828 46564 2884 47404
rect 2940 47394 2996 47404
rect 3164 47460 3220 47470
rect 3164 47366 3220 47404
rect 3500 47458 3556 47470
rect 3500 47406 3502 47458
rect 3554 47406 3556 47458
rect 3500 47348 3556 47406
rect 3500 47068 3556 47292
rect 2716 46562 2884 46564
rect 2716 46510 2718 46562
rect 2770 46510 2884 46562
rect 2716 46508 2884 46510
rect 2716 46498 2772 46508
rect 2604 46284 2772 46340
rect 2380 45714 2436 45724
rect 2492 45780 2548 45790
rect 2492 45778 2660 45780
rect 2492 45726 2494 45778
rect 2546 45726 2660 45778
rect 2492 45724 2660 45726
rect 2492 45714 2548 45724
rect 2156 45500 2548 45556
rect 2380 45332 2436 45342
rect 2044 44942 2046 44994
rect 2098 44942 2100 44994
rect 2044 44660 2100 44942
rect 1932 44604 2100 44660
rect 2268 45106 2324 45118
rect 2268 45054 2270 45106
rect 2322 45054 2324 45106
rect 1820 43764 1876 43774
rect 1708 43708 1820 43764
rect 1820 43698 1876 43708
rect 1820 42754 1876 42766
rect 1820 42702 1822 42754
rect 1874 42702 1876 42754
rect 1708 42420 1764 42430
rect 1708 41970 1764 42364
rect 1708 41918 1710 41970
rect 1762 41918 1764 41970
rect 1708 40628 1764 41918
rect 1596 40572 1764 40628
rect 1596 38948 1652 40572
rect 1708 40402 1764 40414
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 39732 1764 40350
rect 1708 39060 1764 39676
rect 1820 39620 1876 42702
rect 1932 39844 1988 44604
rect 2268 44546 2324 45054
rect 2268 44494 2270 44546
rect 2322 44494 2324 44546
rect 2268 44482 2324 44494
rect 2380 44212 2436 45276
rect 2492 44882 2548 45500
rect 2604 45330 2660 45724
rect 2604 45278 2606 45330
rect 2658 45278 2660 45330
rect 2604 45266 2660 45278
rect 2492 44830 2494 44882
rect 2546 44830 2548 44882
rect 2492 44818 2548 44830
rect 2492 44436 2548 44446
rect 2716 44436 2772 46284
rect 2828 45332 2884 46508
rect 3164 47012 3556 47068
rect 3164 46564 3220 47012
rect 3612 46788 3668 48748
rect 3612 46722 3668 46732
rect 3164 46470 3220 46508
rect 3612 46562 3668 46574
rect 3612 46510 3614 46562
rect 3666 46510 3668 46562
rect 3612 46452 3668 46510
rect 3612 46386 3668 46396
rect 2828 45266 2884 45276
rect 3612 45220 3668 45230
rect 2828 45108 2884 45118
rect 2828 45014 2884 45052
rect 3052 45108 3108 45118
rect 3500 45108 3556 45118
rect 3612 45108 3668 45164
rect 3052 45106 3332 45108
rect 3052 45054 3054 45106
rect 3106 45054 3332 45106
rect 3052 45052 3332 45054
rect 3052 45042 3108 45052
rect 2492 44434 2772 44436
rect 2492 44382 2494 44434
rect 2546 44382 2772 44434
rect 2492 44380 2772 44382
rect 2828 44884 2884 44894
rect 2828 44436 2884 44828
rect 2492 44370 2548 44380
rect 2492 44212 2548 44222
rect 2380 44156 2492 44212
rect 2492 44146 2548 44156
rect 2156 44100 2212 44110
rect 2156 44098 2324 44100
rect 2156 44046 2158 44098
rect 2210 44046 2324 44098
rect 2156 44044 2324 44046
rect 2156 44034 2212 44044
rect 2156 43764 2212 43774
rect 2268 43764 2324 44044
rect 2380 43764 2436 43774
rect 2268 43708 2380 43764
rect 2156 43670 2212 43708
rect 2380 43698 2436 43708
rect 2492 43652 2548 43662
rect 2492 43558 2548 43596
rect 2828 43538 2884 44380
rect 3164 44546 3220 44558
rect 3164 44494 3166 44546
rect 3218 44494 3220 44546
rect 3052 44100 3108 44110
rect 3052 44006 3108 44044
rect 3164 43876 3220 44494
rect 2828 43486 2830 43538
rect 2882 43486 2884 43538
rect 2828 43474 2884 43486
rect 2940 43820 3220 43876
rect 2604 43426 2660 43438
rect 2604 43374 2606 43426
rect 2658 43374 2660 43426
rect 2492 42642 2548 42654
rect 2492 42590 2494 42642
rect 2546 42590 2548 42642
rect 2492 42194 2548 42590
rect 2492 42142 2494 42194
rect 2546 42142 2548 42194
rect 2492 42130 2548 42142
rect 2044 42082 2100 42094
rect 2044 42030 2046 42082
rect 2098 42030 2100 42082
rect 2044 41188 2100 42030
rect 2044 41132 2212 41188
rect 2044 40964 2100 40974
rect 2044 40870 2100 40908
rect 2044 40514 2100 40526
rect 2044 40462 2046 40514
rect 2098 40462 2100 40514
rect 2044 40404 2100 40462
rect 2044 40338 2100 40348
rect 2044 39844 2100 39854
rect 1932 39788 2044 39844
rect 2044 39778 2100 39788
rect 1820 39618 1988 39620
rect 1820 39566 1822 39618
rect 1874 39566 1988 39618
rect 1820 39564 1988 39566
rect 1820 39554 1876 39564
rect 1820 39060 1876 39070
rect 1708 39004 1820 39060
rect 1820 38994 1876 39004
rect 1596 38892 1764 38948
rect 1708 38836 1764 38892
rect 1820 38836 1876 38846
rect 1708 38834 1876 38836
rect 1708 38782 1822 38834
rect 1874 38782 1876 38834
rect 1708 38780 1876 38782
rect 1820 38770 1876 38780
rect 1820 37268 1876 37278
rect 1932 37268 1988 39564
rect 1820 37266 1988 37268
rect 1820 37214 1822 37266
rect 1874 37214 1988 37266
rect 1820 37212 1988 37214
rect 1820 37202 1876 37212
rect 1708 37044 1764 37054
rect 1708 36482 1764 36988
rect 1708 36430 1710 36482
rect 1762 36430 1764 36482
rect 1708 36418 1764 36430
rect 1820 35586 1876 35598
rect 1820 35534 1822 35586
rect 1874 35534 1876 35586
rect 1708 34804 1764 34814
rect 1820 34804 1876 35534
rect 1708 34802 1876 34804
rect 1708 34750 1710 34802
rect 1762 34750 1876 34802
rect 1708 34748 1876 34750
rect 1932 35252 1988 37212
rect 2044 36260 2100 36270
rect 2044 36166 2100 36204
rect 1708 34356 1764 34748
rect 1708 34290 1764 34300
rect 1820 34132 1876 34142
rect 1932 34132 1988 35196
rect 1820 34130 1988 34132
rect 1820 34078 1822 34130
rect 1874 34078 1988 34130
rect 1820 34076 1988 34078
rect 2044 34690 2100 34702
rect 2044 34638 2046 34690
rect 2098 34638 2100 34690
rect 1820 34066 1876 34076
rect 2044 33348 2100 34638
rect 2044 33282 2100 33292
rect 1820 32450 1876 32462
rect 1820 32398 1822 32450
rect 1874 32398 1876 32450
rect 1708 31668 1764 31678
rect 1820 31668 1876 32398
rect 2156 31892 2212 41132
rect 2380 40962 2436 40974
rect 2380 40910 2382 40962
rect 2434 40910 2436 40962
rect 2380 40852 2436 40910
rect 2380 40786 2436 40796
rect 2492 40516 2548 40526
rect 2492 40402 2548 40460
rect 2492 40350 2494 40402
rect 2546 40350 2548 40402
rect 2492 40338 2548 40350
rect 2604 40178 2660 43374
rect 2940 42308 2996 43820
rect 3164 43652 3220 43662
rect 2716 42252 2996 42308
rect 2716 41972 2772 42252
rect 2716 41878 2772 41916
rect 2716 41746 2772 41758
rect 2716 41694 2718 41746
rect 2770 41694 2772 41746
rect 2716 41410 2772 41694
rect 2716 41358 2718 41410
rect 2770 41358 2772 41410
rect 2716 41346 2772 41358
rect 2828 40962 2884 40974
rect 2828 40910 2830 40962
rect 2882 40910 2884 40962
rect 2604 40126 2606 40178
rect 2658 40126 2660 40178
rect 2604 40114 2660 40126
rect 2716 40626 2772 40638
rect 2716 40574 2718 40626
rect 2770 40574 2772 40626
rect 2492 39732 2548 39742
rect 2716 39732 2772 40574
rect 2828 40404 2884 40910
rect 2940 40628 2996 42252
rect 3052 43540 3108 43550
rect 3052 42082 3108 43484
rect 3052 42030 3054 42082
rect 3106 42030 3108 42082
rect 3052 42018 3108 42030
rect 3052 41412 3108 41422
rect 3164 41412 3220 43596
rect 3276 42082 3332 45052
rect 3500 45106 3668 45108
rect 3500 45054 3502 45106
rect 3554 45054 3668 45106
rect 3500 45052 3668 45054
rect 3500 45042 3556 45052
rect 3388 44996 3444 45006
rect 3388 44902 3444 44940
rect 3724 44772 3780 49420
rect 4284 49252 4340 49980
rect 4172 49196 4340 49252
rect 4396 49252 4452 50204
rect 4620 49810 4676 49822
rect 4620 49758 4622 49810
rect 4674 49758 4676 49810
rect 4620 49588 4676 49758
rect 5068 49700 5124 51660
rect 5628 51602 5684 51996
rect 5628 51550 5630 51602
rect 5682 51550 5684 51602
rect 5628 51538 5684 51550
rect 5180 51492 5236 51502
rect 5180 51398 5236 51436
rect 5740 51380 5796 52444
rect 5964 52386 6020 52398
rect 5964 52334 5966 52386
rect 6018 52334 6020 52386
rect 5852 52276 5908 52286
rect 5852 52182 5908 52220
rect 5964 51604 6020 52334
rect 6524 52386 6580 58772
rect 6636 57876 6692 57886
rect 6692 57820 6804 57876
rect 6636 57810 6692 57820
rect 6636 57650 6692 57662
rect 6636 57598 6638 57650
rect 6690 57598 6692 57650
rect 6636 55972 6692 57598
rect 6636 55906 6692 55916
rect 6748 56196 6804 57820
rect 6860 57426 6916 57438
rect 6860 57374 6862 57426
rect 6914 57374 6916 57426
rect 6860 56868 6916 57374
rect 6860 56774 6916 56812
rect 6636 55412 6692 55422
rect 6748 55412 6804 56140
rect 6636 55410 6916 55412
rect 6636 55358 6638 55410
rect 6690 55358 6916 55410
rect 6636 55356 6916 55358
rect 6636 55346 6692 55356
rect 6636 54404 6692 54414
rect 6860 54404 6916 55356
rect 6972 54628 7028 59388
rect 7308 59220 7364 59230
rect 7420 59220 7476 59388
rect 7308 59218 7476 59220
rect 7308 59166 7310 59218
rect 7362 59166 7476 59218
rect 7308 59164 7476 59166
rect 7308 59154 7364 59164
rect 7084 58996 7140 59006
rect 7420 58996 7476 59006
rect 7084 58994 7476 58996
rect 7084 58942 7086 58994
rect 7138 58942 7422 58994
rect 7474 58942 7476 58994
rect 7084 58940 7476 58942
rect 7084 58930 7140 58940
rect 7420 58930 7476 58940
rect 7532 58212 7588 60510
rect 7644 60674 7700 60686
rect 7644 60622 7646 60674
rect 7698 60622 7700 60674
rect 7644 58994 7700 60622
rect 7756 59892 7812 61404
rect 8016 61180 8280 61190
rect 8072 61124 8120 61180
rect 8176 61124 8224 61180
rect 8016 61114 8280 61124
rect 7868 60786 7924 60798
rect 7868 60734 7870 60786
rect 7922 60734 7924 60786
rect 7868 60116 7924 60734
rect 8316 60788 8372 60798
rect 8316 60694 8372 60732
rect 7868 60050 7924 60060
rect 8428 60228 8484 62524
rect 7756 59836 7924 59892
rect 7644 58942 7646 58994
rect 7698 58942 7700 58994
rect 7644 58930 7700 58942
rect 7756 59220 7812 59230
rect 7756 58548 7812 59164
rect 7084 58156 7532 58212
rect 7084 57876 7140 58156
rect 7532 58146 7588 58156
rect 7644 58492 7756 58548
rect 7084 57782 7140 57820
rect 7532 57876 7588 57886
rect 7644 57876 7700 58492
rect 7756 58482 7812 58492
rect 7532 57874 7700 57876
rect 7532 57822 7534 57874
rect 7586 57822 7700 57874
rect 7532 57820 7700 57822
rect 7196 57426 7252 57438
rect 7196 57374 7198 57426
rect 7250 57374 7252 57426
rect 7196 55410 7252 57374
rect 7532 57316 7588 57820
rect 7532 57250 7588 57260
rect 7532 56756 7588 56766
rect 7532 56662 7588 56700
rect 7420 55972 7476 55982
rect 7420 55878 7476 55916
rect 7196 55358 7198 55410
rect 7250 55358 7252 55410
rect 7196 55346 7252 55358
rect 7756 55412 7812 55422
rect 7644 55074 7700 55086
rect 7644 55022 7646 55074
rect 7698 55022 7700 55074
rect 6972 54572 7252 54628
rect 6972 54404 7028 54414
rect 6636 54402 6804 54404
rect 6636 54350 6638 54402
rect 6690 54350 6804 54402
rect 6636 54348 6804 54350
rect 6860 54402 7028 54404
rect 6860 54350 6974 54402
rect 7026 54350 7028 54402
rect 6860 54348 7028 54350
rect 6636 54338 6692 54348
rect 6636 53844 6692 53854
rect 6636 52946 6692 53788
rect 6748 53620 6804 54348
rect 6972 54338 7028 54348
rect 7084 54402 7140 54414
rect 7084 54350 7086 54402
rect 7138 54350 7140 54402
rect 6748 53554 6804 53564
rect 6636 52894 6638 52946
rect 6690 52894 6692 52946
rect 6636 52882 6692 52894
rect 7084 52836 7140 54350
rect 6972 52780 7140 52836
rect 6636 52724 6692 52734
rect 6972 52724 7028 52780
rect 6636 52722 7028 52724
rect 6636 52670 6638 52722
rect 6690 52670 7028 52722
rect 6636 52668 7028 52670
rect 6636 52658 6692 52668
rect 6524 52334 6526 52386
rect 6578 52334 6580 52386
rect 6524 52322 6580 52334
rect 6748 52500 6804 52510
rect 6748 52274 6804 52444
rect 6748 52222 6750 52274
rect 6802 52222 6804 52274
rect 6748 52210 6804 52222
rect 7084 52276 7140 52286
rect 7084 52182 7140 52220
rect 6188 52052 6244 52062
rect 6188 51958 6244 51996
rect 5852 51492 5908 51502
rect 5964 51492 6020 51548
rect 5852 51490 6020 51492
rect 5852 51438 5854 51490
rect 5906 51438 6020 51490
rect 5852 51436 6020 51438
rect 5852 51426 5908 51436
rect 5516 51324 5796 51380
rect 6188 51378 6244 51390
rect 6188 51326 6190 51378
rect 6242 51326 6244 51378
rect 5404 51268 5460 51278
rect 5180 50708 5236 50718
rect 5180 50614 5236 50652
rect 5292 49924 5348 49934
rect 5404 49924 5460 51212
rect 5292 49922 5460 49924
rect 5292 49870 5294 49922
rect 5346 49870 5460 49922
rect 5292 49868 5460 49870
rect 5292 49858 5348 49868
rect 5068 49644 5236 49700
rect 4620 49522 4676 49532
rect 4614 49420 4878 49430
rect 4670 49364 4718 49420
rect 4774 49364 4822 49420
rect 4614 49354 4878 49364
rect 3948 49028 4004 49066
rect 4172 49028 4228 49196
rect 4396 49186 4452 49196
rect 5068 49252 5124 49262
rect 4396 49028 4452 49038
rect 4172 48972 4340 49028
rect 3948 48962 4004 48972
rect 4060 48802 4116 48814
rect 4060 48750 4062 48802
rect 4114 48750 4116 48802
rect 3724 44706 3780 44716
rect 3836 48580 3892 48590
rect 3836 44660 3892 48524
rect 4060 47684 4116 48750
rect 4172 48804 4228 48814
rect 4172 48710 4228 48748
rect 4060 47618 4116 47628
rect 4172 48468 4228 48478
rect 3836 44594 3892 44604
rect 3948 47572 4004 47582
rect 3948 44548 4004 47516
rect 4060 46900 4116 46910
rect 4060 45444 4116 46844
rect 4060 45378 4116 45388
rect 4172 45108 4228 48412
rect 4284 47570 4340 48972
rect 4284 47518 4286 47570
rect 4338 47518 4340 47570
rect 4284 47348 4340 47518
rect 4284 47282 4340 47292
rect 3948 44482 4004 44492
rect 4060 45052 4228 45108
rect 4284 46452 4340 46462
rect 4284 45330 4340 46396
rect 4284 45278 4286 45330
rect 4338 45278 4340 45330
rect 3724 44436 3780 44446
rect 3724 44342 3780 44380
rect 3388 44212 3444 44222
rect 3388 44118 3444 44156
rect 3836 44100 3892 44110
rect 3836 43428 3892 44044
rect 3836 43362 3892 43372
rect 3276 42030 3278 42082
rect 3330 42030 3332 42082
rect 3276 41748 3332 42030
rect 3724 41972 3780 41982
rect 3780 41916 3892 41972
rect 3724 41878 3780 41916
rect 3388 41748 3444 41758
rect 3276 41692 3388 41748
rect 3276 41682 3444 41692
rect 3276 41580 3388 41682
rect 3276 41412 3332 41422
rect 3052 41410 3332 41412
rect 3052 41358 3054 41410
rect 3106 41358 3278 41410
rect 3330 41358 3332 41410
rect 3052 41356 3332 41358
rect 3052 40964 3108 41356
rect 3276 41346 3332 41356
rect 3052 40898 3108 40908
rect 3500 41300 3556 41310
rect 3500 40962 3556 41244
rect 3836 41188 3892 41916
rect 3836 41122 3892 41132
rect 3948 41410 4004 41422
rect 3948 41358 3950 41410
rect 4002 41358 4004 41410
rect 3948 41298 4004 41358
rect 3948 41246 3950 41298
rect 4002 41246 4004 41298
rect 3500 40910 3502 40962
rect 3554 40910 3556 40962
rect 2940 40562 2996 40572
rect 3164 40852 3220 40862
rect 3164 40514 3220 40796
rect 3500 40852 3556 40910
rect 3500 40786 3556 40796
rect 3164 40462 3166 40514
rect 3218 40462 3220 40514
rect 2828 40338 2884 40348
rect 2940 40402 2996 40414
rect 2940 40350 2942 40402
rect 2994 40350 2996 40402
rect 2492 39730 2772 39732
rect 2492 39678 2494 39730
rect 2546 39678 2772 39730
rect 2492 39676 2772 39678
rect 2492 39666 2548 39676
rect 2940 39508 2996 40350
rect 3164 40068 3220 40462
rect 3612 40404 3668 40414
rect 3612 40310 3668 40348
rect 3724 40180 3780 40190
rect 3724 40086 3780 40124
rect 3948 40068 4004 41246
rect 4060 40180 4116 45052
rect 4284 44436 4340 45278
rect 4172 44380 4340 44436
rect 4172 43652 4228 44380
rect 4396 44324 4452 48972
rect 4620 48804 4676 48814
rect 4620 48130 4676 48748
rect 4956 48804 5012 48814
rect 5068 48804 5124 49196
rect 4956 48802 5124 48804
rect 4956 48750 4958 48802
rect 5010 48750 5124 48802
rect 4956 48748 5124 48750
rect 4956 48738 5012 48748
rect 4620 48078 4622 48130
rect 4674 48078 4676 48130
rect 4620 48020 4676 48078
rect 4620 47954 4676 47964
rect 4956 48356 5012 48366
rect 4956 48018 5012 48300
rect 4956 47966 4958 48018
rect 5010 47966 5012 48018
rect 4956 47908 5012 47966
rect 4614 47852 4878 47862
rect 4670 47796 4718 47852
rect 4774 47796 4822 47852
rect 4956 47842 5012 47852
rect 4614 47786 4878 47796
rect 5068 47684 5124 48748
rect 4844 47628 5124 47684
rect 4732 47572 4788 47582
rect 4732 47478 4788 47516
rect 4508 47460 4564 47470
rect 4508 46564 4564 47404
rect 4844 47068 4900 47628
rect 4844 47002 4900 47012
rect 4956 47460 5012 47470
rect 4508 46470 4564 46508
rect 4844 46788 4900 46798
rect 4956 46788 5012 47404
rect 5068 47236 5124 47246
rect 5068 46898 5124 47180
rect 5068 46846 5070 46898
rect 5122 46846 5124 46898
rect 5068 46834 5124 46846
rect 4844 46786 5012 46788
rect 4844 46734 4846 46786
rect 4898 46734 5012 46786
rect 4844 46732 5012 46734
rect 5180 46788 5236 49644
rect 5292 49140 5348 49150
rect 5292 48242 5348 49084
rect 5292 48190 5294 48242
rect 5346 48190 5348 48242
rect 5292 48178 5348 48190
rect 5516 48132 5572 51324
rect 5964 51268 6020 51278
rect 5964 51174 6020 51212
rect 6188 51268 6244 51326
rect 6412 51380 6468 51390
rect 6412 51378 6580 51380
rect 6412 51326 6414 51378
rect 6466 51326 6580 51378
rect 6412 51324 6580 51326
rect 6412 51314 6468 51324
rect 6188 51202 6244 51212
rect 6412 51156 6468 51166
rect 5628 51044 5684 51054
rect 5628 50428 5684 50988
rect 5964 50932 6020 50942
rect 5628 50372 5908 50428
rect 5628 49924 5684 49934
rect 5628 49140 5684 49868
rect 5628 49046 5684 49084
rect 5740 48804 5796 48814
rect 5740 48710 5796 48748
rect 5852 48580 5908 50372
rect 5852 48514 5908 48524
rect 5852 48356 5908 48366
rect 5852 48262 5908 48300
rect 5516 48076 5908 48132
rect 5292 48018 5348 48030
rect 5292 47966 5294 48018
rect 5346 47966 5348 48018
rect 5292 47908 5348 47966
rect 5292 47852 5684 47908
rect 5516 47684 5572 47694
rect 5516 47068 5572 47628
rect 4844 46452 4900 46732
rect 5180 46722 5236 46732
rect 5404 47012 5572 47068
rect 5404 46676 5460 47012
rect 5404 46610 5460 46620
rect 5516 46900 5572 46910
rect 5516 46674 5572 46844
rect 5516 46622 5518 46674
rect 5570 46622 5572 46674
rect 5516 46610 5572 46622
rect 4844 46386 4900 46396
rect 5180 46452 5236 46462
rect 5180 46450 5572 46452
rect 5180 46398 5182 46450
rect 5234 46398 5572 46450
rect 5180 46396 5572 46398
rect 5180 46386 5236 46396
rect 4614 46284 4878 46294
rect 4670 46228 4718 46284
rect 4774 46228 4822 46284
rect 4614 46218 4878 46228
rect 4620 46002 4676 46014
rect 4620 45950 4622 46002
rect 4674 45950 4676 46002
rect 4620 45220 4676 45950
rect 5180 45668 5236 45706
rect 5180 45602 5236 45612
rect 5180 45444 5236 45454
rect 5180 45332 5236 45388
rect 5180 45330 5348 45332
rect 5180 45278 5182 45330
rect 5234 45278 5348 45330
rect 5180 45276 5348 45278
rect 5180 45266 5236 45276
rect 4620 45154 4676 45164
rect 4844 44996 4900 45006
rect 4844 44902 4900 44940
rect 4614 44716 4878 44726
rect 4670 44660 4718 44716
rect 4774 44660 4822 44716
rect 4614 44650 4878 44660
rect 4172 43586 4228 43596
rect 4284 44268 4452 44324
rect 4284 42084 4340 44268
rect 4508 44210 4564 44222
rect 4508 44158 4510 44210
rect 4562 44158 4564 44210
rect 4396 44098 4452 44110
rect 4396 44046 4398 44098
rect 4450 44046 4452 44098
rect 4396 43540 4452 44046
rect 4396 43474 4452 43484
rect 4508 43316 4564 44158
rect 5180 44100 5236 44138
rect 5180 44034 5236 44044
rect 5292 43652 5348 45276
rect 5404 43652 5460 43662
rect 5068 43650 5460 43652
rect 5068 43598 5406 43650
rect 5458 43598 5460 43650
rect 5068 43596 5460 43598
rect 4844 43540 4900 43550
rect 4844 43538 5012 43540
rect 4844 43486 4846 43538
rect 4898 43486 5012 43538
rect 4844 43484 5012 43486
rect 4844 43474 4900 43484
rect 4396 43260 4564 43316
rect 4396 42868 4452 43260
rect 4614 43148 4878 43158
rect 4670 43092 4718 43148
rect 4774 43092 4822 43148
rect 4614 43082 4878 43092
rect 4620 42868 4676 42878
rect 4396 42866 4676 42868
rect 4396 42814 4622 42866
rect 4674 42814 4676 42866
rect 4396 42812 4676 42814
rect 4620 42644 4676 42812
rect 4956 42868 5012 43484
rect 4956 42802 5012 42812
rect 5068 42866 5124 43596
rect 5404 43586 5460 43596
rect 5068 42814 5070 42866
rect 5122 42814 5124 42866
rect 4620 42578 4676 42588
rect 4844 42084 4900 42094
rect 4284 42028 4452 42084
rect 4172 41972 4228 41982
rect 4228 41916 4340 41972
rect 4172 41878 4228 41916
rect 4284 40628 4340 41916
rect 4396 41188 4452 42028
rect 4844 41970 4900 42028
rect 5068 41972 5124 42814
rect 5516 42532 5572 46396
rect 5628 44436 5684 47852
rect 5740 47458 5796 47470
rect 5740 47406 5742 47458
rect 5794 47406 5796 47458
rect 5740 47236 5796 47406
rect 5740 47170 5796 47180
rect 5852 47234 5908 48076
rect 5852 47182 5854 47234
rect 5906 47182 5908 47234
rect 5852 47124 5908 47182
rect 5852 47058 5908 47068
rect 5852 46900 5908 46910
rect 5740 45332 5796 45342
rect 5740 45238 5796 45276
rect 5852 44884 5908 46844
rect 5964 45108 6020 50876
rect 6188 50596 6244 50606
rect 6188 50502 6244 50540
rect 6412 50594 6468 51100
rect 6524 50706 6580 51324
rect 7196 51156 7252 54572
rect 7308 54514 7364 54526
rect 7308 54462 7310 54514
rect 7362 54462 7364 54514
rect 7308 53844 7364 54462
rect 7308 53778 7364 53788
rect 7644 53508 7700 55022
rect 7644 53442 7700 53452
rect 7644 52834 7700 52846
rect 7644 52782 7646 52834
rect 7698 52782 7700 52834
rect 7644 52612 7700 52782
rect 7308 52556 7644 52612
rect 7308 51602 7364 52556
rect 7644 52546 7700 52556
rect 7532 52388 7588 52398
rect 7532 52162 7588 52332
rect 7532 52110 7534 52162
rect 7586 52110 7588 52162
rect 7532 52098 7588 52110
rect 7756 51828 7812 55356
rect 7308 51550 7310 51602
rect 7362 51550 7364 51602
rect 7308 51538 7364 51550
rect 7644 51772 7812 51828
rect 7196 51090 7252 51100
rect 7644 50820 7700 51772
rect 7756 51604 7812 51614
rect 7756 51510 7812 51548
rect 7868 51044 7924 59836
rect 8016 59612 8280 59622
rect 8072 59556 8120 59612
rect 8176 59556 8224 59612
rect 8016 59546 8280 59556
rect 8016 58044 8280 58054
rect 8072 57988 8120 58044
rect 8176 57988 8224 58044
rect 8016 57978 8280 57988
rect 8092 57876 8148 57886
rect 8428 57876 8484 60172
rect 8540 60116 8596 60126
rect 8540 59444 8596 60060
rect 8540 59378 8596 59388
rect 8652 57988 8708 68012
rect 8876 67060 8932 67070
rect 8764 67058 8932 67060
rect 8764 67006 8878 67058
rect 8930 67006 8932 67058
rect 8764 67004 8932 67006
rect 8764 66946 8820 67004
rect 8876 66994 8932 67004
rect 8764 66894 8766 66946
rect 8818 66894 8820 66946
rect 8764 66882 8820 66894
rect 8876 66836 8932 66846
rect 8764 65380 8820 65390
rect 8876 65380 8932 66780
rect 8764 65378 8932 65380
rect 8764 65326 8766 65378
rect 8818 65326 8932 65378
rect 8764 65324 8932 65326
rect 8764 65314 8820 65324
rect 8876 63812 8932 65324
rect 8988 66500 9044 66510
rect 8988 64820 9044 66444
rect 8988 64726 9044 64764
rect 9212 64372 9268 68012
rect 9548 66500 9604 68574
rect 9660 67844 9716 70702
rect 9772 70644 9828 71710
rect 9772 70578 9828 70588
rect 9772 70420 9828 70430
rect 9772 70326 9828 70364
rect 9660 67778 9716 67788
rect 9660 67620 9716 67630
rect 9660 67526 9716 67564
rect 9660 66948 9716 66958
rect 9660 66854 9716 66892
rect 9548 66386 9604 66444
rect 9548 66334 9550 66386
rect 9602 66334 9604 66386
rect 9548 66322 9604 66334
rect 9884 65716 9940 73724
rect 9996 72324 10052 74060
rect 10108 75010 10500 75012
rect 10108 74958 10222 75010
rect 10274 74958 10500 75010
rect 10108 74956 10500 74958
rect 10108 74338 10164 74956
rect 10220 74946 10276 74956
rect 10332 74788 10388 74798
rect 10108 74286 10110 74338
rect 10162 74286 10164 74338
rect 10108 73554 10164 74286
rect 10108 73502 10110 73554
rect 10162 73502 10164 73554
rect 10108 72660 10164 73502
rect 10108 72594 10164 72604
rect 10220 74786 10388 74788
rect 10220 74734 10334 74786
rect 10386 74734 10388 74786
rect 10220 74732 10388 74734
rect 9996 71204 10052 72268
rect 10108 72434 10164 72446
rect 10108 72382 10110 72434
rect 10162 72382 10164 72434
rect 10108 71988 10164 72382
rect 10108 71922 10164 71932
rect 10220 71762 10276 74732
rect 10332 74722 10388 74732
rect 10444 74226 10500 74956
rect 10444 74174 10446 74226
rect 10498 74174 10500 74226
rect 10444 74162 10500 74174
rect 10556 73948 10612 76636
rect 10668 76468 10724 76478
rect 10668 76466 10836 76468
rect 10668 76414 10670 76466
rect 10722 76414 10836 76466
rect 10668 76412 10836 76414
rect 10668 76402 10724 76412
rect 10780 75348 10836 76412
rect 10892 75572 10948 85652
rect 12012 85586 12068 85596
rect 12124 86434 12180 86446
rect 12124 86382 12126 86434
rect 12178 86382 12180 86434
rect 11418 85484 11682 85494
rect 11474 85428 11522 85484
rect 11578 85428 11626 85484
rect 11418 85418 11682 85428
rect 11452 84978 11508 84990
rect 12124 84980 12180 86382
rect 11452 84926 11454 84978
rect 11506 84926 11508 84978
rect 11452 84420 11508 84926
rect 11452 84354 11508 84364
rect 11788 84924 12180 84980
rect 11788 84418 11844 84924
rect 12348 84868 12404 88060
rect 11788 84366 11790 84418
rect 11842 84366 11844 84418
rect 11788 84354 11844 84366
rect 11900 84812 12404 84868
rect 11116 84308 11172 84318
rect 11116 84214 11172 84252
rect 11418 83916 11682 83926
rect 11474 83860 11522 83916
rect 11578 83860 11626 83916
rect 11418 83850 11682 83860
rect 11564 83300 11620 83310
rect 11228 83076 11284 83086
rect 11116 82964 11172 82974
rect 11116 82870 11172 82908
rect 11228 82962 11284 83020
rect 11228 82910 11230 82962
rect 11282 82910 11284 82962
rect 11228 82898 11284 82910
rect 11564 82962 11620 83244
rect 11564 82910 11566 82962
rect 11618 82910 11620 82962
rect 11564 82898 11620 82910
rect 11340 82740 11396 82750
rect 11116 82738 11396 82740
rect 11116 82686 11342 82738
rect 11394 82686 11396 82738
rect 11116 82684 11396 82686
rect 11116 82404 11172 82684
rect 11340 82674 11396 82684
rect 11116 82348 11284 82404
rect 11228 82178 11284 82348
rect 11418 82348 11682 82358
rect 11474 82292 11522 82348
rect 11578 82292 11626 82348
rect 11418 82282 11682 82292
rect 11228 82126 11230 82178
rect 11282 82126 11284 82178
rect 11116 81732 11172 81742
rect 11004 81730 11172 81732
rect 11004 81678 11118 81730
rect 11170 81678 11172 81730
rect 11004 81676 11172 81678
rect 11004 81620 11060 81676
rect 11116 81666 11172 81676
rect 11004 80946 11060 81564
rect 11228 81284 11284 82126
rect 11564 81732 11620 81742
rect 11564 81396 11620 81676
rect 11900 81396 11956 84812
rect 12348 83634 12404 83646
rect 12348 83582 12350 83634
rect 12402 83582 12404 83634
rect 12348 82738 12404 83582
rect 12348 82686 12350 82738
rect 12402 82686 12404 82738
rect 12348 82674 12404 82686
rect 12124 82516 12180 82526
rect 11564 81330 11620 81340
rect 11788 81394 11956 81396
rect 11788 81342 11902 81394
rect 11954 81342 11956 81394
rect 11788 81340 11956 81342
rect 11340 81284 11396 81294
rect 11228 81228 11340 81284
rect 11340 81218 11396 81228
rect 11004 80894 11006 80946
rect 11058 80894 11060 80946
rect 11004 78932 11060 80894
rect 11116 80948 11172 80958
rect 11116 80854 11172 80892
rect 11418 80780 11682 80790
rect 11474 80724 11522 80780
rect 11578 80724 11626 80780
rect 11418 80714 11682 80724
rect 11676 79604 11732 79614
rect 11788 79604 11844 81340
rect 11900 81330 11956 81340
rect 12012 81730 12068 81742
rect 12012 81678 12014 81730
rect 12066 81678 12068 81730
rect 11732 79548 11844 79604
rect 12012 79604 12068 81678
rect 11676 79510 11732 79548
rect 12012 79538 12068 79548
rect 12012 79380 12068 79390
rect 11418 79212 11682 79222
rect 11474 79156 11522 79212
rect 11578 79156 11626 79212
rect 11418 79146 11682 79156
rect 11004 78866 11060 78876
rect 11228 78930 11284 78942
rect 11228 78878 11230 78930
rect 11282 78878 11284 78930
rect 11004 78708 11060 78718
rect 11004 78258 11060 78652
rect 11004 78206 11006 78258
rect 11058 78206 11060 78258
rect 11004 78194 11060 78206
rect 11228 77028 11284 78878
rect 12012 78930 12068 79324
rect 12012 78878 12014 78930
rect 12066 78878 12068 78930
rect 11418 77644 11682 77654
rect 11474 77588 11522 77644
rect 11578 77588 11626 77644
rect 11418 77578 11682 77588
rect 11116 76692 11172 76702
rect 11116 76598 11172 76636
rect 11228 76690 11284 76972
rect 11228 76638 11230 76690
rect 11282 76638 11284 76690
rect 11228 76626 11284 76638
rect 11900 77140 11956 77150
rect 11900 76690 11956 77084
rect 11900 76638 11902 76690
rect 11954 76638 11956 76690
rect 11900 76626 11956 76638
rect 11788 76468 11844 76478
rect 11004 76244 11060 76254
rect 11004 76150 11060 76188
rect 11418 76076 11682 76086
rect 11474 76020 11522 76076
rect 11578 76020 11626 76076
rect 11418 76010 11682 76020
rect 11788 75908 11844 76412
rect 11676 75852 11844 75908
rect 11004 75572 11060 75582
rect 10892 75516 11004 75572
rect 11004 75506 11060 75516
rect 10780 75292 11396 75348
rect 11004 75124 11060 75134
rect 11228 75124 11284 75134
rect 11004 75122 11228 75124
rect 11004 75070 11006 75122
rect 11058 75070 11228 75122
rect 11004 75068 11228 75070
rect 11004 75058 11060 75068
rect 11228 75030 11284 75068
rect 11340 75122 11396 75292
rect 11340 75070 11342 75122
rect 11394 75070 11396 75122
rect 11340 75058 11396 75070
rect 11452 74900 11508 74910
rect 11452 74806 11508 74844
rect 11676 74676 11732 75852
rect 11900 75794 11956 75806
rect 11900 75742 11902 75794
rect 11954 75742 11956 75794
rect 11228 74620 11732 74676
rect 11788 74898 11844 74910
rect 11788 74846 11790 74898
rect 11842 74846 11844 74898
rect 10892 74002 10948 74014
rect 10892 73950 10894 74002
rect 10946 73950 10948 74002
rect 10556 73892 10724 73948
rect 10220 71710 10222 71762
rect 10274 71710 10276 71762
rect 10220 71698 10276 71710
rect 10444 72212 10500 72222
rect 10444 71874 10500 72156
rect 10556 71988 10612 71998
rect 10556 71894 10612 71932
rect 10444 71822 10446 71874
rect 10498 71822 10500 71874
rect 9996 71148 10164 71204
rect 9996 70978 10052 70990
rect 9996 70926 9998 70978
rect 10050 70926 10052 70978
rect 9996 70420 10052 70926
rect 9996 70354 10052 70364
rect 9996 70196 10052 70206
rect 10108 70196 10164 71148
rect 10444 70980 10500 71822
rect 10668 71204 10724 73892
rect 10892 73556 10948 73950
rect 10668 71138 10724 71148
rect 10780 71764 10836 71774
rect 10780 70980 10836 71708
rect 10444 70914 10500 70924
rect 10668 70924 10836 70980
rect 10444 70756 10500 70766
rect 10668 70756 10724 70924
rect 10444 70754 10724 70756
rect 10444 70702 10446 70754
rect 10498 70702 10724 70754
rect 10444 70700 10724 70702
rect 10780 70756 10836 70766
rect 10444 70644 10500 70700
rect 10444 70578 10500 70588
rect 10220 70420 10276 70430
rect 10668 70420 10724 70430
rect 10220 70326 10276 70364
rect 10332 70364 10668 70420
rect 9996 70194 10164 70196
rect 9996 70142 9998 70194
rect 10050 70142 10164 70194
rect 9996 70140 10164 70142
rect 10220 70196 10276 70206
rect 10332 70196 10388 70364
rect 10668 70354 10724 70364
rect 10220 70194 10388 70196
rect 10220 70142 10222 70194
rect 10274 70142 10388 70194
rect 10220 70140 10388 70142
rect 9996 69188 10052 70140
rect 10220 70130 10276 70140
rect 9996 69122 10052 69132
rect 10444 69188 10500 69198
rect 10444 69094 10500 69132
rect 10332 68516 10388 68526
rect 10332 68514 10500 68516
rect 10332 68462 10334 68514
rect 10386 68462 10500 68514
rect 10332 68460 10500 68462
rect 10332 68450 10388 68460
rect 10444 67954 10500 68460
rect 10444 67902 10446 67954
rect 10498 67902 10500 67954
rect 10444 67890 10500 67902
rect 10220 67842 10276 67854
rect 10220 67790 10222 67842
rect 10274 67790 10276 67842
rect 9996 67620 10052 67630
rect 10220 67620 10276 67790
rect 10668 67732 10724 67742
rect 10668 67638 10724 67676
rect 9996 67618 10276 67620
rect 9996 67566 9998 67618
rect 10050 67566 10276 67618
rect 9996 67564 10276 67566
rect 9996 67554 10052 67564
rect 9212 64306 9268 64316
rect 9324 65660 9940 65716
rect 8876 63718 8932 63756
rect 8988 63924 9044 63934
rect 8764 62804 8820 62814
rect 8764 62578 8820 62748
rect 8764 62526 8766 62578
rect 8818 62526 8820 62578
rect 8764 62356 8820 62526
rect 8764 62290 8820 62300
rect 8988 61572 9044 63868
rect 8988 61570 9156 61572
rect 8988 61518 8990 61570
rect 9042 61518 9156 61570
rect 8988 61516 9156 61518
rect 8988 61506 9044 61516
rect 8988 60788 9044 60798
rect 8988 60676 9044 60732
rect 8876 60674 9044 60676
rect 8876 60622 8990 60674
rect 9042 60622 9044 60674
rect 8876 60620 9044 60622
rect 8876 58324 8932 60620
rect 8988 60610 9044 60620
rect 8988 60228 9044 60238
rect 8988 60114 9044 60172
rect 8988 60062 8990 60114
rect 9042 60062 9044 60114
rect 8988 60050 9044 60062
rect 9100 59332 9156 61516
rect 9100 59266 9156 59276
rect 8876 58258 8932 58268
rect 9100 58436 9156 58446
rect 8988 57988 9044 57998
rect 8652 57932 8988 57988
rect 8092 57874 8484 57876
rect 8092 57822 8094 57874
rect 8146 57822 8484 57874
rect 8092 57820 8484 57822
rect 8540 57876 8596 57886
rect 8092 57426 8148 57820
rect 8540 57782 8596 57820
rect 8988 57874 9044 57932
rect 8988 57822 8990 57874
rect 9042 57822 9044 57874
rect 8988 57810 9044 57822
rect 8092 57374 8094 57426
rect 8146 57374 8148 57426
rect 8092 57362 8148 57374
rect 8428 56756 8484 56766
rect 8016 56476 8280 56486
rect 8072 56420 8120 56476
rect 8176 56420 8224 56476
rect 8016 56410 8280 56420
rect 8428 56306 8484 56700
rect 8428 56254 8430 56306
rect 8482 56254 8484 56306
rect 8428 56242 8484 56254
rect 8652 56420 8708 56430
rect 8652 56194 8708 56364
rect 8988 56308 9044 56318
rect 8652 56142 8654 56194
rect 8706 56142 8708 56194
rect 8316 56084 8372 56094
rect 8316 56082 8484 56084
rect 8316 56030 8318 56082
rect 8370 56030 8484 56082
rect 8316 56028 8484 56030
rect 8316 56018 8372 56028
rect 8092 55970 8148 55982
rect 8092 55918 8094 55970
rect 8146 55918 8148 55970
rect 8092 55860 8148 55918
rect 8092 55794 8148 55804
rect 7980 55412 8036 55422
rect 7980 55318 8036 55356
rect 8428 55074 8484 56028
rect 8652 55412 8708 56142
rect 8876 56196 8932 56206
rect 8876 56102 8932 56140
rect 8652 55346 8708 55356
rect 8876 55412 8932 55422
rect 8988 55412 9044 56252
rect 8876 55410 9044 55412
rect 8876 55358 8878 55410
rect 8930 55358 9044 55410
rect 8876 55356 9044 55358
rect 8876 55346 8932 55356
rect 8428 55022 8430 55074
rect 8482 55022 8484 55074
rect 8016 54908 8280 54918
rect 8072 54852 8120 54908
rect 8176 54852 8224 54908
rect 8016 54842 8280 54852
rect 8428 54572 8484 55022
rect 8428 54516 8708 54572
rect 8204 54402 8260 54414
rect 8204 54350 8206 54402
rect 8258 54350 8260 54402
rect 8204 54180 8260 54350
rect 8540 54402 8596 54414
rect 8540 54350 8542 54402
rect 8594 54350 8596 54402
rect 8540 54292 8596 54350
rect 8204 54114 8260 54124
rect 8428 54236 8540 54292
rect 8016 53340 8280 53350
rect 8072 53284 8120 53340
rect 8176 53284 8224 53340
rect 8016 53274 8280 53284
rect 8092 52834 8148 52846
rect 8092 52782 8094 52834
rect 8146 52782 8148 52834
rect 8092 52500 8148 52782
rect 8092 52434 8148 52444
rect 8204 52722 8260 52734
rect 8204 52670 8206 52722
rect 8258 52670 8260 52722
rect 8204 52274 8260 52670
rect 8204 52222 8206 52274
rect 8258 52222 8260 52274
rect 8204 52210 8260 52222
rect 8428 52276 8484 54236
rect 8540 54226 8596 54236
rect 8428 52210 8484 52220
rect 8540 53844 8596 53854
rect 8428 52052 8484 52062
rect 8016 51772 8280 51782
rect 8072 51716 8120 51772
rect 8176 51716 8224 51772
rect 8016 51706 8280 51716
rect 8428 51378 8484 51996
rect 8540 51716 8596 53788
rect 8652 53732 8708 54516
rect 9100 54404 9156 58380
rect 9212 58324 9268 58334
rect 9212 58230 9268 58268
rect 8988 54402 9156 54404
rect 8988 54350 9102 54402
rect 9154 54350 9156 54402
rect 8988 54348 9156 54350
rect 8764 53732 8820 53742
rect 8652 53730 8820 53732
rect 8652 53678 8766 53730
rect 8818 53678 8820 53730
rect 8652 53676 8820 53678
rect 8764 53620 8820 53676
rect 8988 53732 9044 54348
rect 9100 54338 9156 54348
rect 9212 54852 9268 54862
rect 8988 53666 9044 53676
rect 9100 54068 9156 54078
rect 9212 54068 9268 54796
rect 9156 54012 9268 54068
rect 9100 53730 9156 54012
rect 9100 53678 9102 53730
rect 9154 53678 9156 53730
rect 9100 53666 9156 53678
rect 8764 53554 8820 53564
rect 8988 53506 9044 53518
rect 8988 53454 8990 53506
rect 9042 53454 9044 53506
rect 8652 53396 8708 53406
rect 8652 53170 8708 53340
rect 8652 53118 8654 53170
rect 8706 53118 8708 53170
rect 8652 53106 8708 53118
rect 8988 52722 9044 53454
rect 9100 53284 9156 53294
rect 9100 53170 9156 53228
rect 9100 53118 9102 53170
rect 9154 53118 9156 53170
rect 9100 53106 9156 53118
rect 8988 52670 8990 52722
rect 9042 52670 9044 52722
rect 8988 52658 9044 52670
rect 9212 53060 9268 53070
rect 9212 52724 9268 53004
rect 9212 52658 9268 52668
rect 8988 51828 9044 51838
rect 8764 51716 8820 51726
rect 8540 51660 8764 51716
rect 8764 51650 8820 51660
rect 8988 51602 9044 51772
rect 8988 51550 8990 51602
rect 9042 51550 9044 51602
rect 8988 51492 9044 51550
rect 8988 51426 9044 51436
rect 8428 51326 8430 51378
rect 8482 51326 8484 51378
rect 8428 51314 8484 51326
rect 8764 51380 8820 51390
rect 8764 51286 8820 51324
rect 8204 51268 8260 51278
rect 8204 51174 8260 51212
rect 8876 51266 8932 51278
rect 8876 51214 8878 51266
rect 8930 51214 8932 51266
rect 7868 50978 7924 50988
rect 8652 51044 8708 51054
rect 7196 50764 7700 50820
rect 6524 50654 6526 50706
rect 6578 50654 6580 50706
rect 6524 50642 6580 50654
rect 6860 50708 6916 50718
rect 6412 50542 6414 50594
rect 6466 50542 6468 50594
rect 6412 50428 6468 50542
rect 6636 50596 6692 50606
rect 6636 50594 6804 50596
rect 6636 50542 6638 50594
rect 6690 50542 6804 50594
rect 6636 50540 6804 50542
rect 6636 50530 6692 50540
rect 6748 50484 6804 50540
rect 6412 50372 6692 50428
rect 6748 50418 6804 50428
rect 6860 50482 6916 50652
rect 6860 50430 6862 50482
rect 6914 50430 6916 50482
rect 6860 50428 6916 50430
rect 6860 50372 7028 50428
rect 6300 50036 6356 50046
rect 6188 49588 6244 49598
rect 6188 48466 6244 49532
rect 6188 48414 6190 48466
rect 6242 48414 6244 48466
rect 6188 48402 6244 48414
rect 6300 48244 6356 49980
rect 6524 49812 6580 49822
rect 6524 49138 6580 49756
rect 6524 49086 6526 49138
rect 6578 49086 6580 49138
rect 6524 49074 6580 49086
rect 6188 48188 6356 48244
rect 6412 48804 6468 48814
rect 6076 48018 6132 48030
rect 6076 47966 6078 48018
rect 6130 47966 6132 48018
rect 6076 45666 6132 47966
rect 6076 45614 6078 45666
rect 6130 45614 6132 45666
rect 6076 45444 6132 45614
rect 6188 45556 6244 48188
rect 6300 46564 6356 46574
rect 6300 46470 6356 46508
rect 6412 46228 6468 48748
rect 6524 48580 6580 48590
rect 6524 47796 6580 48524
rect 6636 48130 6692 50372
rect 6636 48078 6638 48130
rect 6690 48078 6692 48130
rect 6636 48018 6692 48078
rect 6636 47966 6638 48018
rect 6690 47966 6692 48018
rect 6636 47954 6692 47966
rect 6748 50260 6804 50270
rect 6524 47740 6692 47796
rect 6412 46162 6468 46172
rect 6412 45780 6468 45790
rect 6412 45686 6468 45724
rect 6188 45490 6244 45500
rect 6524 45668 6580 45678
rect 6076 45378 6132 45388
rect 5964 45042 6020 45052
rect 6188 44994 6244 45006
rect 6188 44942 6190 44994
rect 6242 44942 6244 44994
rect 6188 44884 6244 44942
rect 5852 44882 6244 44884
rect 5852 44830 6190 44882
rect 6242 44830 6244 44882
rect 5852 44828 6244 44830
rect 6188 44818 6244 44828
rect 6300 44996 6356 45006
rect 6188 44548 6244 44558
rect 6188 44454 6244 44492
rect 5628 44380 6020 44436
rect 4844 41918 4846 41970
rect 4898 41918 4900 41970
rect 4844 41906 4900 41918
rect 4956 41916 5068 41972
rect 4614 41580 4878 41590
rect 4670 41524 4718 41580
rect 4774 41524 4822 41580
rect 4614 41514 4878 41524
rect 4844 41300 4900 41310
rect 4956 41300 5012 41916
rect 5068 41906 5124 41916
rect 5404 42476 5572 42532
rect 5628 44212 5684 44222
rect 4844 41298 4956 41300
rect 4844 41246 4846 41298
rect 4898 41246 4956 41298
rect 4844 41244 4956 41246
rect 4844 41234 4900 41244
rect 4956 41206 5012 41244
rect 4396 41132 4788 41188
rect 4732 41076 4788 41132
rect 4732 41020 5012 41076
rect 4284 40402 4340 40572
rect 4284 40350 4286 40402
rect 4338 40350 4340 40402
rect 4284 40338 4340 40350
rect 4396 40964 4452 40974
rect 4060 40124 4340 40180
rect 3164 40002 3220 40012
rect 3836 40012 4004 40068
rect 2940 39452 3444 39508
rect 2268 39060 2324 39070
rect 2268 38966 2324 39004
rect 3388 39058 3444 39452
rect 3388 39006 3390 39058
rect 3442 39006 3444 39058
rect 3388 38994 3444 39006
rect 3500 39060 3556 39070
rect 3500 38946 3556 39004
rect 3500 38894 3502 38946
rect 3554 38894 3556 38946
rect 3500 38882 3556 38894
rect 3612 38948 3668 38958
rect 2380 38276 2436 38286
rect 2380 38182 2436 38220
rect 2380 38052 2436 38062
rect 2380 37958 2436 37996
rect 3388 38052 3444 38062
rect 3388 37958 3444 37996
rect 2716 37940 2772 37950
rect 2940 37940 2996 37950
rect 2716 37938 2884 37940
rect 2716 37886 2718 37938
rect 2770 37886 2884 37938
rect 2716 37884 2884 37886
rect 2716 37874 2772 37884
rect 2492 37826 2548 37838
rect 2492 37774 2494 37826
rect 2546 37774 2548 37826
rect 2492 37378 2548 37774
rect 2492 37326 2494 37378
rect 2546 37326 2548 37378
rect 2492 37314 2548 37326
rect 2492 37044 2548 37054
rect 2828 37044 2884 37884
rect 2940 37846 2996 37884
rect 2828 36988 3220 37044
rect 2492 36594 2548 36988
rect 3164 36706 3220 36988
rect 3164 36654 3166 36706
rect 3218 36654 3220 36706
rect 3164 36642 3220 36654
rect 3276 36708 3332 36718
rect 2492 36542 2494 36594
rect 2546 36542 2548 36594
rect 2492 36530 2548 36542
rect 3276 36594 3332 36652
rect 3276 36542 3278 36594
rect 3330 36542 3332 36594
rect 3276 36530 3332 36542
rect 2940 35028 2996 35038
rect 2940 34934 2996 34972
rect 2828 34916 2884 34926
rect 2716 34914 2884 34916
rect 2716 34862 2830 34914
rect 2882 34862 2884 34914
rect 2716 34860 2884 34862
rect 2492 34018 2548 34030
rect 2492 33966 2494 34018
rect 2546 33966 2548 34018
rect 2380 33572 2436 33582
rect 2380 33348 2436 33516
rect 2156 31826 2212 31836
rect 2268 33346 2436 33348
rect 2268 33294 2382 33346
rect 2434 33294 2436 33346
rect 2268 33292 2436 33294
rect 1764 31612 1876 31668
rect 2044 31780 2100 31790
rect 2044 31666 2100 31724
rect 2044 31614 2046 31666
rect 2098 31614 2100 31666
rect 1708 31574 1764 31612
rect 2044 31602 2100 31614
rect 1820 30994 1876 31006
rect 1820 30942 1822 30994
rect 1874 30942 1876 30994
rect 1708 29426 1764 29438
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 28980 1764 29374
rect 1708 28644 1764 28924
rect 1708 28578 1764 28588
rect 1820 28084 1876 30942
rect 2044 30212 2100 30222
rect 2268 30212 2324 33292
rect 2380 33282 2436 33292
rect 2492 33124 2548 33966
rect 2604 33460 2660 33470
rect 2604 33366 2660 33404
rect 2716 33348 2772 34860
rect 2828 34850 2884 34860
rect 3500 34916 3556 34926
rect 3500 34822 3556 34860
rect 3388 34804 3444 34814
rect 2940 34802 3444 34804
rect 2940 34750 3390 34802
rect 3442 34750 3444 34802
rect 2940 34748 3444 34750
rect 2716 33282 2772 33292
rect 2828 33348 2884 33358
rect 2940 33348 2996 34748
rect 3388 34738 3444 34748
rect 3388 33572 3444 33582
rect 2828 33346 2996 33348
rect 2828 33294 2830 33346
rect 2882 33294 2996 33346
rect 2828 33292 2996 33294
rect 3276 33516 3388 33572
rect 2828 33282 2884 33292
rect 3052 33236 3108 33246
rect 3052 33234 3220 33236
rect 3052 33182 3054 33234
rect 3106 33182 3220 33234
rect 3052 33180 3220 33182
rect 3052 33170 3108 33180
rect 2604 33124 2660 33134
rect 2492 33122 2660 33124
rect 2492 33070 2606 33122
rect 2658 33070 2660 33122
rect 2492 33068 2660 33070
rect 2604 33058 2660 33068
rect 2604 32788 2660 32798
rect 2492 32732 2604 32788
rect 2492 32002 2548 32732
rect 2604 32694 2660 32732
rect 3052 32788 3108 32798
rect 3052 32694 3108 32732
rect 3164 32338 3220 33180
rect 3276 33124 3332 33516
rect 3388 33506 3444 33516
rect 3500 33460 3556 33470
rect 3500 33366 3556 33404
rect 3388 33348 3444 33358
rect 3388 33254 3444 33292
rect 3276 33068 3556 33124
rect 3500 32786 3556 33068
rect 3500 32734 3502 32786
rect 3554 32734 3556 32786
rect 3500 32722 3556 32734
rect 3164 32286 3166 32338
rect 3218 32286 3220 32338
rect 3164 32274 3220 32286
rect 3500 32338 3556 32350
rect 3500 32286 3502 32338
rect 3554 32286 3556 32338
rect 2492 31950 2494 32002
rect 2546 31950 2548 32002
rect 2492 31938 2548 31950
rect 3388 32004 3444 32014
rect 3388 31890 3444 31948
rect 3388 31838 3390 31890
rect 3442 31838 3444 31890
rect 3388 31826 3444 31838
rect 2828 31780 2884 31790
rect 2828 31686 2884 31724
rect 3500 31668 3556 32286
rect 3388 31612 3556 31668
rect 2604 31554 2660 31566
rect 3276 31556 3332 31566
rect 2604 31502 2606 31554
rect 2658 31502 2660 31554
rect 1932 30210 2324 30212
rect 1932 30158 2046 30210
rect 2098 30158 2270 30210
rect 2322 30158 2324 30210
rect 1932 30156 2324 30158
rect 1932 28756 1988 30156
rect 2044 30146 2100 30156
rect 2268 30146 2324 30156
rect 2492 30882 2548 30894
rect 2492 30830 2494 30882
rect 2546 30830 2548 30882
rect 2492 29988 2548 30830
rect 2604 30434 2660 31502
rect 2604 30382 2606 30434
rect 2658 30382 2660 30434
rect 2604 30370 2660 30382
rect 2828 31554 3332 31556
rect 2828 31502 3278 31554
rect 3330 31502 3332 31554
rect 2828 31500 3332 31502
rect 2828 30210 2884 31500
rect 3276 31490 3332 31500
rect 2828 30158 2830 30210
rect 2882 30158 2884 30210
rect 2828 30146 2884 30158
rect 3052 30100 3108 30110
rect 3388 30100 3444 31612
rect 3052 30098 3444 30100
rect 3052 30046 3054 30098
rect 3106 30046 3444 30098
rect 3052 30044 3444 30046
rect 3500 30434 3556 30446
rect 3500 30382 3502 30434
rect 3554 30382 3556 30434
rect 3052 30034 3108 30044
rect 2604 29988 2660 29998
rect 2492 29986 2660 29988
rect 2492 29934 2606 29986
rect 2658 29934 2660 29986
rect 2492 29932 2660 29934
rect 2604 29922 2660 29932
rect 2044 29540 2100 29550
rect 2044 29538 2212 29540
rect 2044 29486 2046 29538
rect 2098 29486 2212 29538
rect 2044 29484 2212 29486
rect 2044 29474 2100 29484
rect 2044 28866 2100 28878
rect 2044 28814 2046 28866
rect 2098 28814 2100 28866
rect 2044 28756 2100 28814
rect 1932 28754 2100 28756
rect 1932 28702 2046 28754
rect 2098 28702 2100 28754
rect 1932 28700 2100 28702
rect 2044 28690 2100 28700
rect 1820 27858 1876 28028
rect 1820 27806 1822 27858
rect 1874 27806 1876 27858
rect 1820 27794 1876 27806
rect 2156 27860 2212 29484
rect 2828 29426 2884 29438
rect 2828 29374 2830 29426
rect 2882 29374 2884 29426
rect 2492 29316 2548 29326
rect 2492 29222 2548 29260
rect 2156 27794 2212 27804
rect 2268 28866 2324 28878
rect 2268 28814 2270 28866
rect 2322 28814 2324 28866
rect 2268 28644 2324 28814
rect 2716 28756 2772 28766
rect 2716 28662 2772 28700
rect 2380 28644 2436 28654
rect 2268 28642 2436 28644
rect 2268 28590 2382 28642
rect 2434 28590 2436 28642
rect 2268 28588 2436 28590
rect 1708 26962 1764 26974
rect 1708 26910 1710 26962
rect 1762 26910 1764 26962
rect 1708 26852 1764 26910
rect 2268 26908 2324 28588
rect 2380 28578 2436 28588
rect 2604 28644 2660 28654
rect 2380 28420 2436 28430
rect 2380 28418 2548 28420
rect 2380 28366 2382 28418
rect 2434 28366 2548 28418
rect 2380 28364 2548 28366
rect 2380 28354 2436 28364
rect 2492 27970 2548 28364
rect 2492 27918 2494 27970
rect 2546 27918 2548 27970
rect 2492 27906 2548 27918
rect 2492 27188 2548 27198
rect 2604 27188 2660 28588
rect 2828 28084 2884 29374
rect 3164 29316 3220 30044
rect 3500 29316 3556 30382
rect 3612 30212 3668 38892
rect 3836 38052 3892 40012
rect 4060 39844 4116 39854
rect 3724 37996 3892 38052
rect 3948 39788 4060 39844
rect 3948 39058 4004 39788
rect 4060 39778 4116 39788
rect 3948 39006 3950 39058
rect 4002 39006 4004 39058
rect 3948 38948 4004 39006
rect 3948 38052 4004 38892
rect 3724 36484 3780 37996
rect 3724 35922 3780 36428
rect 3836 37828 3892 37838
rect 3836 36260 3892 37772
rect 3948 36596 4004 37996
rect 4172 38052 4228 38062
rect 3948 36502 4004 36540
rect 4060 37156 4116 37166
rect 3948 36260 4004 36270
rect 3836 36204 3948 36260
rect 3724 35870 3726 35922
rect 3778 35870 3780 35922
rect 3724 33570 3780 35870
rect 3836 36036 3892 36046
rect 3836 34356 3892 35980
rect 3836 34290 3892 34300
rect 3724 33518 3726 33570
rect 3778 33518 3780 33570
rect 3724 32788 3780 33518
rect 3780 32732 3892 32788
rect 3724 32722 3780 32732
rect 3612 30156 3780 30212
rect 3612 29988 3668 29998
rect 3612 29894 3668 29932
rect 3612 29540 3668 29550
rect 3612 29446 3668 29484
rect 3500 29260 3668 29316
rect 2940 28644 2996 28654
rect 2940 28550 2996 28588
rect 3164 28532 3220 29260
rect 3500 28756 3556 28766
rect 3500 28662 3556 28700
rect 3164 28530 3332 28532
rect 3164 28478 3166 28530
rect 3218 28478 3332 28530
rect 3164 28476 3332 28478
rect 3164 28466 3220 28476
rect 2940 28084 2996 28094
rect 2828 28028 2940 28084
rect 2940 28018 2996 28028
rect 2492 27186 2660 27188
rect 2492 27134 2494 27186
rect 2546 27134 2660 27186
rect 2492 27132 2660 27134
rect 2828 27188 2884 27198
rect 2492 27122 2548 27132
rect 1708 26292 1764 26796
rect 2044 26850 2100 26862
rect 2044 26798 2046 26850
rect 2098 26798 2100 26850
rect 1708 26226 1764 26236
rect 1932 26404 1988 26414
rect 1820 23938 1876 23950
rect 1820 23886 1822 23938
rect 1874 23886 1876 23938
rect 1820 23604 1876 23886
rect 1708 23380 1764 23390
rect 1708 23154 1764 23324
rect 1708 23102 1710 23154
rect 1762 23102 1764 23154
rect 1708 22148 1764 23102
rect 1820 22372 1876 23548
rect 1932 22484 1988 26348
rect 2044 25508 2100 26798
rect 2044 25442 2100 25452
rect 2156 26852 2324 26908
rect 2156 25396 2212 26852
rect 2828 26516 2884 27132
rect 2940 27074 2996 27086
rect 2940 27022 2942 27074
rect 2994 27022 2996 27074
rect 2940 26852 2996 27022
rect 2940 26786 2996 26796
rect 3276 26852 3332 28476
rect 3612 28530 3668 29260
rect 3612 28478 3614 28530
rect 3666 28478 3668 28530
rect 3612 28466 3668 28478
rect 3724 28196 3780 30156
rect 3500 28140 3780 28196
rect 3836 28866 3892 32732
rect 3948 32452 4004 36204
rect 4060 35698 4116 37100
rect 4060 35646 4062 35698
rect 4114 35646 4116 35698
rect 4060 35252 4116 35646
rect 4060 35186 4116 35196
rect 3948 32338 4004 32396
rect 3948 32286 3950 32338
rect 4002 32286 4004 32338
rect 3948 32274 4004 32286
rect 4172 32116 4228 37996
rect 3948 32060 4228 32116
rect 3948 30212 4004 32060
rect 4060 31892 4116 31902
rect 4060 31778 4116 31836
rect 4060 31726 4062 31778
rect 4114 31726 4116 31778
rect 4060 30434 4116 31726
rect 4172 31554 4228 31566
rect 4172 31502 4174 31554
rect 4226 31502 4228 31554
rect 4172 31220 4228 31502
rect 4172 31154 4228 31164
rect 4060 30382 4062 30434
rect 4114 30382 4116 30434
rect 4060 30370 4116 30382
rect 3948 30146 4004 30156
rect 4284 30100 4340 40124
rect 4396 39956 4452 40908
rect 4614 40012 4878 40022
rect 4670 39956 4718 40012
rect 4774 39956 4822 40012
rect 4614 39946 4878 39956
rect 4396 39890 4452 39900
rect 4396 39732 4452 39742
rect 4396 39058 4452 39676
rect 4396 39006 4398 39058
rect 4450 39006 4452 39058
rect 4396 37828 4452 39006
rect 4620 39730 4676 39742
rect 4620 39678 4622 39730
rect 4674 39678 4676 39730
rect 4620 39060 4676 39678
rect 4620 38994 4676 39004
rect 4614 38444 4878 38454
rect 4670 38388 4718 38444
rect 4774 38388 4822 38444
rect 4614 38378 4878 38388
rect 4396 37762 4452 37772
rect 4396 37380 4452 37390
rect 4396 36484 4452 37324
rect 4956 37380 5012 41020
rect 5068 40292 5124 40302
rect 5068 40290 5236 40292
rect 5068 40238 5070 40290
rect 5122 40238 5236 40290
rect 5068 40236 5236 40238
rect 5068 40226 5124 40236
rect 5068 39732 5124 39742
rect 5068 39638 5124 39676
rect 5180 39284 5236 40236
rect 5180 39218 5236 39228
rect 5068 38948 5124 38958
rect 5068 38854 5124 38892
rect 5292 38948 5348 38958
rect 4956 37314 5012 37324
rect 4620 37154 4676 37166
rect 4620 37102 4622 37154
rect 4674 37102 4676 37154
rect 4620 37044 4676 37102
rect 5068 37156 5124 37166
rect 5068 37062 5124 37100
rect 4732 37044 4788 37054
rect 4620 36988 4732 37044
rect 4732 36978 4788 36988
rect 4614 36876 4878 36886
rect 4670 36820 4718 36876
rect 4774 36820 4822 36876
rect 4614 36810 4878 36820
rect 5068 36594 5124 36606
rect 5068 36542 5070 36594
rect 5122 36542 5124 36594
rect 4732 36484 4788 36494
rect 4396 36428 4564 36484
rect 4396 36260 4452 36270
rect 4396 36166 4452 36204
rect 4508 35476 4564 36428
rect 4732 36390 4788 36428
rect 5068 36484 5124 36542
rect 5068 36418 5124 36428
rect 5180 36596 5236 36606
rect 4956 36372 5012 36382
rect 4956 36278 5012 36316
rect 4956 36148 5012 36158
rect 4844 35812 4900 35822
rect 4844 35718 4900 35756
rect 4396 35420 4564 35476
rect 4396 33348 4452 35420
rect 4614 35308 4878 35318
rect 4670 35252 4718 35308
rect 4774 35252 4822 35308
rect 4614 35242 4878 35252
rect 4844 35140 4900 35150
rect 4844 35026 4900 35084
rect 4844 34974 4846 35026
rect 4898 34974 4900 35026
rect 4844 34962 4900 34974
rect 4620 34916 4676 34926
rect 4620 34018 4676 34860
rect 4620 33966 4622 34018
rect 4674 33966 4676 34018
rect 4620 33954 4676 33966
rect 4614 33740 4878 33750
rect 4670 33684 4718 33740
rect 4774 33684 4822 33740
rect 4614 33674 4878 33684
rect 4844 33460 4900 33470
rect 4396 33292 4564 33348
rect 4396 33124 4452 33134
rect 4396 33030 4452 33068
rect 4508 32788 4564 33292
rect 4396 32732 4564 32788
rect 4844 33122 4900 33404
rect 4956 33348 5012 36092
rect 5180 34130 5236 36540
rect 5180 34078 5182 34130
rect 5234 34078 5236 34130
rect 5180 33572 5236 34078
rect 5180 33506 5236 33516
rect 5180 33348 5236 33358
rect 4956 33292 5180 33348
rect 5180 33282 5236 33292
rect 4844 33070 4846 33122
rect 4898 33070 4900 33122
rect 4396 30212 4452 32732
rect 4844 32452 4900 33070
rect 4844 32386 4900 32396
rect 4614 32172 4878 32182
rect 4670 32116 4718 32172
rect 4774 32116 4822 32172
rect 4614 32106 4878 32116
rect 4620 32004 4676 32014
rect 4620 30882 4676 31948
rect 4732 31780 4788 31790
rect 4732 31686 4788 31724
rect 5068 31668 5124 31678
rect 5068 31666 5236 31668
rect 5068 31614 5070 31666
rect 5122 31614 5236 31666
rect 5068 31612 5236 31614
rect 5068 31602 5124 31612
rect 5180 31556 5236 31612
rect 5180 31490 5236 31500
rect 5068 31332 5124 31342
rect 5068 31218 5124 31276
rect 5068 31166 5070 31218
rect 5122 31166 5124 31218
rect 5068 31154 5124 31166
rect 4620 30830 4622 30882
rect 4674 30830 4676 30882
rect 4620 30818 4676 30830
rect 4614 30604 4878 30614
rect 4670 30548 4718 30604
rect 4774 30548 4822 30604
rect 4614 30538 4878 30548
rect 4732 30436 4788 30446
rect 4396 30156 4564 30212
rect 4060 30044 4340 30100
rect 3948 29986 4004 29998
rect 3948 29934 3950 29986
rect 4002 29934 4004 29986
rect 3948 29876 4004 29934
rect 3948 29810 4004 29820
rect 3836 28814 3838 28866
rect 3890 28814 3892 28866
rect 3388 26852 3444 26862
rect 3276 26850 3444 26852
rect 3276 26798 3390 26850
rect 3442 26798 3444 26850
rect 3276 26796 3444 26798
rect 2492 26514 2884 26516
rect 2492 26462 2830 26514
rect 2882 26462 2884 26514
rect 2492 26460 2884 26462
rect 2492 25844 2548 26460
rect 2828 26450 2884 26460
rect 2268 25788 2548 25844
rect 2268 25618 2324 25788
rect 2492 25730 2548 25788
rect 2492 25678 2494 25730
rect 2546 25678 2548 25730
rect 2492 25666 2548 25678
rect 2268 25566 2270 25618
rect 2322 25566 2324 25618
rect 2268 25554 2324 25566
rect 3276 25620 3332 26796
rect 3388 26786 3444 26796
rect 3388 26404 3444 26414
rect 3388 26310 3444 26348
rect 3500 25732 3556 28140
rect 3836 28084 3892 28814
rect 3612 28028 3892 28084
rect 3612 27188 3668 28028
rect 4060 27972 4116 30044
rect 4396 29988 4452 29998
rect 4396 29894 4452 29932
rect 4508 29764 4564 30156
rect 4732 29876 4788 30380
rect 5068 30436 5124 30446
rect 5068 30434 5236 30436
rect 5068 30382 5070 30434
rect 5122 30382 5236 30434
rect 5068 30380 5236 30382
rect 5068 30370 5124 30380
rect 5180 30324 5236 30380
rect 5180 30258 5236 30268
rect 5068 30212 5124 30222
rect 5068 30118 5124 30156
rect 4732 29810 4788 29820
rect 5180 29988 5236 29998
rect 4396 29708 4564 29764
rect 4284 29428 4340 29438
rect 4284 28756 4340 29372
rect 4284 28662 4340 28700
rect 4172 28644 4228 28654
rect 4172 28550 4228 28588
rect 3612 27122 3668 27132
rect 3724 27916 4116 27972
rect 4284 28532 4340 28542
rect 2716 25508 2772 25518
rect 2268 25396 2324 25406
rect 2156 25340 2268 25396
rect 2044 24724 2100 24734
rect 2268 24724 2324 25340
rect 2716 25394 2772 25452
rect 2716 25342 2718 25394
rect 2770 25342 2772 25394
rect 2716 25330 2772 25342
rect 2604 25282 2660 25294
rect 2604 25230 2606 25282
rect 2658 25230 2660 25282
rect 2380 24948 2436 24958
rect 2380 24946 2548 24948
rect 2380 24894 2382 24946
rect 2434 24894 2548 24946
rect 2380 24892 2548 24894
rect 2380 24882 2436 24892
rect 2380 24724 2436 24734
rect 2044 24722 2436 24724
rect 2044 24670 2046 24722
rect 2098 24670 2382 24722
rect 2434 24670 2436 24722
rect 2044 24668 2436 24670
rect 2044 24658 2100 24668
rect 2044 23380 2100 23390
rect 2044 23286 2100 23324
rect 1932 22428 2324 22484
rect 1820 22370 1988 22372
rect 1820 22318 1822 22370
rect 1874 22318 1988 22370
rect 1820 22316 1988 22318
rect 1820 22306 1876 22316
rect 1820 22148 1876 22158
rect 1708 22092 1820 22148
rect 1820 22082 1876 22092
rect 1820 21586 1876 21598
rect 1820 21534 1822 21586
rect 1874 21534 1876 21586
rect 1820 20916 1876 21534
rect 1820 20822 1876 20860
rect 1820 19236 1876 19246
rect 1932 19236 1988 22316
rect 2044 21698 2100 21710
rect 2044 21646 2046 21698
rect 2098 21646 2100 21698
rect 2044 20804 2100 21646
rect 2044 20738 2100 20748
rect 1820 19234 1988 19236
rect 1820 19182 1822 19234
rect 1874 19182 1988 19234
rect 1820 19180 1988 19182
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18228 1764 18398
rect 1708 18162 1764 18172
rect 1820 16882 1876 19180
rect 2268 18788 2324 22428
rect 2380 21588 2436 24668
rect 2492 24050 2548 24892
rect 2604 24498 2660 25230
rect 2940 24724 2996 24734
rect 2940 24630 2996 24668
rect 3164 24724 3220 24734
rect 3276 24724 3332 25564
rect 3164 24722 3332 24724
rect 3164 24670 3166 24722
rect 3218 24670 3332 24722
rect 3164 24668 3332 24670
rect 3388 25676 3556 25732
rect 2604 24446 2606 24498
rect 2658 24446 2660 24498
rect 2604 24434 2660 24446
rect 2492 23998 2494 24050
rect 2546 23998 2548 24050
rect 2492 23986 2548 23998
rect 3164 23548 3220 24668
rect 2716 23492 3220 23548
rect 2716 23042 2772 23492
rect 3164 23380 3220 23390
rect 3388 23380 3444 25676
rect 3500 25508 3556 25518
rect 3500 25414 3556 25452
rect 3612 24836 3668 24846
rect 3612 24742 3668 24780
rect 3500 24724 3556 24734
rect 3500 24630 3556 24668
rect 3724 23548 3780 27916
rect 3836 27188 3892 27198
rect 3836 27094 3892 27132
rect 4284 27186 4340 28476
rect 4284 27134 4286 27186
rect 4338 27134 4340 27186
rect 4284 26404 4340 27134
rect 4284 26338 4340 26348
rect 4060 25508 4116 25518
rect 4060 25414 4116 25452
rect 4396 24948 4452 29708
rect 4614 29036 4878 29046
rect 4670 28980 4718 29036
rect 4774 28980 4822 29036
rect 4614 28970 4878 28980
rect 4620 28756 4676 28766
rect 4620 27746 4676 28700
rect 5180 28754 5236 29932
rect 5180 28702 5182 28754
rect 5234 28702 5236 28754
rect 5180 28690 5236 28702
rect 5068 28084 5124 28094
rect 5068 27990 5124 28028
rect 4620 27694 4622 27746
rect 4674 27694 4676 27746
rect 4620 27682 4676 27694
rect 4614 27468 4878 27478
rect 4670 27412 4718 27468
rect 4774 27412 4822 27468
rect 4614 27402 4878 27412
rect 5068 27188 5124 27198
rect 5068 27094 5124 27132
rect 5292 26908 5348 38892
rect 5404 33906 5460 42476
rect 5628 42420 5684 44156
rect 5852 44212 5908 44222
rect 5852 44118 5908 44156
rect 5516 42364 5684 42420
rect 5740 44098 5796 44110
rect 5740 44046 5742 44098
rect 5794 44046 5796 44098
rect 5516 41076 5572 42364
rect 5740 42084 5796 44046
rect 5740 42018 5796 42028
rect 5628 41300 5684 41310
rect 5684 41244 5796 41300
rect 5628 41234 5684 41244
rect 5740 41188 5796 41244
rect 5852 41188 5908 41198
rect 5740 41186 5908 41188
rect 5740 41134 5854 41186
rect 5906 41134 5908 41186
rect 5740 41132 5908 41134
rect 5852 41122 5908 41132
rect 5516 41020 5796 41076
rect 5516 40628 5572 40638
rect 5516 40068 5572 40572
rect 5516 39058 5572 40012
rect 5628 39844 5684 39854
rect 5628 39618 5684 39788
rect 5628 39566 5630 39618
rect 5682 39566 5684 39618
rect 5628 39554 5684 39566
rect 5628 39394 5684 39406
rect 5628 39342 5630 39394
rect 5682 39342 5684 39394
rect 5628 39284 5684 39342
rect 5628 39218 5684 39228
rect 5516 39006 5518 39058
rect 5570 39006 5572 39058
rect 5516 37268 5572 39006
rect 5740 38668 5796 41020
rect 5964 39842 6020 44380
rect 6300 44212 6356 44940
rect 6524 44548 6580 45612
rect 6636 45332 6692 47740
rect 6748 47458 6804 50204
rect 6860 49140 6916 49150
rect 6860 48356 6916 49084
rect 6972 49028 7028 50372
rect 6972 48962 7028 48972
rect 7084 49812 7140 49822
rect 7084 48804 7140 49756
rect 6860 48290 6916 48300
rect 6972 48748 7140 48804
rect 6748 47406 6750 47458
rect 6802 47406 6804 47458
rect 6748 47348 6804 47406
rect 6748 47282 6804 47292
rect 6860 46564 6916 46574
rect 6860 46002 6916 46508
rect 6860 45950 6862 46002
rect 6914 45950 6916 46002
rect 6860 45938 6916 45950
rect 6748 45778 6804 45790
rect 6748 45726 6750 45778
rect 6802 45726 6804 45778
rect 6748 45668 6804 45726
rect 6748 45602 6804 45612
rect 6972 45444 7028 48748
rect 7084 48130 7140 48142
rect 7084 48078 7086 48130
rect 7138 48078 7140 48130
rect 7084 47908 7140 48078
rect 7084 47842 7140 47852
rect 7084 47124 7140 47134
rect 7084 46116 7140 47068
rect 7084 46050 7140 46060
rect 6972 45378 7028 45388
rect 7084 45778 7140 45790
rect 7084 45726 7086 45778
rect 7138 45726 7140 45778
rect 6636 44660 6692 45276
rect 7084 45332 7140 45726
rect 7196 45444 7252 50764
rect 7308 50596 7364 50606
rect 7308 50502 7364 50540
rect 7868 50596 7924 50606
rect 7532 50484 7588 50494
rect 7420 50372 7588 50428
rect 7420 49698 7476 50372
rect 7868 50036 7924 50540
rect 8092 50482 8148 50494
rect 8092 50430 8094 50482
rect 8146 50430 8148 50482
rect 8092 50428 8148 50430
rect 8092 50372 8596 50428
rect 8428 50260 8484 50270
rect 8016 50204 8280 50214
rect 8072 50148 8120 50204
rect 8176 50148 8224 50204
rect 8016 50138 8280 50148
rect 8092 50036 8148 50046
rect 7868 50034 8148 50036
rect 7868 49982 8094 50034
rect 8146 49982 8148 50034
rect 7868 49980 8148 49982
rect 8092 49970 8148 49980
rect 7420 49646 7422 49698
rect 7474 49646 7476 49698
rect 7420 49634 7476 49646
rect 8204 49924 8260 49934
rect 7420 49250 7476 49262
rect 7420 49198 7422 49250
rect 7474 49198 7476 49250
rect 7420 49138 7476 49198
rect 7420 49086 7422 49138
rect 7474 49086 7476 49138
rect 7420 49074 7476 49086
rect 7868 49252 7924 49262
rect 7868 49138 7924 49196
rect 7868 49086 7870 49138
rect 7922 49086 7924 49138
rect 7868 49074 7924 49086
rect 8204 49250 8260 49868
rect 8204 49198 8206 49250
rect 8258 49198 8260 49250
rect 8204 49138 8260 49198
rect 8204 49086 8206 49138
rect 8258 49086 8260 49138
rect 8204 49074 8260 49086
rect 8428 49810 8484 50204
rect 8540 50034 8596 50372
rect 8540 49982 8542 50034
rect 8594 49982 8596 50034
rect 8540 49970 8596 49982
rect 8428 49758 8430 49810
rect 8482 49758 8484 49810
rect 8428 49140 8484 49758
rect 8652 49812 8708 50988
rect 8652 49718 8708 49756
rect 8764 50260 8820 50270
rect 7308 49028 7364 49038
rect 7308 46116 7364 48972
rect 8016 48636 8280 48646
rect 8072 48580 8120 48636
rect 8176 48580 8224 48636
rect 8016 48570 8280 48580
rect 7532 48468 7588 48478
rect 8428 48468 8484 49084
rect 8652 49252 8708 49262
rect 8652 49138 8708 49196
rect 8652 49086 8654 49138
rect 8706 49086 8708 49138
rect 8652 49074 8708 49086
rect 7532 48374 7588 48412
rect 8316 48412 8484 48468
rect 8316 48244 8372 48412
rect 8316 48150 8372 48188
rect 8540 48356 8596 48366
rect 8540 48242 8596 48300
rect 8540 48190 8542 48242
rect 8594 48190 8596 48242
rect 7420 48132 7476 48142
rect 7420 47570 7476 48076
rect 8092 48130 8148 48142
rect 8092 48078 8094 48130
rect 8146 48078 8148 48130
rect 8092 47684 8148 48078
rect 8428 48132 8484 48142
rect 8428 48038 8484 48076
rect 8204 47684 8260 47694
rect 8092 47628 8204 47684
rect 8204 47618 8260 47628
rect 7420 47518 7422 47570
rect 7474 47518 7476 47570
rect 7420 47506 7476 47518
rect 8016 47068 8280 47078
rect 8072 47012 8120 47068
rect 8176 47012 8224 47068
rect 8540 47068 8596 48190
rect 8540 47012 8708 47068
rect 8016 47002 8280 47012
rect 8428 46562 8484 46574
rect 8428 46510 8430 46562
rect 8482 46510 8484 46562
rect 8428 46228 8484 46510
rect 7308 46050 7364 46060
rect 8204 46172 8484 46228
rect 7308 45892 7364 45902
rect 7868 45892 7924 45902
rect 7308 45890 7924 45892
rect 7308 45838 7310 45890
rect 7362 45838 7870 45890
rect 7922 45838 7924 45890
rect 7308 45836 7924 45838
rect 7308 45826 7364 45836
rect 7868 45826 7924 45836
rect 7980 45892 8036 45902
rect 7980 45798 8036 45836
rect 8204 45892 8260 46172
rect 7756 45666 7812 45678
rect 7756 45614 7758 45666
rect 7810 45614 7812 45666
rect 7756 45556 7812 45614
rect 8204 45668 8260 45836
rect 8316 45892 8372 45902
rect 8316 45890 8484 45892
rect 8316 45838 8318 45890
rect 8370 45838 8484 45890
rect 8316 45836 8484 45838
rect 8316 45826 8372 45836
rect 8204 45602 8260 45612
rect 8428 45780 8484 45836
rect 8428 45556 8484 45724
rect 7756 45490 7812 45500
rect 8016 45500 8280 45510
rect 8072 45444 8120 45500
rect 8176 45444 8224 45500
rect 8428 45490 8484 45500
rect 8016 45434 8280 45444
rect 7196 45378 7252 45388
rect 7084 45266 7140 45276
rect 8428 45332 8484 45342
rect 7644 45218 7700 45230
rect 7644 45166 7646 45218
rect 7698 45166 7700 45218
rect 7644 45108 7700 45166
rect 7644 45052 7924 45108
rect 6748 44994 6804 45006
rect 6748 44942 6750 44994
rect 6802 44942 6804 44994
rect 6748 44884 6804 44942
rect 7196 44996 7252 45034
rect 7196 44930 7252 44940
rect 7532 44996 7588 45006
rect 7588 44940 7700 44996
rect 7532 44930 7588 44940
rect 6748 44818 6804 44828
rect 6748 44660 6804 44670
rect 6636 44604 6748 44660
rect 6748 44594 6804 44604
rect 7532 44660 7588 44670
rect 6860 44548 6916 44558
rect 6524 44492 6692 44548
rect 6300 44146 6356 44156
rect 6412 44322 6468 44334
rect 6412 44270 6414 44322
rect 6466 44270 6468 44322
rect 6188 44100 6244 44110
rect 6076 42868 6132 42878
rect 6076 42774 6132 42812
rect 6188 42644 6244 44044
rect 6412 43540 6468 44270
rect 6412 43474 6468 43484
rect 5964 39790 5966 39842
rect 6018 39790 6020 39842
rect 5964 39778 6020 39790
rect 6076 42588 6244 42644
rect 6524 42754 6580 42766
rect 6524 42702 6526 42754
rect 6578 42702 6580 42754
rect 6076 38948 6132 42588
rect 6524 41188 6580 42702
rect 6524 41122 6580 41132
rect 6300 41076 6356 41086
rect 6300 40982 6356 41020
rect 6188 40962 6244 40974
rect 6188 40910 6190 40962
rect 6242 40910 6244 40962
rect 6188 39618 6244 40910
rect 6524 40516 6580 40526
rect 6188 39566 6190 39618
rect 6242 39566 6244 39618
rect 6188 39554 6244 39566
rect 6412 39732 6468 39742
rect 6412 39618 6468 39676
rect 6412 39566 6414 39618
rect 6466 39566 6468 39618
rect 6412 39554 6468 39566
rect 6076 38882 6132 38892
rect 5516 37202 5572 37212
rect 5628 38612 5796 38668
rect 5628 36820 5684 38612
rect 5404 33854 5406 33906
rect 5458 33854 5460 33906
rect 5404 33842 5460 33854
rect 5516 36764 5684 36820
rect 5740 38500 5796 38510
rect 5180 26852 5348 26908
rect 5404 33348 5460 33358
rect 5404 31556 5460 33292
rect 4956 26292 5012 26302
rect 4956 26198 5012 26236
rect 4614 25900 4878 25910
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4614 25834 4878 25844
rect 5068 25620 5124 25630
rect 5068 25526 5124 25564
rect 4620 25396 4676 25406
rect 4620 25302 4676 25340
rect 5180 25060 5236 26852
rect 5404 26740 5460 31500
rect 5516 30884 5572 36764
rect 5628 36596 5684 36606
rect 5628 36482 5684 36540
rect 5628 36430 5630 36482
rect 5682 36430 5684 36482
rect 5628 36418 5684 36430
rect 5628 36258 5684 36270
rect 5628 36206 5630 36258
rect 5682 36206 5684 36258
rect 5628 35812 5684 36206
rect 5628 35746 5684 35756
rect 5740 34468 5796 38444
rect 6188 38050 6244 38062
rect 6188 37998 6190 38050
rect 6242 37998 6244 38050
rect 5852 37828 5908 37838
rect 6188 37828 6244 37998
rect 5852 37826 6244 37828
rect 5852 37774 5854 37826
rect 5906 37774 6244 37826
rect 5852 37772 6244 37774
rect 5852 37268 5908 37772
rect 6412 37492 6468 37502
rect 6412 37398 6468 37436
rect 5852 37202 5908 37212
rect 5964 37156 6020 37166
rect 5964 37062 6020 37100
rect 5852 37042 5908 37054
rect 5852 36990 5854 37042
rect 5906 36990 5908 37042
rect 5852 36708 5908 36990
rect 5852 36652 6132 36708
rect 5964 36484 6020 36494
rect 5964 36390 6020 36428
rect 6076 36482 6132 36652
rect 6076 36430 6078 36482
rect 6130 36430 6132 36482
rect 6076 36418 6132 36430
rect 6412 36370 6468 36382
rect 6412 36318 6414 36370
rect 6466 36318 6468 36370
rect 6412 36260 6468 36318
rect 6412 36194 6468 36204
rect 5516 30818 5572 30828
rect 5628 34412 5796 34468
rect 5628 31220 5684 34412
rect 6412 34356 6468 34366
rect 5740 34354 6468 34356
rect 5740 34302 6414 34354
rect 6466 34302 6468 34354
rect 5740 34300 6468 34302
rect 6524 34356 6580 40460
rect 6636 38164 6692 44492
rect 6748 44324 6804 44334
rect 6748 44230 6804 44268
rect 6860 44322 6916 44492
rect 6860 44270 6862 44322
rect 6914 44270 6916 44322
rect 6860 44258 6916 44270
rect 7308 44324 7364 44334
rect 6972 44098 7028 44110
rect 6972 44046 6974 44098
rect 7026 44046 7028 44098
rect 6748 43988 6804 43998
rect 6748 38388 6804 43932
rect 6972 42532 7028 44046
rect 7196 42980 7252 42990
rect 7196 42866 7252 42924
rect 7196 42814 7198 42866
rect 7250 42814 7252 42866
rect 7196 42802 7252 42814
rect 6860 41860 6916 41870
rect 6860 41186 6916 41804
rect 6972 41858 7028 42476
rect 6972 41806 6974 41858
rect 7026 41806 7028 41858
rect 6972 41794 7028 41806
rect 6860 41134 6862 41186
rect 6914 41134 6916 41186
rect 6860 41122 6916 41134
rect 7196 41076 7252 41086
rect 7196 40292 7252 41020
rect 7308 40962 7364 44268
rect 7532 44100 7588 44604
rect 7644 44324 7700 44940
rect 7644 44258 7700 44268
rect 7756 44882 7812 44894
rect 7756 44830 7758 44882
rect 7810 44830 7812 44882
rect 7756 44322 7812 44830
rect 7868 44548 7924 45052
rect 7868 44482 7924 44492
rect 7980 44996 8036 45006
rect 7980 44436 8036 44940
rect 7980 44370 8036 44380
rect 8428 44434 8484 45276
rect 8428 44382 8430 44434
rect 8482 44382 8484 44434
rect 8428 44370 8484 44382
rect 8540 44994 8596 45006
rect 8540 44942 8542 44994
rect 8594 44942 8596 44994
rect 8540 44882 8596 44942
rect 8652 44996 8708 47012
rect 8652 44930 8708 44940
rect 8540 44830 8542 44882
rect 8594 44830 8596 44882
rect 7756 44270 7758 44322
rect 7810 44270 7812 44322
rect 7756 44258 7812 44270
rect 7868 44212 7924 44222
rect 7532 44044 7812 44100
rect 7756 42756 7812 44044
rect 7756 42690 7812 42700
rect 7756 41970 7812 41982
rect 7756 41918 7758 41970
rect 7810 41918 7812 41970
rect 7532 41858 7588 41870
rect 7532 41806 7534 41858
rect 7586 41806 7588 41858
rect 7532 41748 7588 41806
rect 7532 41682 7588 41692
rect 7308 40910 7310 40962
rect 7362 40910 7364 40962
rect 7308 40852 7364 40910
rect 7308 40786 7364 40796
rect 7644 41188 7700 41198
rect 7196 40290 7364 40292
rect 7196 40238 7198 40290
rect 7250 40238 7364 40290
rect 7196 40236 7364 40238
rect 7196 40226 7252 40236
rect 7196 40068 7252 40078
rect 7196 39730 7252 40012
rect 7308 39842 7364 40236
rect 7644 40068 7700 41132
rect 7756 40740 7812 41918
rect 7756 40674 7812 40684
rect 7756 40516 7812 40526
rect 7868 40516 7924 44156
rect 8016 43932 8280 43942
rect 8072 43876 8120 43932
rect 8176 43876 8224 43932
rect 8016 43866 8280 43876
rect 8540 43540 8596 44830
rect 8764 44436 8820 50204
rect 8876 49810 8932 51214
rect 8876 49758 8878 49810
rect 8930 49758 8932 49810
rect 8876 49746 8932 49758
rect 9100 51268 9156 51278
rect 9100 49138 9156 51212
rect 9100 49086 9102 49138
rect 9154 49086 9156 49138
rect 9100 48916 9156 49086
rect 9100 48850 9156 48860
rect 8876 48242 8932 48254
rect 8876 48190 8878 48242
rect 8930 48190 8932 48242
rect 8876 48132 8932 48190
rect 9212 48132 9268 48142
rect 8876 48076 9212 48132
rect 9212 48066 9268 48076
rect 9212 47908 9268 47918
rect 9100 47684 9156 47694
rect 8988 46564 9044 46574
rect 8876 46508 8988 46564
rect 8876 44882 8932 46508
rect 8988 46470 9044 46508
rect 8988 46004 9044 46014
rect 9100 46004 9156 47628
rect 8988 46002 9156 46004
rect 8988 45950 8990 46002
rect 9042 45950 9156 46002
rect 8988 45948 9156 45950
rect 8988 45938 9044 45948
rect 9212 45892 9268 47852
rect 9212 45826 9268 45836
rect 9212 45444 9268 45454
rect 9100 45108 9156 45146
rect 9100 45042 9156 45052
rect 8876 44830 8878 44882
rect 8930 44830 8932 44882
rect 8876 44818 8932 44830
rect 8988 44996 9044 45006
rect 8876 44436 8932 44446
rect 8764 44380 8876 44436
rect 8876 44370 8932 44380
rect 8652 44322 8708 44334
rect 8652 44270 8654 44322
rect 8706 44270 8708 44322
rect 8652 44100 8708 44270
rect 8652 44034 8708 44044
rect 8988 44210 9044 44940
rect 9212 44660 9268 45388
rect 8988 44158 8990 44210
rect 9042 44158 9044 44210
rect 8540 43474 8596 43484
rect 8652 43876 8708 43886
rect 8540 42980 8596 42990
rect 8016 42364 8280 42374
rect 8072 42308 8120 42364
rect 8176 42308 8224 42364
rect 8016 42298 8280 42308
rect 8316 42196 8372 42206
rect 8204 42140 8316 42196
rect 8092 41972 8148 41982
rect 8092 41188 8148 41916
rect 8204 41970 8260 42140
rect 8316 42130 8372 42140
rect 8540 42194 8596 42924
rect 8540 42142 8542 42194
rect 8594 42142 8596 42194
rect 8540 42130 8596 42142
rect 8204 41918 8206 41970
rect 8258 41918 8260 41970
rect 8204 41906 8260 41918
rect 8540 41970 8596 41982
rect 8540 41918 8542 41970
rect 8594 41918 8596 41970
rect 8092 41122 8148 41132
rect 8428 41074 8484 41086
rect 8428 41022 8430 41074
rect 8482 41022 8484 41074
rect 8016 40796 8280 40806
rect 8072 40740 8120 40796
rect 8176 40740 8224 40796
rect 8016 40730 8280 40740
rect 8428 40626 8484 41022
rect 8428 40574 8430 40626
rect 8482 40574 8484 40626
rect 8428 40562 8484 40574
rect 7812 40460 7924 40516
rect 8204 40516 8260 40526
rect 7756 40450 7812 40460
rect 7868 40292 7924 40302
rect 8204 40292 8260 40460
rect 7868 40290 8260 40292
rect 7868 40238 7870 40290
rect 7922 40238 8260 40290
rect 7868 40236 8260 40238
rect 7868 40226 7924 40236
rect 7756 40068 7812 40078
rect 7644 40012 7756 40068
rect 7756 40002 7812 40012
rect 7308 39790 7310 39842
rect 7362 39790 7364 39842
rect 7308 39778 7364 39790
rect 7868 39842 7924 39854
rect 7868 39790 7870 39842
rect 7922 39790 7924 39842
rect 7196 39678 7198 39730
rect 7250 39678 7252 39730
rect 7196 39666 7252 39678
rect 7756 39394 7812 39406
rect 7756 39342 7758 39394
rect 7810 39342 7812 39394
rect 7756 38948 7812 39342
rect 7756 38882 7812 38892
rect 7644 38836 7700 38846
rect 6748 38322 6804 38332
rect 7420 38388 7476 38398
rect 6636 38108 6916 38164
rect 6860 37492 6916 38108
rect 6972 37940 7028 37950
rect 6972 37938 7364 37940
rect 6972 37886 6974 37938
rect 7026 37886 7364 37938
rect 6972 37884 7364 37886
rect 6972 37874 7028 37884
rect 7196 37716 7252 37726
rect 6860 37490 7140 37492
rect 6860 37438 6862 37490
rect 6914 37438 7140 37490
rect 6860 37436 7140 37438
rect 6860 37426 6916 37436
rect 7084 37266 7140 37436
rect 7084 37214 7086 37266
rect 7138 37214 7140 37266
rect 6972 36932 7028 36942
rect 6860 36708 6916 36718
rect 6748 36482 6804 36494
rect 6748 36430 6750 36482
rect 6802 36430 6804 36482
rect 6748 36372 6804 36430
rect 6748 36306 6804 36316
rect 6748 36148 6804 36158
rect 6524 34300 6692 34356
rect 5740 34242 5796 34300
rect 6412 34290 6468 34300
rect 5740 34190 5742 34242
rect 5794 34190 5796 34242
rect 5740 34178 5796 34190
rect 5964 34130 6020 34142
rect 5964 34078 5966 34130
rect 6018 34078 6020 34130
rect 5852 34018 5908 34030
rect 5852 33966 5854 34018
rect 5906 33966 5908 34018
rect 5852 33460 5908 33966
rect 5964 33684 6020 34078
rect 6524 34018 6580 34030
rect 6524 33966 6526 34018
rect 6578 33966 6580 34018
rect 6524 33796 6580 33966
rect 6524 33730 6580 33740
rect 5964 33618 6020 33628
rect 6412 33460 6468 33470
rect 5852 33458 6468 33460
rect 5852 33406 6414 33458
rect 6466 33406 6468 33458
rect 5852 33404 6468 33406
rect 6412 33394 6468 33404
rect 5740 33348 5796 33358
rect 5740 33346 5908 33348
rect 5740 33294 5742 33346
rect 5794 33294 5908 33346
rect 5740 33292 5908 33294
rect 5740 33282 5796 33292
rect 5852 31780 5908 33292
rect 6300 32452 6356 32462
rect 6300 31780 6356 32396
rect 5852 31778 6356 31780
rect 5852 31726 5854 31778
rect 5906 31726 6302 31778
rect 6354 31726 6356 31778
rect 5852 31724 6356 31726
rect 5852 31332 5908 31724
rect 5852 31266 5908 31276
rect 5740 31220 5796 31230
rect 5628 31218 5796 31220
rect 5628 31166 5742 31218
rect 5794 31166 5796 31218
rect 5628 31164 5796 31166
rect 5628 30996 5684 31164
rect 5740 31154 5796 31164
rect 5628 30212 5684 30940
rect 5852 30434 5908 30446
rect 5852 30382 5854 30434
rect 5906 30382 5908 30434
rect 5852 30324 5908 30382
rect 5852 30258 5908 30268
rect 5516 30210 5684 30212
rect 5516 30158 5630 30210
rect 5682 30158 5684 30210
rect 5516 30156 5684 30158
rect 5516 29988 5572 30156
rect 5628 30146 5684 30156
rect 5740 30212 5796 30222
rect 5516 29922 5572 29932
rect 5628 29986 5684 29998
rect 5628 29934 5630 29986
rect 5682 29934 5684 29986
rect 5628 29540 5684 29934
rect 5628 29474 5684 29484
rect 5740 29314 5796 30156
rect 6076 29428 6132 31724
rect 6300 31714 6356 31724
rect 6300 31220 6356 31230
rect 6300 31126 6356 31164
rect 6636 31108 6692 34300
rect 6748 33460 6804 36092
rect 6748 33394 6804 33404
rect 6860 32116 6916 36652
rect 6972 35586 7028 36876
rect 6972 35534 6974 35586
rect 7026 35534 7028 35586
rect 6972 35522 7028 35534
rect 7084 35364 7140 37214
rect 6972 35308 7140 35364
rect 6972 32676 7028 35308
rect 7196 35252 7252 37660
rect 7308 37490 7364 37884
rect 7308 37438 7310 37490
rect 7362 37438 7364 37490
rect 7308 37426 7364 37438
rect 7420 37492 7476 38332
rect 7420 37426 7476 37436
rect 7532 37828 7588 37838
rect 7532 37380 7588 37772
rect 7532 37286 7588 37324
rect 7420 37268 7476 37278
rect 7420 35922 7476 37212
rect 7420 35870 7422 35922
rect 7474 35870 7476 35922
rect 7420 35858 7476 35870
rect 7084 35196 7252 35252
rect 7084 35028 7140 35196
rect 7084 33684 7140 34972
rect 7196 34356 7252 34366
rect 7196 34262 7252 34300
rect 7532 34020 7588 34030
rect 7084 33618 7140 33628
rect 7420 33964 7532 34020
rect 6972 32610 7028 32620
rect 6860 32060 7364 32116
rect 6972 31668 7028 31678
rect 7196 31668 7252 31678
rect 6972 31666 7140 31668
rect 6972 31614 6974 31666
rect 7026 31614 7140 31666
rect 6972 31612 7140 31614
rect 6972 31602 7028 31612
rect 7084 31218 7140 31612
rect 7084 31166 7086 31218
rect 7138 31166 7140 31218
rect 7084 31154 7140 31166
rect 7196 31220 7252 31612
rect 6524 31052 6692 31108
rect 7196 31106 7252 31164
rect 7196 31054 7198 31106
rect 7250 31054 7252 31106
rect 6412 30884 6468 30894
rect 6412 30210 6468 30828
rect 6412 30158 6414 30210
rect 6466 30158 6468 30210
rect 6412 30146 6468 30158
rect 5740 29262 5742 29314
rect 5794 29262 5796 29314
rect 5740 29250 5796 29262
rect 5964 29426 6132 29428
rect 5964 29374 6078 29426
rect 6130 29374 6132 29426
rect 5964 29372 6132 29374
rect 5964 28866 6020 29372
rect 6076 29362 6132 29372
rect 6188 30100 6244 30110
rect 5964 28814 5966 28866
rect 6018 28814 6020 28866
rect 5964 28754 6020 28814
rect 5964 28702 5966 28754
rect 6018 28702 6020 28754
rect 5964 28084 6020 28702
rect 6020 28028 6132 28084
rect 5964 28018 6020 28028
rect 5852 27860 5908 27870
rect 5628 27188 5684 27198
rect 5628 27094 5684 27132
rect 5852 27076 5908 27804
rect 5852 26962 5908 27020
rect 5852 26910 5854 26962
rect 5906 26910 5908 26962
rect 5852 26898 5908 26910
rect 5964 27186 6020 27198
rect 5964 27134 5966 27186
rect 6018 27134 6020 27186
rect 5404 26684 5908 26740
rect 5740 25506 5796 25518
rect 5740 25454 5742 25506
rect 5794 25454 5796 25506
rect 5740 25396 5796 25454
rect 5740 25330 5796 25340
rect 5628 25284 5684 25294
rect 5068 25004 5236 25060
rect 5516 25282 5684 25284
rect 5516 25230 5630 25282
rect 5682 25230 5684 25282
rect 5516 25228 5684 25230
rect 3164 23286 3220 23324
rect 3276 23324 3444 23380
rect 3500 23492 3780 23548
rect 3836 24892 4452 24948
rect 4508 24948 4564 24958
rect 2716 22990 2718 23042
rect 2770 22990 2772 23042
rect 2492 22258 2548 22270
rect 2492 22206 2494 22258
rect 2546 22206 2548 22258
rect 2492 21812 2548 22206
rect 2716 22036 2772 22990
rect 2716 21970 2772 21980
rect 3052 22930 3108 22942
rect 3052 22878 3054 22930
rect 3106 22878 3108 22930
rect 2716 21812 2772 21822
rect 2492 21810 2772 21812
rect 2492 21758 2718 21810
rect 2770 21758 2772 21810
rect 2492 21756 2772 21758
rect 2716 21746 2772 21756
rect 2716 21588 2772 21598
rect 2380 21586 2772 21588
rect 2380 21534 2718 21586
rect 2770 21534 2772 21586
rect 2380 21532 2772 21534
rect 2380 21252 2436 21262
rect 2380 20914 2436 21196
rect 2380 20862 2382 20914
rect 2434 20862 2436 20914
rect 2380 20850 2436 20862
rect 2492 20244 2548 20254
rect 2380 20242 2548 20244
rect 2380 20190 2494 20242
rect 2546 20190 2548 20242
rect 2380 20188 2548 20190
rect 2380 19348 2436 20188
rect 2492 20178 2548 20188
rect 2604 20018 2660 21532
rect 2716 21522 2772 21532
rect 3052 21586 3108 22878
rect 3276 22932 3332 23324
rect 3388 23156 3444 23166
rect 3500 23156 3556 23492
rect 3836 23266 3892 24892
rect 4060 24724 4116 24734
rect 4060 24164 4116 24668
rect 4508 24722 4564 24892
rect 4508 24670 4510 24722
rect 4562 24670 4564 24722
rect 4508 24658 4564 24670
rect 4956 24948 5012 24958
rect 4614 24332 4878 24342
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4614 24266 4878 24276
rect 4060 24098 4116 24108
rect 4620 24164 4676 24174
rect 4620 24050 4676 24108
rect 4620 23998 4622 24050
rect 4674 23998 4676 24050
rect 4620 23986 4676 23998
rect 4956 23604 5012 24892
rect 5068 23940 5124 25004
rect 5516 24948 5572 25228
rect 5628 25218 5684 25228
rect 5180 24892 5572 24948
rect 5740 24948 5796 24958
rect 5180 24834 5236 24892
rect 5180 24782 5182 24834
rect 5234 24782 5236 24834
rect 5180 24770 5236 24782
rect 5740 24050 5796 24892
rect 5740 23998 5742 24050
rect 5794 23998 5796 24050
rect 5740 23986 5796 23998
rect 5068 23884 5348 23940
rect 5068 23714 5124 23726
rect 5068 23662 5070 23714
rect 5122 23662 5124 23714
rect 5068 23604 5124 23662
rect 5012 23548 5124 23604
rect 4956 23538 5012 23548
rect 4620 23380 4676 23390
rect 4620 23286 4676 23324
rect 3836 23214 3838 23266
rect 3890 23214 3892 23266
rect 3388 23154 3668 23156
rect 3388 23102 3390 23154
rect 3442 23102 3668 23154
rect 3388 23100 3668 23102
rect 3388 23090 3444 23100
rect 3276 22876 3444 22932
rect 3276 22260 3332 22270
rect 3276 21698 3332 22204
rect 3276 21646 3278 21698
rect 3330 21646 3332 21698
rect 3276 21634 3332 21646
rect 3052 21534 3054 21586
rect 3106 21534 3108 21586
rect 3052 21522 3108 21534
rect 3052 21252 3108 21262
rect 3052 21026 3108 21196
rect 3052 20974 3054 21026
rect 3106 20974 3108 21026
rect 2604 19966 2606 20018
rect 2658 19966 2660 20018
rect 2492 19348 2548 19358
rect 2380 19346 2548 19348
rect 2380 19294 2494 19346
rect 2546 19294 2548 19346
rect 2380 19292 2548 19294
rect 2492 19282 2548 19292
rect 1820 16830 1822 16882
rect 1874 16830 1876 16882
rect 1820 16818 1876 16830
rect 1932 18732 2324 18788
rect 1820 16098 1876 16110
rect 1820 16046 1822 16098
rect 1874 16046 1876 16098
rect 1820 15540 1876 16046
rect 1820 15446 1876 15484
rect 1820 12962 1876 12974
rect 1820 12910 1822 12962
rect 1874 12910 1876 12962
rect 1708 12852 1764 12862
rect 1708 12178 1764 12796
rect 1708 12126 1710 12178
rect 1762 12126 1764 12178
rect 1708 8372 1764 12126
rect 1820 10836 1876 12910
rect 1820 9826 1876 10780
rect 1820 9774 1822 9826
rect 1874 9774 1876 9826
rect 1820 9762 1876 9774
rect 1932 9156 1988 18732
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 2044 17668 2100 18510
rect 2604 18564 2660 19966
rect 2716 20804 2772 20814
rect 2716 20020 2772 20748
rect 2940 20578 2996 20590
rect 2940 20526 2942 20578
rect 2994 20526 2996 20578
rect 2716 19954 2772 19964
rect 2828 20020 2884 20030
rect 2940 20020 2996 20526
rect 3052 20356 3108 20974
rect 3388 20804 3444 22876
rect 3500 22036 3556 22046
rect 3500 21586 3556 21980
rect 3500 21534 3502 21586
rect 3554 21534 3556 21586
rect 3500 21028 3556 21534
rect 3612 21924 3668 23100
rect 3724 22930 3780 22942
rect 3724 22878 3726 22930
rect 3778 22878 3780 22930
rect 3724 22260 3780 22878
rect 3836 22596 3892 23214
rect 4508 23156 4564 23166
rect 4508 23062 4564 23100
rect 4614 22764 4878 22774
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4614 22698 4878 22708
rect 3836 22530 3892 22540
rect 4620 22596 4676 22606
rect 4620 22482 4676 22540
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 4620 22418 4676 22430
rect 3724 22194 3780 22204
rect 4396 22148 4452 22158
rect 3612 21868 4004 21924
rect 3612 21252 3668 21868
rect 3948 21810 4004 21868
rect 3948 21758 3950 21810
rect 4002 21758 4004 21810
rect 3948 21746 4004 21758
rect 4396 21810 4452 22092
rect 4396 21758 4398 21810
rect 4450 21758 4452 21810
rect 4396 21746 4452 21758
rect 5068 22146 5124 23548
rect 5068 22094 5070 22146
rect 5122 22094 5124 22146
rect 5068 21586 5124 22094
rect 5068 21534 5070 21586
rect 5122 21534 5124 21586
rect 3612 21186 3668 21196
rect 4614 21196 4878 21206
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4614 21130 4878 21140
rect 3500 20972 3780 21028
rect 3500 20804 3556 20814
rect 3612 20804 3668 20814
rect 3388 20802 3668 20804
rect 3388 20750 3502 20802
rect 3554 20750 3614 20802
rect 3666 20750 3668 20802
rect 3388 20748 3668 20750
rect 3500 20738 3556 20748
rect 3612 20738 3668 20748
rect 3388 20580 3444 20590
rect 3052 20290 3108 20300
rect 3164 20578 3444 20580
rect 3164 20526 3390 20578
rect 3442 20526 3444 20578
rect 3164 20524 3444 20526
rect 3052 20132 3108 20142
rect 3164 20132 3220 20524
rect 3388 20514 3444 20524
rect 3388 20356 3444 20366
rect 3052 20130 3220 20132
rect 3052 20078 3054 20130
rect 3106 20078 3220 20130
rect 3052 20076 3220 20078
rect 3276 20132 3332 20142
rect 3052 20066 3108 20076
rect 3276 20038 3332 20076
rect 2828 20018 2996 20020
rect 2828 19966 2830 20018
rect 2882 19966 2996 20018
rect 2828 19964 2996 19966
rect 2828 19954 2884 19964
rect 3388 19796 3444 20300
rect 3276 19740 3444 19796
rect 3500 20132 3556 20142
rect 3724 20132 3780 20972
rect 4284 21026 4340 21038
rect 4284 20974 4286 21026
rect 4338 20974 4340 21026
rect 3948 20580 4004 20590
rect 3556 20076 3780 20132
rect 3836 20578 4004 20580
rect 3836 20526 3950 20578
rect 4002 20526 4004 20578
rect 3836 20524 4004 20526
rect 3276 18676 3332 19740
rect 3500 19684 3556 20076
rect 2492 18338 2548 18350
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 2492 18228 2548 18286
rect 2492 18162 2548 18172
rect 2044 17602 2100 17612
rect 2492 16772 2548 16782
rect 2380 16770 2548 16772
rect 2380 16718 2494 16770
rect 2546 16718 2548 16770
rect 2380 16716 2548 16718
rect 2044 15876 2100 15886
rect 2380 15876 2436 16716
rect 2492 16706 2548 16716
rect 2604 16098 2660 18508
rect 2604 16046 2606 16098
rect 2658 16046 2660 16098
rect 2492 15876 2548 15886
rect 2044 15874 2324 15876
rect 2044 15822 2046 15874
rect 2098 15822 2324 15874
rect 2044 15820 2324 15822
rect 2380 15874 2548 15876
rect 2380 15822 2494 15874
rect 2546 15822 2548 15874
rect 2380 15820 2548 15822
rect 2044 15810 2100 15820
rect 2044 15204 2100 15214
rect 2044 15092 2212 15148
rect 2044 14980 2100 14990
rect 2044 14642 2100 14924
rect 2044 14590 2046 14642
rect 2098 14590 2100 14642
rect 2044 14578 2100 14590
rect 2156 14532 2212 15092
rect 2268 14756 2324 15820
rect 2492 15810 2548 15820
rect 2604 15204 2660 16046
rect 2604 15138 2660 15148
rect 2716 18674 3332 18676
rect 2716 18622 3278 18674
rect 3330 18622 3332 18674
rect 2716 18620 3332 18622
rect 2716 17890 2772 18620
rect 3276 18610 3332 18620
rect 3388 19628 3556 19684
rect 3836 19908 3892 20524
rect 3948 20514 4004 20524
rect 3948 20020 4004 20030
rect 3948 19926 4004 19964
rect 3388 18004 3444 19628
rect 3836 18564 3892 19852
rect 4284 19460 4340 20974
rect 4844 21026 4900 21038
rect 4844 20974 4846 21026
rect 4898 20974 4900 21026
rect 4844 20914 4900 20974
rect 4844 20862 4846 20914
rect 4898 20862 4900 20914
rect 4844 20850 4900 20862
rect 5068 20916 5124 21534
rect 4396 20578 4452 20590
rect 4396 20526 4398 20578
rect 4450 20526 4452 20578
rect 4396 20132 4452 20526
rect 4396 20066 4452 20076
rect 4956 19908 5012 19918
rect 4508 19796 4564 19834
rect 4956 19814 5012 19852
rect 4508 19730 4564 19740
rect 4614 19628 4878 19638
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4614 19562 4878 19572
rect 4284 19404 4676 19460
rect 4620 19346 4676 19404
rect 4620 19294 4622 19346
rect 4674 19294 4676 19346
rect 4620 19282 4676 19294
rect 3836 18498 3892 18508
rect 5068 19010 5124 20860
rect 5068 18958 5070 19010
rect 5122 18958 5124 19010
rect 3724 18452 3780 18462
rect 2716 17838 2718 17890
rect 2770 17838 2772 17890
rect 2716 15876 2772 17838
rect 3276 17948 3444 18004
rect 3500 18396 3724 18452
rect 2940 17668 2996 17678
rect 2940 17554 2996 17612
rect 2940 17502 2942 17554
rect 2994 17502 2996 17554
rect 2940 17490 2996 17502
rect 2828 17442 2884 17454
rect 2828 17390 2830 17442
rect 2882 17390 2884 17442
rect 2828 16322 2884 17390
rect 2828 16270 2830 16322
rect 2882 16270 2884 16322
rect 2828 16258 2884 16270
rect 3052 17444 3108 17454
rect 3052 16098 3108 17388
rect 3052 16046 3054 16098
rect 3106 16046 3108 16098
rect 3052 16034 3108 16046
rect 3276 15986 3332 17948
rect 3500 17778 3556 18396
rect 3724 18358 3780 18396
rect 4396 18452 4452 18462
rect 3500 17726 3502 17778
rect 3554 17726 3556 17778
rect 3500 17714 3556 17726
rect 4172 17668 4228 17678
rect 4172 17574 4228 17612
rect 3388 17444 3444 17454
rect 3388 17350 3444 17388
rect 4396 16772 4452 18396
rect 4956 18340 5012 18350
rect 4614 18060 4878 18070
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4614 17994 4878 18004
rect 4732 17444 4788 17454
rect 4956 17444 5012 18284
rect 4732 17442 5012 17444
rect 4732 17390 4734 17442
rect 4786 17390 5012 17442
rect 4732 17388 5012 17390
rect 4732 17378 4788 17388
rect 4620 16772 4676 16782
rect 4396 16770 4676 16772
rect 4396 16718 4622 16770
rect 4674 16718 4676 16770
rect 4396 16716 4676 16718
rect 4620 16706 4676 16716
rect 4614 16492 4878 16502
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4614 16426 4878 16436
rect 3276 15934 3278 15986
rect 3330 15934 3332 15986
rect 2716 15820 3108 15876
rect 2268 14690 2324 14700
rect 2380 14980 2436 14990
rect 2268 14532 2324 14542
rect 2156 14530 2324 14532
rect 2156 14478 2270 14530
rect 2322 14478 2324 14530
rect 2156 14476 2324 14478
rect 2044 12290 2100 12302
rect 2044 12238 2046 12290
rect 2098 12238 2100 12290
rect 2044 11396 2100 12238
rect 2156 11396 2212 14476
rect 2268 14466 2324 14476
rect 2268 13972 2324 13982
rect 2268 13878 2324 13916
rect 2380 13636 2436 14924
rect 2716 14980 2772 15820
rect 3052 15538 3108 15820
rect 3052 15486 3054 15538
rect 3106 15486 3108 15538
rect 3052 15474 3108 15486
rect 2716 14914 2772 14924
rect 3164 15092 3220 15102
rect 3276 15092 3332 15934
rect 3724 15876 3780 15886
rect 3500 15874 3780 15876
rect 3500 15822 3726 15874
rect 3778 15822 3780 15874
rect 3500 15820 3780 15822
rect 3500 15538 3556 15820
rect 3724 15810 3780 15820
rect 4172 15874 4228 15886
rect 4172 15822 4174 15874
rect 4226 15822 4228 15874
rect 3500 15486 3502 15538
rect 3554 15486 3556 15538
rect 3500 15204 3556 15486
rect 3500 15138 3556 15148
rect 3836 15204 3892 15214
rect 3164 15090 3332 15092
rect 3164 15038 3166 15090
rect 3218 15038 3332 15090
rect 3164 15036 3332 15038
rect 2492 14532 2548 14542
rect 2492 13860 2548 14476
rect 2604 14532 2660 14542
rect 2604 14530 2772 14532
rect 2604 14478 2606 14530
rect 2658 14478 2772 14530
rect 2604 14476 2772 14478
rect 2604 14466 2660 14476
rect 2492 13794 2548 13804
rect 2604 14306 2660 14318
rect 2604 14254 2606 14306
rect 2658 14254 2660 14306
rect 2492 13636 2548 13646
rect 2380 13634 2548 13636
rect 2380 13582 2494 13634
rect 2546 13582 2548 13634
rect 2380 13580 2548 13582
rect 2380 12404 2436 13580
rect 2492 13570 2548 13580
rect 2492 13076 2548 13086
rect 2604 13076 2660 14254
rect 2716 14084 2772 14476
rect 2828 14420 2884 14430
rect 2828 14326 2884 14364
rect 3052 14420 3108 14430
rect 3164 14420 3220 15036
rect 3612 14530 3668 14542
rect 3612 14478 3614 14530
rect 3666 14478 3668 14530
rect 3052 14418 3220 14420
rect 3052 14366 3054 14418
rect 3106 14366 3220 14418
rect 3052 14364 3220 14366
rect 3276 14420 3332 14430
rect 2716 14028 2884 14084
rect 2716 13860 2772 13870
rect 2716 13766 2772 13804
rect 2828 13634 2884 14028
rect 2828 13582 2830 13634
rect 2882 13582 2884 13634
rect 2828 13570 2884 13582
rect 3052 13636 3108 14364
rect 3276 13970 3332 14364
rect 3276 13918 3278 13970
rect 3330 13918 3332 13970
rect 3276 13906 3332 13918
rect 3388 13972 3444 13982
rect 3388 13636 3444 13916
rect 3612 13860 3668 14478
rect 3612 13794 3668 13804
rect 3052 13580 3220 13636
rect 2492 13074 2660 13076
rect 2492 13022 2494 13074
rect 2546 13022 2660 13074
rect 2492 13020 2660 13022
rect 2492 13010 2548 13020
rect 2380 12290 2436 12348
rect 2604 12292 2660 12302
rect 2380 12238 2382 12290
rect 2434 12238 2436 12290
rect 2380 12226 2436 12238
rect 2492 12290 2660 12292
rect 2492 12238 2606 12290
rect 2658 12238 2660 12290
rect 2492 12236 2660 12238
rect 2492 11844 2548 12236
rect 2604 12226 2660 12236
rect 2716 12180 2772 12190
rect 2380 11788 2548 11844
rect 2604 12066 2660 12078
rect 2604 12014 2606 12066
rect 2658 12014 2660 12066
rect 2268 11396 2324 11406
rect 2156 11394 2324 11396
rect 2156 11342 2270 11394
rect 2322 11342 2324 11394
rect 2156 11340 2324 11342
rect 2044 11330 2100 11340
rect 2044 11172 2100 11182
rect 2044 11078 2100 11116
rect 2268 10948 2324 11340
rect 2268 10882 2324 10892
rect 2156 10836 2212 10846
rect 2156 10724 2212 10780
rect 2268 10724 2324 10734
rect 2156 10722 2324 10724
rect 2156 10670 2270 10722
rect 2322 10670 2324 10722
rect 2156 10668 2324 10670
rect 1932 9090 1988 9100
rect 2044 10276 2100 10286
rect 1820 8372 1876 8382
rect 1708 8370 1876 8372
rect 1708 8318 1822 8370
rect 1874 8318 1876 8370
rect 1708 8316 1876 8318
rect 1820 8306 1876 8316
rect 2044 7698 2100 10220
rect 2156 8930 2212 8942
rect 2156 8878 2158 8930
rect 2210 8878 2212 8930
rect 2156 8372 2212 8878
rect 2156 8306 2212 8316
rect 2268 8258 2324 10668
rect 2380 10276 2436 11788
rect 2604 11618 2660 12014
rect 2604 11566 2606 11618
rect 2658 11566 2660 11618
rect 2604 11554 2660 11566
rect 2604 11172 2660 11182
rect 2380 10210 2436 10220
rect 2492 11170 2660 11172
rect 2492 11118 2606 11170
rect 2658 11118 2660 11170
rect 2492 11116 2660 11118
rect 2492 9938 2548 11116
rect 2604 11106 2660 11116
rect 2492 9886 2494 9938
rect 2546 9886 2548 9938
rect 2492 9874 2548 9886
rect 2604 10948 2660 10958
rect 2380 9156 2436 9166
rect 2380 9062 2436 9100
rect 2604 8484 2660 10892
rect 2716 10164 2772 12124
rect 3052 12180 3108 12190
rect 3052 12086 3108 12124
rect 3164 11788 3220 13580
rect 3388 13542 3444 13580
rect 3388 12292 3444 12302
rect 3388 12290 3556 12292
rect 3388 12238 3390 12290
rect 3442 12238 3556 12290
rect 3388 12236 3556 12238
rect 3388 12226 3444 12236
rect 3164 11732 3332 11788
rect 3276 11508 3332 11732
rect 3052 11452 3332 11508
rect 3052 11394 3108 11452
rect 3052 11342 3054 11394
rect 3106 11342 3108 11394
rect 3052 11330 3108 11342
rect 2828 11284 2884 11294
rect 2828 11190 2884 11228
rect 2716 10098 2772 10108
rect 2604 8418 2660 8428
rect 3164 9154 3220 11452
rect 3388 11394 3444 11406
rect 3388 11342 3390 11394
rect 3442 11342 3444 11394
rect 3388 10276 3444 11342
rect 3500 11396 3556 12236
rect 3500 11330 3556 11340
rect 3388 10210 3444 10220
rect 3164 9102 3166 9154
rect 3218 9102 3220 9154
rect 2268 8206 2270 8258
rect 2322 8206 2324 8258
rect 2268 8194 2324 8206
rect 2828 8372 2884 8382
rect 2044 7646 2046 7698
rect 2098 7646 2100 7698
rect 2044 7634 2100 7646
rect 2828 7698 2884 8316
rect 3164 8372 3220 9102
rect 3164 8306 3220 8316
rect 3724 8372 3780 8382
rect 2828 7646 2830 7698
rect 2882 7646 2884 7698
rect 2828 7588 2884 7646
rect 2940 8146 2996 8158
rect 2940 8094 2942 8146
rect 2994 8094 2996 8146
rect 2940 7700 2996 8094
rect 3724 7700 3780 8316
rect 2940 7634 2996 7644
rect 3388 7698 3780 7700
rect 3388 7646 3726 7698
rect 3778 7646 3780 7698
rect 3388 7644 3780 7646
rect 2828 7522 2884 7532
rect 1708 7476 1764 7486
rect 1708 7382 1764 7420
rect 2492 7476 2548 7486
rect 2492 6802 2548 7420
rect 2492 6750 2494 6802
rect 2546 6750 2548 6802
rect 2492 6738 2548 6750
rect 3276 7474 3332 7486
rect 3276 7422 3278 7474
rect 3330 7422 3332 7474
rect 3276 6580 3332 7422
rect 3388 6802 3444 7644
rect 3724 7634 3780 7644
rect 3836 7476 3892 15148
rect 3948 15204 4004 15214
rect 4172 15204 4228 15822
rect 3948 15202 4228 15204
rect 3948 15150 3950 15202
rect 4002 15150 4228 15202
rect 3948 15148 4228 15150
rect 4396 15202 4452 15214
rect 4396 15150 4398 15202
rect 4450 15150 4452 15202
rect 4396 15148 4452 15150
rect 3948 15090 4004 15148
rect 3948 15038 3950 15090
rect 4002 15038 4004 15090
rect 3948 15026 4004 15038
rect 4284 15092 4452 15148
rect 4172 14306 4228 14318
rect 4172 14254 4174 14306
rect 4226 14254 4228 14306
rect 4172 13634 4228 14254
rect 4172 13582 4174 13634
rect 4226 13582 4228 13634
rect 4172 13524 4228 13582
rect 4172 13458 4228 13468
rect 4060 12404 4116 12414
rect 3948 11620 4004 11630
rect 3948 11526 4004 11564
rect 4060 11284 4116 12348
rect 4284 12180 4340 15092
rect 4614 14924 4878 14934
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4614 14858 4878 14868
rect 4620 14420 4676 14430
rect 4620 14326 4676 14364
rect 4956 14420 5012 17388
rect 5068 17106 5124 18958
rect 5180 18450 5236 18462
rect 5180 18398 5182 18450
rect 5234 18398 5236 18450
rect 5180 17780 5236 18398
rect 5180 17714 5236 17724
rect 5068 17054 5070 17106
rect 5122 17054 5124 17106
rect 5068 17042 5124 17054
rect 5180 16884 5236 16894
rect 4956 14354 5012 14364
rect 5068 16828 5180 16884
rect 5068 14644 5124 16828
rect 5180 16818 5236 16828
rect 5292 16770 5348 23884
rect 5852 23548 5908 26684
rect 5964 25730 6020 27134
rect 5964 25678 5966 25730
rect 6018 25678 6020 25730
rect 5964 25666 6020 25678
rect 6076 26402 6132 28028
rect 6076 26350 6078 26402
rect 6130 26350 6132 26402
rect 6076 24948 6132 26350
rect 6188 26404 6244 30044
rect 6412 28866 6468 28878
rect 6412 28814 6414 28866
rect 6466 28814 6468 28866
rect 6412 28754 6468 28814
rect 6412 28702 6414 28754
rect 6466 28702 6468 28754
rect 6412 28690 6468 28702
rect 6524 28084 6580 31052
rect 7196 31042 7252 31054
rect 6972 30994 7028 31006
rect 6972 30942 6974 30994
rect 7026 30942 7028 30994
rect 6636 30884 6692 30894
rect 6972 30884 7028 30942
rect 6692 30828 7028 30884
rect 6636 30790 6692 30828
rect 6748 30324 6804 30334
rect 6748 28756 6804 30268
rect 6860 30324 6916 30828
rect 7308 30324 7364 32060
rect 7420 30548 7476 33964
rect 7532 33926 7588 33964
rect 7644 31332 7700 38780
rect 7868 37492 7924 39790
rect 8092 39732 8148 39742
rect 8204 39732 8260 40236
rect 8092 39730 8260 39732
rect 8092 39678 8094 39730
rect 8146 39678 8260 39730
rect 8092 39676 8260 39678
rect 8428 40402 8484 40414
rect 8428 40350 8430 40402
rect 8482 40350 8484 40402
rect 8428 40292 8484 40350
rect 8092 39666 8148 39676
rect 8016 39228 8280 39238
rect 8072 39172 8120 39228
rect 8176 39172 8224 39228
rect 8016 39162 8280 39172
rect 8428 38948 8484 40236
rect 8540 40404 8596 41918
rect 8540 39730 8596 40348
rect 8540 39678 8542 39730
rect 8594 39678 8596 39730
rect 8540 39666 8596 39678
rect 8540 38948 8596 38958
rect 8428 38892 8540 38948
rect 8540 38882 8596 38892
rect 8652 38668 8708 43820
rect 8988 41972 9044 44158
rect 8876 41970 9044 41972
rect 8876 41918 8990 41970
rect 9042 41918 9044 41970
rect 8876 41916 9044 41918
rect 8764 40178 8820 40190
rect 8764 40126 8766 40178
rect 8818 40126 8820 40178
rect 8764 39842 8820 40126
rect 8764 39790 8766 39842
rect 8818 39790 8820 39842
rect 8764 39778 8820 39790
rect 8540 38612 8708 38668
rect 8428 38164 8484 38174
rect 8016 37660 8280 37670
rect 8072 37604 8120 37660
rect 8176 37604 8224 37660
rect 8016 37594 8280 37604
rect 8204 37492 8260 37502
rect 7868 37436 8148 37492
rect 7756 37380 7812 37390
rect 7756 37378 8036 37380
rect 7756 37326 7758 37378
rect 7810 37326 8036 37378
rect 7756 37324 8036 37326
rect 7756 37314 7812 37324
rect 7980 37268 8036 37324
rect 7980 37202 8036 37212
rect 8092 36260 8148 37436
rect 8204 37044 8260 37436
rect 8428 37490 8484 38108
rect 8428 37438 8430 37490
rect 8482 37438 8484 37490
rect 8428 37426 8484 37438
rect 8316 37268 8372 37278
rect 8316 37174 8372 37212
rect 8204 36978 8260 36988
rect 8204 36820 8260 36830
rect 8204 36482 8260 36764
rect 8204 36430 8206 36482
rect 8258 36430 8260 36482
rect 8204 36418 8260 36430
rect 8428 36484 8484 36494
rect 8540 36484 8596 38612
rect 8764 37492 8820 37502
rect 8652 37380 8708 37390
rect 8652 36594 8708 37324
rect 8764 37266 8820 37436
rect 8764 37214 8766 37266
rect 8818 37214 8820 37266
rect 8764 37202 8820 37214
rect 8652 36542 8654 36594
rect 8706 36542 8708 36594
rect 8652 36530 8708 36542
rect 8428 36482 8596 36484
rect 8428 36430 8430 36482
rect 8482 36430 8596 36482
rect 8428 36428 8596 36430
rect 8428 36418 8484 36428
rect 7868 36204 8148 36260
rect 7868 35924 7924 36204
rect 8016 36092 8280 36102
rect 8072 36036 8120 36092
rect 8176 36036 8224 36092
rect 8016 36026 8280 36036
rect 8540 35924 8596 36428
rect 8876 36484 8932 41916
rect 8988 41906 9044 41916
rect 9100 44604 9268 44660
rect 8988 40404 9044 40414
rect 8988 39730 9044 40348
rect 8988 39678 8990 39730
rect 9042 39678 9044 39730
rect 8988 39666 9044 39678
rect 9100 38668 9156 44604
rect 9324 44548 9380 65660
rect 9660 65490 9716 65502
rect 9660 65438 9662 65490
rect 9714 65438 9716 65490
rect 9436 64820 9492 64830
rect 9436 63028 9492 64764
rect 9660 63924 9716 65438
rect 10220 64596 10276 67564
rect 10780 67060 10836 70700
rect 10892 70418 10948 73500
rect 11116 72660 11172 72670
rect 11004 71876 11060 71886
rect 11116 71876 11172 72604
rect 11228 72212 11284 74620
rect 11418 74508 11682 74518
rect 11474 74452 11522 74508
rect 11578 74452 11626 74508
rect 11418 74442 11682 74452
rect 11788 74452 11844 74846
rect 11900 74900 11956 75742
rect 11900 74834 11956 74844
rect 11788 74386 11844 74396
rect 11900 74564 11956 74574
rect 11788 74228 11844 74238
rect 11676 74004 11732 74042
rect 11676 73938 11732 73948
rect 11418 72940 11682 72950
rect 11474 72884 11522 72940
rect 11578 72884 11626 72940
rect 11418 72874 11682 72884
rect 11788 72324 11844 74172
rect 11228 72146 11284 72156
rect 11340 72268 11844 72324
rect 11340 71876 11396 72268
rect 11676 72100 11732 72110
rect 11676 71986 11732 72044
rect 11676 71934 11678 71986
rect 11730 71934 11732 71986
rect 11676 71922 11732 71934
rect 11788 71988 11844 72268
rect 11788 71922 11844 71932
rect 11564 71876 11620 71886
rect 11116 71820 11284 71876
rect 11340 71820 11508 71876
rect 11004 71782 11060 71820
rect 11228 71204 11284 71820
rect 11452 71762 11508 71820
rect 11564 71782 11620 71820
rect 11452 71710 11454 71762
rect 11506 71710 11508 71762
rect 11452 71698 11508 71710
rect 11418 71372 11682 71382
rect 11474 71316 11522 71372
rect 11578 71316 11626 71372
rect 11418 71306 11682 71316
rect 11228 71148 11396 71204
rect 11228 70980 11284 70990
rect 11228 70886 11284 70924
rect 10892 70366 10894 70418
rect 10946 70366 10948 70418
rect 10892 70308 10948 70366
rect 11340 70420 11396 71148
rect 11340 70326 11396 70364
rect 11788 70644 11844 70654
rect 10892 70242 10948 70252
rect 11418 69804 11682 69814
rect 11474 69748 11522 69804
rect 11578 69748 11626 69804
rect 11418 69738 11682 69748
rect 11788 69634 11844 70588
rect 11900 70308 11956 74508
rect 12012 70868 12068 78878
rect 12124 78818 12180 82460
rect 12460 81730 12516 89852
rect 12572 89796 12628 92652
rect 12684 92642 12740 92652
rect 12796 92372 12852 92382
rect 12684 91588 12740 91598
rect 12684 91474 12740 91532
rect 12684 91422 12686 91474
rect 12738 91422 12740 91474
rect 12684 91410 12740 91422
rect 12796 91362 12852 92316
rect 13580 92260 13636 93884
rect 13916 93874 13972 93884
rect 13692 93716 13748 93726
rect 13692 92930 13748 93660
rect 14028 93492 14084 93502
rect 13692 92878 13694 92930
rect 13746 92878 13748 92930
rect 13692 92866 13748 92878
rect 13804 93268 13860 93278
rect 13580 92194 13636 92204
rect 13468 92034 13524 92046
rect 13468 91982 13470 92034
rect 13522 91982 13524 92034
rect 12796 91310 12798 91362
rect 12850 91310 12852 91362
rect 12796 91298 12852 91310
rect 12908 91476 12964 91486
rect 12908 91250 12964 91420
rect 12908 91198 12910 91250
rect 12962 91198 12964 91250
rect 12908 91186 12964 91198
rect 13356 91138 13412 91150
rect 13356 91086 13358 91138
rect 13410 91086 13412 91138
rect 12684 90580 12740 90590
rect 12684 90486 12740 90524
rect 13356 90580 13412 91086
rect 13468 90804 13524 91982
rect 13580 91476 13636 91486
rect 13580 91250 13636 91420
rect 13580 91198 13582 91250
rect 13634 91198 13636 91250
rect 13580 91186 13636 91198
rect 13692 91252 13748 91262
rect 13692 91158 13748 91196
rect 13468 90738 13524 90748
rect 12908 90466 12964 90478
rect 12908 90414 12910 90466
rect 12962 90414 12964 90466
rect 12908 90020 12964 90414
rect 13356 90466 13412 90524
rect 13356 90414 13358 90466
rect 13410 90414 13412 90466
rect 13356 90402 13412 90414
rect 13468 90578 13524 90590
rect 13468 90526 13470 90578
rect 13522 90526 13524 90578
rect 12908 89954 12964 89964
rect 13468 90020 13524 90526
rect 13804 90132 13860 93212
rect 14028 93044 14084 93436
rect 13916 92988 14084 93044
rect 13916 92818 13972 92988
rect 13916 92766 13918 92818
rect 13970 92766 13972 92818
rect 13916 92754 13972 92766
rect 14028 92818 14084 92830
rect 14028 92766 14030 92818
rect 14082 92766 14084 92818
rect 14028 92484 14084 92766
rect 14028 92418 14084 92428
rect 14028 90692 14084 90702
rect 14140 90692 14196 94670
rect 14252 93940 14308 95788
rect 14364 95778 14420 95788
rect 14588 95396 14644 97468
rect 14820 97244 15084 97254
rect 14876 97188 14924 97244
rect 14980 97188 15028 97244
rect 14820 97178 15084 97188
rect 14700 96796 15092 96852
rect 14700 96180 14756 96796
rect 15036 96738 15092 96796
rect 15036 96686 15038 96738
rect 15090 96686 15092 96738
rect 15036 96674 15092 96686
rect 15148 96850 15204 96862
rect 15148 96798 15150 96850
rect 15202 96798 15204 96850
rect 15148 96628 15204 96798
rect 15148 96562 15204 96572
rect 14700 96086 14756 96124
rect 15372 96404 15428 96414
rect 15484 96404 15540 99036
rect 15596 98418 15652 100604
rect 15596 98366 15598 98418
rect 15650 98366 15652 98418
rect 15596 98354 15652 98366
rect 15596 97636 15652 97646
rect 15596 96516 15652 97580
rect 15708 96962 15764 105868
rect 15820 104356 15876 105982
rect 15932 105588 15988 106206
rect 16268 106146 16324 107772
rect 16716 107826 16772 107996
rect 16716 107774 16718 107826
rect 16770 107774 16772 107826
rect 16716 107762 16772 107774
rect 16828 107828 16884 107838
rect 16828 106482 16884 107772
rect 16828 106430 16830 106482
rect 16882 106430 16884 106482
rect 16828 106418 16884 106430
rect 16268 106094 16270 106146
rect 16322 106094 16324 106146
rect 16268 105812 16324 106094
rect 16492 106036 16548 106046
rect 16492 105942 16548 105980
rect 16268 105756 16548 105812
rect 16380 105588 16436 105598
rect 15932 105586 16436 105588
rect 15932 105534 16382 105586
rect 16434 105534 16436 105586
rect 15932 105532 16436 105534
rect 16380 105522 16436 105532
rect 15820 104290 15876 104300
rect 16044 104244 16100 104254
rect 15932 98196 15988 98206
rect 15932 97636 15988 98140
rect 15932 97542 15988 97580
rect 15708 96910 15710 96962
rect 15762 96910 15764 96962
rect 15708 96740 15764 96910
rect 15708 96684 15988 96740
rect 15596 96450 15652 96460
rect 15820 96516 15876 96526
rect 15428 96348 15540 96404
rect 14812 96066 14868 96078
rect 14812 96014 14814 96066
rect 14866 96014 14868 96066
rect 14812 95956 14868 96014
rect 14812 95890 14868 95900
rect 15372 95954 15428 96348
rect 15372 95902 15374 95954
rect 15426 95902 15428 95954
rect 15372 95890 15428 95902
rect 15596 96292 15652 96302
rect 15260 95844 15316 95854
rect 15148 95788 15260 95844
rect 14820 95676 15084 95686
rect 14876 95620 14924 95676
rect 14980 95620 15028 95676
rect 14820 95610 15084 95620
rect 14812 95508 14868 95518
rect 15148 95508 15204 95788
rect 15260 95778 15316 95788
rect 14588 95340 14756 95396
rect 14476 95282 14532 95294
rect 14476 95230 14478 95282
rect 14530 95230 14532 95282
rect 14364 95060 14420 95070
rect 14364 94610 14420 95004
rect 14364 94558 14366 94610
rect 14418 94558 14420 94610
rect 14364 94164 14420 94558
rect 14364 94098 14420 94108
rect 14364 93940 14420 93950
rect 14252 93938 14420 93940
rect 14252 93886 14366 93938
rect 14418 93886 14420 93938
rect 14252 93884 14420 93886
rect 14364 93874 14420 93884
rect 14252 93716 14308 93726
rect 14252 93622 14308 93660
rect 14476 93268 14532 95230
rect 14700 95282 14756 95340
rect 14700 95230 14702 95282
rect 14754 95230 14756 95282
rect 14700 95218 14756 95230
rect 14588 95170 14644 95182
rect 14588 95118 14590 95170
rect 14642 95118 14644 95170
rect 14588 95060 14644 95118
rect 14588 95004 14756 95060
rect 14700 94500 14756 95004
rect 14700 94434 14756 94444
rect 14588 94386 14644 94398
rect 14588 94334 14590 94386
rect 14642 94334 14644 94386
rect 14588 93940 14644 94334
rect 14812 94276 14868 95452
rect 15036 95452 15204 95508
rect 15596 95506 15652 96236
rect 15820 96180 15876 96460
rect 15708 96124 15876 96180
rect 15708 95842 15764 96124
rect 15932 96066 15988 96684
rect 15932 96014 15934 96066
rect 15986 96014 15988 96066
rect 15932 96002 15988 96014
rect 15708 95790 15710 95842
rect 15762 95790 15764 95842
rect 15708 95778 15764 95790
rect 15820 95844 15876 95854
rect 15820 95750 15876 95788
rect 15596 95454 15598 95506
rect 15650 95454 15652 95506
rect 15036 95394 15092 95452
rect 15596 95442 15652 95454
rect 15932 95732 15988 95742
rect 15036 95342 15038 95394
rect 15090 95342 15092 95394
rect 15036 95330 15092 95342
rect 15932 95394 15988 95676
rect 15932 95342 15934 95394
rect 15986 95342 15988 95394
rect 15372 95282 15428 95294
rect 15372 95230 15374 95282
rect 15426 95230 15428 95282
rect 15372 95172 15428 95230
rect 15596 95284 15652 95294
rect 15596 95190 15652 95228
rect 15372 95106 15428 95116
rect 15932 95060 15988 95342
rect 15932 94994 15988 95004
rect 16044 94948 16100 104188
rect 16492 103236 16548 105756
rect 17164 104020 17220 108668
rect 17388 108658 17444 108668
rect 17276 108386 17332 108398
rect 17276 108334 17278 108386
rect 17330 108334 17332 108386
rect 17276 106036 17332 108334
rect 17500 108386 17556 108398
rect 17500 108334 17502 108386
rect 17554 108334 17556 108386
rect 17500 108164 17556 108334
rect 17500 108098 17556 108108
rect 17388 107940 17444 107950
rect 17388 107938 17556 107940
rect 17388 107886 17390 107938
rect 17442 107886 17556 107938
rect 17388 107884 17556 107886
rect 17388 107874 17444 107884
rect 17500 106258 17556 107884
rect 17500 106206 17502 106258
rect 17554 106206 17556 106258
rect 17500 106194 17556 106206
rect 17388 106036 17444 106046
rect 17276 105980 17388 106036
rect 17164 103954 17220 103964
rect 16492 103170 16548 103180
rect 16828 103908 16884 103918
rect 16156 103122 16212 103134
rect 16156 103070 16158 103122
rect 16210 103070 16212 103122
rect 16156 95508 16212 103070
rect 16828 102450 16884 103852
rect 17388 103348 17444 105980
rect 17612 105588 17668 116956
rect 17724 116452 17780 116462
rect 17836 116452 17892 117742
rect 18396 117234 18452 117246
rect 18396 117182 18398 117234
rect 18450 117182 18452 117234
rect 18396 117012 18452 117182
rect 18396 116956 18676 117012
rect 18222 116844 18486 116854
rect 18278 116788 18326 116844
rect 18382 116788 18430 116844
rect 18222 116778 18486 116788
rect 18620 116562 18676 116956
rect 18620 116510 18622 116562
rect 18674 116510 18676 116562
rect 17780 116396 17892 116452
rect 18396 116452 18452 116462
rect 18620 116452 18676 116510
rect 18452 116396 18676 116452
rect 17724 116358 17780 116396
rect 18396 116386 18452 116396
rect 18396 115668 18452 115678
rect 18620 115668 18676 116396
rect 18396 115666 18676 115668
rect 18396 115614 18398 115666
rect 18450 115614 18676 115666
rect 18396 115612 18676 115614
rect 18396 115602 18452 115612
rect 18222 115276 18486 115286
rect 18278 115220 18326 115276
rect 18382 115220 18430 115276
rect 18222 115210 18486 115220
rect 18620 114996 18676 115612
rect 18060 114884 18116 114894
rect 18060 114790 18116 114828
rect 18508 114660 18564 114670
rect 18620 114660 18676 114940
rect 18508 114658 18676 114660
rect 18508 114606 18510 114658
rect 18562 114606 18676 114658
rect 18508 114604 18676 114606
rect 18508 114268 18564 114604
rect 19292 114268 19348 119600
rect 19404 118018 19460 118030
rect 19404 117966 19406 118018
rect 19458 117966 19460 118018
rect 19404 117012 19460 117966
rect 20076 118018 20132 118030
rect 20076 117966 20078 118018
rect 20130 117966 20132 118018
rect 20076 117234 20132 117966
rect 20860 117796 20916 117806
rect 20076 117182 20078 117234
rect 20130 117182 20132 117234
rect 19516 117012 19572 117022
rect 19404 117010 19908 117012
rect 19404 116958 19518 117010
rect 19570 116958 19908 117010
rect 19404 116956 19908 116958
rect 19516 116946 19572 116956
rect 19852 116562 19908 116956
rect 19852 116510 19854 116562
rect 19906 116510 19908 116562
rect 19740 115892 19796 115902
rect 19852 115892 19908 116510
rect 19740 115890 19908 115892
rect 19740 115838 19742 115890
rect 19794 115838 19908 115890
rect 19740 115836 19908 115838
rect 19740 115826 19796 115836
rect 19852 114994 19908 115836
rect 19852 114942 19854 114994
rect 19906 114942 19908 114994
rect 19852 114268 19908 114942
rect 18172 114212 18564 114268
rect 18732 114212 19348 114268
rect 19516 114212 19908 114268
rect 20076 115666 20132 117182
rect 20748 117794 20916 117796
rect 20748 117742 20862 117794
rect 20914 117742 20916 117794
rect 20748 117740 20916 117742
rect 20748 117234 20804 117740
rect 20860 117730 20916 117740
rect 20748 117182 20750 117234
rect 20802 117182 20804 117234
rect 20300 116228 20356 116238
rect 20748 116228 20804 117182
rect 20300 116226 20916 116228
rect 20300 116174 20302 116226
rect 20354 116174 20750 116226
rect 20802 116174 20916 116226
rect 20300 116172 20916 116174
rect 20300 116162 20356 116172
rect 20748 116162 20804 116172
rect 20076 115614 20078 115666
rect 20130 115614 20132 115666
rect 20076 114884 20132 115614
rect 20076 114324 20132 114828
rect 18172 114100 18228 114212
rect 18060 114098 18228 114100
rect 18060 114046 18174 114098
rect 18226 114046 18228 114098
rect 18060 114044 18228 114046
rect 18060 111748 18116 114044
rect 18172 114034 18228 114044
rect 18222 113708 18486 113718
rect 18278 113652 18326 113708
rect 18382 113652 18430 113708
rect 18222 113642 18486 113652
rect 18620 113316 18676 113326
rect 18620 113222 18676 113260
rect 18222 112140 18486 112150
rect 18278 112084 18326 112140
rect 18382 112084 18430 112140
rect 18222 112074 18486 112084
rect 18172 111748 18228 111758
rect 18060 111692 18172 111748
rect 18172 110962 18228 111692
rect 18172 110910 18174 110962
rect 18226 110910 18228 110962
rect 18172 110898 18228 110910
rect 18222 110572 18486 110582
rect 18278 110516 18326 110572
rect 18382 110516 18430 110572
rect 18222 110506 18486 110516
rect 18732 109508 18788 114212
rect 19516 113874 19572 114212
rect 19516 113822 19518 113874
rect 19570 113822 19572 113874
rect 19180 113316 19236 113326
rect 19180 112530 19236 113260
rect 19180 112478 19182 112530
rect 19234 112478 19236 112530
rect 19180 112466 19236 112478
rect 19292 113316 19348 113326
rect 19516 113316 19572 113822
rect 19292 113314 19572 113316
rect 19292 113262 19294 113314
rect 19346 113262 19572 113314
rect 19292 113260 19572 113262
rect 20076 114098 20132 114268
rect 20076 114046 20078 114098
rect 20130 114046 20132 114098
rect 20076 113316 20132 114046
rect 19292 112532 19348 113260
rect 18956 111748 19012 111758
rect 19292 111748 19348 112476
rect 19964 112532 20020 112542
rect 19964 112438 20020 112476
rect 19012 111746 19572 111748
rect 19012 111694 19294 111746
rect 19346 111694 19572 111746
rect 19012 111692 19572 111694
rect 18956 111654 19012 111692
rect 19292 111682 19348 111692
rect 19516 110740 19572 111692
rect 20076 110964 20132 113260
rect 20860 115666 20916 116172
rect 20860 115614 20862 115666
rect 20914 115614 20916 115666
rect 20860 114098 20916 115614
rect 20860 114046 20862 114098
rect 20914 114046 20916 114098
rect 20860 113092 20916 114046
rect 20748 113090 20916 113092
rect 20748 113038 20862 113090
rect 20914 113038 20916 113090
rect 20748 113036 20916 113038
rect 20748 110964 20804 113036
rect 20860 113026 20916 113036
rect 20076 110870 20132 110908
rect 20636 110962 20804 110964
rect 20636 110910 20750 110962
rect 20802 110910 20804 110962
rect 20636 110908 20804 110910
rect 19516 110738 19908 110740
rect 19516 110686 19518 110738
rect 19570 110686 19908 110738
rect 19516 110684 19908 110686
rect 19516 110674 19572 110684
rect 19852 110292 19908 110684
rect 19852 110290 20132 110292
rect 19852 110238 19854 110290
rect 19906 110238 20132 110290
rect 19852 110236 20132 110238
rect 19852 110226 19908 110236
rect 18620 109452 18788 109508
rect 19404 109954 19460 109966
rect 19404 109902 19406 109954
rect 19458 109902 19460 109954
rect 18172 109284 18228 109294
rect 17836 109282 18228 109284
rect 17836 109230 18174 109282
rect 18226 109230 18228 109282
rect 17836 109228 18228 109230
rect 17836 108610 17892 109228
rect 18172 109218 18228 109228
rect 18222 109004 18486 109014
rect 18278 108948 18326 109004
rect 18382 108948 18430 109004
rect 18222 108938 18486 108948
rect 17836 108558 17838 108610
rect 17890 108558 17892 108610
rect 17724 107826 17780 107838
rect 17724 107774 17726 107826
rect 17778 107774 17780 107826
rect 17724 107044 17780 107774
rect 17724 106978 17780 106988
rect 17724 106820 17780 106830
rect 17724 106726 17780 106764
rect 17612 105522 17668 105532
rect 17612 104578 17668 104590
rect 17612 104526 17614 104578
rect 17666 104526 17668 104578
rect 17500 103796 17556 103806
rect 17500 103702 17556 103740
rect 17500 103348 17556 103358
rect 17388 103346 17556 103348
rect 17388 103294 17502 103346
rect 17554 103294 17556 103346
rect 17388 103292 17556 103294
rect 17500 103282 17556 103292
rect 16828 102398 16830 102450
rect 16882 102398 16884 102450
rect 16828 102386 16884 102398
rect 17276 103122 17332 103134
rect 17276 103070 17278 103122
rect 17330 103070 17332 103122
rect 16716 99204 16772 99214
rect 16604 97634 16660 97646
rect 16604 97582 16606 97634
rect 16658 97582 16660 97634
rect 16492 97300 16548 97310
rect 16380 97188 16436 97198
rect 16380 96852 16436 97132
rect 16268 96738 16324 96750
rect 16268 96686 16270 96738
rect 16322 96686 16324 96738
rect 16268 96292 16324 96686
rect 16268 96226 16324 96236
rect 16380 96066 16436 96796
rect 16492 96850 16548 97244
rect 16492 96798 16494 96850
rect 16546 96798 16548 96850
rect 16492 96786 16548 96798
rect 16380 96014 16382 96066
rect 16434 96014 16436 96066
rect 16380 96002 16436 96014
rect 16604 96068 16660 97582
rect 16716 97522 16772 99148
rect 16716 97470 16718 97522
rect 16770 97470 16772 97522
rect 16716 97458 16772 97470
rect 17276 97468 17332 103070
rect 17612 102452 17668 104526
rect 17500 101780 17556 101790
rect 17612 101780 17668 102396
rect 17500 101778 17668 101780
rect 17500 101726 17502 101778
rect 17554 101726 17668 101778
rect 17500 101724 17668 101726
rect 17724 103122 17780 103134
rect 17724 103070 17726 103122
rect 17778 103070 17780 103122
rect 17500 101714 17556 101724
rect 17500 100772 17556 100782
rect 17052 97412 17332 97468
rect 17388 98980 17444 98990
rect 17388 97748 17444 98924
rect 17500 98196 17556 100716
rect 17500 98140 17668 98196
rect 17388 97522 17444 97692
rect 17388 97470 17390 97522
rect 17442 97470 17444 97522
rect 16604 96002 16660 96012
rect 16716 97076 16772 97086
rect 16940 97076 16996 97086
rect 16716 96180 16772 97020
rect 16828 97020 16940 97076
rect 16828 96738 16884 97020
rect 16940 97010 16996 97020
rect 16828 96686 16830 96738
rect 16882 96686 16884 96738
rect 16828 96674 16884 96686
rect 16716 95732 16772 96124
rect 16716 95666 16772 95676
rect 16268 95508 16324 95518
rect 16156 95452 16268 95508
rect 16268 95394 16324 95452
rect 16828 95508 16884 95518
rect 16828 95414 16884 95452
rect 16268 95342 16270 95394
rect 16322 95342 16324 95394
rect 16268 95330 16324 95342
rect 16380 95284 16436 95294
rect 16044 94892 16324 94948
rect 14924 94836 14980 94846
rect 14980 94780 15092 94836
rect 14924 94770 14980 94780
rect 15036 94500 15092 94780
rect 15596 94500 15652 94510
rect 14588 93874 14644 93884
rect 14700 94220 14868 94276
rect 14924 94386 14980 94398
rect 14924 94334 14926 94386
rect 14978 94334 14980 94386
rect 14924 94276 14980 94334
rect 15036 94386 15092 94444
rect 15036 94334 15038 94386
rect 15090 94334 15092 94386
rect 15036 94322 15092 94334
rect 15372 94498 15652 94500
rect 15372 94446 15598 94498
rect 15650 94446 15652 94498
rect 15372 94444 15652 94446
rect 15260 94276 15316 94286
rect 14588 93716 14644 93726
rect 14700 93716 14756 94220
rect 14924 94210 14980 94220
rect 15148 94274 15316 94276
rect 15148 94222 15262 94274
rect 15314 94222 15316 94274
rect 15148 94220 15316 94222
rect 14820 94108 15084 94118
rect 14876 94052 14924 94108
rect 14980 94052 15028 94108
rect 14820 94042 15084 94052
rect 15148 93826 15204 94220
rect 15260 94210 15316 94220
rect 15148 93774 15150 93826
rect 15202 93774 15204 93826
rect 15148 93762 15204 93774
rect 15260 94052 15316 94062
rect 15260 93938 15316 93996
rect 15260 93886 15262 93938
rect 15314 93886 15316 93938
rect 14588 93714 14756 93716
rect 14588 93662 14590 93714
rect 14642 93662 14756 93714
rect 14588 93660 14756 93662
rect 14812 93714 14868 93726
rect 14812 93662 14814 93714
rect 14866 93662 14868 93714
rect 14588 93650 14644 93660
rect 14476 93202 14532 93212
rect 14588 92932 14644 92942
rect 14476 92930 14644 92932
rect 14476 92878 14590 92930
rect 14642 92878 14644 92930
rect 14476 92876 14644 92878
rect 14364 92820 14420 92830
rect 14364 92036 14420 92764
rect 14364 91970 14420 91980
rect 14476 91812 14532 92876
rect 14588 92866 14644 92876
rect 14812 92708 14868 93662
rect 15260 93380 15316 93886
rect 14924 93324 15316 93380
rect 14924 93154 14980 93324
rect 14924 93102 14926 93154
rect 14978 93102 14980 93154
rect 14924 93090 14980 93102
rect 14700 92652 14868 92708
rect 14252 91756 14532 91812
rect 14588 92260 14644 92270
rect 14252 91588 14308 91756
rect 14252 91250 14308 91532
rect 14588 91588 14644 92204
rect 14588 91474 14644 91532
rect 14588 91422 14590 91474
rect 14642 91422 14644 91474
rect 14588 91410 14644 91422
rect 14252 91198 14254 91250
rect 14306 91198 14308 91250
rect 14252 91186 14308 91198
rect 14700 91140 14756 92652
rect 14820 92540 15084 92550
rect 14876 92484 14924 92540
rect 14980 92484 15028 92540
rect 14820 92474 15084 92484
rect 15372 91476 15428 94444
rect 15596 94434 15652 94444
rect 15932 94500 15988 94510
rect 15708 94276 15764 94286
rect 15708 94274 15876 94276
rect 15708 94222 15710 94274
rect 15762 94222 15876 94274
rect 15708 94220 15876 94222
rect 15708 94210 15764 94220
rect 15484 93828 15540 93838
rect 15484 93826 15764 93828
rect 15484 93774 15486 93826
rect 15538 93774 15764 93826
rect 15484 93772 15764 93774
rect 15484 93762 15540 93772
rect 15708 93714 15764 93772
rect 15708 93662 15710 93714
rect 15762 93662 15764 93714
rect 15708 93650 15764 93662
rect 15820 93492 15876 94220
rect 15932 93828 15988 94444
rect 16156 94500 16212 94510
rect 16156 94406 16212 94444
rect 15932 93762 15988 93772
rect 16044 94276 16100 94286
rect 16044 93714 16100 94220
rect 16268 93938 16324 94892
rect 16380 94498 16436 95228
rect 16380 94446 16382 94498
rect 16434 94446 16436 94498
rect 16380 94434 16436 94446
rect 16492 95060 16548 95070
rect 16492 94388 16548 95004
rect 16604 94612 16660 94622
rect 16604 94610 16996 94612
rect 16604 94558 16606 94610
rect 16658 94558 16996 94610
rect 16604 94556 16996 94558
rect 16604 94546 16660 94556
rect 16940 94498 16996 94556
rect 16940 94446 16942 94498
rect 16994 94446 16996 94498
rect 16940 94434 16996 94446
rect 16716 94388 16772 94398
rect 16492 94386 16772 94388
rect 16492 94334 16718 94386
rect 16770 94334 16772 94386
rect 16492 94332 16772 94334
rect 16716 94322 16772 94332
rect 16268 93886 16270 93938
rect 16322 93886 16324 93938
rect 16268 93874 16324 93886
rect 16380 94052 16436 94062
rect 16380 93938 16436 93996
rect 16380 93886 16382 93938
rect 16434 93886 16436 93938
rect 16380 93874 16436 93886
rect 16044 93662 16046 93714
rect 16098 93662 16100 93714
rect 16044 93650 16100 93662
rect 16156 93714 16212 93726
rect 16156 93662 16158 93714
rect 16210 93662 16212 93714
rect 15932 93492 15988 93502
rect 15820 93436 15932 93492
rect 15932 93426 15988 93436
rect 15596 93268 15652 93278
rect 15596 93042 15652 93212
rect 15596 92990 15598 93042
rect 15650 92990 15652 93042
rect 15596 92978 15652 92990
rect 16156 93044 16212 93662
rect 15932 92820 15988 92830
rect 15596 92148 15652 92158
rect 15372 91410 15428 91420
rect 15484 92036 15540 92046
rect 15484 91364 15540 91980
rect 15484 91270 15540 91308
rect 14700 91074 14756 91084
rect 14820 90972 15084 90982
rect 14876 90916 14924 90972
rect 14980 90916 15028 90972
rect 14820 90906 15084 90916
rect 15484 90804 15540 90814
rect 14700 90692 14756 90702
rect 14028 90690 14756 90692
rect 14028 90638 14030 90690
rect 14082 90638 14702 90690
rect 14754 90638 14756 90690
rect 14028 90636 14756 90638
rect 14028 90626 14084 90636
rect 13804 90076 13972 90132
rect 13468 89954 13524 89964
rect 13580 89908 13636 89918
rect 12684 89796 12740 89806
rect 12572 89740 12684 89796
rect 12684 89730 12740 89740
rect 13580 89794 13636 89852
rect 13916 89906 13972 90076
rect 13916 89854 13918 89906
rect 13970 89854 13972 89906
rect 13916 89842 13972 89854
rect 14588 89908 14644 90636
rect 14700 90626 14756 90636
rect 14924 90692 14980 90702
rect 14924 90598 14980 90636
rect 15148 90580 15204 90590
rect 15148 90486 15204 90524
rect 15372 90578 15428 90590
rect 15372 90526 15374 90578
rect 15426 90526 15428 90578
rect 15372 90468 15428 90526
rect 15260 90412 15372 90468
rect 13580 89742 13582 89794
rect 13634 89742 13636 89794
rect 13580 89730 13636 89742
rect 13804 89796 13860 89806
rect 13692 89572 13748 89582
rect 13356 88900 13412 88910
rect 12908 88338 12964 88350
rect 12908 88286 12910 88338
rect 12962 88286 12964 88338
rect 12908 88228 12964 88286
rect 12908 88162 12964 88172
rect 13244 88116 13300 88126
rect 13020 87556 13076 87566
rect 12572 86660 12628 86670
rect 12572 86658 12852 86660
rect 12572 86606 12574 86658
rect 12626 86606 12852 86658
rect 12572 86604 12852 86606
rect 12572 86594 12628 86604
rect 12796 86100 12852 86604
rect 12572 86044 12852 86100
rect 12572 85090 12628 86044
rect 13020 85708 13076 87500
rect 13244 87330 13300 88060
rect 13356 88004 13412 88844
rect 13468 88228 13524 88238
rect 13468 88134 13524 88172
rect 13356 87948 13524 88004
rect 13244 87278 13246 87330
rect 13298 87278 13300 87330
rect 13244 87220 13300 87278
rect 13244 87154 13300 87164
rect 13468 85874 13524 87948
rect 13468 85822 13470 85874
rect 13522 85822 13524 85874
rect 13468 85810 13524 85822
rect 13580 85988 13636 85998
rect 12572 85038 12574 85090
rect 12626 85038 12628 85090
rect 12572 85026 12628 85038
rect 12908 85652 13076 85708
rect 12796 84980 12852 84990
rect 12796 84886 12852 84924
rect 12908 84978 12964 85652
rect 12908 84926 12910 84978
rect 12962 84926 12964 84978
rect 12908 83410 12964 84926
rect 12908 83358 12910 83410
rect 12962 83358 12964 83410
rect 12572 83300 12628 83310
rect 12572 83206 12628 83244
rect 12796 83300 12852 83310
rect 12796 83206 12852 83244
rect 12908 82964 12964 83358
rect 12908 82898 12964 82908
rect 13468 83300 13524 83310
rect 13580 83300 13636 85932
rect 13692 85876 13748 89516
rect 13804 88900 13860 89740
rect 14588 89794 14644 89852
rect 15036 89908 15092 89918
rect 15036 89814 15092 89852
rect 14588 89742 14590 89794
rect 14642 89742 14644 89794
rect 14028 89684 14084 89694
rect 14028 89590 14084 89628
rect 13804 88834 13860 88844
rect 14028 88452 14084 88462
rect 13804 87556 13860 87566
rect 13804 87462 13860 87500
rect 14028 87442 14084 88396
rect 14028 87390 14030 87442
rect 14082 87390 14084 87442
rect 13916 87332 13972 87342
rect 13916 87238 13972 87276
rect 14028 86660 14084 87390
rect 14476 87442 14532 87454
rect 14476 87390 14478 87442
rect 14530 87390 14532 87442
rect 14252 87332 14308 87342
rect 14308 87276 14420 87332
rect 14252 87266 14308 87276
rect 13692 85810 13748 85820
rect 13916 86604 14084 86660
rect 13916 85708 13972 86604
rect 13524 83244 13636 83300
rect 13692 85652 13972 85708
rect 13468 82626 13524 83244
rect 13468 82574 13470 82626
rect 13522 82574 13524 82626
rect 13468 82562 13524 82574
rect 13692 82348 13748 85652
rect 14364 85204 14420 87276
rect 14476 86660 14532 87390
rect 14588 87444 14644 89742
rect 15260 89794 15316 90412
rect 15372 90402 15428 90412
rect 15484 89906 15540 90748
rect 15484 89854 15486 89906
rect 15538 89854 15540 89906
rect 15484 89842 15540 89854
rect 15596 90578 15652 92092
rect 15932 92036 15988 92764
rect 16156 92484 16212 92988
rect 16380 93716 16436 93726
rect 16380 92820 16436 93660
rect 16380 92754 16436 92764
rect 16492 93492 16548 93502
rect 16492 92930 16548 93436
rect 16492 92878 16494 92930
rect 16546 92878 16548 92930
rect 16156 92418 16212 92428
rect 15932 91970 15988 91980
rect 16268 91588 16324 91598
rect 16044 91364 16100 91374
rect 15708 91362 16100 91364
rect 15708 91310 16046 91362
rect 16098 91310 16100 91362
rect 15708 91308 16100 91310
rect 15708 91252 15764 91308
rect 16044 91298 16100 91308
rect 15708 90804 15764 91196
rect 16268 91028 16324 91532
rect 16380 91252 16436 91262
rect 16492 91252 16548 92878
rect 16604 92820 16660 92830
rect 16940 92820 16996 92830
rect 16604 92818 16940 92820
rect 16604 92766 16606 92818
rect 16658 92766 16940 92818
rect 16604 92764 16940 92766
rect 16604 92754 16660 92764
rect 16940 92726 16996 92764
rect 16828 92596 16884 92606
rect 16828 92370 16884 92540
rect 16828 92318 16830 92370
rect 16882 92318 16884 92370
rect 16828 92306 16884 92318
rect 16380 91250 16548 91252
rect 16380 91198 16382 91250
rect 16434 91198 16548 91250
rect 16380 91196 16548 91198
rect 16828 91364 16884 91374
rect 16828 91250 16884 91308
rect 16828 91198 16830 91250
rect 16882 91198 16884 91250
rect 16380 91186 16436 91196
rect 16268 90972 16436 91028
rect 15708 90802 15876 90804
rect 15708 90750 15710 90802
rect 15762 90750 15876 90802
rect 15708 90748 15876 90750
rect 15708 90738 15764 90748
rect 15596 90526 15598 90578
rect 15650 90526 15652 90578
rect 15260 89742 15262 89794
rect 15314 89742 15316 89794
rect 14812 89682 14868 89694
rect 14812 89630 14814 89682
rect 14866 89630 14868 89682
rect 14812 89572 14868 89630
rect 14812 89506 14868 89516
rect 15260 89684 15316 89742
rect 15596 89684 15652 90526
rect 14820 89404 15084 89414
rect 14876 89348 14924 89404
rect 14980 89348 15028 89404
rect 14820 89338 15084 89348
rect 14700 89012 14756 89022
rect 14700 87668 14756 88956
rect 15148 88788 15204 88798
rect 14820 87836 15084 87846
rect 14876 87780 14924 87836
rect 14980 87780 15028 87836
rect 14820 87770 15084 87780
rect 14700 87602 14756 87612
rect 15148 87666 15204 88732
rect 15148 87614 15150 87666
rect 15202 87614 15204 87666
rect 15148 87602 15204 87614
rect 15036 87556 15092 87566
rect 14700 87444 14756 87454
rect 14588 87442 14756 87444
rect 14588 87390 14702 87442
rect 14754 87390 14756 87442
rect 14588 87388 14756 87390
rect 14700 87378 14756 87388
rect 14924 87442 14980 87454
rect 14924 87390 14926 87442
rect 14978 87390 14980 87442
rect 14924 87220 14980 87390
rect 15036 87444 15092 87500
rect 15260 87554 15316 89628
rect 15484 89628 15652 89684
rect 15708 90020 15764 90030
rect 15708 89794 15764 89964
rect 15708 89742 15710 89794
rect 15762 89742 15764 89794
rect 15260 87502 15262 87554
rect 15314 87502 15316 87554
rect 15260 87490 15316 87502
rect 15372 88900 15428 88910
rect 15036 87388 15204 87444
rect 15036 87220 15092 87230
rect 14924 87164 15036 87220
rect 15036 87154 15092 87164
rect 15036 86772 15092 86782
rect 14476 86604 14644 86660
rect 14476 85204 14532 85214
rect 14364 85202 14532 85204
rect 14364 85150 14478 85202
rect 14530 85150 14532 85202
rect 14364 85148 14532 85150
rect 14476 85138 14532 85148
rect 13804 85090 13860 85102
rect 13804 85038 13806 85090
rect 13858 85038 13860 85090
rect 13804 84308 13860 85038
rect 14028 84980 14084 84990
rect 14028 84530 14084 84924
rect 14028 84478 14030 84530
rect 14082 84478 14084 84530
rect 14028 84466 14084 84478
rect 13804 83300 13860 84252
rect 14364 84420 14420 84430
rect 14364 84308 14420 84364
rect 14476 84308 14532 84318
rect 14364 84306 14532 84308
rect 14364 84254 14478 84306
rect 14530 84254 14532 84306
rect 14364 84252 14532 84254
rect 13916 83300 13972 83310
rect 13804 83298 13972 83300
rect 13804 83246 13918 83298
rect 13970 83246 13972 83298
rect 13804 83244 13972 83246
rect 13692 82292 13860 82348
rect 12460 81678 12462 81730
rect 12514 81678 12516 81730
rect 12236 81170 12292 81182
rect 12236 81118 12238 81170
rect 12290 81118 12292 81170
rect 12236 80498 12292 81118
rect 12236 80446 12238 80498
rect 12290 80446 12292 80498
rect 12236 80434 12292 80446
rect 12460 79044 12516 81678
rect 13020 81732 13076 81742
rect 13580 81732 13636 81742
rect 13020 81730 13300 81732
rect 13020 81678 13022 81730
rect 13074 81678 13300 81730
rect 13020 81676 13300 81678
rect 13020 81666 13076 81676
rect 13020 80162 13076 80174
rect 13020 80110 13022 80162
rect 13074 80110 13076 80162
rect 12684 79714 12740 79726
rect 12684 79662 12686 79714
rect 12738 79662 12740 79714
rect 12684 79604 12740 79662
rect 12684 79538 12740 79548
rect 12460 78978 12516 78988
rect 12124 78766 12126 78818
rect 12178 78766 12180 78818
rect 12124 78754 12180 78766
rect 12236 78932 12292 78942
rect 12236 78818 12292 78876
rect 12236 78766 12238 78818
rect 12290 78766 12292 78818
rect 12124 76466 12180 76478
rect 12124 76414 12126 76466
rect 12178 76414 12180 76466
rect 12124 76356 12180 76414
rect 12124 75684 12180 76300
rect 12124 75618 12180 75628
rect 12124 74452 12180 74462
rect 12124 74226 12180 74396
rect 12124 74174 12126 74226
rect 12178 74174 12180 74226
rect 12124 74162 12180 74174
rect 12236 72884 12292 78766
rect 13020 78820 13076 80110
rect 13132 79490 13188 79502
rect 13132 79438 13134 79490
rect 13186 79438 13188 79490
rect 13132 79380 13188 79438
rect 13132 79314 13188 79324
rect 13020 78754 13076 78764
rect 13244 78932 13300 81676
rect 13020 78596 13076 78606
rect 13020 78502 13076 78540
rect 13020 78034 13076 78046
rect 13020 77982 13022 78034
rect 13074 77982 13076 78034
rect 12908 77364 12964 77374
rect 12572 77362 12964 77364
rect 12572 77310 12910 77362
rect 12962 77310 12964 77362
rect 12572 77308 12964 77310
rect 12348 76466 12404 76478
rect 12348 76414 12350 76466
rect 12402 76414 12404 76466
rect 12348 75796 12404 76414
rect 12460 75796 12516 75806
rect 12348 75794 12516 75796
rect 12348 75742 12462 75794
rect 12514 75742 12516 75794
rect 12348 75740 12516 75742
rect 12460 75730 12516 75740
rect 12572 75682 12628 77308
rect 12908 77298 12964 77308
rect 13020 77140 13076 77982
rect 12572 75630 12574 75682
rect 12626 75630 12628 75682
rect 12348 75458 12404 75470
rect 12348 75406 12350 75458
rect 12402 75406 12404 75458
rect 12348 75124 12404 75406
rect 12348 75030 12404 75068
rect 12572 75012 12628 75630
rect 12796 76916 12852 76926
rect 12796 76244 12852 76860
rect 12796 75684 12852 76188
rect 12908 75684 12964 75694
rect 12796 75682 12964 75684
rect 12796 75630 12910 75682
rect 12962 75630 12964 75682
rect 12796 75628 12964 75630
rect 12908 75618 12964 75628
rect 12572 74946 12628 74956
rect 12460 74900 12516 74910
rect 12348 74452 12404 74462
rect 12348 73948 12404 74396
rect 12460 74226 12516 74844
rect 12796 74786 12852 74798
rect 12796 74734 12798 74786
rect 12850 74734 12852 74786
rect 12572 74674 12628 74686
rect 12572 74622 12574 74674
rect 12626 74622 12628 74674
rect 12572 74338 12628 74622
rect 12796 74564 12852 74734
rect 13020 74564 13076 77084
rect 13132 76916 13188 76926
rect 13132 76690 13188 76860
rect 13132 76638 13134 76690
rect 13186 76638 13188 76690
rect 13132 76626 13188 76638
rect 13244 76580 13300 78876
rect 13468 81730 13636 81732
rect 13468 81678 13582 81730
rect 13634 81678 13636 81730
rect 13468 81676 13636 81678
rect 13468 78484 13524 81676
rect 13580 81666 13636 81676
rect 13692 81732 13748 81742
rect 13468 78418 13524 78428
rect 13580 80388 13636 80398
rect 13692 80388 13748 81676
rect 13580 80386 13748 80388
rect 13580 80334 13582 80386
rect 13634 80334 13748 80386
rect 13580 80332 13748 80334
rect 13580 78260 13636 80332
rect 13580 77924 13636 78204
rect 13244 76514 13300 76524
rect 13468 77922 13636 77924
rect 13468 77870 13582 77922
rect 13634 77870 13636 77922
rect 13468 77868 13636 77870
rect 13468 77252 13524 77868
rect 13580 77858 13636 77868
rect 13692 78820 13748 78830
rect 13692 77924 13748 78764
rect 13804 78484 13860 82292
rect 13916 81732 13972 83244
rect 13916 81666 13972 81676
rect 14028 81730 14084 81742
rect 14028 81678 14030 81730
rect 14082 81678 14084 81730
rect 14028 81620 14084 81678
rect 14084 81564 14196 81620
rect 14028 81554 14084 81564
rect 14028 81058 14084 81070
rect 14028 81006 14030 81058
rect 14082 81006 14084 81058
rect 13916 78932 13972 78942
rect 13916 78818 13972 78876
rect 13916 78766 13918 78818
rect 13970 78766 13972 78818
rect 13916 78754 13972 78766
rect 13804 78428 13972 78484
rect 13692 77858 13748 77868
rect 13468 75796 13524 77196
rect 13580 77138 13636 77150
rect 13580 77086 13582 77138
rect 13634 77086 13636 77138
rect 13580 77028 13636 77086
rect 13580 76962 13636 76972
rect 13692 77026 13748 77038
rect 13692 76974 13694 77026
rect 13746 76974 13748 77026
rect 13468 75684 13524 75740
rect 13580 75684 13636 75694
rect 13468 75682 13636 75684
rect 13468 75630 13582 75682
rect 13634 75630 13636 75682
rect 13468 75628 13636 75630
rect 13580 75460 13636 75628
rect 13580 75394 13636 75404
rect 13580 75012 13636 75022
rect 13580 74918 13636 74956
rect 13244 74900 13300 74910
rect 13692 74900 13748 76974
rect 13916 77028 13972 78428
rect 13916 76962 13972 76972
rect 14028 76468 14084 81006
rect 14140 81060 14196 81564
rect 14140 80994 14196 81004
rect 14252 80948 14308 80958
rect 14252 79042 14308 80892
rect 14364 80612 14420 84252
rect 14476 84242 14532 84252
rect 14476 83524 14532 83534
rect 14476 83430 14532 83468
rect 14588 83522 14644 86604
rect 15036 86658 15092 86716
rect 15036 86606 15038 86658
rect 15090 86606 15092 86658
rect 15036 86594 15092 86606
rect 15036 86436 15092 86474
rect 14588 83470 14590 83522
rect 14642 83470 14644 83522
rect 14588 83458 14644 83470
rect 14700 86380 15036 86436
rect 14476 81732 14532 81742
rect 14476 81638 14532 81676
rect 14364 80546 14420 80556
rect 14252 78990 14254 79042
rect 14306 78990 14308 79042
rect 14252 78978 14308 78990
rect 14364 80274 14420 80286
rect 14364 80222 14366 80274
rect 14418 80222 14420 80274
rect 14252 78818 14308 78830
rect 14252 78766 14254 78818
rect 14306 78766 14308 78818
rect 14252 78484 14308 78766
rect 14364 78596 14420 80222
rect 14700 79156 14756 86380
rect 15036 86370 15092 86380
rect 14820 86268 15084 86278
rect 14876 86212 14924 86268
rect 14980 86212 15028 86268
rect 14820 86202 15084 86212
rect 15148 86100 15204 87388
rect 15372 86884 15428 88844
rect 15484 88116 15540 89628
rect 15708 89124 15764 89742
rect 15820 89684 15876 90748
rect 16268 90468 16324 90478
rect 16156 90466 16324 90468
rect 16156 90414 16270 90466
rect 16322 90414 16324 90466
rect 16156 90412 16324 90414
rect 15820 89682 15988 89684
rect 15820 89630 15822 89682
rect 15874 89630 15988 89682
rect 15820 89628 15988 89630
rect 15820 89618 15876 89628
rect 15708 89030 15764 89068
rect 15820 89236 15876 89246
rect 15820 89122 15876 89180
rect 15820 89070 15822 89122
rect 15874 89070 15876 89122
rect 15820 88340 15876 89070
rect 15932 89066 15988 89628
rect 15932 89014 15934 89066
rect 15986 89014 15988 89066
rect 15932 89002 15988 89014
rect 16156 89012 16212 90412
rect 16268 90402 16324 90412
rect 16380 90468 16436 90972
rect 16380 90402 16436 90412
rect 16604 90468 16660 90478
rect 16604 90374 16660 90412
rect 16828 90020 16884 91198
rect 16828 89954 16884 89964
rect 17052 89908 17108 97412
rect 17388 96850 17444 97470
rect 17500 97634 17556 97646
rect 17500 97582 17502 97634
rect 17554 97582 17556 97634
rect 17500 97076 17556 97582
rect 17500 97010 17556 97020
rect 17388 96798 17390 96850
rect 17442 96798 17444 96850
rect 17388 96786 17444 96798
rect 17500 96852 17556 96862
rect 17500 96628 17556 96796
rect 17388 96572 17556 96628
rect 17276 95508 17332 95518
rect 17164 94276 17220 94286
rect 17164 94182 17220 94220
rect 17276 93156 17332 95452
rect 17388 95172 17444 96572
rect 17612 96292 17668 98140
rect 17724 97746 17780 103070
rect 17836 102340 17892 108558
rect 17948 108836 18004 108846
rect 17948 107828 18004 108780
rect 18508 108610 18564 108622
rect 18508 108558 18510 108610
rect 18562 108558 18564 108610
rect 18172 108500 18228 108510
rect 18172 108406 18228 108444
rect 18508 108276 18564 108558
rect 18508 108210 18564 108220
rect 18172 107828 18228 107838
rect 17948 107826 18228 107828
rect 17948 107774 18174 107826
rect 18226 107774 18228 107826
rect 17948 107772 18228 107774
rect 18060 107044 18116 107772
rect 18172 107762 18228 107772
rect 18222 107436 18486 107446
rect 18278 107380 18326 107436
rect 18382 107380 18430 107436
rect 18222 107370 18486 107380
rect 18172 107044 18228 107054
rect 18060 107042 18228 107044
rect 18060 106990 18174 107042
rect 18226 106990 18228 107042
rect 18060 106988 18228 106990
rect 18172 106978 18228 106988
rect 18284 106260 18340 106270
rect 18060 106258 18340 106260
rect 18060 106206 18286 106258
rect 18338 106206 18340 106258
rect 18060 106204 18340 106206
rect 18060 105868 18116 106204
rect 18284 106194 18340 106204
rect 17948 105812 18116 105868
rect 18222 105868 18486 105878
rect 18278 105812 18326 105868
rect 18382 105812 18430 105868
rect 17948 104132 18004 105812
rect 18222 105802 18486 105812
rect 18620 104916 18676 109452
rect 18732 109284 18788 109294
rect 18956 109284 19012 109294
rect 19404 109284 19460 109902
rect 20076 109844 20132 110236
rect 20636 109954 20692 110908
rect 20748 110898 20804 110908
rect 20636 109902 20638 109954
rect 20690 109902 20692 109954
rect 20636 109844 20692 109902
rect 20076 109788 20692 109844
rect 19516 109396 19572 109406
rect 19516 109302 19572 109340
rect 18788 109282 19460 109284
rect 18788 109230 18958 109282
rect 19010 109230 19460 109282
rect 18788 109228 19460 109230
rect 19964 109282 20020 109294
rect 19964 109230 19966 109282
rect 20018 109230 20020 109282
rect 19964 109228 20020 109230
rect 18732 108722 18788 109228
rect 18956 109218 19012 109228
rect 18732 108670 18734 108722
rect 18786 108670 18788 108722
rect 18732 108658 18788 108670
rect 19180 108500 19236 109228
rect 19180 108406 19236 108444
rect 19852 109172 20020 109228
rect 19852 108610 19908 109172
rect 19852 108558 19854 108610
rect 19906 108558 19908 108610
rect 19068 108388 19124 108398
rect 19068 108294 19124 108332
rect 19180 107826 19236 107838
rect 19180 107774 19182 107826
rect 19234 107774 19236 107826
rect 18620 104850 18676 104860
rect 18956 107492 19012 107502
rect 18956 106260 19012 107436
rect 19180 107044 19236 107774
rect 19852 107492 19908 108558
rect 19852 107426 19908 107436
rect 20076 108388 20132 109788
rect 20524 109508 20580 109518
rect 20524 109506 20692 109508
rect 20524 109454 20526 109506
rect 20578 109454 20692 109506
rect 20524 109452 20692 109454
rect 20524 109442 20580 109452
rect 20412 109284 20468 109294
rect 20412 108722 20468 109228
rect 20636 109228 20692 109452
rect 20636 109172 20804 109228
rect 20412 108670 20414 108722
rect 20466 108670 20468 108722
rect 20188 108388 20244 108398
rect 20076 108332 20188 108388
rect 20076 107268 20132 108332
rect 20188 108322 20244 108332
rect 19852 107212 20132 107268
rect 19852 107044 19908 107212
rect 20076 107154 20132 107212
rect 20076 107102 20078 107154
rect 20130 107102 20132 107154
rect 20076 107090 20132 107102
rect 19180 107042 19908 107044
rect 19180 106990 19182 107042
rect 19234 106990 19908 107042
rect 19180 106988 19908 106990
rect 19180 106820 19236 106988
rect 19180 106754 19236 106764
rect 19852 106482 19908 106988
rect 19852 106430 19854 106482
rect 19906 106430 19908 106482
rect 19852 106418 19908 106430
rect 19964 107044 20020 107054
rect 18172 104692 18228 104702
rect 17948 104066 18004 104076
rect 18060 104690 18228 104692
rect 18060 104638 18174 104690
rect 18226 104638 18228 104690
rect 18060 104636 18228 104638
rect 18060 103348 18116 104636
rect 18172 104626 18228 104636
rect 18508 104692 18564 104702
rect 18508 104578 18564 104636
rect 18508 104526 18510 104578
rect 18562 104526 18564 104578
rect 18508 104514 18564 104526
rect 18222 104300 18486 104310
rect 18278 104244 18326 104300
rect 18382 104244 18430 104300
rect 18222 104234 18486 104244
rect 18396 104132 18452 104142
rect 18060 103292 18340 103348
rect 17836 102274 17892 102284
rect 17948 103122 18004 103134
rect 17948 103070 17950 103122
rect 18002 103070 18004 103122
rect 17948 100884 18004 103070
rect 17948 100818 18004 100828
rect 18060 99092 18116 103292
rect 18284 103234 18340 103292
rect 18396 103346 18452 104076
rect 18396 103294 18398 103346
rect 18450 103294 18452 103346
rect 18396 103282 18452 103294
rect 18284 103182 18286 103234
rect 18338 103182 18340 103234
rect 18284 103170 18340 103182
rect 18844 103122 18900 103134
rect 18844 103070 18846 103122
rect 18898 103070 18900 103122
rect 18222 102732 18486 102742
rect 18278 102676 18326 102732
rect 18382 102676 18430 102732
rect 18222 102666 18486 102676
rect 18844 102452 18900 103070
rect 18844 102386 18900 102396
rect 18844 101332 18900 101342
rect 18956 101332 19012 106204
rect 19964 105698 20020 106988
rect 19964 105646 19966 105698
rect 20018 105646 20020 105698
rect 19964 105634 20020 105646
rect 20188 106148 20244 106158
rect 20412 106148 20468 108670
rect 20748 108500 20804 109172
rect 20748 108498 20916 108500
rect 20748 108446 20750 108498
rect 20802 108446 20916 108498
rect 20748 108444 20916 108446
rect 20748 108434 20804 108444
rect 20524 108388 20580 108398
rect 20524 108050 20580 108332
rect 20524 107998 20526 108050
rect 20578 107998 20580 108050
rect 20524 107986 20580 107998
rect 20748 107828 20804 107838
rect 20748 107734 20804 107772
rect 20860 107268 20916 108444
rect 21084 108050 21140 119600
rect 21624 117628 21888 117638
rect 21680 117572 21728 117628
rect 21784 117572 21832 117628
rect 21624 117562 21888 117572
rect 22316 117124 22372 117134
rect 22652 117124 22708 117134
rect 22316 117122 22708 117124
rect 22316 117070 22318 117122
rect 22370 117070 22654 117122
rect 22706 117070 22708 117122
rect 22316 117068 22708 117070
rect 21624 116060 21888 116070
rect 21680 116004 21728 116060
rect 21784 116004 21832 116060
rect 21624 115994 21888 116004
rect 22316 115556 22372 117068
rect 22652 117058 22708 117068
rect 22316 115554 22484 115556
rect 22316 115502 22318 115554
rect 22370 115502 22484 115554
rect 22316 115500 22484 115502
rect 22316 115490 22372 115500
rect 21420 114882 21476 114894
rect 21420 114830 21422 114882
rect 21474 114830 21476 114882
rect 21420 114324 21476 114830
rect 22428 114882 22484 115500
rect 22428 114830 22430 114882
rect 22482 114830 22484 114882
rect 22428 114660 22484 114830
rect 22652 115554 22708 115566
rect 22652 115502 22654 115554
rect 22706 115502 22708 115554
rect 22652 114660 22708 115502
rect 22428 114604 22652 114660
rect 21624 114492 21888 114502
rect 21680 114436 21728 114492
rect 21784 114436 21832 114492
rect 21624 114426 21888 114436
rect 21420 114258 21476 114268
rect 22652 113986 22708 114604
rect 22876 114436 22932 119600
rect 22876 114370 22932 114380
rect 23660 114268 23716 119644
rect 24332 119476 24388 119644
rect 24640 119600 24752 120000
rect 25676 119644 26180 119700
rect 24668 119476 24724 119600
rect 24332 119420 24724 119476
rect 25026 118412 25290 118422
rect 25082 118356 25130 118412
rect 25186 118356 25234 118412
rect 25026 118346 25290 118356
rect 25676 117458 25732 119644
rect 26124 119476 26180 119644
rect 26432 119600 26544 120000
rect 28224 119600 28336 120000
rect 26460 119476 26516 119600
rect 26124 119420 26516 119476
rect 25676 117406 25678 117458
rect 25730 117406 25732 117458
rect 25676 117394 25732 117406
rect 24668 117236 24724 117246
rect 24668 117122 24724 117180
rect 25340 117236 25396 117246
rect 25340 117142 25396 117180
rect 24668 117070 24670 117122
rect 24722 117070 24724 117122
rect 23772 114660 23828 114670
rect 24108 114660 24164 114698
rect 23772 114658 24108 114660
rect 23772 114606 23774 114658
rect 23826 114606 24108 114658
rect 23772 114604 24108 114606
rect 23772 114594 23828 114604
rect 24108 114594 24164 114604
rect 22652 113934 22654 113986
rect 22706 113934 22708 113986
rect 22092 113874 22148 113886
rect 22092 113822 22094 113874
rect 22146 113822 22148 113874
rect 22092 113540 22148 113822
rect 22652 113540 22708 113934
rect 22092 113538 22708 113540
rect 22092 113486 22094 113538
rect 22146 113486 22708 113538
rect 22092 113484 22708 113486
rect 23548 114212 23716 114268
rect 24108 114436 24164 114446
rect 24108 114268 24164 114380
rect 24108 114212 24276 114268
rect 22092 113474 22148 113484
rect 21420 113090 21476 113102
rect 21420 113038 21422 113090
rect 21474 113038 21476 113090
rect 21420 112420 21476 113038
rect 21624 112924 21888 112934
rect 21680 112868 21728 112924
rect 21784 112868 21832 112924
rect 21624 112858 21888 112868
rect 21532 112420 21588 112430
rect 21868 112420 21924 112430
rect 22316 112420 22372 113484
rect 23436 113314 23492 113326
rect 23436 113262 23438 113314
rect 23490 113262 23492 113314
rect 21420 112418 22372 112420
rect 21420 112366 21534 112418
rect 21586 112366 21870 112418
rect 21922 112366 22372 112418
rect 21420 112364 22372 112366
rect 21532 112354 21588 112364
rect 21868 112354 21924 112364
rect 21624 111356 21888 111366
rect 21680 111300 21728 111356
rect 21784 111300 21832 111356
rect 21624 111290 21888 111300
rect 21420 110964 21476 110974
rect 21420 110178 21476 110908
rect 21420 110126 21422 110178
rect 21474 110126 21476 110178
rect 21420 109618 21476 110126
rect 22316 110852 22372 112364
rect 22540 112530 22596 112542
rect 22540 112478 22542 112530
rect 22594 112478 22596 112530
rect 22540 111748 22596 112478
rect 23436 112530 23492 113262
rect 23436 112478 23438 112530
rect 23490 112478 23492 112530
rect 23212 111748 23268 111758
rect 22540 111746 23268 111748
rect 22540 111694 23214 111746
rect 23266 111694 23268 111746
rect 22540 111692 23268 111694
rect 22652 110852 22708 110862
rect 22316 110850 22708 110852
rect 22316 110798 22318 110850
rect 22370 110798 22654 110850
rect 22706 110798 22708 110850
rect 22316 110796 22708 110798
rect 22316 110178 22372 110796
rect 22652 110786 22708 110796
rect 22316 110126 22318 110178
rect 22370 110126 22372 110178
rect 21624 109788 21888 109798
rect 21680 109732 21728 109788
rect 21784 109732 21832 109788
rect 21624 109722 21888 109732
rect 21420 109566 21422 109618
rect 21474 109566 21476 109618
rect 21420 109554 21476 109566
rect 21308 109394 21364 109406
rect 21308 109342 21310 109394
rect 21362 109342 21364 109394
rect 21308 108834 21364 109342
rect 22316 109228 22372 110126
rect 21308 108782 21310 108834
rect 21362 108782 21364 108834
rect 21308 108770 21364 108782
rect 22204 109172 22372 109228
rect 22428 109282 22484 109294
rect 22428 109230 22430 109282
rect 22482 109230 22484 109282
rect 21084 107998 21086 108050
rect 21138 107998 21140 108050
rect 21084 107986 21140 107998
rect 21420 108500 21476 108510
rect 21420 107716 21476 108444
rect 21868 108388 21924 108426
rect 21868 108322 21924 108332
rect 22204 108388 22260 109172
rect 22204 108322 22260 108332
rect 22316 108724 22372 108734
rect 22316 108610 22372 108668
rect 22316 108558 22318 108610
rect 22370 108558 22372 108610
rect 21624 108220 21888 108230
rect 21680 108164 21728 108220
rect 21784 108164 21832 108220
rect 21624 108154 21888 108164
rect 22316 107826 22372 108558
rect 22316 107774 22318 107826
rect 22370 107774 22372 107826
rect 21532 107716 21588 107726
rect 21420 107714 21700 107716
rect 21420 107662 21534 107714
rect 21586 107662 21700 107714
rect 21420 107660 21700 107662
rect 21532 107650 21588 107660
rect 21644 107604 21700 107660
rect 21532 107268 21588 107278
rect 20860 107266 21588 107268
rect 20860 107214 21534 107266
rect 21586 107214 21588 107266
rect 20860 107212 21588 107214
rect 21532 107202 21588 107212
rect 21308 107044 21364 107054
rect 21644 107044 21700 107548
rect 21196 107042 21700 107044
rect 21196 106990 21310 107042
rect 21362 106990 21700 107042
rect 21196 106988 21700 106990
rect 22316 107042 22372 107774
rect 22428 107604 22484 109230
rect 23212 108724 23268 111692
rect 23436 111748 23492 112478
rect 23436 111682 23492 111692
rect 23212 108658 23268 108668
rect 22428 107538 22484 107548
rect 23100 108612 23156 108622
rect 23100 107826 23156 108556
rect 23100 107774 23102 107826
rect 23154 107774 23156 107826
rect 22316 106990 22318 107042
rect 22370 106990 22372 107042
rect 21196 106596 21252 106988
rect 21308 106978 21364 106988
rect 21868 106820 21924 106830
rect 21868 106818 22036 106820
rect 21868 106766 21870 106818
rect 21922 106766 22036 106818
rect 21868 106764 22036 106766
rect 21868 106754 21924 106764
rect 20188 106146 20468 106148
rect 20188 106094 20190 106146
rect 20242 106094 20468 106146
rect 20188 106092 20468 106094
rect 20636 106540 21252 106596
rect 21624 106652 21888 106662
rect 21680 106596 21728 106652
rect 21784 106596 21832 106652
rect 21624 106586 21888 106596
rect 20188 105588 20244 106092
rect 20188 105522 20244 105532
rect 20636 105700 20692 106540
rect 21308 106484 21364 106494
rect 21308 106390 21364 106428
rect 21868 106372 21924 106382
rect 21980 106372 22036 106764
rect 22316 106484 22372 106990
rect 23100 107042 23156 107774
rect 23100 106990 23102 107042
rect 23154 106990 23156 107042
rect 22316 106418 22372 106428
rect 22764 106484 22820 106494
rect 23100 106484 23156 106990
rect 22764 106482 23156 106484
rect 22764 106430 22766 106482
rect 22818 106430 23156 106482
rect 22764 106428 23156 106430
rect 22764 106418 22820 106428
rect 21868 106370 22036 106372
rect 21868 106318 21870 106370
rect 21922 106318 22036 106370
rect 21868 106316 22036 106318
rect 21868 106306 21924 106316
rect 22204 106260 22260 106270
rect 22204 106166 22260 106204
rect 20300 105474 20356 105486
rect 20300 105422 20302 105474
rect 20354 105422 20356 105474
rect 20300 105364 20356 105422
rect 20524 105476 20580 105486
rect 20636 105476 20692 105644
rect 22540 106148 22596 106158
rect 22540 105698 22596 106092
rect 23324 106148 23380 106158
rect 23324 106054 23380 106092
rect 22540 105646 22542 105698
rect 22594 105646 22596 105698
rect 22540 105634 22596 105646
rect 23436 106034 23492 106046
rect 23436 105982 23438 106034
rect 23490 105982 23492 106034
rect 22204 105588 22260 105598
rect 20524 105474 20692 105476
rect 20524 105422 20526 105474
rect 20578 105422 20692 105474
rect 20524 105420 20692 105422
rect 20524 105410 20580 105420
rect 19068 104804 19124 104814
rect 19068 104710 19124 104748
rect 20300 104804 20356 105308
rect 20300 104738 20356 104748
rect 18900 101276 19012 101332
rect 19404 104690 19460 104702
rect 19404 104638 19406 104690
rect 19458 104638 19460 104690
rect 19404 101666 19460 104638
rect 19516 103012 19572 103022
rect 20636 103012 20692 105420
rect 19516 103010 19908 103012
rect 19516 102958 19518 103010
rect 19570 102958 19908 103010
rect 19516 102956 19908 102958
rect 19516 102946 19572 102956
rect 19740 102228 19796 102238
rect 19740 102134 19796 102172
rect 19404 101614 19406 101666
rect 19458 101614 19460 101666
rect 18222 101164 18486 101174
rect 18278 101108 18326 101164
rect 18382 101108 18430 101164
rect 18222 101098 18486 101108
rect 18284 100996 18340 101006
rect 18284 99986 18340 100940
rect 18284 99934 18286 99986
rect 18338 99934 18340 99986
rect 18284 99922 18340 99934
rect 18732 100884 18788 100894
rect 18222 99596 18486 99606
rect 18278 99540 18326 99596
rect 18382 99540 18430 99596
rect 18222 99530 18486 99540
rect 18060 99026 18116 99036
rect 18172 99428 18228 99438
rect 17836 98980 17892 98990
rect 17836 98530 17892 98924
rect 17948 98756 18004 98766
rect 18004 98700 18116 98756
rect 17948 98690 18004 98700
rect 18060 98642 18116 98700
rect 18060 98590 18062 98642
rect 18114 98590 18116 98642
rect 18060 98578 18116 98590
rect 18172 98642 18228 99372
rect 18172 98590 18174 98642
rect 18226 98590 18228 98642
rect 18172 98578 18228 98590
rect 18732 98642 18788 100828
rect 18732 98590 18734 98642
rect 18786 98590 18788 98642
rect 18732 98578 18788 98590
rect 18844 99540 18900 101276
rect 19404 100996 19460 101614
rect 19404 100930 19460 100940
rect 18844 98642 18900 99484
rect 19740 100770 19796 100782
rect 19740 100718 19742 100770
rect 19794 100718 19796 100770
rect 19180 99204 19236 99214
rect 19180 99110 19236 99148
rect 19740 99204 19796 100718
rect 19740 99138 19796 99148
rect 19852 99202 19908 102956
rect 20188 102564 20244 102574
rect 20188 102450 20244 102508
rect 20188 102398 20190 102450
rect 20242 102398 20244 102450
rect 20188 102386 20244 102398
rect 20636 102450 20692 102956
rect 20636 102398 20638 102450
rect 20690 102398 20692 102450
rect 20636 102386 20692 102398
rect 20748 105532 21588 105588
rect 20748 102450 20804 105532
rect 21308 105364 21364 105374
rect 21308 105270 21364 105308
rect 21532 105362 21588 105532
rect 22204 105494 22260 105532
rect 22540 105476 22596 105486
rect 22540 105474 22932 105476
rect 22540 105422 22542 105474
rect 22594 105422 22932 105474
rect 22540 105420 22932 105422
rect 22540 105410 22596 105420
rect 21532 105310 21534 105362
rect 21586 105310 21588 105362
rect 21532 105298 21588 105310
rect 21420 105250 21476 105262
rect 21420 105198 21422 105250
rect 21474 105198 21476 105250
rect 21420 103906 21476 105198
rect 21624 105084 21888 105094
rect 21680 105028 21728 105084
rect 21784 105028 21832 105084
rect 21624 105018 21888 105028
rect 21420 103854 21422 103906
rect 21474 103854 21476 103906
rect 21420 103842 21476 103854
rect 22204 104578 22260 104590
rect 22204 104526 22206 104578
rect 22258 104526 22260 104578
rect 21624 103516 21888 103526
rect 21680 103460 21728 103516
rect 21784 103460 21832 103516
rect 21624 103450 21888 103460
rect 22204 103122 22260 104526
rect 22316 104356 22372 104366
rect 22316 103906 22372 104300
rect 22316 103854 22318 103906
rect 22370 103854 22372 103906
rect 22316 103842 22372 103854
rect 22876 103346 22932 105420
rect 23212 105474 23268 105486
rect 23212 105422 23214 105474
rect 23266 105422 23268 105474
rect 23212 105364 23268 105422
rect 23212 105298 23268 105308
rect 23436 104244 23492 105982
rect 23436 104178 23492 104188
rect 22876 103294 22878 103346
rect 22930 103294 22932 103346
rect 22876 103282 22932 103294
rect 23324 103348 23380 103358
rect 23548 103348 23604 114212
rect 24108 113316 24164 113326
rect 24108 113222 24164 113260
rect 24108 111748 24164 111758
rect 24108 111654 24164 111692
rect 23660 110068 23716 110078
rect 23660 110066 23940 110068
rect 23660 110014 23662 110066
rect 23714 110014 23940 110066
rect 23660 110012 23940 110014
rect 23660 110002 23716 110012
rect 23884 109956 23940 110012
rect 23996 109956 24052 109966
rect 23884 109954 24052 109956
rect 23884 109902 23998 109954
rect 24050 109902 24052 109954
rect 23884 109900 24052 109902
rect 23996 108388 24052 109900
rect 23996 108322 24052 108332
rect 23772 106148 23828 106158
rect 23772 106054 23828 106092
rect 23996 106034 24052 106046
rect 23996 105982 23998 106034
rect 24050 105982 24052 106034
rect 23884 105364 23940 105374
rect 23660 105308 23884 105364
rect 23660 104356 23716 105308
rect 23884 105270 23940 105308
rect 23660 104018 23716 104300
rect 23660 103966 23662 104018
rect 23714 103966 23716 104018
rect 23660 103954 23716 103966
rect 23772 104244 23828 104254
rect 23660 103348 23716 103358
rect 23548 103346 23716 103348
rect 23548 103294 23662 103346
rect 23714 103294 23716 103346
rect 23548 103292 23716 103294
rect 23324 103254 23380 103292
rect 23660 103282 23716 103292
rect 22204 103070 22206 103122
rect 22258 103070 22260 103122
rect 22204 103058 22260 103070
rect 22428 103236 22484 103246
rect 21644 103010 21700 103022
rect 21980 103012 22036 103022
rect 21644 102958 21646 103010
rect 21698 102958 21700 103010
rect 21644 102564 21700 102958
rect 20748 102398 20750 102450
rect 20802 102398 20804 102450
rect 20748 102386 20804 102398
rect 21084 102508 21700 102564
rect 21756 103010 22036 103012
rect 21756 102958 21982 103010
rect 22034 102958 22036 103010
rect 21756 102956 22036 102958
rect 21756 102564 21812 102956
rect 21980 102946 22036 102956
rect 22428 102564 22484 103180
rect 22540 103124 22596 103134
rect 22540 103010 22596 103068
rect 22540 102958 22542 103010
rect 22594 102958 22596 103010
rect 22540 102946 22596 102958
rect 22988 103012 23044 103022
rect 22988 102918 23044 102956
rect 23660 103012 23716 103022
rect 22540 102564 22596 102574
rect 22428 102562 22596 102564
rect 22428 102510 22542 102562
rect 22594 102510 22596 102562
rect 22428 102508 22596 102510
rect 20412 102338 20468 102350
rect 20412 102286 20414 102338
rect 20466 102286 20468 102338
rect 19964 102226 20020 102238
rect 19964 102174 19966 102226
rect 20018 102174 20020 102226
rect 19964 99428 20020 102174
rect 20076 100772 20132 100782
rect 20076 100678 20132 100716
rect 19964 99362 20020 99372
rect 20300 100658 20356 100670
rect 20300 100606 20302 100658
rect 20354 100606 20356 100658
rect 19852 99150 19854 99202
rect 19906 99150 19908 99202
rect 19852 99138 19908 99150
rect 20188 99204 20244 99214
rect 20300 99204 20356 100606
rect 20188 99202 20356 99204
rect 20188 99150 20190 99202
rect 20242 99150 20356 99202
rect 20188 99148 20356 99150
rect 20188 99138 20244 99148
rect 19292 99092 19348 99102
rect 19068 98980 19124 98990
rect 18844 98590 18846 98642
rect 18898 98590 18900 98642
rect 18844 98578 18900 98590
rect 18956 98978 19124 98980
rect 18956 98926 19070 98978
rect 19122 98926 19124 98978
rect 18956 98924 19124 98926
rect 17836 98478 17838 98530
rect 17890 98478 17892 98530
rect 17836 98466 17892 98478
rect 17948 98532 18004 98570
rect 17948 98466 18004 98476
rect 18284 98420 18340 98430
rect 18284 98326 18340 98364
rect 18620 98418 18676 98430
rect 18956 98420 19012 98924
rect 19068 98914 19124 98924
rect 19292 98978 19348 99036
rect 19292 98926 19294 98978
rect 19346 98926 19348 98978
rect 18620 98366 18622 98418
rect 18674 98366 18676 98418
rect 18620 98196 18676 98366
rect 18620 98130 18676 98140
rect 18732 98364 19012 98420
rect 19180 98644 19236 98654
rect 19180 98418 19236 98588
rect 19180 98366 19182 98418
rect 19234 98366 19236 98418
rect 18222 98028 18486 98038
rect 18278 97972 18326 98028
rect 18382 97972 18430 98028
rect 18222 97962 18486 97972
rect 17724 97694 17726 97746
rect 17778 97694 17780 97746
rect 17724 97682 17780 97694
rect 18508 97636 18564 97646
rect 18172 97524 18228 97534
rect 17724 97412 17780 97422
rect 17724 97410 17892 97412
rect 17724 97358 17726 97410
rect 17778 97358 17892 97410
rect 17724 97356 17892 97358
rect 17724 97346 17780 97356
rect 17836 96964 17892 97356
rect 17948 97410 18004 97422
rect 17948 97358 17950 97410
rect 18002 97358 18004 97410
rect 17948 97188 18004 97358
rect 17948 97122 18004 97132
rect 18172 97074 18228 97468
rect 18172 97022 18174 97074
rect 18226 97022 18228 97074
rect 18172 97010 18228 97022
rect 18396 97410 18452 97422
rect 18396 97358 18398 97410
rect 18450 97358 18452 97410
rect 18396 97076 18452 97358
rect 18396 97010 18452 97020
rect 18508 97074 18564 97580
rect 18508 97022 18510 97074
rect 18562 97022 18564 97074
rect 18508 97010 18564 97022
rect 18732 97300 18788 98364
rect 19180 98308 19236 98366
rect 17948 96964 18004 96974
rect 17836 96962 18004 96964
rect 17836 96910 17950 96962
rect 18002 96910 18004 96962
rect 17836 96908 18004 96910
rect 17724 96850 17780 96862
rect 17724 96798 17726 96850
rect 17778 96798 17780 96850
rect 17724 96404 17780 96798
rect 17948 96852 18004 96908
rect 17948 96786 18004 96796
rect 18732 96852 18788 97244
rect 18844 98252 19236 98308
rect 18844 97076 18900 98252
rect 19292 97860 19348 98926
rect 19516 98980 19572 98990
rect 19516 98886 19572 98924
rect 20076 98980 20132 98990
rect 20076 98886 20132 98924
rect 20188 98420 20244 98430
rect 20188 98326 20244 98364
rect 19740 98308 19796 98318
rect 19740 98306 19908 98308
rect 19740 98254 19742 98306
rect 19794 98254 19908 98306
rect 19740 98252 19908 98254
rect 19740 98242 19796 98252
rect 19180 97804 19348 97860
rect 18956 97524 19012 97562
rect 18956 97458 19012 97468
rect 18844 97010 18900 97020
rect 18844 96852 18900 96862
rect 18732 96850 18900 96852
rect 18732 96798 18846 96850
rect 18898 96798 18900 96850
rect 18732 96796 18900 96798
rect 17836 96740 17892 96750
rect 17836 96646 17892 96684
rect 18222 96460 18486 96470
rect 18278 96404 18326 96460
rect 18382 96404 18430 96460
rect 17724 96348 18116 96404
rect 18222 96394 18486 96404
rect 18060 96292 18116 96348
rect 18284 96292 18340 96302
rect 17612 96236 18004 96292
rect 18060 96290 18340 96292
rect 18060 96238 18286 96290
rect 18338 96238 18340 96290
rect 18060 96236 18340 96238
rect 17500 96066 17556 96078
rect 17500 96014 17502 96066
rect 17554 96014 17556 96066
rect 17500 95508 17556 96014
rect 17724 96068 17780 96078
rect 17612 95954 17668 95966
rect 17612 95902 17614 95954
rect 17666 95902 17668 95954
rect 17612 95620 17668 95902
rect 17724 95842 17780 96012
rect 17724 95790 17726 95842
rect 17778 95790 17780 95842
rect 17724 95778 17780 95790
rect 17612 95564 17892 95620
rect 17500 95452 17780 95508
rect 17612 95284 17668 95294
rect 17612 95190 17668 95228
rect 17388 94724 17444 95116
rect 17500 95170 17556 95182
rect 17500 95118 17502 95170
rect 17554 95118 17556 95170
rect 17500 94948 17556 95118
rect 17500 94882 17556 94892
rect 17388 94668 17556 94724
rect 17164 93100 17332 93156
rect 17388 94386 17444 94398
rect 17388 94334 17390 94386
rect 17442 94334 17444 94386
rect 17164 92708 17220 93100
rect 17164 92642 17220 92652
rect 17276 92932 17332 92942
rect 17052 89842 17108 89852
rect 17164 92484 17220 92494
rect 16604 89794 16660 89806
rect 16604 89742 16606 89794
rect 16658 89742 16660 89794
rect 16156 88946 16212 88956
rect 16268 89682 16324 89694
rect 16268 89630 16270 89682
rect 16322 89630 16324 89682
rect 16268 88452 16324 89630
rect 16380 89572 16436 89582
rect 16380 89010 16436 89516
rect 16380 88958 16382 89010
rect 16434 88958 16436 89010
rect 16380 88946 16436 88958
rect 16604 89348 16660 89742
rect 16716 89348 16772 89358
rect 16604 89292 16716 89348
rect 15484 88050 15540 88060
rect 15708 88284 15876 88340
rect 15932 88396 16324 88452
rect 15372 86818 15428 86828
rect 15484 87668 15540 87678
rect 15484 86660 15540 87612
rect 15372 86604 15540 86660
rect 15708 86660 15764 88284
rect 15820 87554 15876 87566
rect 15820 87502 15822 87554
rect 15874 87502 15876 87554
rect 15820 86996 15876 87502
rect 15932 87330 15988 88396
rect 15932 87278 15934 87330
rect 15986 87278 15988 87330
rect 15932 87266 15988 87278
rect 16044 88228 16100 88238
rect 16044 87444 16100 88172
rect 16604 88228 16660 89292
rect 16716 89282 16772 89292
rect 16828 89012 16884 89022
rect 16828 88340 16884 88956
rect 17164 88452 17220 92428
rect 17276 91474 17332 92876
rect 17276 91422 17278 91474
rect 17330 91422 17332 91474
rect 17276 91410 17332 91422
rect 17388 90020 17444 94334
rect 17500 94052 17556 94668
rect 17612 94388 17668 94398
rect 17724 94388 17780 95452
rect 17612 94386 17780 94388
rect 17612 94334 17614 94386
rect 17666 94334 17780 94386
rect 17612 94332 17780 94334
rect 17612 94322 17668 94332
rect 17500 93042 17556 93996
rect 17612 93716 17668 93726
rect 17612 93622 17668 93660
rect 17500 92990 17502 93042
rect 17554 92990 17556 93042
rect 17500 92978 17556 92990
rect 17612 93268 17668 93278
rect 17612 92930 17668 93212
rect 17612 92878 17614 92930
rect 17666 92878 17668 92930
rect 17500 92148 17556 92158
rect 17612 92148 17668 92878
rect 17724 92370 17780 94332
rect 17724 92318 17726 92370
rect 17778 92318 17780 92370
rect 17724 92306 17780 92318
rect 17836 92372 17892 95564
rect 17948 95396 18004 96236
rect 18284 96226 18340 96236
rect 18620 96292 18676 96302
rect 18732 96292 18788 96796
rect 18844 96786 18900 96796
rect 18620 96290 18788 96292
rect 18620 96238 18622 96290
rect 18674 96238 18788 96290
rect 18620 96236 18788 96238
rect 18620 96226 18676 96236
rect 18060 96068 18116 96078
rect 18060 96066 18452 96068
rect 18060 96014 18062 96066
rect 18114 96014 18452 96066
rect 18060 96012 18452 96014
rect 18060 96002 18116 96012
rect 18396 95620 18452 96012
rect 18396 95564 18676 95620
rect 18620 95506 18676 95564
rect 18620 95454 18622 95506
rect 18674 95454 18676 95506
rect 18620 95442 18676 95454
rect 18172 95396 18228 95406
rect 17948 95394 18228 95396
rect 17948 95342 18174 95394
rect 18226 95342 18228 95394
rect 17948 95340 18228 95342
rect 18172 95330 18228 95340
rect 18396 95282 18452 95294
rect 18396 95230 18398 95282
rect 18450 95230 18452 95282
rect 18396 95060 18452 95230
rect 18452 95004 18676 95060
rect 18396 94994 18452 95004
rect 18222 94892 18486 94902
rect 18278 94836 18326 94892
rect 18382 94836 18430 94892
rect 18222 94826 18486 94836
rect 18396 94724 18452 94734
rect 18284 94668 18396 94724
rect 18172 94500 18228 94510
rect 18060 94388 18116 94398
rect 18060 94294 18116 94332
rect 18172 94386 18228 94444
rect 18172 94334 18174 94386
rect 18226 94334 18228 94386
rect 18172 94322 18228 94334
rect 18284 94386 18340 94668
rect 18396 94658 18452 94668
rect 18284 94334 18286 94386
rect 18338 94334 18340 94386
rect 18284 94322 18340 94334
rect 17948 94274 18004 94286
rect 17948 94222 17950 94274
rect 18002 94222 18004 94274
rect 17948 93044 18004 94222
rect 18620 94164 18676 95004
rect 18620 94098 18676 94108
rect 18732 94498 18788 96236
rect 19068 96740 19124 96750
rect 18844 95956 18900 95966
rect 18844 95862 18900 95900
rect 18844 95508 18900 95518
rect 19068 95508 19124 96684
rect 18844 95394 18900 95452
rect 18844 95342 18846 95394
rect 18898 95342 18900 95394
rect 18844 95330 18900 95342
rect 18956 95452 19124 95508
rect 18956 95172 19012 95452
rect 18732 94446 18734 94498
rect 18786 94446 18788 94498
rect 18508 93714 18564 93726
rect 18508 93662 18510 93714
rect 18562 93662 18564 93714
rect 18060 93604 18116 93614
rect 18060 93268 18116 93548
rect 18508 93492 18564 93662
rect 18508 93426 18564 93436
rect 18222 93324 18486 93334
rect 18278 93268 18326 93324
rect 18382 93268 18430 93324
rect 18222 93258 18486 93268
rect 18060 93202 18116 93212
rect 17948 92988 18116 93044
rect 17836 92306 17892 92316
rect 17948 92820 18004 92830
rect 17556 92092 17668 92148
rect 17836 92146 17892 92158
rect 17836 92094 17838 92146
rect 17890 92094 17892 92146
rect 17500 92054 17556 92092
rect 17836 91588 17892 92094
rect 17948 92146 18004 92764
rect 17948 92094 17950 92146
rect 18002 92094 18004 92146
rect 17948 92082 18004 92094
rect 17836 91522 17892 91532
rect 18060 91474 18116 92988
rect 18620 92820 18676 92830
rect 18732 92820 18788 94446
rect 18676 92764 18788 92820
rect 18844 95116 19012 95172
rect 19068 95282 19124 95294
rect 19068 95230 19070 95282
rect 19122 95230 19124 95282
rect 19068 95172 19124 95230
rect 18620 92754 18676 92764
rect 18508 92372 18564 92382
rect 18564 92316 18676 92372
rect 18508 92278 18564 92316
rect 18222 91756 18486 91766
rect 18278 91700 18326 91756
rect 18382 91700 18430 91756
rect 18222 91690 18486 91700
rect 18620 91588 18676 92316
rect 18844 92036 18900 95116
rect 19068 95106 19124 95116
rect 19180 94724 19236 97804
rect 19404 97748 19460 97758
rect 18956 94668 19236 94724
rect 19292 97634 19348 97646
rect 19292 97582 19294 97634
rect 19346 97582 19348 97634
rect 18956 92932 19012 94668
rect 19068 94500 19124 94510
rect 19068 94406 19124 94444
rect 19180 94388 19236 94398
rect 19068 93826 19124 93838
rect 19068 93774 19070 93826
rect 19122 93774 19124 93826
rect 19068 93604 19124 93774
rect 19068 93538 19124 93548
rect 19180 93602 19236 94332
rect 19180 93550 19182 93602
rect 19234 93550 19236 93602
rect 19180 93538 19236 93550
rect 19292 93156 19348 97582
rect 18956 92866 19012 92876
rect 19068 93100 19348 93156
rect 18844 91970 18900 91980
rect 18956 92034 19012 92046
rect 18956 91982 18958 92034
rect 19010 91982 19012 92034
rect 18956 91812 19012 91982
rect 18956 91746 19012 91756
rect 18060 91422 18062 91474
rect 18114 91422 18116 91474
rect 18060 91410 18116 91422
rect 18172 91532 18676 91588
rect 18732 91532 19012 91588
rect 18060 91252 18116 91262
rect 18172 91252 18228 91532
rect 18508 91364 18564 91374
rect 18732 91364 18788 91532
rect 18956 91474 19012 91532
rect 18956 91422 18958 91474
rect 19010 91422 19012 91474
rect 18956 91410 19012 91422
rect 18508 91362 18788 91364
rect 18508 91310 18510 91362
rect 18562 91310 18788 91362
rect 18508 91308 18788 91310
rect 18844 91362 18900 91374
rect 18844 91310 18846 91362
rect 18898 91310 18900 91362
rect 18508 91298 18564 91308
rect 18060 91250 18228 91252
rect 18060 91198 18062 91250
rect 18114 91198 18228 91250
rect 18060 91196 18228 91198
rect 18844 91252 18900 91310
rect 18956 91252 19012 91262
rect 18844 91196 18956 91252
rect 18060 91186 18116 91196
rect 18956 91186 19012 91196
rect 17948 91138 18004 91150
rect 17948 91086 17950 91138
rect 18002 91086 18004 91138
rect 17948 91028 18004 91086
rect 18284 91138 18340 91150
rect 18284 91086 18286 91138
rect 18338 91086 18340 91138
rect 17948 90972 18228 91028
rect 18172 90580 18228 90972
rect 18172 90514 18228 90524
rect 17388 89954 17444 89964
rect 17612 90466 17668 90478
rect 17612 90414 17614 90466
rect 17666 90414 17668 90466
rect 17612 89684 17668 90414
rect 17948 90468 18004 90478
rect 17948 90354 18004 90412
rect 18284 90356 18340 91086
rect 18844 90580 18900 90590
rect 17948 90302 17950 90354
rect 18002 90302 18004 90354
rect 17724 89796 17780 89806
rect 17724 89702 17780 89740
rect 17612 89618 17668 89628
rect 17948 89684 18004 90302
rect 18060 90300 18340 90356
rect 18396 90466 18452 90478
rect 18396 90414 18398 90466
rect 18450 90414 18452 90466
rect 18396 90354 18452 90414
rect 18396 90302 18398 90354
rect 18450 90302 18452 90354
rect 18060 89796 18116 90300
rect 18396 90290 18452 90302
rect 18222 90188 18486 90198
rect 18278 90132 18326 90188
rect 18382 90132 18430 90188
rect 18222 90122 18486 90132
rect 18508 90020 18564 90030
rect 18844 90020 18900 90524
rect 18060 89740 18228 89796
rect 17948 89618 18004 89628
rect 18060 89572 18116 89582
rect 18060 89478 18116 89516
rect 17500 89348 17556 89358
rect 17500 89010 17556 89292
rect 18172 89236 18228 89740
rect 18396 89684 18452 89694
rect 18060 89180 18228 89236
rect 18284 89236 18340 89246
rect 17500 88958 17502 89010
rect 17554 88958 17556 89010
rect 17500 88946 17556 88958
rect 17948 89124 18004 89134
rect 17948 89010 18004 89068
rect 17948 88958 17950 89010
rect 18002 88958 18004 89010
rect 17948 88946 18004 88958
rect 17724 88898 17780 88910
rect 17724 88846 17726 88898
rect 17778 88846 17780 88898
rect 17164 88396 17332 88452
rect 16828 88338 16996 88340
rect 16828 88286 16830 88338
rect 16882 88286 16996 88338
rect 16828 88284 16996 88286
rect 16828 88274 16884 88284
rect 16604 88162 16660 88172
rect 16716 88116 16772 88126
rect 16604 87668 16660 87678
rect 16604 87574 16660 87612
rect 16044 87388 16548 87444
rect 16044 87330 16100 87388
rect 16044 87278 16046 87330
rect 16098 87278 16100 87330
rect 16044 87266 16100 87278
rect 16380 87220 16436 87230
rect 16268 87218 16436 87220
rect 16268 87166 16382 87218
rect 16434 87166 16436 87218
rect 16268 87164 16436 87166
rect 16268 86996 16324 87164
rect 16380 87154 16436 87164
rect 15820 86940 16324 86996
rect 15708 86658 16212 86660
rect 15708 86606 15710 86658
rect 15762 86606 16212 86658
rect 15708 86604 16212 86606
rect 15260 86100 15316 86110
rect 15148 86098 15316 86100
rect 15148 86046 15262 86098
rect 15314 86046 15316 86098
rect 15148 86044 15316 86046
rect 15036 85876 15092 85886
rect 15036 85652 15092 85820
rect 15036 85596 15204 85652
rect 14820 84700 15084 84710
rect 14876 84644 14924 84700
rect 14980 84644 15028 84700
rect 14820 84634 15084 84644
rect 14812 84420 14868 84430
rect 14812 83410 14868 84364
rect 14924 83524 14980 83534
rect 14924 83430 14980 83468
rect 14812 83358 14814 83410
rect 14866 83358 14868 83410
rect 14812 83346 14868 83358
rect 14820 83132 15084 83142
rect 14876 83076 14924 83132
rect 14980 83076 15028 83132
rect 14820 83066 15084 83076
rect 14812 81954 14868 81966
rect 14812 81902 14814 81954
rect 14866 81902 14868 81954
rect 14812 81732 14868 81902
rect 14812 81666 14868 81676
rect 14820 81564 15084 81574
rect 14876 81508 14924 81564
rect 14980 81508 15028 81564
rect 14820 81498 15084 81508
rect 14820 79996 15084 80006
rect 14876 79940 14924 79996
rect 14980 79940 15028 79996
rect 14820 79930 15084 79940
rect 15148 79828 15204 85596
rect 15260 83748 15316 86044
rect 15260 83682 15316 83692
rect 15372 84418 15428 86604
rect 15708 86594 15764 86604
rect 15372 84366 15374 84418
rect 15426 84366 15428 84418
rect 15372 82964 15428 84366
rect 15484 86324 15540 86334
rect 15484 85316 15540 86268
rect 15932 85988 15988 85998
rect 15932 85894 15988 85932
rect 16156 85986 16212 86604
rect 16156 85934 16158 85986
rect 16210 85934 16212 85986
rect 15484 84420 15540 85260
rect 16156 84980 16212 85934
rect 16156 84914 16212 84924
rect 15484 84354 15540 84364
rect 16268 84308 16324 86940
rect 16492 86884 16548 87388
rect 16716 87330 16772 88060
rect 16716 87278 16718 87330
rect 16770 87278 16772 87330
rect 16716 87266 16772 87278
rect 16492 86770 16548 86828
rect 16492 86718 16494 86770
rect 16546 86718 16548 86770
rect 16492 86706 16548 86718
rect 16380 86546 16436 86558
rect 16380 86494 16382 86546
rect 16434 86494 16436 86546
rect 16380 85986 16436 86494
rect 16380 85934 16382 85986
rect 16434 85934 16436 85986
rect 16380 85316 16436 85934
rect 16828 85764 16884 85774
rect 16716 85652 16772 85662
rect 16716 85558 16772 85596
rect 16380 85250 16436 85260
rect 16604 85202 16660 85214
rect 16604 85150 16606 85202
rect 16658 85150 16660 85202
rect 16604 85092 16660 85150
rect 16604 85026 16660 85036
rect 16324 84252 16548 84308
rect 16268 84242 16324 84252
rect 15932 83748 15988 83758
rect 15596 83636 15652 83646
rect 15596 83542 15652 83580
rect 15372 82898 15428 82908
rect 15708 83524 15764 83534
rect 15708 82852 15764 83468
rect 15932 83300 15988 83692
rect 16380 83300 16436 83310
rect 15932 83298 16436 83300
rect 15932 83246 15934 83298
rect 15986 83246 16382 83298
rect 16434 83246 16436 83298
rect 15932 83244 16436 83246
rect 15932 83234 15988 83244
rect 15932 82964 15988 82974
rect 15708 82796 15876 82852
rect 15596 82740 15652 82750
rect 15596 82646 15652 82684
rect 15820 82738 15876 82796
rect 15820 82686 15822 82738
rect 15874 82686 15876 82738
rect 15708 82626 15764 82638
rect 15708 82574 15710 82626
rect 15762 82574 15764 82626
rect 15596 82068 15652 82078
rect 15708 82068 15764 82574
rect 15820 82404 15876 82686
rect 15820 82338 15876 82348
rect 15596 82066 15764 82068
rect 15596 82014 15598 82066
rect 15650 82014 15764 82066
rect 15596 82012 15764 82014
rect 15596 82002 15652 82012
rect 15148 79772 15316 79828
rect 14812 79716 14868 79726
rect 14812 79622 14868 79660
rect 14924 79604 14980 79614
rect 14924 79510 14980 79548
rect 14700 79090 14756 79100
rect 14812 78820 14868 78830
rect 14700 78818 14868 78820
rect 14700 78766 14814 78818
rect 14866 78766 14868 78818
rect 14700 78764 14868 78766
rect 14476 78596 14532 78606
rect 14364 78594 14532 78596
rect 14364 78542 14478 78594
rect 14530 78542 14532 78594
rect 14364 78540 14532 78542
rect 14476 78530 14532 78540
rect 14252 78148 14308 78428
rect 14700 78260 14756 78764
rect 14812 78754 14868 78764
rect 14820 78428 15084 78438
rect 14876 78372 14924 78428
rect 14980 78372 15028 78428
rect 14820 78362 15084 78372
rect 14700 78194 14756 78204
rect 14364 78148 14420 78158
rect 14252 78092 14364 78148
rect 14364 78082 14420 78092
rect 15036 77252 15092 77262
rect 15036 77158 15092 77196
rect 14820 76860 15084 76870
rect 14876 76804 14924 76860
rect 14980 76804 15028 76860
rect 14820 76794 15084 76804
rect 14028 76374 14084 76412
rect 15260 76578 15316 79772
rect 15820 79716 15876 79726
rect 15932 79716 15988 82908
rect 16044 82740 16100 83244
rect 16380 83234 16436 83244
rect 16492 82964 16548 84252
rect 16828 84194 16884 85708
rect 16828 84142 16830 84194
rect 16882 84142 16884 84194
rect 16828 84084 16884 84142
rect 16716 84028 16884 84084
rect 16604 83636 16660 83646
rect 16716 83636 16772 84028
rect 16660 83580 16772 83636
rect 16604 83570 16660 83580
rect 16828 83300 16884 83310
rect 16604 82964 16660 82974
rect 16492 82962 16660 82964
rect 16492 82910 16606 82962
rect 16658 82910 16660 82962
rect 16492 82908 16660 82910
rect 16604 82898 16660 82908
rect 16380 82850 16436 82862
rect 16380 82798 16382 82850
rect 16434 82798 16436 82850
rect 16044 82674 16100 82684
rect 16268 82740 16324 82750
rect 16380 82740 16436 82798
rect 16268 82738 16436 82740
rect 16268 82686 16270 82738
rect 16322 82686 16436 82738
rect 16268 82684 16436 82686
rect 16716 82740 16772 82750
rect 16268 82674 16324 82684
rect 16716 82646 16772 82684
rect 15820 79714 15988 79716
rect 15820 79662 15822 79714
rect 15874 79662 15988 79714
rect 15820 79660 15988 79662
rect 16380 82068 16436 82078
rect 15596 78706 15652 78718
rect 15596 78654 15598 78706
rect 15650 78654 15652 78706
rect 15596 78260 15652 78654
rect 15596 78194 15652 78204
rect 15260 76526 15262 76578
rect 15314 76526 15316 76578
rect 15260 76020 15316 76526
rect 15260 75954 15316 75964
rect 14252 75570 14308 75582
rect 14252 75518 14254 75570
rect 14306 75518 14308 75570
rect 14252 75122 14308 75518
rect 15596 75348 15652 75358
rect 14820 75292 15084 75302
rect 14876 75236 14924 75292
rect 14980 75236 15028 75292
rect 14820 75226 15084 75236
rect 14252 75070 14254 75122
rect 14306 75070 14308 75122
rect 14252 75058 14308 75070
rect 15148 75124 15204 75134
rect 14028 74900 14084 74910
rect 13692 74844 13860 74900
rect 13244 74806 13300 74844
rect 13356 74674 13412 74686
rect 13356 74622 13358 74674
rect 13410 74622 13412 74674
rect 13020 74508 13300 74564
rect 12796 74498 12852 74508
rect 12572 74286 12574 74338
rect 12626 74286 12628 74338
rect 12572 74274 12628 74286
rect 12460 74174 12462 74226
rect 12514 74174 12516 74226
rect 12460 74162 12516 74174
rect 12572 74116 12628 74126
rect 12348 73892 12516 73948
rect 12236 72818 12292 72828
rect 12236 72658 12292 72670
rect 12236 72606 12238 72658
rect 12290 72606 12292 72658
rect 12236 72212 12292 72606
rect 12236 72146 12292 72156
rect 12460 71988 12516 73892
rect 12124 71986 12516 71988
rect 12124 71934 12462 71986
rect 12514 71934 12516 71986
rect 12124 71932 12516 71934
rect 12124 71762 12180 71932
rect 12460 71922 12516 71932
rect 12124 71710 12126 71762
rect 12178 71710 12180 71762
rect 12124 71698 12180 71710
rect 12012 70812 12292 70868
rect 11900 70252 12180 70308
rect 11900 70084 11956 70094
rect 11900 69990 11956 70028
rect 11788 69582 11790 69634
rect 11842 69582 11844 69634
rect 11788 69570 11844 69582
rect 11788 69188 11844 69198
rect 11788 69094 11844 69132
rect 12012 68740 12068 68750
rect 11418 68236 11682 68246
rect 11474 68180 11522 68236
rect 11578 68180 11626 68236
rect 11418 68170 11682 68180
rect 10892 67844 10948 67854
rect 11564 67844 11620 67854
rect 10892 67842 11620 67844
rect 10892 67790 10894 67842
rect 10946 67790 11566 67842
rect 11618 67790 11620 67842
rect 10892 67788 11620 67790
rect 10892 67778 10948 67788
rect 11564 67778 11620 67788
rect 11676 67844 11732 67854
rect 11676 67750 11732 67788
rect 12012 67842 12068 68684
rect 12012 67790 12014 67842
rect 12066 67790 12068 67842
rect 11452 67620 11508 67630
rect 11340 67564 11452 67620
rect 11340 67284 11396 67564
rect 11452 67526 11508 67564
rect 10780 66994 10836 67004
rect 10892 67282 11396 67284
rect 10892 67230 11342 67282
rect 11394 67230 11396 67282
rect 10892 67228 11396 67230
rect 10780 66834 10836 66846
rect 10780 66782 10782 66834
rect 10834 66782 10836 66834
rect 10332 65378 10388 65390
rect 10332 65326 10334 65378
rect 10386 65326 10388 65378
rect 10332 64818 10388 65326
rect 10332 64766 10334 64818
rect 10386 64766 10388 64818
rect 10332 64754 10388 64766
rect 10444 64706 10500 64718
rect 10444 64654 10446 64706
rect 10498 64654 10500 64706
rect 10332 64596 10388 64606
rect 10220 64594 10332 64596
rect 10220 64542 10222 64594
rect 10274 64542 10332 64594
rect 10220 64540 10332 64542
rect 10220 64530 10276 64540
rect 9884 64484 9940 64494
rect 9884 64390 9940 64428
rect 9660 63858 9716 63868
rect 10108 63924 10164 63934
rect 10108 63830 10164 63868
rect 9548 63810 9604 63822
rect 9548 63758 9550 63810
rect 9602 63758 9604 63810
rect 9548 63252 9604 63758
rect 9996 63812 10052 63822
rect 9660 63700 9716 63710
rect 9660 63606 9716 63644
rect 9660 63252 9716 63262
rect 9548 63196 9660 63252
rect 9660 63158 9716 63196
rect 9436 62972 9940 63028
rect 9884 62578 9940 62972
rect 9884 62526 9886 62578
rect 9938 62526 9940 62578
rect 9884 62514 9940 62526
rect 9996 62914 10052 63756
rect 10220 63252 10276 63262
rect 10220 63138 10276 63196
rect 10220 63086 10222 63138
rect 10274 63086 10276 63138
rect 10220 63074 10276 63086
rect 9996 62862 9998 62914
rect 10050 62862 10052 62914
rect 9996 62580 10052 62862
rect 10108 62914 10164 62926
rect 10108 62862 10110 62914
rect 10162 62862 10164 62914
rect 10108 62692 10164 62862
rect 10108 62626 10164 62636
rect 9996 62514 10052 62524
rect 10332 62356 10388 64540
rect 10108 62300 10388 62356
rect 10444 64484 10500 64654
rect 10780 64706 10836 66782
rect 10780 64654 10782 64706
rect 10834 64654 10836 64706
rect 10780 64642 10836 64654
rect 9996 61572 10052 61582
rect 9660 61458 9716 61470
rect 9660 61406 9662 61458
rect 9714 61406 9716 61458
rect 9660 61012 9716 61406
rect 9660 60946 9716 60956
rect 9772 60676 9828 60686
rect 9772 60582 9828 60620
rect 9884 59444 9940 59454
rect 9884 59350 9940 59388
rect 9660 59220 9716 59230
rect 9548 58324 9604 58334
rect 9548 57874 9604 58268
rect 9660 58210 9716 59164
rect 9772 59218 9828 59230
rect 9772 59166 9774 59218
rect 9826 59166 9828 59218
rect 9772 58828 9828 59166
rect 9884 58996 9940 59006
rect 9996 58996 10052 61516
rect 9884 58994 10052 58996
rect 9884 58942 9886 58994
rect 9938 58942 10052 58994
rect 9884 58940 10052 58942
rect 10108 60786 10164 62300
rect 10332 61012 10388 61022
rect 10332 60918 10388 60956
rect 10108 60734 10110 60786
rect 10162 60734 10164 60786
rect 10108 60676 10164 60734
rect 10332 60788 10388 60798
rect 10332 60694 10388 60732
rect 9884 58930 9940 58940
rect 9772 58772 10052 58828
rect 9660 58158 9662 58210
rect 9714 58158 9716 58210
rect 9660 58100 9716 58158
rect 9660 58034 9716 58044
rect 9996 58212 10052 58772
rect 10108 58658 10164 60620
rect 10444 60564 10500 64428
rect 10892 64036 10948 67228
rect 11340 67218 11396 67228
rect 11564 67060 11620 67070
rect 12012 67060 12068 67790
rect 11564 66966 11620 67004
rect 11788 67058 12068 67060
rect 11788 67006 12014 67058
rect 12066 67006 12068 67058
rect 11788 67004 12068 67006
rect 11004 66948 11060 66958
rect 11452 66948 11508 66958
rect 11004 66854 11060 66892
rect 11116 66946 11508 66948
rect 11116 66894 11454 66946
rect 11506 66894 11508 66946
rect 11116 66892 11508 66894
rect 11116 66834 11172 66892
rect 11452 66882 11508 66892
rect 11116 66782 11118 66834
rect 11170 66782 11172 66834
rect 11116 66770 11172 66782
rect 11418 66668 11682 66678
rect 11474 66612 11522 66668
rect 11578 66612 11626 66668
rect 11418 66602 11682 66612
rect 11418 65100 11682 65110
rect 11474 65044 11522 65100
rect 11578 65044 11626 65100
rect 11418 65034 11682 65044
rect 11228 64596 11284 64606
rect 11228 64502 11284 64540
rect 10780 63980 10948 64036
rect 10780 63588 10836 63980
rect 10892 63812 10948 63822
rect 10892 63810 11284 63812
rect 10892 63758 10894 63810
rect 10946 63758 11284 63810
rect 10892 63756 11284 63758
rect 10892 63746 10948 63756
rect 10780 63532 10948 63588
rect 10556 63138 10612 63150
rect 10556 63086 10558 63138
rect 10610 63086 10612 63138
rect 10556 62578 10612 63086
rect 10556 62526 10558 62578
rect 10610 62526 10612 62578
rect 10556 61684 10612 62526
rect 10556 61618 10612 61628
rect 10892 60900 10948 63532
rect 11228 63252 11284 63756
rect 11418 63532 11682 63542
rect 11474 63476 11522 63532
rect 11578 63476 11626 63532
rect 11418 63466 11682 63476
rect 11788 63364 11844 67004
rect 12012 66948 12068 67004
rect 12012 66882 12068 66892
rect 11676 63308 11844 63364
rect 12012 63924 12068 63934
rect 11340 63252 11396 63262
rect 11228 63250 11396 63252
rect 11228 63198 11342 63250
rect 11394 63198 11396 63250
rect 11228 63196 11396 63198
rect 11340 63186 11396 63196
rect 11564 63252 11620 63262
rect 11564 63140 11620 63196
rect 11452 63138 11620 63140
rect 11452 63086 11566 63138
rect 11618 63086 11620 63138
rect 11452 63084 11620 63086
rect 11228 63026 11284 63038
rect 11228 62974 11230 63026
rect 11282 62974 11284 63026
rect 11228 62804 11284 62974
rect 11228 62738 11284 62748
rect 11004 62580 11060 62590
rect 11452 62580 11508 63084
rect 11564 63074 11620 63084
rect 11676 62692 11732 63308
rect 11788 63140 11844 63150
rect 11788 63046 11844 63084
rect 11676 62636 11788 62692
rect 11004 62486 11060 62524
rect 11116 62578 11508 62580
rect 11116 62526 11454 62578
rect 11506 62526 11508 62578
rect 11116 62524 11508 62526
rect 11732 62580 11788 62636
rect 11732 62524 11956 62580
rect 11116 60900 11172 62524
rect 11452 62514 11508 62524
rect 11418 61964 11682 61974
rect 11474 61908 11522 61964
rect 11578 61908 11626 61964
rect 11418 61898 11682 61908
rect 11788 61682 11844 61694
rect 11788 61630 11790 61682
rect 11842 61630 11844 61682
rect 11788 61348 11844 61630
rect 11452 60900 11508 60910
rect 10892 60844 11060 60900
rect 11116 60844 11284 60900
rect 10668 60788 10724 60798
rect 10668 60786 10948 60788
rect 10668 60734 10670 60786
rect 10722 60734 10948 60786
rect 10668 60732 10948 60734
rect 10668 60722 10724 60732
rect 10892 60674 10948 60732
rect 10892 60622 10894 60674
rect 10946 60622 10948 60674
rect 10892 60610 10948 60622
rect 10444 60498 10500 60508
rect 10780 60564 10836 60574
rect 10444 59780 10500 59790
rect 10444 59686 10500 59724
rect 10444 59332 10500 59342
rect 10444 59220 10500 59276
rect 10108 58606 10110 58658
rect 10162 58606 10164 58658
rect 10108 58594 10164 58606
rect 10220 59218 10500 59220
rect 10220 59166 10446 59218
rect 10498 59166 10500 59218
rect 10220 59164 10500 59166
rect 10108 58212 10164 58222
rect 9996 58210 10164 58212
rect 9996 58158 10110 58210
rect 10162 58158 10164 58210
rect 9996 58156 10164 58158
rect 9548 57822 9550 57874
rect 9602 57822 9604 57874
rect 9548 57810 9604 57822
rect 9772 57650 9828 57662
rect 9772 57598 9774 57650
rect 9826 57598 9828 57650
rect 9660 57538 9716 57550
rect 9660 57486 9662 57538
rect 9714 57486 9716 57538
rect 9660 57204 9716 57486
rect 9548 57148 9716 57204
rect 9548 56196 9604 57148
rect 9660 56980 9716 56990
rect 9772 56980 9828 57598
rect 9660 56978 9828 56980
rect 9660 56926 9662 56978
rect 9714 56926 9828 56978
rect 9660 56924 9828 56926
rect 9660 56644 9716 56924
rect 9660 56578 9716 56588
rect 9772 56532 9828 56542
rect 9772 56308 9828 56476
rect 9548 56130 9604 56140
rect 9660 56252 9828 56308
rect 9436 55412 9492 55422
rect 9436 55318 9492 55356
rect 9660 55188 9716 56252
rect 9772 56082 9828 56094
rect 9772 56030 9774 56082
rect 9826 56030 9828 56082
rect 9772 55972 9828 56030
rect 9996 56084 10052 58156
rect 10108 58146 10164 58156
rect 10108 57876 10164 57886
rect 10108 57650 10164 57820
rect 10108 57598 10110 57650
rect 10162 57598 10164 57650
rect 10108 57586 10164 57598
rect 10108 56868 10164 56878
rect 10220 56868 10276 59164
rect 10444 59154 10500 59164
rect 10444 58884 10500 58894
rect 10108 56866 10276 56868
rect 10108 56814 10110 56866
rect 10162 56814 10276 56866
rect 10108 56812 10276 56814
rect 10332 58658 10388 58670
rect 10332 58606 10334 58658
rect 10386 58606 10388 58658
rect 10332 57540 10388 58606
rect 10444 57876 10500 58828
rect 10556 58548 10612 58586
rect 10556 58482 10612 58492
rect 10556 58324 10612 58334
rect 10780 58324 10836 60508
rect 10892 59780 10948 59790
rect 11004 59780 11060 60844
rect 11116 60674 11172 60686
rect 11116 60622 11118 60674
rect 11170 60622 11172 60674
rect 11116 60228 11172 60622
rect 11228 60452 11284 60844
rect 11452 60806 11508 60844
rect 11228 60386 11284 60396
rect 11418 60396 11682 60406
rect 11474 60340 11522 60396
rect 11578 60340 11626 60396
rect 11418 60330 11682 60340
rect 11788 60228 11844 61292
rect 11116 60172 11396 60228
rect 11340 60114 11396 60172
rect 11340 60062 11342 60114
rect 11394 60062 11396 60114
rect 11340 60050 11396 60062
rect 11676 60172 11844 60228
rect 11452 60004 11508 60014
rect 11676 60004 11732 60172
rect 11452 60002 11732 60004
rect 11452 59950 11454 60002
rect 11506 59950 11732 60002
rect 11452 59948 11732 59950
rect 11900 60004 11956 62524
rect 12012 62578 12068 63868
rect 12012 62526 12014 62578
rect 12066 62526 12068 62578
rect 12012 62514 12068 62526
rect 12124 61796 12180 70252
rect 12236 70196 12292 70812
rect 12460 70756 12516 70766
rect 12460 70662 12516 70700
rect 12460 70196 12516 70206
rect 12572 70196 12628 74060
rect 13132 73892 13188 73902
rect 13132 73330 13188 73836
rect 13132 73278 13134 73330
rect 13186 73278 13188 73330
rect 13132 73266 13188 73278
rect 12236 70194 12404 70196
rect 12236 70142 12238 70194
rect 12290 70142 12404 70194
rect 12236 70140 12404 70142
rect 12236 70130 12292 70140
rect 12348 69860 12404 70140
rect 12460 70194 12628 70196
rect 12460 70142 12462 70194
rect 12514 70142 12628 70194
rect 12460 70140 12628 70142
rect 12684 72884 12740 72894
rect 12460 70130 12516 70140
rect 12684 70084 12740 72828
rect 12908 72660 12964 72670
rect 12908 72566 12964 72604
rect 12684 69990 12740 70028
rect 12796 72324 12852 72334
rect 12796 69972 12852 72268
rect 12908 71988 12964 71998
rect 12908 71894 12964 71932
rect 13020 71204 13076 71214
rect 12908 70754 12964 70766
rect 12908 70702 12910 70754
rect 12962 70702 12964 70754
rect 12908 70644 12964 70702
rect 12908 70578 12964 70588
rect 13020 70418 13076 71148
rect 13020 70366 13022 70418
rect 13074 70366 13076 70418
rect 13020 70354 13076 70366
rect 13244 71092 13300 74508
rect 13356 73330 13412 74622
rect 13692 74674 13748 74686
rect 13692 74622 13694 74674
rect 13746 74622 13748 74674
rect 13692 74004 13748 74622
rect 13804 74228 13860 74844
rect 14084 74844 14196 74900
rect 14028 74806 14084 74844
rect 13804 74162 13860 74172
rect 14028 74676 14084 74686
rect 14028 74226 14084 74620
rect 14028 74174 14030 74226
rect 14082 74174 14084 74226
rect 14028 74162 14084 74174
rect 14140 74116 14196 74844
rect 14252 74898 14308 74910
rect 14252 74846 14254 74898
rect 14306 74846 14308 74898
rect 14252 74564 14308 74846
rect 14588 74900 14644 74910
rect 14588 74806 14644 74844
rect 14924 74898 14980 74910
rect 14924 74846 14926 74898
rect 14978 74846 14980 74898
rect 14924 74788 14980 74846
rect 15036 74900 15092 74910
rect 15036 74806 15092 74844
rect 14924 74722 14980 74732
rect 14252 74498 14308 74508
rect 14140 74060 14420 74116
rect 13692 73938 13748 73948
rect 13356 73278 13358 73330
rect 13410 73278 13412 73330
rect 13356 73266 13412 73278
rect 13580 73890 13636 73902
rect 13580 73838 13582 73890
rect 13634 73838 13636 73890
rect 13580 73332 13636 73838
rect 14028 73444 14084 73454
rect 14028 73350 14084 73388
rect 13692 73332 13748 73342
rect 13580 73330 13748 73332
rect 13580 73278 13694 73330
rect 13746 73278 13748 73330
rect 13580 73276 13748 73278
rect 13692 73220 13748 73276
rect 13804 73332 13860 73342
rect 13804 73238 13860 73276
rect 14252 73332 14308 73342
rect 13692 73154 13748 73164
rect 13916 73218 13972 73230
rect 13916 73166 13918 73218
rect 13970 73166 13972 73218
rect 13916 72884 13972 73166
rect 13692 72828 13972 72884
rect 13692 72770 13748 72828
rect 14028 72772 14084 72782
rect 13692 72718 13694 72770
rect 13746 72718 13748 72770
rect 13692 72706 13748 72718
rect 13916 72716 14028 72772
rect 13916 72658 13972 72716
rect 14028 72706 14084 72716
rect 14252 72770 14308 73276
rect 14252 72718 14254 72770
rect 14306 72718 14308 72770
rect 14252 72706 14308 72718
rect 13916 72606 13918 72658
rect 13970 72606 13972 72658
rect 13916 72594 13972 72606
rect 13580 72548 13636 72558
rect 13580 72454 13636 72492
rect 14140 72546 14196 72558
rect 14140 72494 14142 72546
rect 14194 72494 14196 72546
rect 14140 72324 14196 72494
rect 14364 72324 14420 74060
rect 14924 74004 14980 74014
rect 15148 74004 15204 75068
rect 15596 74898 15652 75292
rect 15596 74846 15598 74898
rect 15650 74846 15652 74898
rect 15596 74834 15652 74846
rect 15708 74674 15764 74686
rect 15708 74622 15710 74674
rect 15762 74622 15764 74674
rect 15596 74116 15652 74126
rect 15708 74116 15764 74622
rect 15596 74114 15708 74116
rect 15596 74062 15598 74114
rect 15650 74062 15708 74114
rect 15596 74060 15708 74062
rect 15596 74050 15652 74060
rect 14924 74002 15204 74004
rect 14924 73950 14926 74002
rect 14978 73950 15204 74002
rect 14924 73948 15204 73950
rect 14924 73938 14980 73948
rect 14588 73892 14644 73902
rect 14812 73892 14868 73902
rect 14588 73798 14644 73836
rect 14700 73890 14868 73892
rect 14700 73838 14814 73890
rect 14866 73838 14868 73890
rect 14700 73836 14868 73838
rect 14700 73444 14756 73836
rect 14812 73826 14868 73836
rect 15372 73892 15428 73902
rect 14820 73724 15084 73734
rect 14876 73668 14924 73724
rect 14980 73668 15028 73724
rect 14820 73658 15084 73668
rect 14700 73378 14756 73388
rect 15260 73444 15316 73454
rect 14588 73218 14644 73230
rect 14588 73166 14590 73218
rect 14642 73166 14644 73218
rect 14588 72548 14644 73166
rect 14588 72482 14644 72492
rect 15148 73220 15204 73230
rect 15148 72436 15204 73164
rect 14364 72268 14756 72324
rect 14140 72258 14196 72268
rect 14252 72100 14308 72110
rect 13580 71820 14084 71876
rect 13468 71540 13524 71550
rect 13468 71446 13524 71484
rect 13580 71538 13636 71820
rect 13580 71486 13582 71538
rect 13634 71486 13636 71538
rect 13580 71474 13636 71486
rect 13804 71538 13860 71550
rect 13804 71486 13806 71538
rect 13858 71486 13860 71538
rect 13804 71316 13860 71486
rect 13916 71540 13972 71550
rect 13916 71446 13972 71484
rect 13468 71260 13860 71316
rect 13468 71204 13524 71260
rect 14028 71204 14084 71820
rect 14252 71874 14308 72044
rect 14364 71988 14420 71998
rect 14700 71988 14756 72268
rect 14820 72156 15084 72166
rect 14876 72100 14924 72156
rect 14980 72100 15028 72156
rect 14820 72090 15084 72100
rect 15036 71988 15092 71998
rect 14700 71932 14868 71988
rect 14364 71894 14420 71932
rect 14252 71822 14254 71874
rect 14306 71822 14308 71874
rect 14252 71810 14308 71822
rect 14252 71540 14308 71550
rect 14308 71484 14420 71540
rect 14252 71474 14308 71484
rect 13468 71138 13524 71148
rect 13580 71148 13972 71204
rect 14028 71148 14308 71204
rect 12908 70196 12964 70206
rect 12908 70102 12964 70140
rect 13132 70194 13188 70206
rect 13132 70142 13134 70194
rect 13186 70142 13188 70194
rect 12796 69916 13076 69972
rect 12348 69804 12852 69860
rect 12348 69634 12404 69646
rect 12348 69582 12350 69634
rect 12402 69582 12404 69634
rect 12236 69186 12292 69198
rect 12236 69134 12238 69186
rect 12290 69134 12292 69186
rect 12236 68740 12292 69134
rect 12236 68674 12292 68684
rect 12348 64930 12404 69582
rect 12684 69636 12740 69646
rect 12684 69542 12740 69580
rect 12572 69298 12628 69310
rect 12572 69246 12574 69298
rect 12626 69246 12628 69298
rect 12460 68516 12516 68526
rect 12572 68516 12628 69246
rect 12796 68738 12852 69804
rect 12796 68686 12798 68738
rect 12850 68686 12852 68738
rect 12796 68674 12852 68686
rect 12460 68514 12628 68516
rect 12460 68462 12462 68514
rect 12514 68462 12628 68514
rect 12460 68460 12628 68462
rect 12460 67844 12516 68460
rect 12908 67956 12964 67966
rect 12460 67778 12516 67788
rect 12684 67900 12908 67956
rect 12460 67620 12516 67630
rect 12460 67396 12516 67564
rect 12460 65716 12516 67340
rect 12460 65650 12516 65660
rect 12572 67060 12628 67070
rect 12460 65380 12516 65390
rect 12572 65380 12628 67004
rect 12684 66164 12740 67900
rect 12908 67862 12964 67900
rect 13020 67284 13076 69916
rect 13132 69860 13188 70142
rect 13132 69794 13188 69804
rect 13244 69636 13300 71036
rect 13580 71090 13636 71148
rect 13580 71038 13582 71090
rect 13634 71038 13636 71090
rect 13580 70644 13636 71038
rect 13580 70578 13636 70588
rect 13692 70980 13748 70990
rect 13132 69580 13300 69636
rect 13356 70196 13412 70206
rect 13132 67508 13188 69580
rect 13356 69522 13412 70140
rect 13356 69470 13358 69522
rect 13410 69470 13412 69522
rect 13356 69458 13412 69470
rect 13468 70084 13524 70094
rect 13468 69524 13524 70028
rect 13244 69412 13300 69422
rect 13244 69300 13300 69356
rect 13468 69410 13524 69468
rect 13692 69412 13748 70924
rect 13804 70978 13860 70990
rect 13804 70926 13806 70978
rect 13858 70926 13860 70978
rect 13804 70868 13860 70926
rect 13916 70980 13972 71148
rect 14252 71090 14308 71148
rect 14252 71038 14254 71090
rect 14306 71038 14308 71090
rect 14252 71026 14308 71038
rect 13916 70914 13972 70924
rect 14028 70978 14084 70990
rect 14028 70926 14030 70978
rect 14082 70926 14084 70978
rect 13804 70802 13860 70812
rect 14028 70756 14084 70926
rect 14140 70868 14196 70878
rect 14252 70868 14308 70878
rect 14196 70866 14308 70868
rect 14196 70814 14254 70866
rect 14306 70814 14308 70866
rect 14196 70812 14308 70814
rect 14140 70802 14196 70812
rect 14028 70196 14084 70700
rect 14028 70130 14084 70140
rect 14140 70644 14196 70654
rect 13468 69358 13470 69410
rect 13522 69358 13524 69410
rect 13468 69346 13524 69358
rect 13580 69356 13748 69412
rect 14028 69412 14084 69422
rect 13244 69244 13412 69300
rect 13132 67452 13300 67508
rect 13132 67284 13188 67294
rect 13020 67282 13188 67284
rect 13020 67230 13134 67282
rect 13186 67230 13188 67282
rect 13020 67228 13188 67230
rect 13132 67218 13188 67228
rect 13244 66948 13300 67452
rect 12908 66892 13300 66948
rect 12796 66836 12852 66846
rect 12796 66742 12852 66780
rect 12908 66388 12964 66892
rect 13356 66836 13412 69244
rect 13468 68404 13524 68414
rect 13468 67956 13524 68348
rect 13468 67862 13524 67900
rect 13580 67172 13636 69356
rect 13692 69186 13748 69198
rect 13692 69134 13694 69186
rect 13746 69134 13748 69186
rect 13692 68292 13748 69134
rect 13916 69188 13972 69198
rect 13916 69094 13972 69132
rect 14028 68852 14084 69356
rect 13692 68226 13748 68236
rect 13916 68796 14084 68852
rect 12908 66294 12964 66332
rect 13244 66780 13412 66836
rect 13468 67116 13636 67172
rect 13692 67842 13748 67854
rect 13692 67790 13694 67842
rect 13746 67790 13748 67842
rect 12684 66108 12964 66164
rect 12460 65378 12628 65380
rect 12460 65326 12462 65378
rect 12514 65326 12628 65378
rect 12460 65324 12628 65326
rect 12684 65492 12740 65502
rect 12460 65314 12516 65324
rect 12684 65268 12740 65436
rect 12348 64878 12350 64930
rect 12402 64878 12404 64930
rect 12348 64866 12404 64878
rect 12572 65212 12740 65268
rect 12236 63140 12292 63150
rect 12460 63140 12516 63150
rect 12292 63084 12404 63140
rect 12236 63074 12292 63084
rect 12348 63026 12404 63084
rect 12460 63046 12516 63084
rect 12348 62974 12350 63026
rect 12402 62974 12404 63026
rect 12348 62962 12404 62974
rect 12236 62914 12292 62926
rect 12236 62862 12238 62914
rect 12290 62862 12292 62914
rect 12236 62580 12292 62862
rect 12236 62514 12292 62524
rect 12460 62804 12516 62814
rect 12460 62578 12516 62748
rect 12460 62526 12462 62578
rect 12514 62526 12516 62578
rect 12460 62514 12516 62526
rect 12572 62188 12628 65212
rect 12684 64482 12740 64494
rect 12684 64430 12686 64482
rect 12738 64430 12740 64482
rect 12684 63924 12740 64430
rect 12684 63858 12740 63868
rect 12684 62916 12740 62926
rect 12684 62822 12740 62860
rect 12124 61730 12180 61740
rect 12236 62132 12628 62188
rect 12684 62356 12740 62366
rect 12124 61460 12180 61470
rect 12124 61366 12180 61404
rect 12236 61236 12292 62132
rect 12348 61796 12404 61806
rect 12348 61570 12404 61740
rect 12684 61682 12740 62300
rect 12908 62188 12964 66108
rect 13132 65380 13188 65390
rect 13020 64930 13076 64942
rect 13020 64878 13022 64930
rect 13074 64878 13076 64930
rect 13020 64036 13076 64878
rect 13132 64260 13188 65324
rect 13132 64194 13188 64204
rect 13020 63980 13188 64036
rect 13020 63810 13076 63822
rect 13020 63758 13022 63810
rect 13074 63758 13076 63810
rect 13020 63140 13076 63758
rect 13020 63074 13076 63084
rect 13020 62580 13076 62590
rect 13020 62486 13076 62524
rect 13132 62356 13188 63980
rect 12684 61630 12686 61682
rect 12738 61630 12740 61682
rect 12684 61618 12740 61630
rect 12796 62132 12964 62188
rect 13020 62300 13188 62356
rect 12348 61518 12350 61570
rect 12402 61518 12404 61570
rect 12348 61506 12404 61518
rect 12348 61348 12404 61358
rect 12572 61348 12628 61358
rect 12404 61346 12628 61348
rect 12404 61294 12574 61346
rect 12626 61294 12628 61346
rect 12404 61292 12628 61294
rect 12348 61282 12404 61292
rect 12572 61282 12628 61292
rect 12684 61348 12740 61358
rect 12684 61254 12740 61292
rect 11452 59938 11508 59948
rect 11900 59910 11956 59948
rect 12124 61180 12292 61236
rect 11228 59780 11284 59790
rect 10892 59778 11284 59780
rect 10892 59726 10894 59778
rect 10946 59726 11230 59778
rect 11282 59726 11284 59778
rect 10892 59724 11284 59726
rect 10892 58436 10948 59724
rect 11228 59714 11284 59724
rect 11228 59106 11284 59118
rect 11228 59054 11230 59106
rect 11282 59054 11284 59106
rect 11228 58548 11284 59054
rect 11900 58996 11956 59006
rect 11418 58828 11682 58838
rect 11474 58772 11522 58828
rect 11578 58772 11626 58828
rect 11418 58762 11682 58772
rect 11788 58660 11844 58670
rect 11788 58566 11844 58604
rect 11452 58548 11508 58558
rect 11228 58546 11508 58548
rect 11228 58494 11454 58546
rect 11506 58494 11508 58546
rect 11228 58492 11508 58494
rect 11452 58482 11508 58492
rect 11900 58436 11956 58940
rect 10892 58370 10948 58380
rect 11788 58380 11956 58436
rect 12012 58434 12068 58446
rect 12012 58382 12014 58434
rect 12066 58382 12068 58434
rect 10612 58268 10836 58324
rect 11340 58324 11396 58334
rect 11564 58324 11620 58334
rect 10556 58258 10612 58268
rect 11340 58230 11396 58268
rect 11452 58322 11620 58324
rect 11452 58270 11566 58322
rect 11618 58270 11620 58322
rect 11452 58268 11620 58270
rect 11004 58212 11060 58222
rect 11004 58118 11060 58156
rect 10444 57820 10948 57876
rect 10668 57652 10724 57690
rect 10108 56532 10164 56812
rect 10108 56466 10164 56476
rect 10220 56644 10276 56654
rect 10220 56194 10276 56588
rect 10220 56142 10222 56194
rect 10274 56142 10276 56194
rect 10220 56130 10276 56142
rect 10332 56196 10388 57484
rect 10332 56130 10388 56140
rect 10556 57596 10668 57652
rect 9996 56082 10164 56084
rect 9996 56030 9998 56082
rect 10050 56030 10164 56082
rect 9996 56028 10164 56030
rect 9996 56018 10052 56028
rect 9772 55906 9828 55916
rect 9660 54514 9716 55132
rect 10108 55860 10164 56028
rect 10444 56082 10500 56094
rect 10444 56030 10446 56082
rect 10498 56030 10500 56082
rect 10332 55972 10388 55982
rect 10332 55878 10388 55916
rect 9884 55074 9940 55086
rect 9884 55022 9886 55074
rect 9938 55022 9940 55074
rect 9884 54964 9940 55022
rect 9996 54964 10052 54974
rect 9884 54908 9996 54964
rect 9996 54898 10052 54908
rect 10108 54740 10164 55804
rect 10444 55860 10500 56030
rect 10444 55794 10500 55804
rect 9660 54462 9662 54514
rect 9714 54462 9716 54514
rect 9660 53844 9716 54462
rect 9660 53778 9716 53788
rect 9996 54684 10164 54740
rect 10220 55522 10276 55534
rect 10220 55470 10222 55522
rect 10274 55470 10276 55522
rect 10220 55074 10276 55470
rect 10220 55022 10222 55074
rect 10274 55022 10276 55074
rect 9436 53620 9492 53630
rect 9996 53620 10052 54684
rect 10220 54292 10276 55022
rect 10556 54852 10612 57596
rect 10668 57586 10724 57596
rect 10780 56980 10836 56990
rect 10780 56886 10836 56924
rect 10892 56308 10948 57820
rect 11340 57652 11396 57662
rect 11452 57652 11508 58268
rect 11564 58258 11620 58268
rect 11396 57596 11508 57652
rect 11340 57586 11396 57596
rect 11116 57540 11172 57550
rect 11116 57446 11172 57484
rect 11564 57538 11620 57550
rect 11564 57486 11566 57538
rect 11618 57486 11620 57538
rect 10892 56082 10948 56252
rect 10892 56030 10894 56082
rect 10946 56030 10948 56082
rect 10892 56018 10948 56030
rect 11004 57426 11060 57438
rect 11004 57374 11006 57426
rect 11058 57374 11060 57426
rect 10892 55860 10948 55870
rect 10892 55766 10948 55804
rect 10668 55076 10724 55086
rect 10668 54982 10724 55020
rect 10556 54786 10612 54796
rect 10332 54516 10388 54526
rect 10332 54514 10724 54516
rect 10332 54462 10334 54514
rect 10386 54462 10724 54514
rect 10332 54460 10724 54462
rect 10332 54450 10388 54460
rect 10220 54236 10388 54292
rect 10220 53844 10276 53854
rect 9436 53618 9828 53620
rect 9436 53566 9438 53618
rect 9490 53566 9828 53618
rect 9436 53564 9828 53566
rect 9436 53554 9492 53564
rect 9548 53172 9604 53182
rect 9436 53116 9548 53172
rect 9604 53116 9716 53172
rect 9436 51828 9492 53116
rect 9548 53106 9604 53116
rect 9660 53058 9716 53116
rect 9772 53170 9828 53564
rect 9996 53554 10052 53564
rect 10108 53788 10220 53844
rect 9772 53118 9774 53170
rect 9826 53118 9828 53170
rect 9772 53106 9828 53118
rect 9660 53006 9662 53058
rect 9714 53006 9716 53058
rect 9660 52994 9716 53006
rect 9884 52946 9940 52958
rect 9884 52894 9886 52946
rect 9938 52894 9940 52946
rect 9884 52276 9940 52894
rect 9884 52210 9940 52220
rect 10108 52388 10164 53788
rect 10220 53750 10276 53788
rect 10220 53060 10276 53070
rect 10220 52946 10276 53004
rect 10220 52894 10222 52946
rect 10274 52894 10276 52946
rect 10220 52882 10276 52894
rect 10332 52724 10388 54236
rect 10556 54180 10612 54190
rect 9436 49140 9492 51772
rect 9548 51716 9604 51726
rect 9548 49922 9604 51660
rect 10108 51490 10164 52332
rect 10220 52668 10388 52724
rect 10444 53732 10500 53742
rect 10444 52722 10500 53676
rect 10556 53618 10612 54124
rect 10668 53842 10724 54460
rect 10668 53790 10670 53842
rect 10722 53790 10724 53842
rect 10668 53778 10724 53790
rect 10556 53566 10558 53618
rect 10610 53566 10612 53618
rect 10556 52948 10612 53566
rect 10780 53730 10836 53742
rect 10780 53678 10782 53730
rect 10834 53678 10836 53730
rect 10780 53508 10836 53678
rect 10780 53442 10836 53452
rect 10556 52882 10612 52892
rect 10892 52834 10948 52846
rect 10892 52782 10894 52834
rect 10946 52782 10948 52834
rect 10444 52670 10446 52722
rect 10498 52670 10500 52722
rect 10220 51940 10276 52668
rect 10332 52276 10388 52286
rect 10332 52182 10388 52220
rect 10220 51884 10388 51940
rect 10108 51438 10110 51490
rect 10162 51438 10164 51490
rect 10108 51426 10164 51438
rect 9996 51380 10052 51390
rect 9996 50708 10052 51324
rect 10220 50708 10276 50718
rect 9996 50706 10276 50708
rect 9996 50654 10222 50706
rect 10274 50654 10276 50706
rect 9996 50652 10276 50654
rect 9996 50034 10052 50652
rect 10220 50642 10276 50652
rect 10332 50260 10388 51884
rect 10332 50194 10388 50204
rect 9996 49982 9998 50034
rect 10050 49982 10052 50034
rect 9996 49970 10052 49982
rect 9548 49870 9550 49922
rect 9602 49870 9604 49922
rect 9548 49858 9604 49870
rect 9772 49810 9828 49822
rect 9772 49758 9774 49810
rect 9826 49758 9828 49810
rect 9772 49588 9828 49758
rect 10108 49812 10164 49822
rect 9772 49522 9828 49532
rect 9884 49698 9940 49710
rect 9884 49646 9886 49698
rect 9938 49646 9940 49698
rect 9548 49140 9604 49150
rect 9436 49138 9604 49140
rect 9436 49086 9550 49138
rect 9602 49086 9604 49138
rect 9436 49084 9604 49086
rect 9436 48468 9492 48478
rect 9436 46114 9492 48412
rect 9548 48466 9604 49084
rect 9548 48414 9550 48466
rect 9602 48414 9604 48466
rect 9548 47908 9604 48414
rect 9772 48242 9828 48254
rect 9772 48190 9774 48242
rect 9826 48190 9828 48242
rect 9660 48132 9716 48142
rect 9660 48038 9716 48076
rect 9548 47842 9604 47852
rect 9548 47572 9604 47582
rect 9772 47572 9828 48190
rect 9548 47570 9828 47572
rect 9548 47518 9550 47570
rect 9602 47518 9828 47570
rect 9548 47516 9828 47518
rect 9548 47460 9604 47516
rect 9548 47394 9604 47404
rect 9884 47236 9940 49646
rect 9996 48802 10052 48814
rect 9996 48750 9998 48802
rect 10050 48750 10052 48802
rect 9996 48692 10052 48750
rect 9996 48626 10052 48636
rect 9996 48468 10052 48478
rect 9996 48374 10052 48412
rect 9996 48020 10052 48030
rect 9996 47346 10052 47964
rect 10108 47908 10164 49756
rect 10444 48468 10500 52670
rect 10668 52724 10724 52734
rect 10668 52386 10724 52668
rect 10892 52724 10948 52782
rect 10892 52658 10948 52668
rect 11004 52612 11060 57374
rect 11564 57426 11620 57486
rect 11564 57374 11566 57426
rect 11618 57374 11620 57426
rect 11564 57362 11620 57374
rect 11418 57260 11682 57270
rect 11474 57204 11522 57260
rect 11578 57204 11626 57260
rect 11418 57194 11682 57204
rect 11788 56306 11844 58380
rect 12012 58100 12068 58382
rect 12012 58034 12068 58044
rect 11900 57650 11956 57662
rect 11900 57598 11902 57650
rect 11954 57598 11956 57650
rect 11900 57540 11956 57598
rect 11900 57474 11956 57484
rect 12012 57538 12068 57550
rect 12012 57486 12014 57538
rect 12066 57486 12068 57538
rect 12012 56980 12068 57486
rect 12012 56914 12068 56924
rect 11788 56254 11790 56306
rect 11842 56254 11844 56306
rect 11788 56242 11844 56254
rect 11900 56644 11956 56654
rect 11900 56306 11956 56588
rect 11900 56254 11902 56306
rect 11954 56254 11956 56306
rect 11900 56242 11956 56254
rect 11228 56196 11284 56206
rect 11228 56102 11284 56140
rect 11452 56196 11508 56206
rect 11452 55860 11508 56140
rect 11676 56082 11732 56094
rect 11676 56030 11678 56082
rect 11730 56030 11732 56082
rect 11676 55860 11732 56030
rect 12012 56084 12068 56094
rect 12124 56084 12180 61180
rect 12348 60788 12404 60798
rect 12348 60674 12404 60732
rect 12348 60622 12350 60674
rect 12402 60622 12404 60674
rect 12236 57988 12292 57998
rect 12236 57650 12292 57932
rect 12236 57598 12238 57650
rect 12290 57598 12292 57650
rect 12236 57204 12292 57598
rect 12236 57138 12292 57148
rect 12236 56532 12292 56542
rect 12236 56194 12292 56476
rect 12236 56142 12238 56194
rect 12290 56142 12292 56194
rect 12236 56130 12292 56142
rect 12012 56082 12180 56084
rect 12012 56030 12014 56082
rect 12066 56030 12180 56082
rect 12012 56028 12180 56030
rect 12012 56018 12068 56028
rect 11676 55804 11844 55860
rect 11452 55794 11508 55804
rect 11418 55692 11682 55702
rect 11474 55636 11522 55692
rect 11578 55636 11626 55692
rect 11418 55626 11682 55636
rect 11340 55524 11396 55534
rect 11228 55188 11284 55198
rect 11340 55188 11396 55468
rect 11676 55524 11732 55534
rect 11788 55524 11844 55804
rect 11676 55522 11844 55524
rect 11676 55470 11678 55522
rect 11730 55470 11844 55522
rect 11676 55468 11844 55470
rect 11676 55458 11732 55468
rect 11228 55186 11396 55188
rect 11228 55134 11230 55186
rect 11282 55134 11396 55186
rect 11228 55132 11396 55134
rect 11564 55188 11620 55198
rect 11228 55122 11284 55132
rect 11564 55094 11620 55132
rect 12012 55188 12068 55226
rect 12012 55122 12068 55132
rect 12012 54964 12068 54974
rect 12124 54964 12180 56028
rect 12068 54908 12180 54964
rect 11418 54124 11682 54134
rect 11474 54068 11522 54124
rect 11578 54068 11626 54124
rect 11418 54058 11682 54068
rect 11900 54068 11956 54078
rect 11116 53844 11172 53854
rect 11116 53730 11172 53788
rect 11788 53844 11844 53854
rect 11788 53750 11844 53788
rect 11116 53678 11118 53730
rect 11170 53678 11172 53730
rect 11116 53666 11172 53678
rect 11228 53732 11284 53742
rect 11228 53170 11284 53676
rect 11900 53730 11956 54012
rect 11900 53678 11902 53730
rect 11954 53678 11956 53730
rect 11900 53666 11956 53678
rect 11228 53118 11230 53170
rect 11282 53118 11284 53170
rect 11228 53106 11284 53118
rect 11676 53506 11732 53518
rect 11676 53454 11678 53506
rect 11730 53454 11732 53506
rect 11116 53060 11172 53070
rect 11116 52948 11172 53004
rect 11116 52892 11284 52948
rect 11228 52612 11284 52892
rect 11340 52724 11396 52734
rect 11676 52724 11732 53454
rect 11788 53508 11844 53518
rect 12012 53508 12068 54908
rect 12348 54516 12404 60622
rect 12460 60788 12516 60798
rect 12796 60788 12852 62132
rect 12460 60786 12852 60788
rect 12460 60734 12462 60786
rect 12514 60734 12852 60786
rect 12460 60732 12852 60734
rect 12460 59778 12516 60732
rect 12908 60676 12964 60686
rect 12460 59726 12462 59778
rect 12514 59726 12516 59778
rect 12460 57988 12516 59726
rect 12796 60620 12908 60676
rect 12572 58660 12628 58670
rect 12572 58548 12628 58604
rect 12684 58548 12740 58558
rect 12572 58546 12740 58548
rect 12572 58494 12686 58546
rect 12738 58494 12740 58546
rect 12572 58492 12740 58494
rect 12684 58482 12740 58492
rect 12572 58324 12628 58334
rect 12572 58230 12628 58268
rect 12796 58212 12852 60620
rect 12908 60610 12964 60620
rect 12908 60340 12964 60350
rect 12908 60114 12964 60284
rect 12908 60062 12910 60114
rect 12962 60062 12964 60114
rect 12908 60050 12964 60062
rect 12908 58996 12964 59006
rect 12908 58434 12964 58940
rect 13020 58548 13076 62300
rect 13020 58482 13076 58492
rect 13132 61348 13188 61358
rect 12908 58382 12910 58434
rect 12962 58382 12964 58434
rect 12908 58370 12964 58382
rect 12796 58156 13076 58212
rect 12460 57922 12516 57932
rect 13020 57874 13076 58156
rect 13020 57822 13022 57874
rect 13074 57822 13076 57874
rect 13020 57810 13076 57822
rect 13132 57764 13188 61292
rect 12460 57650 12516 57662
rect 12460 57598 12462 57650
rect 12514 57598 12516 57650
rect 12460 56980 12516 57598
rect 12460 56914 12516 56924
rect 12684 57204 12740 57214
rect 12572 56084 12628 56094
rect 12572 55990 12628 56028
rect 12236 54460 12404 54516
rect 12460 55522 12516 55534
rect 12460 55470 12462 55522
rect 12514 55470 12516 55522
rect 11844 53452 11956 53508
rect 11788 53442 11844 53452
rect 11340 52722 11732 52724
rect 11340 52670 11342 52722
rect 11394 52670 11732 52722
rect 11340 52668 11732 52670
rect 11788 53284 11844 53294
rect 11340 52658 11396 52668
rect 11004 52556 11172 52612
rect 10668 52334 10670 52386
rect 10722 52334 10724 52386
rect 10668 52322 10724 52334
rect 11004 52388 11060 52398
rect 11004 52294 11060 52332
rect 10556 52276 10612 52286
rect 10556 51716 10612 52220
rect 10556 51660 10948 51716
rect 10668 51492 10724 51502
rect 10556 50708 10612 50718
rect 10556 49922 10612 50652
rect 10668 50706 10724 51436
rect 10668 50654 10670 50706
rect 10722 50654 10724 50706
rect 10668 50642 10724 50654
rect 10556 49870 10558 49922
rect 10610 49870 10612 49922
rect 10556 49858 10612 49870
rect 10668 50036 10724 50046
rect 10892 50036 10948 51660
rect 11116 51604 11172 52556
rect 11228 52274 11284 52556
rect 11418 52556 11682 52566
rect 11474 52500 11522 52556
rect 11578 52500 11626 52556
rect 11418 52490 11682 52500
rect 11228 52222 11230 52274
rect 11282 52222 11284 52274
rect 11228 52210 11284 52222
rect 11788 52164 11844 53228
rect 11900 53058 11956 53452
rect 12012 53442 12068 53452
rect 12124 53506 12180 53518
rect 12124 53454 12126 53506
rect 12178 53454 12180 53506
rect 12124 53396 12180 53454
rect 12124 53330 12180 53340
rect 12124 53060 12180 53070
rect 11900 53006 11902 53058
rect 11954 53006 11956 53058
rect 11900 52994 11956 53006
rect 12012 53004 12124 53060
rect 12012 52388 12068 53004
rect 12124 52966 12180 53004
rect 11116 50706 11172 51548
rect 11676 52108 11844 52164
rect 11900 52332 12068 52388
rect 11676 51156 11732 52108
rect 11676 51090 11732 51100
rect 11418 50988 11682 50998
rect 11474 50932 11522 50988
rect 11578 50932 11626 50988
rect 11418 50922 11682 50932
rect 11900 50820 11956 52332
rect 12012 52162 12068 52174
rect 12012 52110 12014 52162
rect 12066 52110 12068 52162
rect 12012 51156 12068 52110
rect 12124 52164 12180 52174
rect 12124 52070 12180 52108
rect 12012 51090 12068 51100
rect 11116 50654 11118 50706
rect 11170 50654 11172 50706
rect 11004 50036 11060 50046
rect 10892 50034 11060 50036
rect 10892 49982 11006 50034
rect 11058 49982 11060 50034
rect 10892 49980 11060 49982
rect 10556 48804 10612 48814
rect 10556 48710 10612 48748
rect 10444 48402 10500 48412
rect 10668 48132 10724 49980
rect 11004 49970 11060 49980
rect 10780 49810 10836 49822
rect 10780 49758 10782 49810
rect 10834 49758 10836 49810
rect 10780 49588 10836 49758
rect 11004 49700 11060 49710
rect 11004 49606 11060 49644
rect 11116 49588 11172 50654
rect 11452 50764 11956 50820
rect 11452 50594 11508 50764
rect 12236 50596 12292 54460
rect 12460 54404 12516 55470
rect 12572 55412 12628 55422
rect 12572 55318 12628 55356
rect 12348 54402 12516 54404
rect 12348 54350 12462 54402
rect 12514 54350 12516 54402
rect 12348 54348 12516 54350
rect 12348 54068 12404 54348
rect 12460 54338 12516 54348
rect 12684 54180 12740 57148
rect 12796 57092 12852 57102
rect 12796 56082 12852 57036
rect 12908 56978 12964 56990
rect 12908 56926 12910 56978
rect 12962 56926 12964 56978
rect 12908 56532 12964 56926
rect 12908 56466 12964 56476
rect 13132 56306 13188 57708
rect 13132 56254 13134 56306
rect 13186 56254 13188 56306
rect 13132 56242 13188 56254
rect 13244 56196 13300 66780
rect 13468 66276 13524 67116
rect 13580 66948 13636 66958
rect 13692 66948 13748 67790
rect 13916 67620 13972 68796
rect 14028 68628 14084 68638
rect 14028 68534 14084 68572
rect 14028 67730 14084 67742
rect 14028 67678 14030 67730
rect 14082 67678 14084 67730
rect 14028 67620 14084 67678
rect 13972 67564 14084 67620
rect 13916 67554 13972 67564
rect 14028 67396 14084 67406
rect 14140 67396 14196 70588
rect 14252 70082 14308 70812
rect 14364 70532 14420 71484
rect 14476 71204 14532 71214
rect 14476 70978 14532 71148
rect 14476 70926 14478 70978
rect 14530 70926 14532 70978
rect 14476 70914 14532 70926
rect 14812 70756 14868 71932
rect 14924 71540 14980 71550
rect 14924 71202 14980 71484
rect 14924 71150 14926 71202
rect 14978 71150 14980 71202
rect 14924 70980 14980 71150
rect 15036 71204 15092 71932
rect 15148 71988 15204 72380
rect 15260 72434 15316 73388
rect 15260 72382 15262 72434
rect 15314 72382 15316 72434
rect 15260 72324 15316 72382
rect 15260 72258 15316 72268
rect 15372 72212 15428 73836
rect 15596 73890 15652 73902
rect 15596 73838 15598 73890
rect 15650 73838 15652 73890
rect 15596 73556 15652 73838
rect 15148 71986 15316 71988
rect 15148 71934 15150 71986
rect 15202 71934 15316 71986
rect 15148 71932 15316 71934
rect 15148 71922 15204 71932
rect 15148 71204 15204 71214
rect 15036 71202 15204 71204
rect 15036 71150 15150 71202
rect 15202 71150 15204 71202
rect 15036 71148 15204 71150
rect 15148 71138 15204 71148
rect 14924 70914 14980 70924
rect 15260 71092 15316 71932
rect 15372 71540 15428 72156
rect 15484 73108 15540 73118
rect 15484 71764 15540 73052
rect 15596 72884 15652 73500
rect 15596 72818 15652 72828
rect 15596 72548 15652 72558
rect 15708 72548 15764 74060
rect 15820 73444 15876 79660
rect 16380 79604 16436 82012
rect 16604 81282 16660 81294
rect 16604 81230 16606 81282
rect 16658 81230 16660 81282
rect 16604 81172 16660 81230
rect 16492 80948 16548 80958
rect 16492 80854 16548 80892
rect 16492 80500 16548 80510
rect 16604 80500 16660 81116
rect 16492 80498 16660 80500
rect 16492 80446 16494 80498
rect 16546 80446 16660 80498
rect 16492 80444 16660 80446
rect 16828 81282 16884 83244
rect 16940 82068 16996 88284
rect 16940 82002 16996 82012
rect 17052 87892 17108 87902
rect 17052 85652 17108 87836
rect 17276 87332 17332 88396
rect 17724 88340 17780 88846
rect 17276 87266 17332 87276
rect 17388 88284 17780 88340
rect 18060 88340 18116 89180
rect 18172 89012 18228 89022
rect 18284 89012 18340 89180
rect 18172 89010 18340 89012
rect 18172 88958 18174 89010
rect 18226 88958 18340 89010
rect 18172 88956 18340 88958
rect 18172 88946 18228 88956
rect 18396 88900 18452 89628
rect 18396 88834 18452 88844
rect 18508 88788 18564 89964
rect 18620 90018 18900 90020
rect 18620 89966 18846 90018
rect 18898 89966 18900 90018
rect 18620 89964 18900 89966
rect 18620 89236 18676 89964
rect 18844 89954 18900 89964
rect 18620 89142 18676 89180
rect 18844 89236 18900 89246
rect 19068 89236 19124 93100
rect 19180 92932 19236 92942
rect 19404 92932 19460 97692
rect 19852 97524 19908 98252
rect 19516 97188 19572 97198
rect 19516 96290 19572 97132
rect 19628 96740 19684 96750
rect 19852 96740 19908 97468
rect 19964 97860 20020 97870
rect 19964 97522 20020 97804
rect 20076 97636 20132 97646
rect 20076 97542 20132 97580
rect 19964 97470 19966 97522
rect 20018 97470 20020 97522
rect 19964 97458 20020 97470
rect 20188 96964 20244 96974
rect 20188 96870 20244 96908
rect 19628 96738 19796 96740
rect 19628 96686 19630 96738
rect 19682 96686 19796 96738
rect 19628 96684 19796 96686
rect 19628 96674 19684 96684
rect 19516 96238 19518 96290
rect 19570 96238 19572 96290
rect 19516 96226 19572 96238
rect 19740 96292 19796 96684
rect 19852 96674 19908 96684
rect 19628 95956 19684 95966
rect 19516 95058 19572 95070
rect 19516 95006 19518 95058
rect 19570 95006 19572 95058
rect 19516 94724 19572 95006
rect 19516 94658 19572 94668
rect 19628 94610 19684 95900
rect 19740 94724 19796 96236
rect 20188 96628 20244 96638
rect 19852 96068 19908 96078
rect 19852 96066 20020 96068
rect 19852 96014 19854 96066
rect 19906 96014 20020 96066
rect 19852 96012 20020 96014
rect 19852 96002 19908 96012
rect 19740 94658 19796 94668
rect 19852 95844 19908 95854
rect 19852 95058 19908 95788
rect 19852 95006 19854 95058
rect 19906 95006 19908 95058
rect 19628 94558 19630 94610
rect 19682 94558 19684 94610
rect 19236 92876 19348 92932
rect 19404 92876 19572 92932
rect 19180 92866 19236 92876
rect 19292 92708 19348 92876
rect 19404 92708 19460 92718
rect 19292 92706 19460 92708
rect 19292 92654 19406 92706
rect 19458 92654 19460 92706
rect 19292 92652 19460 92654
rect 19404 92642 19460 92652
rect 19404 92484 19460 92494
rect 19292 92036 19348 92046
rect 19180 91924 19236 91934
rect 19180 91362 19236 91868
rect 19180 91310 19182 91362
rect 19234 91310 19236 91362
rect 19180 91298 19236 91310
rect 19292 90804 19348 91980
rect 19404 91362 19460 92428
rect 19404 91310 19406 91362
rect 19458 91310 19460 91362
rect 19404 91298 19460 91310
rect 19404 90804 19460 90814
rect 19292 90748 19404 90804
rect 19404 90710 19460 90748
rect 18844 89234 19124 89236
rect 18844 89182 18846 89234
rect 18898 89182 19124 89234
rect 18844 89180 19124 89182
rect 19292 89570 19348 89582
rect 19292 89518 19294 89570
rect 19346 89518 19348 89570
rect 18844 89170 18900 89180
rect 18732 89012 18788 89022
rect 18956 89012 19012 89022
rect 18732 89010 18900 89012
rect 18732 88958 18734 89010
rect 18786 88958 18900 89010
rect 18732 88956 18900 88958
rect 18732 88946 18788 88956
rect 18844 88788 18900 88956
rect 18956 89010 19124 89012
rect 18956 88958 18958 89010
rect 19010 88958 19124 89010
rect 18956 88956 19124 88958
rect 18956 88946 19012 88956
rect 18956 88788 19012 88798
rect 18508 88732 18788 88788
rect 18844 88732 18956 88788
rect 18222 88620 18486 88630
rect 18278 88564 18326 88620
rect 18382 88564 18430 88620
rect 18222 88554 18486 88564
rect 18060 88284 18340 88340
rect 17276 86658 17332 86670
rect 17276 86606 17278 86658
rect 17330 86606 17332 86658
rect 17276 85988 17332 86606
rect 17276 85922 17332 85932
rect 17052 84420 17108 85596
rect 17388 85314 17444 88284
rect 18284 88226 18340 88284
rect 18284 88174 18286 88226
rect 18338 88174 18340 88226
rect 18284 88162 18340 88174
rect 17724 88116 17780 88126
rect 17724 88022 17780 88060
rect 18060 88116 18116 88126
rect 18060 88022 18116 88060
rect 18508 88116 18564 88126
rect 18508 88022 18564 88060
rect 18620 88114 18676 88126
rect 18620 88062 18622 88114
rect 18674 88062 18676 88114
rect 17612 88004 17668 88014
rect 17500 87668 17556 87678
rect 17500 87574 17556 87612
rect 17388 85262 17390 85314
rect 17442 85262 17444 85314
rect 17388 85250 17444 85262
rect 17612 85202 17668 87948
rect 18620 87892 18676 88062
rect 18620 87826 18676 87836
rect 18396 87442 18452 87454
rect 18396 87390 18398 87442
rect 18450 87390 18452 87442
rect 17836 87332 17892 87342
rect 18396 87332 18452 87390
rect 18396 87276 18676 87332
rect 17836 87238 17892 87276
rect 18060 87218 18116 87230
rect 18060 87166 18062 87218
rect 18114 87166 18116 87218
rect 17948 86884 18004 86894
rect 17612 85150 17614 85202
rect 17666 85150 17668 85202
rect 17612 85138 17668 85150
rect 17836 85762 17892 85774
rect 17836 85710 17838 85762
rect 17890 85710 17892 85762
rect 17164 84980 17220 84990
rect 17612 84980 17668 84990
rect 17836 84980 17892 85710
rect 17948 85708 18004 86828
rect 18060 86548 18116 87166
rect 18222 87052 18486 87062
rect 18278 86996 18326 87052
rect 18382 86996 18430 87052
rect 18222 86986 18486 86996
rect 18620 86660 18676 87276
rect 18620 86594 18676 86604
rect 18060 86492 18228 86548
rect 18172 85764 18228 86492
rect 18732 86436 18788 88732
rect 18956 88722 19012 88732
rect 18844 87780 18900 87790
rect 18844 87666 18900 87724
rect 18844 87614 18846 87666
rect 18898 87614 18900 87666
rect 18844 87602 18900 87614
rect 18956 86884 19012 86894
rect 18956 86790 19012 86828
rect 18844 86436 18900 86446
rect 18732 86434 18900 86436
rect 18732 86382 18846 86434
rect 18898 86382 18900 86434
rect 18732 86380 18900 86382
rect 18844 86370 18900 86380
rect 19068 86212 19124 88956
rect 19180 89010 19236 89022
rect 19180 88958 19182 89010
rect 19234 88958 19236 89010
rect 19180 88788 19236 88958
rect 19292 89012 19348 89518
rect 19292 88946 19348 88956
rect 19404 88788 19460 88798
rect 19180 88786 19460 88788
rect 19180 88734 19406 88786
rect 19458 88734 19460 88786
rect 19180 88732 19460 88734
rect 19404 88722 19460 88732
rect 19516 88564 19572 92876
rect 19628 92372 19684 94558
rect 19740 94388 19796 94398
rect 19852 94388 19908 95006
rect 19796 94332 19908 94388
rect 19740 94322 19796 94332
rect 19628 92306 19684 92316
rect 19740 94164 19796 94174
rect 19740 92930 19796 94108
rect 19964 93042 20020 96012
rect 20076 95956 20132 95966
rect 20076 95862 20132 95900
rect 20076 95732 20132 95742
rect 20076 95394 20132 95676
rect 20076 95342 20078 95394
rect 20130 95342 20132 95394
rect 20076 95330 20132 95342
rect 20188 95172 20244 96572
rect 19964 92990 19966 93042
rect 20018 92990 20020 93042
rect 19964 92978 20020 92990
rect 20076 95116 20244 95172
rect 19740 92878 19742 92930
rect 19794 92878 19796 92930
rect 19740 92484 19796 92878
rect 19852 92932 19908 92942
rect 19852 92820 19908 92876
rect 19964 92820 20020 92830
rect 19852 92818 20020 92820
rect 19852 92766 19966 92818
rect 20018 92766 20020 92818
rect 19852 92764 20020 92766
rect 19964 92754 20020 92764
rect 19628 91252 19684 91262
rect 19628 89794 19684 91196
rect 19740 90580 19796 92428
rect 19964 90804 20020 90814
rect 19964 90710 20020 90748
rect 20076 90690 20132 95116
rect 20300 93714 20356 93726
rect 20300 93662 20302 93714
rect 20354 93662 20356 93714
rect 20300 93604 20356 93662
rect 20300 93538 20356 93548
rect 20412 93044 20468 102286
rect 20972 102340 21028 102350
rect 20748 100546 20804 100558
rect 20748 100494 20750 100546
rect 20802 100494 20804 100546
rect 20636 99540 20692 99550
rect 20636 99314 20692 99484
rect 20636 99262 20638 99314
rect 20690 99262 20692 99314
rect 20636 99250 20692 99262
rect 20748 99092 20804 100494
rect 20748 99026 20804 99036
rect 20860 98530 20916 98542
rect 20860 98478 20862 98530
rect 20914 98478 20916 98530
rect 20524 98196 20580 98206
rect 20524 98194 20804 98196
rect 20524 98142 20526 98194
rect 20578 98142 20804 98194
rect 20524 98140 20804 98142
rect 20524 98130 20580 98140
rect 20636 97410 20692 97422
rect 20636 97358 20638 97410
rect 20690 97358 20692 97410
rect 20524 96628 20580 96638
rect 20524 96534 20580 96572
rect 20636 96180 20692 97358
rect 20636 96114 20692 96124
rect 20636 95956 20692 95966
rect 20636 95862 20692 95900
rect 20524 95508 20580 95518
rect 20524 95414 20580 95452
rect 20748 93940 20804 98140
rect 20860 97636 20916 98478
rect 20860 96962 20916 97580
rect 20860 96910 20862 96962
rect 20914 96910 20916 96962
rect 20860 96068 20916 96910
rect 20860 96002 20916 96012
rect 20748 93874 20804 93884
rect 20972 94612 21028 102284
rect 21084 99204 21140 102508
rect 21532 102340 21588 102350
rect 21756 102340 21812 102508
rect 22540 102498 22596 102508
rect 22764 102452 22820 102462
rect 22820 102396 23044 102452
rect 22764 102358 22820 102396
rect 21532 102338 21812 102340
rect 21532 102286 21534 102338
rect 21586 102286 21812 102338
rect 21532 102284 21812 102286
rect 21868 102340 21924 102350
rect 21532 102274 21588 102284
rect 21868 102246 21924 102284
rect 21308 102116 21364 102126
rect 21196 102114 21364 102116
rect 21196 102062 21310 102114
rect 21362 102062 21364 102114
rect 21196 102060 21364 102062
rect 21196 100098 21252 102060
rect 21308 102050 21364 102060
rect 21420 102114 21476 102126
rect 21420 102062 21422 102114
rect 21474 102062 21476 102114
rect 21196 100046 21198 100098
rect 21250 100046 21252 100098
rect 21196 100034 21252 100046
rect 21308 101556 21364 101566
rect 21308 100882 21364 101500
rect 21308 100830 21310 100882
rect 21362 100830 21364 100882
rect 21084 95844 21140 99148
rect 21308 99204 21364 100830
rect 21420 100660 21476 102062
rect 22204 102114 22260 102126
rect 22204 102062 22206 102114
rect 22258 102062 22260 102114
rect 21624 101948 21888 101958
rect 21680 101892 21728 101948
rect 21784 101892 21832 101948
rect 21624 101882 21888 101892
rect 22204 101554 22260 102062
rect 22204 101502 22206 101554
rect 22258 101502 22260 101554
rect 22204 101490 22260 101502
rect 21868 100772 21924 100782
rect 21924 100716 22036 100772
rect 21868 100706 21924 100716
rect 21420 100594 21476 100604
rect 21624 100380 21888 100390
rect 21680 100324 21728 100380
rect 21784 100324 21832 100380
rect 21624 100314 21888 100324
rect 21980 99764 22036 100716
rect 21868 99708 22036 99764
rect 22316 99988 22372 99998
rect 22876 99988 22932 99998
rect 21532 99204 21588 99214
rect 21308 99202 21588 99204
rect 21308 99150 21534 99202
rect 21586 99150 21588 99202
rect 21308 99148 21588 99150
rect 21196 98532 21252 98542
rect 21196 98438 21252 98476
rect 21308 96962 21364 99148
rect 21532 99138 21588 99148
rect 21756 99204 21812 99214
rect 21756 99110 21812 99148
rect 21868 99202 21924 99708
rect 22316 99426 22372 99932
rect 22316 99374 22318 99426
rect 22370 99374 22372 99426
rect 22316 99362 22372 99374
rect 22764 99986 22932 99988
rect 22764 99934 22878 99986
rect 22930 99934 22932 99986
rect 22764 99932 22932 99934
rect 21868 99150 21870 99202
rect 21922 99150 21924 99202
rect 21868 99138 21924 99150
rect 21980 99092 22036 99102
rect 21624 98812 21888 98822
rect 21680 98756 21728 98812
rect 21784 98756 21832 98812
rect 21624 98746 21888 98756
rect 21868 98644 21924 98654
rect 21868 98550 21924 98588
rect 21868 98196 21924 98206
rect 21868 97746 21924 98140
rect 21868 97694 21870 97746
rect 21922 97694 21924 97746
rect 21868 97682 21924 97694
rect 21980 97860 22036 99036
rect 22764 98980 22820 99932
rect 22876 99922 22932 99932
rect 22764 98642 22820 98924
rect 22764 98590 22766 98642
rect 22818 98590 22820 98642
rect 22764 98578 22820 98590
rect 22876 99202 22932 99214
rect 22876 99150 22878 99202
rect 22930 99150 22932 99202
rect 21420 97524 21476 97534
rect 21420 97430 21476 97468
rect 21624 97244 21888 97254
rect 21680 97188 21728 97244
rect 21784 97188 21832 97244
rect 21624 97178 21888 97188
rect 21308 96910 21310 96962
rect 21362 96910 21364 96962
rect 21308 96852 21364 96910
rect 21308 96786 21364 96796
rect 21868 96292 21924 96302
rect 21980 96292 22036 97804
rect 22204 98532 22260 98542
rect 22204 97636 22260 98476
rect 22316 98306 22372 98318
rect 22316 98254 22318 98306
rect 22370 98254 22372 98306
rect 22316 98194 22372 98254
rect 22316 98142 22318 98194
rect 22370 98142 22372 98194
rect 22316 98130 22372 98142
rect 22540 97748 22596 97758
rect 22876 97748 22932 99150
rect 22596 97692 22932 97748
rect 22540 97654 22596 97692
rect 22092 96852 22148 96862
rect 22092 96758 22148 96796
rect 21868 96290 22036 96292
rect 21868 96238 21870 96290
rect 21922 96238 22036 96290
rect 21868 96236 22036 96238
rect 22092 96292 22148 96302
rect 22204 96292 22260 97580
rect 22876 97524 22932 97562
rect 22876 97458 22932 97468
rect 22652 96964 22708 96974
rect 22652 96962 22820 96964
rect 22652 96910 22654 96962
rect 22706 96910 22820 96962
rect 22652 96908 22820 96910
rect 22652 96898 22708 96908
rect 22092 96290 22260 96292
rect 22092 96238 22094 96290
rect 22146 96238 22260 96290
rect 22092 96236 22260 96238
rect 22764 96290 22820 96908
rect 22764 96238 22766 96290
rect 22818 96238 22820 96290
rect 21868 96226 21924 96236
rect 22092 96226 22148 96236
rect 22764 96226 22820 96238
rect 22316 96066 22372 96078
rect 22316 96014 22318 96066
rect 22370 96014 22372 96066
rect 21084 95778 21140 95788
rect 21644 95954 21700 95966
rect 21644 95902 21646 95954
rect 21698 95902 21700 95954
rect 21644 95844 21700 95902
rect 22316 95956 22372 96014
rect 22316 95890 22372 95900
rect 21644 95778 21700 95788
rect 21624 95676 21888 95686
rect 21680 95620 21728 95676
rect 21784 95620 21832 95676
rect 21624 95610 21888 95620
rect 20972 93938 21028 94556
rect 21756 94556 22036 94612
rect 20972 93886 20974 93938
rect 21026 93886 21028 93938
rect 20972 93874 21028 93886
rect 21196 94498 21252 94510
rect 21196 94446 21198 94498
rect 21250 94446 21252 94498
rect 20524 93716 20580 93726
rect 20524 93622 20580 93660
rect 20412 92988 20916 93044
rect 20412 92818 20468 92830
rect 20412 92766 20414 92818
rect 20466 92766 20468 92818
rect 20188 92708 20244 92718
rect 20188 92614 20244 92652
rect 20412 92370 20468 92766
rect 20412 92318 20414 92370
rect 20466 92318 20468 92370
rect 20412 92306 20468 92318
rect 20636 92708 20692 92718
rect 20300 92260 20356 92270
rect 20300 91252 20356 92204
rect 20636 92258 20692 92652
rect 20636 92206 20638 92258
rect 20690 92206 20692 92258
rect 20636 92194 20692 92206
rect 20748 92484 20804 92494
rect 20748 92146 20804 92428
rect 20748 92094 20750 92146
rect 20802 92094 20804 92146
rect 20748 92082 20804 92094
rect 20300 90916 20356 91196
rect 20300 90860 20692 90916
rect 20076 90638 20078 90690
rect 20130 90638 20132 90690
rect 20076 90626 20132 90638
rect 19740 90486 19796 90524
rect 20188 90580 20244 90590
rect 20188 90578 20356 90580
rect 20188 90526 20190 90578
rect 20242 90526 20356 90578
rect 20188 90524 20356 90526
rect 20188 90514 20244 90524
rect 20188 90356 20244 90366
rect 20188 89796 20244 90300
rect 19628 89742 19630 89794
rect 19682 89742 19684 89794
rect 19628 89348 19684 89742
rect 20076 89794 20244 89796
rect 20076 89742 20190 89794
rect 20242 89742 20244 89794
rect 20076 89740 20244 89742
rect 19964 89684 20020 89694
rect 19964 89590 20020 89628
rect 19628 89282 19684 89292
rect 19740 89570 19796 89582
rect 19740 89518 19742 89570
rect 19794 89518 19796 89570
rect 19628 88898 19684 88910
rect 19628 88846 19630 88898
rect 19682 88846 19684 88898
rect 19628 88788 19684 88846
rect 19628 88722 19684 88732
rect 19740 88786 19796 89518
rect 20076 89348 20132 89740
rect 20188 89730 20244 89740
rect 19740 88734 19742 88786
rect 19794 88734 19796 88786
rect 19740 88722 19796 88734
rect 19852 89292 20132 89348
rect 19404 88508 19572 88564
rect 19292 88228 19348 88238
rect 19292 88134 19348 88172
rect 19180 88116 19236 88126
rect 19180 88022 19236 88060
rect 19404 87668 19460 88508
rect 19180 86660 19236 86670
rect 19180 86566 19236 86604
rect 18844 86156 19124 86212
rect 17948 85652 18116 85708
rect 18172 85698 18228 85708
rect 18732 85876 18788 85886
rect 18060 85316 18116 85652
rect 18222 85484 18486 85494
rect 18278 85428 18326 85484
rect 18382 85428 18430 85484
rect 18222 85418 18486 85428
rect 18172 85316 18228 85326
rect 18060 85314 18228 85316
rect 18060 85262 18174 85314
rect 18226 85262 18228 85314
rect 18060 85260 18228 85262
rect 18172 85250 18228 85260
rect 17164 84978 17892 84980
rect 17164 84926 17166 84978
rect 17218 84926 17614 84978
rect 17666 84926 17892 84978
rect 17164 84924 17892 84926
rect 17164 84914 17220 84924
rect 17612 84914 17668 84924
rect 16828 81230 16830 81282
rect 16882 81230 16884 81282
rect 16492 80434 16548 80444
rect 16268 79602 16436 79604
rect 16268 79550 16382 79602
rect 16434 79550 16436 79602
rect 16268 79548 16436 79550
rect 15932 75348 15988 75358
rect 15932 75122 15988 75292
rect 15932 75070 15934 75122
rect 15986 75070 15988 75122
rect 15932 75058 15988 75070
rect 16044 74676 16100 74686
rect 16044 74002 16100 74620
rect 16268 74674 16324 79548
rect 16380 79538 16436 79548
rect 16604 79604 16660 79614
rect 16492 76468 16548 76478
rect 16380 75794 16436 75806
rect 16380 75742 16382 75794
rect 16434 75742 16436 75794
rect 16380 75124 16436 75742
rect 16380 75058 16436 75068
rect 16380 74900 16436 74910
rect 16492 74900 16548 76412
rect 16380 74898 16548 74900
rect 16380 74846 16382 74898
rect 16434 74846 16548 74898
rect 16380 74844 16548 74846
rect 16380 74834 16436 74844
rect 16268 74622 16270 74674
rect 16322 74622 16324 74674
rect 16268 74610 16324 74622
rect 16492 74676 16548 74844
rect 16492 74610 16548 74620
rect 16044 73950 16046 74002
rect 16098 73950 16100 74002
rect 16044 73938 16100 73950
rect 15820 73378 15876 73388
rect 15932 73330 15988 73342
rect 15932 73278 15934 73330
rect 15986 73278 15988 73330
rect 15820 73220 15876 73230
rect 15932 73220 15988 73278
rect 15876 73164 15988 73220
rect 16380 73220 16436 73230
rect 16380 73218 16548 73220
rect 16380 73166 16382 73218
rect 16434 73166 16548 73218
rect 16380 73164 16548 73166
rect 15820 73154 15876 73164
rect 16380 73154 16436 73164
rect 15596 72546 15764 72548
rect 15596 72494 15598 72546
rect 15650 72494 15764 72546
rect 15596 72492 15764 72494
rect 16268 72660 16324 72670
rect 15596 72324 15652 72492
rect 15932 72436 15988 72446
rect 15988 72380 16100 72436
rect 15932 72370 15988 72380
rect 15596 72258 15652 72268
rect 16044 71988 16100 72380
rect 16268 72434 16324 72604
rect 16380 72548 16436 72558
rect 16380 72454 16436 72492
rect 16268 72382 16270 72434
rect 16322 72382 16324 72434
rect 16268 72370 16324 72382
rect 15932 71932 16100 71988
rect 16380 72100 16436 72110
rect 15484 71698 15540 71708
rect 15708 71764 15764 71774
rect 15708 71670 15764 71708
rect 15932 71762 15988 71932
rect 16380 71874 16436 72044
rect 16492 71988 16548 73164
rect 16492 71922 16548 71932
rect 16380 71822 16382 71874
rect 16434 71822 16436 71874
rect 16380 71810 16436 71822
rect 16156 71764 16212 71774
rect 15932 71710 15934 71762
rect 15986 71710 15988 71762
rect 15932 71698 15988 71710
rect 16044 71762 16212 71764
rect 16044 71710 16158 71762
rect 16210 71710 16212 71762
rect 16044 71708 16212 71710
rect 15484 71540 15540 71550
rect 15428 71538 15540 71540
rect 15428 71486 15486 71538
rect 15538 71486 15540 71538
rect 15428 71484 15540 71486
rect 15372 71446 15428 71484
rect 15484 71474 15540 71484
rect 16044 71316 16100 71708
rect 16156 71698 16212 71708
rect 16268 71652 16324 71662
rect 16492 71652 16548 71662
rect 16268 71650 16436 71652
rect 16268 71598 16270 71650
rect 16322 71598 16436 71650
rect 16268 71596 16436 71598
rect 16268 71586 16324 71596
rect 15596 71260 16100 71316
rect 16156 71540 16212 71550
rect 15372 71092 15428 71102
rect 15260 71090 15428 71092
rect 15260 71038 15374 71090
rect 15426 71038 15428 71090
rect 15260 71036 15428 71038
rect 15260 70756 15316 71036
rect 15372 71026 15428 71036
rect 14700 70700 14868 70756
rect 15148 70700 15316 70756
rect 15484 70868 15540 70878
rect 14588 70532 14644 70542
rect 14364 70476 14532 70532
rect 14252 70030 14254 70082
rect 14306 70030 14308 70082
rect 14252 70018 14308 70030
rect 14252 68516 14308 68526
rect 14252 68514 14420 68516
rect 14252 68462 14254 68514
rect 14306 68462 14420 68514
rect 14252 68460 14420 68462
rect 14252 68450 14308 68460
rect 14084 67340 14196 67396
rect 14028 67282 14084 67340
rect 14028 67230 14030 67282
rect 14082 67230 14084 67282
rect 14028 67218 14084 67230
rect 13580 66946 13748 66948
rect 13580 66894 13582 66946
rect 13634 66894 13748 66946
rect 13580 66892 13748 66894
rect 13580 66500 13636 66892
rect 13580 66434 13636 66444
rect 13804 66276 13860 66286
rect 13468 66182 13524 66220
rect 13580 66220 13804 66276
rect 13580 65714 13636 66220
rect 13804 66210 13860 66220
rect 14252 66276 14308 66286
rect 14252 66182 14308 66220
rect 13580 65662 13582 65714
rect 13634 65662 13636 65714
rect 13580 65650 13636 65662
rect 13692 66052 13748 66062
rect 13468 65604 13524 65614
rect 13468 65510 13524 65548
rect 13580 64484 13636 64494
rect 13468 64482 13636 64484
rect 13468 64430 13582 64482
rect 13634 64430 13636 64482
rect 13468 64428 13636 64430
rect 13356 63924 13412 63934
rect 13468 63924 13524 64428
rect 13580 64418 13636 64428
rect 13580 64148 13636 64158
rect 13692 64148 13748 65996
rect 13804 65490 13860 65502
rect 13804 65438 13806 65490
rect 13858 65438 13860 65490
rect 13804 65380 13860 65438
rect 13804 65314 13860 65324
rect 14028 65490 14084 65502
rect 14028 65438 14030 65490
rect 14082 65438 14084 65490
rect 14028 65380 14084 65438
rect 14364 65492 14420 68460
rect 14476 68292 14532 70476
rect 14588 68852 14644 70476
rect 14700 69188 14756 70700
rect 14820 70588 15084 70598
rect 14876 70532 14924 70588
rect 14980 70532 15028 70588
rect 14820 70522 15084 70532
rect 15036 70306 15092 70318
rect 15036 70254 15038 70306
rect 15090 70254 15092 70306
rect 15036 70084 15092 70254
rect 15148 70196 15204 70700
rect 15148 70130 15204 70140
rect 15260 70194 15316 70206
rect 15260 70142 15262 70194
rect 15314 70142 15316 70194
rect 15260 70084 15316 70142
rect 15484 70196 15540 70812
rect 15596 70754 15652 71260
rect 16044 70980 16100 70990
rect 15596 70702 15598 70754
rect 15650 70702 15652 70754
rect 15596 70644 15652 70702
rect 15596 70578 15652 70588
rect 15708 70754 15764 70766
rect 15708 70702 15710 70754
rect 15762 70702 15764 70754
rect 15596 70196 15652 70206
rect 15484 70194 15652 70196
rect 15484 70142 15598 70194
rect 15650 70142 15652 70194
rect 15484 70140 15652 70142
rect 15260 70028 15540 70084
rect 15036 69524 15092 70028
rect 15484 69972 15540 70028
rect 15092 69468 15428 69524
rect 15036 69430 15092 69468
rect 14812 69412 14868 69422
rect 14812 69318 14868 69356
rect 15260 69300 15316 69310
rect 15260 69206 15316 69244
rect 14700 69122 14756 69132
rect 14820 69020 15084 69030
rect 14876 68964 14924 69020
rect 14980 68964 15028 69020
rect 14820 68954 15084 68964
rect 14924 68852 14980 68862
rect 14588 68850 14980 68852
rect 14588 68798 14926 68850
rect 14978 68798 14980 68850
rect 14588 68796 14980 68798
rect 14588 68628 14644 68796
rect 14924 68786 14980 68796
rect 15372 68850 15428 69468
rect 15484 68964 15540 69916
rect 15596 69188 15652 70140
rect 15708 69412 15764 70702
rect 15820 70754 15876 70766
rect 15820 70702 15822 70754
rect 15874 70702 15876 70754
rect 15820 69972 15876 70702
rect 15820 69906 15876 69916
rect 15932 70306 15988 70318
rect 15932 70254 15934 70306
rect 15986 70254 15988 70306
rect 15932 69524 15988 70254
rect 16044 70084 16100 70924
rect 16156 70868 16212 71484
rect 16380 70980 16436 71596
rect 16380 70914 16436 70924
rect 16268 70868 16324 70878
rect 16156 70866 16324 70868
rect 16156 70814 16270 70866
rect 16322 70814 16324 70866
rect 16156 70812 16324 70814
rect 16268 70802 16324 70812
rect 16492 70588 16548 71596
rect 16380 70532 16548 70588
rect 16044 70028 16324 70084
rect 15932 69458 15988 69468
rect 15820 69412 15876 69422
rect 15708 69410 15876 69412
rect 15708 69358 15822 69410
rect 15874 69358 15876 69410
rect 15708 69356 15876 69358
rect 15820 69346 15876 69356
rect 16268 69410 16324 70028
rect 16268 69358 16270 69410
rect 16322 69358 16324 69410
rect 16268 69346 16324 69358
rect 16156 69300 16212 69310
rect 15596 69122 15652 69132
rect 15932 69244 16156 69300
rect 15596 68964 15652 68974
rect 15484 68908 15596 68964
rect 15596 68898 15652 68908
rect 15372 68798 15374 68850
rect 15426 68798 15428 68850
rect 15372 68786 15428 68798
rect 15820 68740 15876 68750
rect 14588 68562 14644 68572
rect 15708 68684 15820 68740
rect 14476 67618 14532 68236
rect 14476 67566 14478 67618
rect 14530 67566 14532 67618
rect 14476 65828 14532 67566
rect 14820 67452 15084 67462
rect 14876 67396 14924 67452
rect 14980 67396 15028 67452
rect 14820 67386 15084 67396
rect 15260 66946 15316 66958
rect 15260 66894 15262 66946
rect 15314 66894 15316 66946
rect 15260 66388 15316 66894
rect 15708 66948 15764 68684
rect 15820 68674 15876 68684
rect 15820 67172 15876 67182
rect 15932 67172 15988 69244
rect 16156 69234 16212 69244
rect 16268 69188 16324 69198
rect 15820 67170 15988 67172
rect 15820 67118 15822 67170
rect 15874 67118 15988 67170
rect 15820 67116 15988 67118
rect 16044 68628 16100 68638
rect 16044 67954 16100 68572
rect 16044 67902 16046 67954
rect 16098 67902 16100 67954
rect 15820 67106 15876 67116
rect 16044 67060 16100 67902
rect 16156 67060 16212 67070
rect 16044 67058 16212 67060
rect 16044 67006 16158 67058
rect 16210 67006 16212 67058
rect 16044 67004 16212 67006
rect 16156 66994 16212 67004
rect 15708 66892 15988 66948
rect 15484 66836 15540 66846
rect 15484 66742 15540 66780
rect 14820 65884 15084 65894
rect 14876 65828 14924 65884
rect 14980 65828 15028 65884
rect 14820 65818 15084 65828
rect 14476 65762 14532 65772
rect 14700 65716 14756 65726
rect 15260 65716 15316 66332
rect 15932 65716 15988 66892
rect 16268 66836 16324 69132
rect 16380 67060 16436 70532
rect 16492 69522 16548 69534
rect 16492 69470 16494 69522
rect 16546 69470 16548 69522
rect 16492 67396 16548 69470
rect 16492 67330 16548 67340
rect 16380 67004 16548 67060
rect 14700 65714 15316 65716
rect 14700 65662 14702 65714
rect 14754 65662 15316 65714
rect 14700 65660 15316 65662
rect 15372 65714 15988 65716
rect 15372 65662 15934 65714
rect 15986 65662 15988 65714
rect 15372 65660 15988 65662
rect 14700 65650 14756 65660
rect 14476 65604 14532 65614
rect 14476 65510 14532 65548
rect 14364 65426 14420 65436
rect 14588 65492 14644 65502
rect 15148 65492 15204 65502
rect 15372 65492 15428 65660
rect 15932 65650 15988 65660
rect 16044 66780 16324 66836
rect 16380 66836 16436 66846
rect 14588 65490 14868 65492
rect 14588 65438 14590 65490
rect 14642 65438 14868 65490
rect 14588 65436 14868 65438
rect 14588 65426 14644 65436
rect 14028 65314 14084 65324
rect 14812 65380 14868 65436
rect 15148 65490 15428 65492
rect 15148 65438 15150 65490
rect 15202 65438 15428 65490
rect 15148 65436 15428 65438
rect 15484 65492 15540 65502
rect 15148 65426 15204 65436
rect 14812 65314 14868 65324
rect 15484 65378 15540 65436
rect 15484 65326 15486 65378
rect 15538 65326 15540 65378
rect 15484 65266 15540 65326
rect 15484 65214 15486 65266
rect 15538 65214 15540 65266
rect 15484 65202 15540 65214
rect 15596 64820 15652 64830
rect 14252 64484 14308 64494
rect 14252 64390 14308 64428
rect 14820 64316 15084 64326
rect 14876 64260 14924 64316
rect 14980 64260 15028 64316
rect 14820 64250 15084 64260
rect 13580 64146 13748 64148
rect 13580 64094 13582 64146
rect 13634 64094 13748 64146
rect 13580 64092 13748 64094
rect 13580 64082 13636 64092
rect 13412 63868 13524 63924
rect 13692 63924 13748 64092
rect 13916 63924 13972 63934
rect 13692 63922 13972 63924
rect 13692 63870 13918 63922
rect 13970 63870 13972 63922
rect 13692 63868 13972 63870
rect 13356 62580 13412 63868
rect 13916 63858 13972 63868
rect 14700 63812 14756 63822
rect 14700 63810 15092 63812
rect 14700 63758 14702 63810
rect 14754 63758 15092 63810
rect 14700 63756 15092 63758
rect 14700 63746 14756 63756
rect 13916 63700 13972 63710
rect 13468 63140 13524 63150
rect 13468 63046 13524 63084
rect 13916 63140 13972 63644
rect 14924 63588 14980 63598
rect 14476 63364 14532 63374
rect 14476 63250 14532 63308
rect 14476 63198 14478 63250
rect 14530 63198 14532 63250
rect 14476 63186 14532 63198
rect 14924 63250 14980 63532
rect 14924 63198 14926 63250
rect 14978 63198 14980 63250
rect 14924 63140 14980 63198
rect 15036 63252 15092 63756
rect 15484 63364 15540 63374
rect 15148 63308 15428 63364
rect 15148 63252 15204 63308
rect 15036 63196 15204 63252
rect 15372 63250 15428 63308
rect 15372 63198 15374 63250
rect 15426 63198 15428 63250
rect 15372 63186 15428 63198
rect 15260 63140 15316 63150
rect 14924 63138 15316 63140
rect 14924 63086 15262 63138
rect 15314 63086 15316 63138
rect 14924 63084 15316 63086
rect 13580 62916 13636 62926
rect 13580 62914 13860 62916
rect 13580 62862 13582 62914
rect 13634 62862 13860 62914
rect 13580 62860 13860 62862
rect 13580 62850 13636 62860
rect 13580 62580 13636 62590
rect 13356 62578 13636 62580
rect 13356 62526 13582 62578
rect 13634 62526 13636 62578
rect 13356 62524 13636 62526
rect 13580 62514 13636 62524
rect 13804 62244 13860 62860
rect 13916 62692 13972 63084
rect 15260 63074 15316 63084
rect 15484 63138 15540 63308
rect 15484 63086 15486 63138
rect 15538 63086 15540 63138
rect 15484 63074 15540 63086
rect 14028 62916 14084 62926
rect 15596 62916 15652 64764
rect 15820 63476 15876 63486
rect 15820 63138 15876 63420
rect 15820 63086 15822 63138
rect 15874 63086 15876 63138
rect 15820 63074 15876 63086
rect 14028 62822 14084 62860
rect 15484 62860 15652 62916
rect 14820 62748 15084 62758
rect 14876 62692 14924 62748
rect 14980 62692 15028 62748
rect 14820 62682 15084 62692
rect 13916 62626 13972 62636
rect 14476 62466 14532 62478
rect 14476 62414 14478 62466
rect 14530 62414 14532 62466
rect 14364 62356 14420 62366
rect 14364 62262 14420 62300
rect 13804 62188 14196 62244
rect 14476 62188 14532 62414
rect 13580 61796 13636 61806
rect 13580 61682 13636 61740
rect 13580 61630 13582 61682
rect 13634 61630 13636 61682
rect 13580 61618 13636 61630
rect 14140 61570 14196 62188
rect 14364 62132 14532 62188
rect 14700 62354 14756 62366
rect 14700 62302 14702 62354
rect 14754 62302 14756 62354
rect 14364 61908 14420 62132
rect 14364 61842 14420 61852
rect 14140 61518 14142 61570
rect 14194 61518 14196 61570
rect 14140 61506 14196 61518
rect 14476 61794 14532 61806
rect 14476 61742 14478 61794
rect 14530 61742 14532 61794
rect 13916 61460 13972 61470
rect 14476 61460 14532 61742
rect 13804 60898 13860 60910
rect 13804 60846 13806 60898
rect 13858 60846 13860 60898
rect 13804 60788 13860 60846
rect 13804 60722 13860 60732
rect 13916 60674 13972 61404
rect 14252 61404 14532 61460
rect 14140 61348 14196 61358
rect 13916 60622 13918 60674
rect 13970 60622 13972 60674
rect 13916 60610 13972 60622
rect 14028 60788 14084 60798
rect 13692 60228 13748 60238
rect 13468 60004 13524 60014
rect 13692 60004 13748 60172
rect 13468 60002 13748 60004
rect 13468 59950 13470 60002
rect 13522 59950 13748 60002
rect 13468 59948 13748 59950
rect 13468 59938 13524 59948
rect 13580 59778 13636 59790
rect 13580 59726 13582 59778
rect 13634 59726 13636 59778
rect 13356 59108 13412 59118
rect 13580 59108 13636 59726
rect 13356 59106 13636 59108
rect 13356 59054 13358 59106
rect 13410 59054 13636 59106
rect 13356 59052 13636 59054
rect 13356 58996 13412 59052
rect 13356 58930 13412 58940
rect 13692 58828 13748 59948
rect 13804 60004 13860 60014
rect 14028 60004 14084 60732
rect 14140 60786 14196 61292
rect 14140 60734 14142 60786
rect 14194 60734 14196 60786
rect 14140 60722 14196 60734
rect 14252 60452 14308 61404
rect 14700 61012 14756 62302
rect 15372 62356 15428 62366
rect 15372 62130 15428 62300
rect 15372 62078 15374 62130
rect 15426 62078 15428 62130
rect 15372 62066 15428 62078
rect 14924 61572 14980 61582
rect 14924 61478 14980 61516
rect 15260 61572 15316 61582
rect 15260 61478 15316 61516
rect 14820 61180 15084 61190
rect 14876 61124 14924 61180
rect 14980 61124 15028 61180
rect 14820 61114 15084 61124
rect 14700 60956 14868 61012
rect 14252 60386 14308 60396
rect 14364 60788 14420 60798
rect 14364 60226 14420 60732
rect 14364 60174 14366 60226
rect 14418 60174 14420 60226
rect 14364 60162 14420 60174
rect 14252 60116 14308 60126
rect 13804 60002 13972 60004
rect 13804 59950 13806 60002
rect 13858 59950 13972 60002
rect 13804 59948 13972 59950
rect 14028 59948 14196 60004
rect 13804 59938 13860 59948
rect 13916 59892 13972 59948
rect 13916 59826 13972 59836
rect 13804 59780 13860 59790
rect 13804 59442 13860 59724
rect 13804 59390 13806 59442
rect 13858 59390 13860 59442
rect 13804 59378 13860 59390
rect 14028 59780 14084 59790
rect 14028 58996 14084 59724
rect 14140 59218 14196 59948
rect 14252 60002 14308 60060
rect 14252 59950 14254 60002
rect 14306 59950 14308 60002
rect 14252 59938 14308 59950
rect 14364 60004 14420 60014
rect 14140 59166 14142 59218
rect 14194 59166 14196 59218
rect 14140 59154 14196 59166
rect 14028 58940 14308 58996
rect 13580 58772 13636 58782
rect 13692 58772 14196 58828
rect 13580 58210 13636 58716
rect 13804 58548 13860 58558
rect 13580 58158 13582 58210
rect 13634 58158 13636 58210
rect 13468 57876 13524 57886
rect 13468 57782 13524 57820
rect 13580 57428 13636 58158
rect 13580 57362 13636 57372
rect 13692 58492 13804 58548
rect 13692 57204 13748 58492
rect 13804 58482 13860 58492
rect 14028 58324 14084 58334
rect 14028 58230 14084 58268
rect 12796 56030 12798 56082
rect 12850 56030 12852 56082
rect 12796 55524 12852 56030
rect 12908 56084 12964 56094
rect 12908 55990 12964 56028
rect 13020 56082 13076 56094
rect 13020 56030 13022 56082
rect 13074 56030 13076 56082
rect 12796 55458 12852 55468
rect 12908 55748 12964 55758
rect 12908 55074 12964 55692
rect 13020 55522 13076 56030
rect 13020 55470 13022 55522
rect 13074 55470 13076 55522
rect 13020 55458 13076 55470
rect 12908 55022 12910 55074
rect 12962 55022 12964 55074
rect 12796 54628 12852 54638
rect 12796 54534 12852 54572
rect 12348 54002 12404 54012
rect 12460 54124 12740 54180
rect 12348 53620 12404 53630
rect 12348 52612 12404 53564
rect 12348 52546 12404 52556
rect 11452 50542 11454 50594
rect 11506 50542 11508 50594
rect 11452 50036 11508 50542
rect 11564 50540 12292 50596
rect 12348 52050 12404 52062
rect 12348 51998 12350 52050
rect 12402 51998 12404 52050
rect 11564 50482 11620 50540
rect 11564 50430 11566 50482
rect 11618 50430 11620 50482
rect 11564 50418 11620 50430
rect 11452 49970 11508 49980
rect 11900 50036 11956 50046
rect 11228 49812 11284 49822
rect 11228 49718 11284 49756
rect 11900 49812 11956 49980
rect 11900 49746 11956 49756
rect 11116 49532 11844 49588
rect 10780 49522 10836 49532
rect 11418 49420 11682 49430
rect 10780 49364 10836 49374
rect 11474 49364 11522 49420
rect 11578 49364 11626 49420
rect 10836 49308 10948 49364
rect 11418 49354 11682 49364
rect 10780 49298 10836 49308
rect 10892 49138 10948 49308
rect 11340 49252 11396 49262
rect 11788 49252 11844 49532
rect 10892 49086 10894 49138
rect 10946 49086 10948 49138
rect 10892 49074 10948 49086
rect 11116 49140 11172 49150
rect 11004 48916 11060 48926
rect 10892 48244 10948 48254
rect 10780 48132 10836 48142
rect 10668 48076 10780 48132
rect 10780 48038 10836 48076
rect 10108 47842 10164 47852
rect 10332 47796 10388 47806
rect 10220 47684 10276 47694
rect 10220 47458 10276 47628
rect 10332 47570 10388 47740
rect 10556 47796 10612 47806
rect 10556 47684 10612 47740
rect 10556 47628 10724 47684
rect 10332 47518 10334 47570
rect 10386 47518 10388 47570
rect 10332 47506 10388 47518
rect 10220 47406 10222 47458
rect 10274 47406 10276 47458
rect 10220 47394 10276 47406
rect 10556 47460 10612 47470
rect 10668 47460 10724 47628
rect 10556 47458 10724 47460
rect 10556 47406 10558 47458
rect 10610 47406 10724 47458
rect 10556 47404 10724 47406
rect 10556 47394 10612 47404
rect 9996 47294 9998 47346
rect 10050 47294 10052 47346
rect 9996 47282 10052 47294
rect 10108 47348 10164 47358
rect 9772 47180 9940 47236
rect 9772 47068 9828 47180
rect 9996 47068 10052 47078
rect 9772 47012 9940 47068
rect 9436 46062 9438 46114
rect 9490 46062 9492 46114
rect 9436 46050 9492 46062
rect 9436 45892 9492 45902
rect 9884 45892 9940 47012
rect 9996 46898 10052 47012
rect 9996 46846 9998 46898
rect 10050 46846 10052 46898
rect 9996 46834 10052 46846
rect 10108 46564 10164 47292
rect 10444 47348 10500 47358
rect 10444 47254 10500 47292
rect 10780 47348 10836 47358
rect 10668 47236 10724 47246
rect 10332 47124 10388 47134
rect 10332 46900 10388 47068
rect 10108 46498 10164 46508
rect 10220 46844 10388 46900
rect 10556 47124 10612 47134
rect 9436 45798 9492 45836
rect 9772 45836 9940 45892
rect 9996 46114 10052 46126
rect 9996 46062 9998 46114
rect 10050 46062 10052 46114
rect 9436 45556 9492 45566
rect 9436 44996 9492 45500
rect 9772 45444 9828 45836
rect 9884 45668 9940 45678
rect 9996 45668 10052 46062
rect 9884 45666 10052 45668
rect 9884 45614 9886 45666
rect 9938 45614 10052 45666
rect 9884 45612 10052 45614
rect 9884 45602 9940 45612
rect 9996 45444 10052 45612
rect 10220 45444 10276 46844
rect 10332 46674 10388 46686
rect 10332 46622 10334 46674
rect 10386 46622 10388 46674
rect 10332 46564 10388 46622
rect 10332 46498 10388 46508
rect 10332 46114 10388 46126
rect 10332 46062 10334 46114
rect 10386 46062 10388 46114
rect 10332 46002 10388 46062
rect 10332 45950 10334 46002
rect 10386 45950 10388 46002
rect 10332 45938 10388 45950
rect 10444 45668 10500 45678
rect 9996 45388 10164 45444
rect 10220 45388 10388 45444
rect 9772 45378 9828 45388
rect 10108 45332 10164 45388
rect 10108 45276 10276 45332
rect 9548 45220 9604 45230
rect 9548 45126 9604 45164
rect 9772 45106 9828 45118
rect 9772 45054 9774 45106
rect 9826 45054 9828 45106
rect 9436 44940 9604 44996
rect 8988 38612 9156 38668
rect 9212 44492 9380 44548
rect 9436 44548 9492 44558
rect 8988 37940 9044 38612
rect 9100 38164 9156 38174
rect 9100 38070 9156 38108
rect 8988 37884 9156 37940
rect 8876 36482 9044 36484
rect 8876 36430 8878 36482
rect 8930 36430 9044 36482
rect 8876 36428 9044 36430
rect 8876 36418 8932 36428
rect 8652 36260 8708 36270
rect 8652 36258 8820 36260
rect 8652 36206 8654 36258
rect 8706 36206 8820 36258
rect 8652 36204 8820 36206
rect 8652 36194 8708 36204
rect 7868 35868 8148 35924
rect 7868 35700 7924 35710
rect 7756 34804 7812 34814
rect 7756 34710 7812 34748
rect 7868 34580 7924 35644
rect 8092 34914 8148 35868
rect 8428 35868 8540 35924
rect 8092 34862 8094 34914
rect 8146 34862 8148 34914
rect 8092 34850 8148 34862
rect 8316 34916 8372 34926
rect 8428 34916 8484 35868
rect 8540 35830 8596 35868
rect 8764 35812 8820 36204
rect 8652 35028 8708 35038
rect 8652 34934 8708 34972
rect 8316 34914 8484 34916
rect 8316 34862 8318 34914
rect 8370 34862 8484 34914
rect 8316 34860 8484 34862
rect 8316 34850 8372 34860
rect 7756 34524 7924 34580
rect 8016 34524 8280 34534
rect 7756 33908 7812 34524
rect 8072 34468 8120 34524
rect 8176 34468 8224 34524
rect 8016 34458 8280 34468
rect 8428 34356 8484 34860
rect 8652 34804 8708 34814
rect 8652 34710 8708 34748
rect 8428 34290 8484 34300
rect 8540 34690 8596 34702
rect 8540 34638 8542 34690
rect 8594 34638 8596 34690
rect 7868 34132 7924 34142
rect 7868 34038 7924 34076
rect 8092 34132 8148 34142
rect 8092 34038 8148 34076
rect 8316 34130 8372 34142
rect 8316 34078 8318 34130
rect 8370 34078 8372 34130
rect 8204 34018 8260 34030
rect 8204 33966 8206 34018
rect 8258 33966 8260 34018
rect 7756 33852 7924 33908
rect 7644 31266 7700 31276
rect 7756 33684 7812 33694
rect 7644 31108 7700 31118
rect 7532 30996 7588 31006
rect 7532 30902 7588 30940
rect 7532 30772 7588 30782
rect 7644 30772 7700 31052
rect 7532 30770 7700 30772
rect 7532 30718 7534 30770
rect 7586 30718 7700 30770
rect 7532 30716 7700 30718
rect 7532 30706 7588 30716
rect 7420 30492 7588 30548
rect 6860 30322 7252 30324
rect 6860 30270 6862 30322
rect 6914 30270 7252 30322
rect 6860 30268 7252 30270
rect 6860 30258 6916 30268
rect 6860 29876 6916 29886
rect 6860 29538 6916 29820
rect 6860 29486 6862 29538
rect 6914 29486 6916 29538
rect 6860 29474 6916 29486
rect 7084 29540 7140 30268
rect 7196 30210 7252 30268
rect 7196 30158 7198 30210
rect 7250 30158 7252 30210
rect 7196 30146 7252 30158
rect 7308 30212 7364 30268
rect 7420 30212 7476 30222
rect 7308 30210 7476 30212
rect 7308 30158 7422 30210
rect 7474 30158 7476 30210
rect 7308 30156 7476 30158
rect 7420 30146 7476 30156
rect 7308 29986 7364 29998
rect 7308 29934 7310 29986
rect 7362 29934 7364 29986
rect 7196 29876 7252 29886
rect 7308 29876 7364 29934
rect 7252 29820 7364 29876
rect 7196 29810 7252 29820
rect 6860 28756 6916 28766
rect 6748 28700 6860 28756
rect 7084 28756 7140 29484
rect 7308 28756 7364 28766
rect 7084 28754 7364 28756
rect 7084 28702 7310 28754
rect 7362 28702 7364 28754
rect 7084 28700 7364 28702
rect 6860 28662 6916 28700
rect 7308 28690 7364 28700
rect 7532 28532 7588 30492
rect 7644 30324 7700 30334
rect 7644 30230 7700 30268
rect 7756 30100 7812 33628
rect 7868 30884 7924 33852
rect 8204 33460 8260 33966
rect 8316 34020 8372 34078
rect 8316 33954 8372 33964
rect 8428 34130 8484 34142
rect 8428 34078 8430 34130
rect 8482 34078 8484 34130
rect 8428 33908 8484 34078
rect 8428 33842 8484 33852
rect 8540 33684 8596 34638
rect 8540 33618 8596 33628
rect 8652 33796 8708 33806
rect 8204 33394 8260 33404
rect 8540 33460 8596 33470
rect 8652 33460 8708 33740
rect 8540 33458 8708 33460
rect 8540 33406 8542 33458
rect 8594 33406 8708 33458
rect 8540 33404 8708 33406
rect 8540 33394 8596 33404
rect 8016 32956 8280 32966
rect 8072 32900 8120 32956
rect 8176 32900 8224 32956
rect 8016 32890 8280 32900
rect 8764 32788 8820 35756
rect 8988 35922 9044 36428
rect 8988 35870 8990 35922
rect 9042 35870 9044 35922
rect 8988 34804 9044 35870
rect 8988 34354 9044 34748
rect 9100 34468 9156 37884
rect 9100 34402 9156 34412
rect 8988 34302 8990 34354
rect 9042 34302 9044 34354
rect 8988 33908 9044 34302
rect 8988 33570 9044 33852
rect 8988 33518 8990 33570
rect 9042 33518 9044 33570
rect 8988 33506 9044 33518
rect 9100 34132 9156 34142
rect 9100 33458 9156 34076
rect 9100 33406 9102 33458
rect 9154 33406 9156 33458
rect 9100 33394 9156 33406
rect 8764 32722 8820 32732
rect 8764 32452 8820 32490
rect 8764 32386 8820 32396
rect 8764 32228 8820 32238
rect 8016 31388 8280 31398
rect 8072 31332 8120 31388
rect 8176 31332 8224 31388
rect 8016 31322 8280 31332
rect 7980 31108 8036 31118
rect 8204 31108 8260 31118
rect 8036 31106 8260 31108
rect 8036 31054 8206 31106
rect 8258 31054 8260 31106
rect 8036 31052 8260 31054
rect 7980 31042 8036 31052
rect 8204 31042 8260 31052
rect 8428 30996 8484 31006
rect 8428 30902 8484 30940
rect 8092 30884 8148 30894
rect 7868 30828 8092 30884
rect 7868 30548 7924 30558
rect 7868 30210 7924 30492
rect 8092 30436 8148 30828
rect 8092 30324 8148 30380
rect 8428 30436 8484 30446
rect 8316 30324 8372 30334
rect 8092 30322 8372 30324
rect 8092 30270 8318 30322
rect 8370 30270 8372 30322
rect 8092 30268 8372 30270
rect 7868 30158 7870 30210
rect 7922 30158 7924 30210
rect 7868 30146 7924 30158
rect 7196 28476 7588 28532
rect 7644 30044 7812 30100
rect 6636 28084 6692 28094
rect 6412 28082 6692 28084
rect 6412 28030 6638 28082
rect 6690 28030 6692 28082
rect 6412 28028 6692 28030
rect 6412 27188 6468 28028
rect 6636 28018 6692 28028
rect 6412 27094 6468 27132
rect 6860 27300 6916 27310
rect 6860 27186 6916 27244
rect 6860 27134 6862 27186
rect 6914 27134 6916 27186
rect 6860 27122 6916 27134
rect 6748 27076 6804 27086
rect 6748 26982 6804 27020
rect 7196 26908 7252 28476
rect 6188 26338 6244 26348
rect 6300 26850 6356 26862
rect 6300 26798 6302 26850
rect 6354 26798 6356 26850
rect 6188 25508 6244 25518
rect 6300 25508 6356 26798
rect 7084 26852 7252 26908
rect 7308 27188 7364 27198
rect 6188 25506 6356 25508
rect 6188 25454 6190 25506
rect 6242 25454 6356 25506
rect 6188 25452 6356 25454
rect 6412 25620 6468 25630
rect 6412 25506 6468 25564
rect 6412 25454 6414 25506
rect 6466 25454 6468 25506
rect 6188 25442 6244 25452
rect 6412 25442 6468 25454
rect 6636 25508 6692 25518
rect 6076 23938 6132 24892
rect 6076 23886 6078 23938
rect 6130 23886 6132 23938
rect 6076 23874 6132 23886
rect 5852 23492 6020 23548
rect 5516 23042 5572 23054
rect 5516 22990 5518 23042
rect 5570 22990 5572 23042
rect 5516 22596 5572 22990
rect 5516 22530 5572 22540
rect 5852 21474 5908 21486
rect 5852 21422 5854 21474
rect 5906 21422 5908 21474
rect 5852 21026 5908 21422
rect 5852 20974 5854 21026
rect 5906 20974 5908 21026
rect 5852 20962 5908 20974
rect 5964 20692 6020 23492
rect 6636 23268 6692 25452
rect 6860 23826 6916 23838
rect 6860 23774 6862 23826
rect 6914 23774 6916 23826
rect 6860 23380 6916 23774
rect 6972 23380 7028 23390
rect 6860 23378 7028 23380
rect 6860 23326 6974 23378
rect 7026 23326 7028 23378
rect 6860 23324 7028 23326
rect 6972 23314 7028 23324
rect 6636 23174 6692 23212
rect 6188 23044 6244 23054
rect 6300 23044 6356 23054
rect 6188 23042 6300 23044
rect 6188 22990 6190 23042
rect 6242 22990 6300 23042
rect 6188 22988 6300 22990
rect 6188 22978 6244 22988
rect 6188 20692 6244 20702
rect 5964 20636 6188 20692
rect 6188 20598 6244 20636
rect 5740 20578 5796 20590
rect 5740 20526 5742 20578
rect 5794 20526 5796 20578
rect 5740 20356 5796 20526
rect 6300 20356 6356 22988
rect 6860 21364 6916 21374
rect 6412 21026 6468 21038
rect 6412 20974 6414 21026
rect 6466 20974 6468 21026
rect 6412 20580 6468 20974
rect 6860 21026 6916 21308
rect 6860 20974 6862 21026
rect 6914 20974 6916 21026
rect 6860 20962 6916 20974
rect 7084 20916 7140 26852
rect 7196 25506 7252 25518
rect 7196 25454 7198 25506
rect 7250 25454 7252 25506
rect 7196 25284 7252 25454
rect 7196 25218 7252 25228
rect 7308 24610 7364 27132
rect 7644 26908 7700 30044
rect 8316 29988 8372 30268
rect 8428 30322 8484 30380
rect 8428 30270 8430 30322
rect 8482 30270 8484 30322
rect 8428 30258 8484 30270
rect 8316 29922 8372 29932
rect 8540 29986 8596 29998
rect 8540 29934 8542 29986
rect 8594 29934 8596 29986
rect 8540 29876 8596 29934
rect 8016 29820 8280 29830
rect 8072 29764 8120 29820
rect 8176 29764 8224 29820
rect 8540 29810 8596 29820
rect 8016 29754 8280 29764
rect 8540 29092 8596 29102
rect 8428 29036 8540 29092
rect 7756 28756 7812 28766
rect 7756 27188 7812 28700
rect 8016 28252 8280 28262
rect 8072 28196 8120 28252
rect 8176 28196 8224 28252
rect 8016 28186 8280 28196
rect 7756 27094 7812 27132
rect 8092 27860 8148 27870
rect 8092 27018 8148 27804
rect 8092 26966 8094 27018
rect 8146 26966 8148 27018
rect 8316 27188 8372 27198
rect 8316 27074 8372 27132
rect 8316 27022 8318 27074
rect 8370 27022 8372 27074
rect 8316 27010 8372 27022
rect 8092 26954 8148 26966
rect 7308 24558 7310 24610
rect 7362 24558 7364 24610
rect 7308 24546 7364 24558
rect 7420 26852 7700 26908
rect 8204 26852 8260 26862
rect 7196 23154 7252 23166
rect 7196 23102 7198 23154
rect 7250 23102 7252 23154
rect 7196 23044 7252 23102
rect 7196 22978 7252 22988
rect 7308 22932 7364 22942
rect 7308 22838 7364 22876
rect 6972 20860 7140 20916
rect 7196 21140 7252 21150
rect 6636 20802 6692 20814
rect 6636 20750 6638 20802
rect 6690 20750 6692 20802
rect 6524 20580 6580 20590
rect 6412 20578 6580 20580
rect 6412 20526 6526 20578
rect 6578 20526 6580 20578
rect 6412 20524 6580 20526
rect 6524 20514 6580 20524
rect 6636 20356 6692 20750
rect 5740 20300 6692 20356
rect 6636 20244 6692 20300
rect 6636 20178 6692 20188
rect 5404 20132 5460 20142
rect 5404 20038 5460 20076
rect 6412 19348 6468 19358
rect 6972 19348 7028 20860
rect 7084 20692 7140 20702
rect 7084 20598 7140 20636
rect 6076 19236 6132 19246
rect 6412 19236 6468 19292
rect 6860 19292 7028 19348
rect 7196 20242 7252 21084
rect 7420 21028 7476 26852
rect 7868 26850 8260 26852
rect 7868 26798 8206 26850
rect 8258 26798 8260 26850
rect 7868 26796 8260 26798
rect 7868 25618 7924 26796
rect 8204 26786 8260 26796
rect 8016 26684 8280 26694
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8016 26618 8280 26628
rect 7868 25566 7870 25618
rect 7922 25566 7924 25618
rect 7868 25554 7924 25566
rect 8016 25116 8280 25126
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8016 25050 8280 25060
rect 7756 24948 7812 24958
rect 7756 24854 7812 24892
rect 8016 23548 8280 23558
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8016 23482 8280 23492
rect 7532 23268 7588 23278
rect 7532 23174 7588 23212
rect 7756 23156 7812 23166
rect 7756 23154 7924 23156
rect 7756 23102 7758 23154
rect 7810 23102 7924 23154
rect 7756 23100 7924 23102
rect 7756 23090 7812 23100
rect 7420 20962 7476 20972
rect 7868 22148 7924 23100
rect 8316 23042 8372 23054
rect 8316 22990 8318 23042
rect 8370 22990 8372 23042
rect 8204 22930 8260 22942
rect 8204 22878 8206 22930
rect 8258 22878 8260 22930
rect 8204 22596 8260 22878
rect 8316 22932 8372 22990
rect 8316 22866 8372 22876
rect 8204 22530 8260 22540
rect 7980 22148 8036 22158
rect 7868 22146 8036 22148
rect 7868 22094 7982 22146
rect 8034 22094 8036 22146
rect 7868 22092 8036 22094
rect 7308 20692 7364 20702
rect 7308 20598 7364 20636
rect 7756 20692 7812 20702
rect 7868 20692 7924 22092
rect 7980 22082 8036 22092
rect 8016 21980 8280 21990
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8016 21914 8280 21924
rect 8428 21924 8484 29036
rect 8540 29026 8596 29036
rect 8540 27412 8596 27422
rect 8540 27298 8596 27356
rect 8540 27246 8542 27298
rect 8594 27246 8596 27298
rect 8540 27234 8596 27246
rect 8764 26852 8820 32172
rect 9100 31890 9156 31902
rect 9100 31838 9102 31890
rect 9154 31838 9156 31890
rect 9100 30996 9156 31838
rect 9100 30930 9156 30940
rect 8876 30884 8932 30894
rect 8876 30790 8932 30828
rect 9212 30436 9268 44492
rect 9324 42980 9380 42990
rect 9324 42866 9380 42924
rect 9324 42814 9326 42866
rect 9378 42814 9380 42866
rect 9324 42802 9380 42814
rect 9100 30380 9268 30436
rect 9324 37044 9380 37054
rect 9324 36594 9380 36988
rect 9324 36542 9326 36594
rect 9378 36542 9380 36594
rect 8988 30100 9044 30110
rect 8988 29876 9044 30044
rect 8988 29314 9044 29820
rect 8988 29262 8990 29314
rect 9042 29262 9044 29314
rect 8988 29250 9044 29262
rect 8988 27860 9044 27870
rect 8988 27766 9044 27804
rect 8876 27748 8932 27758
rect 8876 27074 8932 27692
rect 8876 27022 8878 27074
rect 8930 27022 8932 27074
rect 8876 27010 8932 27022
rect 9100 26908 9156 30380
rect 9324 30324 9380 36542
rect 9212 30268 9380 30324
rect 9212 27636 9268 30268
rect 9324 30100 9380 30110
rect 9324 30006 9380 30044
rect 9212 27570 9268 27580
rect 9212 27300 9268 27310
rect 9268 27244 9380 27300
rect 9212 27234 9268 27244
rect 9100 26852 9268 26908
rect 8652 26796 8820 26852
rect 8652 23492 8708 26796
rect 8988 25284 9044 25294
rect 8988 24948 9044 25228
rect 8652 23426 8708 23436
rect 8764 24946 9044 24948
rect 8764 24894 8990 24946
rect 9042 24894 9044 24946
rect 8764 24892 9044 24894
rect 8652 23268 8708 23278
rect 8540 23266 8708 23268
rect 8540 23214 8654 23266
rect 8706 23214 8708 23266
rect 8540 23212 8708 23214
rect 8540 23154 8596 23212
rect 8652 23202 8708 23212
rect 8540 23102 8542 23154
rect 8594 23102 8596 23154
rect 8540 23090 8596 23102
rect 8652 22596 8708 22606
rect 8428 21868 8596 21924
rect 7980 21700 8036 21710
rect 7980 21474 8036 21644
rect 8428 21700 8484 21710
rect 8428 21606 8484 21644
rect 7980 21422 7982 21474
rect 8034 21422 8036 21474
rect 7980 21410 8036 21422
rect 8316 21364 8372 21374
rect 8316 21270 8372 21308
rect 8204 20916 8260 20926
rect 8204 20822 8260 20860
rect 7812 20636 7924 20692
rect 7756 20598 7812 20636
rect 8016 20412 8280 20422
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8016 20346 8280 20356
rect 7196 20190 7198 20242
rect 7250 20190 7252 20242
rect 7196 19348 7252 20190
rect 8316 19908 8372 19918
rect 6076 19142 6132 19180
rect 6188 19234 6468 19236
rect 6188 19182 6414 19234
rect 6466 19182 6468 19234
rect 6188 19180 6468 19182
rect 5964 19012 6020 19022
rect 5964 18562 6020 18956
rect 5964 18510 5966 18562
rect 6018 18510 6020 18562
rect 5964 18498 6020 18510
rect 5740 17780 5796 17790
rect 5740 17666 5796 17724
rect 5740 17614 5742 17666
rect 5794 17614 5796 17666
rect 5740 17602 5796 17614
rect 6076 16884 6132 16922
rect 6188 16884 6244 19180
rect 6412 19170 6468 19180
rect 6636 19236 6692 19246
rect 6524 19012 6580 19022
rect 6524 18918 6580 18956
rect 6636 18564 6692 19180
rect 6300 18508 6636 18564
rect 6300 17332 6356 18508
rect 6636 18498 6692 18508
rect 6636 17780 6692 17790
rect 6412 17556 6468 17566
rect 6412 17554 6580 17556
rect 6412 17502 6414 17554
rect 6466 17502 6580 17554
rect 6412 17500 6580 17502
rect 6412 17490 6468 17500
rect 6300 17276 6468 17332
rect 6300 16884 6356 16894
rect 6132 16882 6356 16884
rect 6132 16830 6302 16882
rect 6354 16830 6356 16882
rect 6132 16828 6356 16830
rect 6076 16818 6132 16828
rect 6300 16818 6356 16828
rect 5292 16718 5294 16770
rect 5346 16718 5348 16770
rect 5292 16706 5348 16718
rect 5628 16772 5684 16782
rect 5628 16678 5684 16716
rect 6076 16658 6132 16670
rect 6076 16606 6078 16658
rect 6130 16606 6132 16658
rect 6076 15538 6132 16606
rect 6076 15486 6078 15538
rect 6130 15486 6132 15538
rect 6076 15428 6132 15486
rect 6076 15362 6132 15372
rect 6188 15316 6244 15326
rect 5628 15204 5684 15242
rect 5628 15138 5684 15148
rect 5068 14530 5124 14588
rect 5068 14478 5070 14530
rect 5122 14478 5124 14530
rect 4508 13748 4564 13758
rect 4396 13746 4564 13748
rect 4396 13694 4510 13746
rect 4562 13694 4564 13746
rect 4396 13692 4564 13694
rect 4396 12180 4452 13692
rect 4508 13682 4564 13692
rect 4956 13636 5012 13646
rect 4614 13356 4878 13366
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4614 13290 4878 13300
rect 4620 13076 4676 13086
rect 4956 13076 5012 13580
rect 4620 13074 5012 13076
rect 4620 13022 4622 13074
rect 4674 13022 5012 13074
rect 4620 13020 5012 13022
rect 5068 13076 5124 14478
rect 5516 14644 5572 14654
rect 5516 14530 5572 14588
rect 5516 14478 5518 14530
rect 5570 14478 5572 14530
rect 5516 14466 5572 14478
rect 6188 14530 6244 15260
rect 6188 14478 6190 14530
rect 6242 14478 6244 14530
rect 6188 14466 6244 14478
rect 5964 14420 6020 14430
rect 6020 14364 6132 14420
rect 5964 14326 6020 14364
rect 5740 14308 5796 14318
rect 5628 14306 5796 14308
rect 5628 14254 5742 14306
rect 5794 14254 5796 14306
rect 5628 14252 5796 14254
rect 5628 13972 5684 14252
rect 5740 14242 5796 14252
rect 5852 14308 5908 14318
rect 5292 13916 5684 13972
rect 5292 13858 5348 13916
rect 5292 13806 5294 13858
rect 5346 13806 5348 13858
rect 5292 13794 5348 13806
rect 5516 13076 5572 13086
rect 5068 13074 5516 13076
rect 5068 13022 5070 13074
rect 5122 13022 5516 13074
rect 5068 13020 5516 13022
rect 4620 13010 4676 13020
rect 5068 13010 5124 13020
rect 5516 12962 5572 13020
rect 5516 12910 5518 12962
rect 5570 12910 5572 12962
rect 5516 12898 5572 12910
rect 5740 12738 5796 12750
rect 5740 12686 5742 12738
rect 5794 12686 5796 12738
rect 5740 12404 5796 12686
rect 5180 12348 5796 12404
rect 5180 12290 5236 12348
rect 5180 12238 5182 12290
rect 5234 12238 5236 12290
rect 5180 12226 5236 12238
rect 4508 12180 4564 12190
rect 4396 12178 4564 12180
rect 4396 12126 4510 12178
rect 4562 12126 4564 12178
rect 4396 12124 4564 12126
rect 4284 12114 4340 12124
rect 4508 11956 4564 12124
rect 4508 11900 5012 11956
rect 4956 11844 5012 11900
rect 4614 11788 4878 11798
rect 4956 11788 5348 11844
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4614 11722 4878 11732
rect 4508 11396 4564 11406
rect 4284 11284 4340 11294
rect 4060 11282 4340 11284
rect 4060 11230 4286 11282
rect 4338 11230 4340 11282
rect 4060 11228 4340 11230
rect 4284 11172 4340 11228
rect 4284 11106 4340 11116
rect 4396 11170 4452 11182
rect 4396 11118 4398 11170
rect 4450 11118 4452 11170
rect 4396 10948 4452 11118
rect 4284 10892 4452 10948
rect 4508 11170 4564 11340
rect 4956 11284 5012 11294
rect 4956 11190 5012 11228
rect 5068 11282 5124 11294
rect 5068 11230 5070 11282
rect 5122 11230 5124 11282
rect 4508 11118 4510 11170
rect 4562 11118 4564 11170
rect 3388 6750 3390 6802
rect 3442 6750 3444 6802
rect 3388 6738 3444 6750
rect 3500 7420 3892 7476
rect 3948 9156 4004 9166
rect 3388 6580 3444 6590
rect 3276 6524 3388 6580
rect 3388 6514 3444 6524
rect 2044 6356 2100 6366
rect 1708 5122 1764 5134
rect 1708 5070 1710 5122
rect 1762 5070 1764 5122
rect 1708 4788 1764 5070
rect 2044 5010 2100 6300
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 2492 5122 2548 5134
rect 2492 5070 2494 5122
rect 2546 5070 2548 5122
rect 1708 4722 1764 4732
rect 2492 4788 2548 5070
rect 2492 4722 2548 4732
rect 3500 3388 3556 7420
rect 3836 6468 3892 6478
rect 3948 6468 4004 9100
rect 4284 7252 4340 10892
rect 4508 10836 4564 11118
rect 4396 10780 4564 10836
rect 5068 10836 5124 11230
rect 4396 9042 4452 10780
rect 4614 10220 4878 10230
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4614 10154 4878 10164
rect 5068 10164 5124 10780
rect 5068 10098 5124 10108
rect 5180 11284 5236 11294
rect 4844 10052 4900 10062
rect 4620 9996 4844 10052
rect 4508 9940 4564 9950
rect 4508 9154 4564 9884
rect 4620 9938 4676 9996
rect 4844 9986 4900 9996
rect 4620 9886 4622 9938
rect 4674 9886 4676 9938
rect 4620 9874 4676 9886
rect 5068 9604 5124 9614
rect 5180 9604 5236 11228
rect 5292 11172 5348 11788
rect 5852 11396 5908 14252
rect 5964 13524 6020 13534
rect 5964 12850 6020 13468
rect 5964 12798 5966 12850
rect 6018 12798 6020 12850
rect 5964 12404 6020 12798
rect 5964 12338 6020 12348
rect 5852 11330 5908 11340
rect 6076 11396 6132 14364
rect 6188 12852 6244 12862
rect 6188 12758 6244 12796
rect 6412 11732 6468 17276
rect 6524 17106 6580 17500
rect 6524 17054 6526 17106
rect 6578 17054 6580 17106
rect 6524 17042 6580 17054
rect 6524 15540 6580 15550
rect 6524 15446 6580 15484
rect 6412 11666 6468 11676
rect 6636 14530 6692 17724
rect 6748 16882 6804 16894
rect 6748 16830 6750 16882
rect 6802 16830 6804 16882
rect 6748 16772 6804 16830
rect 6748 16706 6804 16716
rect 6860 15540 6916 19292
rect 7196 19282 7252 19292
rect 8204 19906 8372 19908
rect 8204 19854 8318 19906
rect 8370 19854 8372 19906
rect 8204 19852 8372 19854
rect 7756 19236 7812 19246
rect 8204 19236 8260 19852
rect 8316 19842 8372 19852
rect 8540 19236 8596 21868
rect 8652 21698 8708 22540
rect 8652 21646 8654 21698
rect 8706 21646 8708 21698
rect 8652 21634 8708 21646
rect 8652 20804 8708 20814
rect 8652 20710 8708 20748
rect 8652 19348 8708 19358
rect 8764 19348 8820 24892
rect 8988 24882 9044 24892
rect 9100 24724 9156 24734
rect 8876 24668 9100 24724
rect 8876 24052 8932 24668
rect 9100 24658 9156 24668
rect 8988 24076 9044 24088
rect 8988 24052 8990 24076
rect 8876 24024 8990 24052
rect 9042 24024 9044 24076
rect 8876 23996 9044 24024
rect 8876 23266 8932 23996
rect 9212 23940 9268 26852
rect 8988 23884 9268 23940
rect 8988 23492 9044 23884
rect 9212 23716 9268 23726
rect 9324 23716 9380 27244
rect 9436 23828 9492 44492
rect 9548 43764 9604 44940
rect 9660 44772 9716 44782
rect 9660 44434 9716 44716
rect 9660 44382 9662 44434
rect 9714 44382 9716 44434
rect 9660 44370 9716 44382
rect 9772 44212 9828 45054
rect 9996 45106 10052 45118
rect 9996 45054 9998 45106
rect 10050 45054 10052 45106
rect 9772 44146 9828 44156
rect 9884 44994 9940 45006
rect 9884 44942 9886 44994
rect 9938 44942 9940 44994
rect 9548 43708 9828 43764
rect 9660 43428 9716 43438
rect 9660 43334 9716 43372
rect 9660 43204 9716 43214
rect 9660 42980 9716 43148
rect 9660 42754 9716 42924
rect 9660 42702 9662 42754
rect 9714 42702 9716 42754
rect 9660 42690 9716 42702
rect 9548 42308 9604 42318
rect 9548 41748 9604 42252
rect 9548 40292 9604 41692
rect 9548 40226 9604 40236
rect 9660 40290 9716 40302
rect 9660 40238 9662 40290
rect 9714 40238 9716 40290
rect 9548 40068 9604 40078
rect 9548 39394 9604 40012
rect 9660 39842 9716 40238
rect 9660 39790 9662 39842
rect 9714 39790 9716 39842
rect 9660 39778 9716 39790
rect 9548 39342 9550 39394
rect 9602 39342 9604 39394
rect 9548 39172 9604 39342
rect 9548 39106 9604 39116
rect 9772 38668 9828 43708
rect 9884 43652 9940 44942
rect 9996 44546 10052 45054
rect 10108 45106 10164 45118
rect 10108 45054 10110 45106
rect 10162 45054 10164 45106
rect 10108 44996 10164 45054
rect 10108 44930 10164 44940
rect 9996 44494 9998 44546
rect 10050 44494 10052 44546
rect 9996 44482 10052 44494
rect 10108 44436 10164 44446
rect 10220 44436 10276 45276
rect 10108 44434 10276 44436
rect 10108 44382 10110 44434
rect 10162 44382 10276 44434
rect 10108 44380 10276 44382
rect 10108 44370 10164 44380
rect 10108 43652 10164 43662
rect 9884 43650 10164 43652
rect 9884 43598 10110 43650
rect 10162 43598 10164 43650
rect 9884 43596 10164 43598
rect 10108 43586 10164 43596
rect 9996 43426 10052 43438
rect 9996 43374 9998 43426
rect 10050 43374 10052 43426
rect 9996 43092 10052 43374
rect 10332 43092 10388 45388
rect 10444 44322 10500 45612
rect 10444 44270 10446 44322
rect 10498 44270 10500 44322
rect 10444 44258 10500 44270
rect 10556 43876 10612 47068
rect 10668 44548 10724 47180
rect 10780 46114 10836 47292
rect 10892 47012 10948 48188
rect 11004 47682 11060 48860
rect 11004 47630 11006 47682
rect 11058 47630 11060 47682
rect 11004 47618 11060 47630
rect 11116 47572 11172 49084
rect 11340 49138 11396 49196
rect 11340 49086 11342 49138
rect 11394 49086 11396 49138
rect 11340 49074 11396 49086
rect 11676 49196 11844 49252
rect 11900 49586 11956 49598
rect 11900 49534 11902 49586
rect 11954 49534 11956 49586
rect 11228 48468 11284 48478
rect 11284 48412 11396 48468
rect 11228 48402 11284 48412
rect 11340 48354 11396 48412
rect 11340 48302 11342 48354
rect 11394 48302 11396 48354
rect 11340 48290 11396 48302
rect 11676 48020 11732 49196
rect 11788 49028 11844 49038
rect 11788 48934 11844 48972
rect 11788 48692 11844 48702
rect 11788 48466 11844 48636
rect 11788 48414 11790 48466
rect 11842 48414 11844 48466
rect 11788 48402 11844 48414
rect 11788 48020 11844 48030
rect 11676 48018 11844 48020
rect 11676 47966 11790 48018
rect 11842 47966 11844 48018
rect 11676 47964 11844 47966
rect 11788 47954 11844 47964
rect 11418 47852 11682 47862
rect 11474 47796 11522 47852
rect 11578 47796 11626 47852
rect 11418 47786 11682 47796
rect 11452 47684 11508 47694
rect 11228 47572 11284 47582
rect 11116 47570 11284 47572
rect 11116 47518 11230 47570
rect 11282 47518 11284 47570
rect 11116 47516 11284 47518
rect 11228 47506 11284 47516
rect 11340 47348 11396 47358
rect 10892 46946 10948 46956
rect 11228 47292 11340 47348
rect 10780 46062 10782 46114
rect 10834 46062 10836 46114
rect 10780 46002 10836 46062
rect 10780 45950 10782 46002
rect 10834 45950 10836 46002
rect 10780 45938 10836 45950
rect 10892 46788 10948 46798
rect 10668 44482 10724 44492
rect 10780 44884 10836 44894
rect 10780 44436 10836 44828
rect 10892 44772 10948 46732
rect 11116 46562 11172 46574
rect 11116 46510 11118 46562
rect 11170 46510 11172 46562
rect 11116 46004 11172 46510
rect 11228 46116 11284 47292
rect 11340 47282 11396 47292
rect 11452 46564 11508 47628
rect 11564 47682 11620 47694
rect 11564 47630 11566 47682
rect 11618 47630 11620 47682
rect 11564 47570 11620 47630
rect 11900 47572 11956 49534
rect 12012 49028 12068 50540
rect 12236 50372 12292 50382
rect 12236 49922 12292 50316
rect 12236 49870 12238 49922
rect 12290 49870 12292 49922
rect 12236 49140 12292 49870
rect 12348 49812 12404 51998
rect 12460 50932 12516 54124
rect 12908 54068 12964 55022
rect 12684 54012 12964 54068
rect 13132 54514 13188 54526
rect 13132 54462 13134 54514
rect 13186 54462 13188 54514
rect 13132 54404 13188 54462
rect 12572 53730 12628 53742
rect 12572 53678 12574 53730
rect 12626 53678 12628 53730
rect 12572 53284 12628 53678
rect 12684 53396 12740 54012
rect 12908 53844 12964 53854
rect 12908 53750 12964 53788
rect 13132 53732 13188 54348
rect 13132 53666 13188 53676
rect 13244 54402 13300 56140
rect 13468 57148 13748 57204
rect 13916 57540 13972 57550
rect 14140 57540 14196 58772
rect 13916 57538 14196 57540
rect 13916 57486 13918 57538
rect 13970 57486 14196 57538
rect 13916 57484 14196 57486
rect 13468 56866 13524 57148
rect 13916 57092 13972 57484
rect 14252 57428 14308 58940
rect 14364 58324 14420 59948
rect 14588 60002 14644 60014
rect 14588 59950 14590 60002
rect 14642 59950 14644 60002
rect 14476 59330 14532 59342
rect 14476 59278 14478 59330
rect 14530 59278 14532 59330
rect 14476 58884 14532 59278
rect 14476 58818 14532 58828
rect 14364 58258 14420 58268
rect 14476 58660 14532 58670
rect 14476 58210 14532 58604
rect 14588 58658 14644 59950
rect 14812 59890 14868 60956
rect 14924 60898 14980 60910
rect 14924 60846 14926 60898
rect 14978 60846 14980 60898
rect 14924 60564 14980 60846
rect 15260 60564 15316 60574
rect 14980 60508 15204 60564
rect 14924 60498 14980 60508
rect 14812 59838 14814 59890
rect 14866 59838 14868 59890
rect 14812 59826 14868 59838
rect 14820 59612 15084 59622
rect 14876 59556 14924 59612
rect 14980 59556 15028 59612
rect 14820 59546 15084 59556
rect 14812 59444 14868 59454
rect 14588 58606 14590 58658
rect 14642 58606 14644 58658
rect 14588 58594 14644 58606
rect 14700 59332 14756 59342
rect 14476 58158 14478 58210
rect 14530 58158 14532 58210
rect 13916 57026 13972 57036
rect 14028 57372 14308 57428
rect 14364 58100 14420 58110
rect 13580 56980 13636 56990
rect 13580 56886 13636 56924
rect 13804 56980 13860 56990
rect 13468 56814 13470 56866
rect 13522 56814 13524 56866
rect 13468 55412 13524 56814
rect 13692 56642 13748 56654
rect 13692 56590 13694 56642
rect 13746 56590 13748 56642
rect 13692 56532 13748 56590
rect 13692 56466 13748 56476
rect 13580 56194 13636 56206
rect 13580 56142 13582 56194
rect 13634 56142 13636 56194
rect 13580 55522 13636 56142
rect 13692 56084 13748 56094
rect 13692 55990 13748 56028
rect 13580 55470 13582 55522
rect 13634 55470 13636 55522
rect 13580 55458 13636 55470
rect 13468 55346 13524 55356
rect 13244 54350 13246 54402
rect 13298 54350 13300 54402
rect 12684 53330 12740 53340
rect 12796 53506 12852 53518
rect 13244 53508 13300 54350
rect 13580 55300 13636 55310
rect 13580 55074 13636 55244
rect 13580 55022 13582 55074
rect 13634 55022 13636 55074
rect 13580 54292 13636 55022
rect 13580 54226 13636 54236
rect 13804 53844 13860 56924
rect 13916 56420 13972 56430
rect 13916 55860 13972 56364
rect 13916 55794 13972 55804
rect 14028 55524 14084 57372
rect 14364 57316 14420 58044
rect 14364 57250 14420 57260
rect 14140 56866 14196 56878
rect 14140 56814 14142 56866
rect 14194 56814 14196 56866
rect 14140 55748 14196 56814
rect 14476 56308 14532 58158
rect 14588 58436 14644 58446
rect 14588 57538 14644 58380
rect 14588 57486 14590 57538
rect 14642 57486 14644 57538
rect 14588 57428 14644 57486
rect 14588 57362 14644 57372
rect 14588 56980 14644 56990
rect 14588 56886 14644 56924
rect 14364 56252 14532 56308
rect 14364 55860 14420 56252
rect 14476 56084 14532 56094
rect 14700 56084 14756 59276
rect 14812 59330 14868 59388
rect 14812 59278 14814 59330
rect 14866 59278 14868 59330
rect 14812 59266 14868 59278
rect 15036 59220 15092 59230
rect 14924 58658 14980 58670
rect 14924 58606 14926 58658
rect 14978 58606 14980 58658
rect 14924 58546 14980 58606
rect 15036 58660 15092 59164
rect 15036 58594 15092 58604
rect 14924 58494 14926 58546
rect 14978 58494 14980 58546
rect 14924 58212 14980 58494
rect 15148 58436 15204 60508
rect 15148 58370 15204 58380
rect 15260 58212 15316 60508
rect 15372 60340 15428 60350
rect 15372 58324 15428 60284
rect 15484 60228 15540 62860
rect 15596 62356 15652 62366
rect 15596 61796 15652 62300
rect 16044 62356 16100 66780
rect 16380 66742 16436 66780
rect 16380 66388 16436 66398
rect 16380 66294 16436 66332
rect 16380 66052 16436 66062
rect 16380 65378 16436 65996
rect 16380 65326 16382 65378
rect 16434 65326 16436 65378
rect 16156 65266 16212 65278
rect 16156 65214 16158 65266
rect 16210 65214 16212 65266
rect 16156 63138 16212 65214
rect 16380 63588 16436 65326
rect 16492 64036 16548 67004
rect 16604 66948 16660 79548
rect 16828 78372 16884 81230
rect 16828 78306 16884 78316
rect 16940 81732 16996 81742
rect 16828 75796 16884 75806
rect 16828 75702 16884 75740
rect 16828 74900 16884 74910
rect 16828 74806 16884 74844
rect 16716 73218 16772 73230
rect 16716 73166 16718 73218
rect 16770 73166 16772 73218
rect 16716 72660 16772 73166
rect 16716 72212 16772 72604
rect 16716 72146 16772 72156
rect 16716 71204 16772 71214
rect 16716 70756 16772 71148
rect 16828 70980 16884 70990
rect 16828 70886 16884 70924
rect 16716 70690 16772 70700
rect 16716 69524 16772 69534
rect 16716 69076 16772 69468
rect 16940 69412 16996 81676
rect 17052 80612 17108 84364
rect 17612 84308 17668 84318
rect 17612 83524 17668 84252
rect 17612 83468 17780 83524
rect 17052 80546 17108 80556
rect 17164 83298 17220 83310
rect 17164 83246 17166 83298
rect 17218 83246 17220 83298
rect 17164 80948 17220 83246
rect 17612 83300 17668 83310
rect 17612 83206 17668 83244
rect 17500 82964 17556 82974
rect 17500 82870 17556 82908
rect 17164 78036 17220 80892
rect 16940 69346 16996 69356
rect 17052 77980 17220 78036
rect 17276 82404 17332 82414
rect 17332 82348 17444 82404
rect 17276 82292 17444 82348
rect 16828 69300 16884 69310
rect 16828 69206 16884 69244
rect 16716 69020 16884 69076
rect 16716 68852 16772 68862
rect 16716 67170 16772 68796
rect 16828 68850 16884 69020
rect 16828 68798 16830 68850
rect 16882 68798 16884 68850
rect 16828 68786 16884 68798
rect 16716 67118 16718 67170
rect 16770 67118 16772 67170
rect 16716 67106 16772 67118
rect 16940 68404 16996 68414
rect 16604 66892 16772 66948
rect 16492 63970 16548 63980
rect 16604 64484 16660 64494
rect 16380 63532 16548 63588
rect 16268 63476 16324 63486
rect 16268 63250 16324 63420
rect 16268 63198 16270 63250
rect 16322 63198 16324 63250
rect 16268 63186 16324 63198
rect 16380 63364 16436 63374
rect 16156 63086 16158 63138
rect 16210 63086 16212 63138
rect 16156 63074 16212 63086
rect 16380 63138 16436 63308
rect 16380 63086 16382 63138
rect 16434 63086 16436 63138
rect 16380 63074 16436 63086
rect 16044 62290 16100 62300
rect 16268 62916 16324 62926
rect 16268 62466 16324 62860
rect 16268 62414 16270 62466
rect 16322 62414 16324 62466
rect 15820 62242 15876 62254
rect 15820 62190 15822 62242
rect 15874 62190 15876 62242
rect 15820 62132 15876 62190
rect 15820 62066 15876 62076
rect 16044 62130 16100 62142
rect 16044 62078 16046 62130
rect 16098 62078 16100 62130
rect 15596 61730 15652 61740
rect 16044 61570 16100 62078
rect 16044 61518 16046 61570
rect 16098 61518 16100 61570
rect 15484 60162 15540 60172
rect 15820 61012 15876 61022
rect 15820 59332 15876 60956
rect 16044 60116 16100 61518
rect 16156 61458 16212 61470
rect 16156 61406 16158 61458
rect 16210 61406 16212 61458
rect 16156 61236 16212 61406
rect 16156 61170 16212 61180
rect 16268 61460 16324 62414
rect 16268 60340 16324 61404
rect 16380 60786 16436 60798
rect 16380 60734 16382 60786
rect 16434 60734 16436 60786
rect 16380 60676 16436 60734
rect 16380 60610 16436 60620
rect 16268 60274 16324 60284
rect 15596 59330 15876 59332
rect 15596 59278 15822 59330
rect 15874 59278 15876 59330
rect 15596 59276 15876 59278
rect 15484 59218 15540 59230
rect 15484 59166 15486 59218
rect 15538 59166 15540 59218
rect 15484 58772 15540 59166
rect 15484 58706 15540 58716
rect 15596 58884 15652 59276
rect 15820 59266 15876 59276
rect 15932 60060 16100 60116
rect 15596 58546 15652 58828
rect 15596 58494 15598 58546
rect 15650 58494 15652 58546
rect 15596 58482 15652 58494
rect 15708 58994 15764 59006
rect 15708 58942 15710 58994
rect 15762 58942 15764 58994
rect 15372 58268 15540 58324
rect 14924 58156 15204 58212
rect 15260 58156 15428 58212
rect 14820 58044 15084 58054
rect 14876 57988 14924 58044
rect 14980 57988 15028 58044
rect 14820 57978 15084 57988
rect 15148 57876 15204 58156
rect 15036 57820 15204 57876
rect 15260 57988 15316 57998
rect 15036 56756 15092 57820
rect 15148 57652 15204 57662
rect 15260 57652 15316 57932
rect 15148 57650 15316 57652
rect 15148 57598 15150 57650
rect 15202 57598 15316 57650
rect 15148 57596 15316 57598
rect 15148 57586 15204 57596
rect 15372 56868 15428 58156
rect 15484 57762 15540 58268
rect 15484 57710 15486 57762
rect 15538 57710 15540 57762
rect 15484 57204 15540 57710
rect 15484 57138 15540 57148
rect 15596 57650 15652 57662
rect 15596 57598 15598 57650
rect 15650 57598 15652 57650
rect 15372 56802 15428 56812
rect 15596 56756 15652 57598
rect 15036 56642 15092 56700
rect 15036 56590 15038 56642
rect 15090 56590 15092 56642
rect 15036 56578 15092 56590
rect 15484 56754 15652 56756
rect 15484 56702 15598 56754
rect 15650 56702 15652 56754
rect 15484 56700 15652 56702
rect 14820 56476 15084 56486
rect 14876 56420 14924 56476
rect 14980 56420 15028 56476
rect 14820 56410 15084 56420
rect 15484 56308 15540 56700
rect 15596 56690 15652 56700
rect 15372 56252 15540 56308
rect 15036 56196 15092 56206
rect 15036 56102 15092 56140
rect 14812 56084 14868 56094
rect 14476 56082 14644 56084
rect 14476 56030 14478 56082
rect 14530 56030 14644 56082
rect 14476 56028 14644 56030
rect 14700 56082 14868 56084
rect 14700 56030 14814 56082
rect 14866 56030 14868 56082
rect 14700 56028 14868 56030
rect 14476 56018 14532 56028
rect 14364 55804 14532 55860
rect 14140 55682 14196 55692
rect 14028 55468 14196 55524
rect 14028 55188 14084 55198
rect 14028 55074 14084 55132
rect 14028 55022 14030 55074
rect 14082 55022 14084 55074
rect 13916 53844 13972 53854
rect 13804 53842 13972 53844
rect 13804 53790 13918 53842
rect 13970 53790 13972 53842
rect 13804 53788 13972 53790
rect 12796 53454 12798 53506
rect 12850 53454 12852 53506
rect 12572 53218 12628 53228
rect 12796 53060 12852 53454
rect 12684 53004 12852 53060
rect 13020 53452 13300 53508
rect 12572 52946 12628 52958
rect 12572 52894 12574 52946
rect 12626 52894 12628 52946
rect 12572 52500 12628 52894
rect 12572 52434 12628 52444
rect 12572 50932 12628 50942
rect 12460 50876 12572 50932
rect 12572 50866 12628 50876
rect 12684 50594 12740 53004
rect 12796 52836 12852 52846
rect 12796 52834 12964 52836
rect 12796 52782 12798 52834
rect 12850 52782 12964 52834
rect 12796 52780 12964 52782
rect 12796 52770 12852 52780
rect 12460 50538 12516 50550
rect 12460 50486 12462 50538
rect 12514 50486 12516 50538
rect 12684 50542 12686 50594
rect 12738 50542 12740 50594
rect 12684 50530 12740 50542
rect 12796 52612 12852 52622
rect 12460 50484 12516 50486
rect 12796 50428 12852 52556
rect 12460 50418 12516 50428
rect 12572 50372 12852 50428
rect 12460 49812 12516 49822
rect 12348 49810 12516 49812
rect 12348 49758 12462 49810
rect 12514 49758 12516 49810
rect 12348 49756 12516 49758
rect 12236 49074 12292 49084
rect 12124 49028 12180 49038
rect 12012 49026 12180 49028
rect 12012 48974 12126 49026
rect 12178 48974 12180 49026
rect 12012 48972 12180 48974
rect 12124 48962 12180 48972
rect 12348 49028 12404 49038
rect 12460 49028 12516 49756
rect 12572 49140 12628 50372
rect 12684 49812 12740 49822
rect 12684 49810 12852 49812
rect 12684 49758 12686 49810
rect 12738 49758 12852 49810
rect 12684 49756 12852 49758
rect 12684 49746 12740 49756
rect 12572 49084 12740 49140
rect 12404 48972 12516 49028
rect 12348 48934 12404 48972
rect 12572 48916 12628 48926
rect 12572 48822 12628 48860
rect 12236 48804 12292 48814
rect 12236 48466 12292 48748
rect 12684 48692 12740 49084
rect 12796 48916 12852 49756
rect 12796 48850 12852 48860
rect 12236 48414 12238 48466
rect 12290 48414 12292 48466
rect 12236 48402 12292 48414
rect 12348 48636 12740 48692
rect 11564 47518 11566 47570
rect 11618 47518 11620 47570
rect 11564 47506 11620 47518
rect 11788 47516 11956 47572
rect 12124 48018 12180 48030
rect 12124 47966 12126 48018
rect 12178 47966 12180 48018
rect 11788 47124 11844 47516
rect 12012 47460 12068 47470
rect 11788 47058 11844 47068
rect 11900 47404 12012 47460
rect 11900 47012 11956 47404
rect 12012 47394 12068 47404
rect 12124 47460 12180 47966
rect 12236 47460 12292 47470
rect 12124 47404 12236 47460
rect 12012 47236 12068 47246
rect 12124 47236 12180 47404
rect 12236 47394 12292 47404
rect 12068 47180 12180 47236
rect 12012 47142 12068 47180
rect 11900 46956 12068 47012
rect 11452 46498 11508 46508
rect 11418 46284 11682 46294
rect 11474 46228 11522 46284
rect 11578 46228 11626 46284
rect 11418 46218 11682 46228
rect 12012 46116 12068 46956
rect 11228 46060 11396 46116
rect 11116 45948 11284 46004
rect 11228 45890 11284 45948
rect 11228 45838 11230 45890
rect 11282 45838 11284 45890
rect 11228 45826 11284 45838
rect 11116 45780 11172 45790
rect 11116 45686 11172 45724
rect 11340 45332 11396 46060
rect 11788 46060 12068 46116
rect 11452 45778 11508 45790
rect 11452 45726 11454 45778
rect 11506 45726 11508 45778
rect 11452 45556 11508 45726
rect 11676 45780 11732 45790
rect 11676 45686 11732 45724
rect 11452 45490 11508 45500
rect 11452 45332 11508 45342
rect 11228 45330 11508 45332
rect 11228 45278 11454 45330
rect 11506 45278 11508 45330
rect 11228 45276 11508 45278
rect 11004 44996 11060 45006
rect 11228 44996 11284 45276
rect 11452 45266 11508 45276
rect 11004 44994 11284 44996
rect 11004 44942 11006 44994
rect 11058 44942 11284 44994
rect 11004 44940 11284 44942
rect 11004 44930 11060 44940
rect 10892 44716 11172 44772
rect 10668 44324 10724 44334
rect 10780 44324 10836 44380
rect 10668 44322 10836 44324
rect 10668 44270 10670 44322
rect 10722 44270 10836 44322
rect 10668 44268 10836 44270
rect 10668 44258 10724 44268
rect 10556 43810 10612 43820
rect 10780 44098 10836 44110
rect 10780 44046 10782 44098
rect 10834 44046 10836 44098
rect 10444 43652 10500 43662
rect 10444 43650 10724 43652
rect 10444 43598 10446 43650
rect 10498 43598 10724 43650
rect 10444 43596 10724 43598
rect 10444 43586 10500 43596
rect 9996 43036 10276 43092
rect 10220 42756 10276 43036
rect 10332 43026 10388 43036
rect 10668 42868 10724 43596
rect 10780 43538 10836 44046
rect 10780 43486 10782 43538
rect 10834 43486 10836 43538
rect 10780 43474 10836 43486
rect 10892 44098 10948 44110
rect 10892 44046 10894 44098
rect 10946 44046 10948 44098
rect 10892 43204 10948 44046
rect 11004 44098 11060 44110
rect 11004 44046 11006 44098
rect 11058 44046 11060 44098
rect 11004 43876 11060 44046
rect 11004 43810 11060 43820
rect 11004 43652 11060 43662
rect 11004 43558 11060 43596
rect 10892 43138 10948 43148
rect 10780 42868 10836 42878
rect 10668 42866 10836 42868
rect 10668 42814 10782 42866
rect 10834 42814 10836 42866
rect 10668 42812 10836 42814
rect 10780 42802 10836 42812
rect 10220 42700 10388 42756
rect 9996 42642 10052 42654
rect 9996 42590 9998 42642
rect 10050 42590 10052 42642
rect 9884 42530 9940 42542
rect 9884 42478 9886 42530
rect 9938 42478 9940 42530
rect 9884 42196 9940 42478
rect 9996 42308 10052 42590
rect 9996 42242 10052 42252
rect 9884 42130 9940 42140
rect 10220 41970 10276 41982
rect 10220 41918 10222 41970
rect 10274 41918 10276 41970
rect 9884 41860 9940 41870
rect 9884 41766 9940 41804
rect 10220 41748 10276 41918
rect 10332 41970 10388 42700
rect 10444 42642 10500 42654
rect 10444 42590 10446 42642
rect 10498 42590 10500 42642
rect 10444 42532 10500 42590
rect 10780 42644 10836 42654
rect 10444 42466 10500 42476
rect 10668 42530 10724 42542
rect 10668 42478 10670 42530
rect 10722 42478 10724 42530
rect 10668 42308 10724 42478
rect 10332 41918 10334 41970
rect 10386 41918 10388 41970
rect 10332 41906 10388 41918
rect 10444 42252 10724 42308
rect 10444 41972 10500 42252
rect 10780 42196 10836 42588
rect 10668 42140 10836 42196
rect 10892 42530 10948 42542
rect 10892 42478 10894 42530
rect 10946 42478 10948 42530
rect 10556 42084 10612 42094
rect 10668 42084 10724 42140
rect 10556 42082 10724 42084
rect 10556 42030 10558 42082
rect 10610 42030 10724 42082
rect 10556 42028 10724 42030
rect 10556 42018 10612 42028
rect 10444 41906 10500 41916
rect 10780 41970 10836 41982
rect 10780 41918 10782 41970
rect 10834 41918 10836 41970
rect 10780 41860 10836 41918
rect 10220 41692 10724 41748
rect 9996 41300 10052 41310
rect 9884 40404 9940 40414
rect 9996 40404 10052 41244
rect 10556 41300 10612 41310
rect 10556 41206 10612 41244
rect 10332 40852 10388 40862
rect 10332 40626 10388 40796
rect 10332 40574 10334 40626
rect 10386 40574 10388 40626
rect 10332 40562 10388 40574
rect 10668 40628 10724 41692
rect 10780 40852 10836 41804
rect 10892 41300 10948 42478
rect 11004 42532 11060 42542
rect 11004 42438 11060 42476
rect 11116 42308 11172 44716
rect 11418 44716 11682 44726
rect 11474 44660 11522 44716
rect 11578 44660 11626 44716
rect 11418 44650 11682 44660
rect 11788 44548 11844 46060
rect 12348 46004 12404 48636
rect 12684 48468 12740 48478
rect 12908 48468 12964 52780
rect 13020 52274 13076 53452
rect 13692 53058 13748 53070
rect 13692 53006 13694 53058
rect 13746 53006 13748 53058
rect 13692 52948 13748 53006
rect 13692 52882 13748 52892
rect 13580 52834 13636 52846
rect 13580 52782 13582 52834
rect 13634 52782 13636 52834
rect 13580 52612 13636 52782
rect 13580 52546 13636 52556
rect 13692 52724 13748 52734
rect 13020 52222 13022 52274
rect 13074 52222 13076 52274
rect 13020 52210 13076 52222
rect 13356 52388 13412 52398
rect 13244 50932 13300 50942
rect 13132 50708 13188 50718
rect 13020 50484 13076 50494
rect 13020 50390 13076 50428
rect 13020 49810 13076 49822
rect 13020 49758 13022 49810
rect 13074 49758 13076 49810
rect 13020 48804 13076 49758
rect 13020 48738 13076 48748
rect 13132 48468 13188 50652
rect 12908 48412 13076 48468
rect 12012 45948 12404 46004
rect 12460 47684 12516 47694
rect 12460 47570 12516 47628
rect 12460 47518 12462 47570
rect 12514 47518 12516 47570
rect 12460 46004 12516 47518
rect 11900 45892 11956 45902
rect 11900 45330 11956 45836
rect 11900 45278 11902 45330
rect 11954 45278 11956 45330
rect 11900 44882 11956 45278
rect 11900 44830 11902 44882
rect 11954 44830 11956 44882
rect 11900 44818 11956 44830
rect 12012 44548 12068 45948
rect 12460 45938 12516 45948
rect 12236 45780 12292 45790
rect 12236 45686 12292 45724
rect 12124 45668 12180 45678
rect 12124 44772 12180 45612
rect 12348 45666 12404 45678
rect 12572 45668 12628 45678
rect 12348 45614 12350 45666
rect 12402 45614 12404 45666
rect 12348 45220 12404 45614
rect 12348 45154 12404 45164
rect 12460 45666 12628 45668
rect 12460 45614 12574 45666
rect 12626 45614 12628 45666
rect 12460 45612 12628 45614
rect 12348 44994 12404 45006
rect 12348 44942 12350 44994
rect 12402 44942 12404 44994
rect 12348 44882 12404 44942
rect 12348 44830 12350 44882
rect 12402 44830 12404 44882
rect 12348 44818 12404 44830
rect 12124 44706 12180 44716
rect 11788 44492 11956 44548
rect 12012 44492 12404 44548
rect 11340 44436 11396 44446
rect 11396 44380 11508 44436
rect 11340 44370 11396 44380
rect 11340 43540 11396 43550
rect 11340 43446 11396 43484
rect 11452 43316 11508 44380
rect 10892 41234 10948 41244
rect 11004 42252 11172 42308
rect 11228 43260 11508 43316
rect 11676 44324 11732 44334
rect 11676 43316 11732 44268
rect 11788 44098 11844 44110
rect 11788 44046 11790 44098
rect 11842 44046 11844 44098
rect 11788 43540 11844 44046
rect 11788 43474 11844 43484
rect 11676 43260 11844 43316
rect 10780 40786 10836 40796
rect 10892 40740 10948 40750
rect 10780 40628 10836 40638
rect 10668 40626 10836 40628
rect 10668 40574 10782 40626
rect 10834 40574 10836 40626
rect 10668 40572 10836 40574
rect 9884 40402 10164 40404
rect 9884 40350 9886 40402
rect 9938 40350 10164 40402
rect 9884 40348 10164 40350
rect 9884 40338 9940 40348
rect 10108 40292 10164 40348
rect 10108 40236 10276 40292
rect 10220 40180 10276 40236
rect 10220 40124 10388 40180
rect 10108 40068 10164 40078
rect 9996 39618 10052 39630
rect 9996 39566 9998 39618
rect 10050 39566 10052 39618
rect 9996 39172 10052 39566
rect 9996 39106 10052 39116
rect 10108 39058 10164 40012
rect 10108 39006 10110 39058
rect 10162 39006 10164 39058
rect 10108 38994 10164 39006
rect 9660 38612 9828 38668
rect 10332 38668 10388 40124
rect 10668 39844 10724 40572
rect 10780 40562 10836 40572
rect 10892 40404 10948 40684
rect 10668 39778 10724 39788
rect 10780 40348 10948 40404
rect 10780 39730 10836 40348
rect 10780 39678 10782 39730
rect 10834 39678 10836 39730
rect 10780 39666 10836 39678
rect 10892 39172 10948 39182
rect 10892 39058 10948 39116
rect 10892 39006 10894 39058
rect 10946 39006 10948 39058
rect 10892 38994 10948 39006
rect 11004 38836 11060 42252
rect 11228 42196 11284 43260
rect 11418 43148 11682 43158
rect 11474 43092 11522 43148
rect 11578 43092 11626 43148
rect 11418 43082 11682 43092
rect 11788 42980 11844 43260
rect 11676 42924 11844 42980
rect 11564 42532 11620 42542
rect 11564 42438 11620 42476
rect 11228 42130 11284 42140
rect 11676 42084 11732 42924
rect 11676 41990 11732 42028
rect 11418 41580 11682 41590
rect 11474 41524 11522 41580
rect 11578 41524 11626 41580
rect 11418 41514 11682 41524
rect 11788 41300 11844 41310
rect 11788 41206 11844 41244
rect 11340 40962 11396 40974
rect 11340 40910 11342 40962
rect 11394 40910 11396 40962
rect 11228 40852 11284 40862
rect 11340 40852 11396 40910
rect 11284 40796 11396 40852
rect 11228 40786 11284 40796
rect 11564 40740 11620 40750
rect 11228 40628 11284 40638
rect 11116 40516 11172 40526
rect 11116 40422 11172 40460
rect 11228 40292 11284 40572
rect 11564 40626 11620 40684
rect 11564 40574 11566 40626
rect 11618 40574 11620 40626
rect 11564 40562 11620 40574
rect 11340 40402 11396 40414
rect 11340 40350 11342 40402
rect 11394 40350 11396 40402
rect 11340 40292 11396 40350
rect 11788 40404 11844 40414
rect 11788 40310 11844 40348
rect 11116 40236 11396 40292
rect 11116 39060 11172 40236
rect 11676 40180 11732 40190
rect 11676 40178 11844 40180
rect 11676 40126 11678 40178
rect 11730 40126 11844 40178
rect 11676 40124 11844 40126
rect 11676 40114 11732 40124
rect 11788 40068 11844 40124
rect 11418 40012 11682 40022
rect 11474 39956 11522 40012
rect 11578 39956 11626 40012
rect 11788 40002 11844 40012
rect 11418 39946 11682 39956
rect 11676 39844 11732 39854
rect 11340 39060 11396 39070
rect 11116 39058 11396 39060
rect 11116 39006 11342 39058
rect 11394 39006 11396 39058
rect 11116 39004 11396 39006
rect 11340 38994 11396 39004
rect 11676 38948 11732 39788
rect 11676 38892 11844 38948
rect 10892 38780 11060 38836
rect 10332 38612 10612 38668
rect 9660 38276 9716 38612
rect 9660 37492 9716 38220
rect 10108 38164 10164 38174
rect 10108 38050 10164 38108
rect 10108 37998 10110 38050
rect 10162 37998 10164 38050
rect 10108 37986 10164 37998
rect 10556 38050 10612 38612
rect 10556 37998 10558 38050
rect 10610 37998 10612 38050
rect 10556 37986 10612 37998
rect 10780 38052 10836 38062
rect 10780 37958 10836 37996
rect 10332 37826 10388 37838
rect 10332 37774 10334 37826
rect 10386 37774 10388 37826
rect 10332 37604 10388 37774
rect 10332 37538 10388 37548
rect 10444 37826 10500 37838
rect 10444 37774 10446 37826
rect 10498 37774 10500 37826
rect 9660 37398 9716 37436
rect 10108 37380 10164 37390
rect 10108 37286 10164 37324
rect 9996 37268 10052 37278
rect 10332 37268 10388 37278
rect 9996 37174 10052 37212
rect 10220 37266 10388 37268
rect 10220 37214 10334 37266
rect 10386 37214 10388 37266
rect 10220 37212 10388 37214
rect 10444 37268 10500 37774
rect 10556 37268 10612 37278
rect 10444 37266 10612 37268
rect 10444 37214 10558 37266
rect 10610 37214 10612 37266
rect 10444 37212 10612 37214
rect 9996 36594 10052 36606
rect 9996 36542 9998 36594
rect 10050 36542 10052 36594
rect 9996 36372 10052 36542
rect 9996 36306 10052 36316
rect 10108 35924 10164 35934
rect 10108 35830 10164 35868
rect 9660 35812 9716 35822
rect 9660 35718 9716 35756
rect 10220 35308 10276 37212
rect 10332 37202 10388 37212
rect 10556 37202 10612 37212
rect 10444 36932 10500 36942
rect 9884 35252 10276 35308
rect 10332 35588 10388 35598
rect 9548 34804 9604 34814
rect 9772 34804 9828 34814
rect 9548 34802 9772 34804
rect 9548 34750 9550 34802
rect 9602 34750 9772 34802
rect 9548 34748 9772 34750
rect 9548 34738 9604 34748
rect 9772 34710 9828 34748
rect 9884 34356 9940 35252
rect 10108 34916 10164 34926
rect 10108 34822 10164 34860
rect 10332 34802 10388 35532
rect 10444 34916 10500 36876
rect 10444 34850 10500 34860
rect 10556 36820 10612 36830
rect 10332 34750 10334 34802
rect 10386 34750 10388 34802
rect 10108 34690 10164 34702
rect 10108 34638 10110 34690
rect 10162 34638 10164 34690
rect 10108 34580 10164 34638
rect 10108 34514 10164 34524
rect 9660 34300 9940 34356
rect 9548 34130 9604 34142
rect 9548 34078 9550 34130
rect 9602 34078 9604 34130
rect 9548 33796 9604 34078
rect 9548 33730 9604 33740
rect 9548 33570 9604 33582
rect 9548 33518 9550 33570
rect 9602 33518 9604 33570
rect 9548 33458 9604 33518
rect 9548 33406 9550 33458
rect 9602 33406 9604 33458
rect 9548 33394 9604 33406
rect 9660 33012 9716 34300
rect 9772 34132 9828 34142
rect 9772 33570 9828 34076
rect 9996 34130 10052 34142
rect 9996 34078 9998 34130
rect 10050 34078 10052 34130
rect 9772 33518 9774 33570
rect 9826 33518 9828 33570
rect 9772 33506 9828 33518
rect 9884 34018 9940 34030
rect 9884 33966 9886 34018
rect 9938 33966 9940 34018
rect 9884 33236 9940 33966
rect 9884 33170 9940 33180
rect 9996 34020 10052 34078
rect 9660 32956 9940 33012
rect 9772 32004 9828 32014
rect 9660 31948 9772 32004
rect 9548 31666 9604 31678
rect 9548 31614 9550 31666
rect 9602 31614 9604 31666
rect 9548 30996 9604 31614
rect 9548 30930 9604 30940
rect 9548 30324 9604 30334
rect 9660 30324 9716 31948
rect 9772 31938 9828 31948
rect 9884 31892 9940 32956
rect 9996 32228 10052 33964
rect 10108 34130 10164 34142
rect 10108 34078 10110 34130
rect 10162 34078 10164 34130
rect 10108 33908 10164 34078
rect 10108 33842 10164 33852
rect 10332 33908 10388 34750
rect 10556 34356 10612 36764
rect 10780 35588 10836 35598
rect 10780 35494 10836 35532
rect 10780 35028 10836 35038
rect 10668 34914 10724 34926
rect 10668 34862 10670 34914
rect 10722 34862 10724 34914
rect 10668 34580 10724 34862
rect 10780 34802 10836 34972
rect 10780 34750 10782 34802
rect 10834 34750 10836 34802
rect 10780 34738 10836 34750
rect 10668 34514 10724 34524
rect 10332 33842 10388 33852
rect 10444 34300 10612 34356
rect 10108 33570 10164 33582
rect 10444 33572 10500 34300
rect 10556 34130 10612 34142
rect 10556 34078 10558 34130
rect 10610 34078 10612 34130
rect 10556 33908 10612 34078
rect 10780 34130 10836 34142
rect 10780 34078 10782 34130
rect 10834 34078 10836 34130
rect 10556 33842 10612 33852
rect 10668 34018 10724 34030
rect 10668 33966 10670 34018
rect 10722 33966 10724 34018
rect 10108 33518 10110 33570
rect 10162 33518 10164 33570
rect 10108 33458 10164 33518
rect 10108 33406 10110 33458
rect 10162 33406 10164 33458
rect 10108 33394 10164 33406
rect 10220 33516 10500 33572
rect 10668 33572 10724 33966
rect 9996 32162 10052 32172
rect 10220 32900 10276 33516
rect 10668 33506 10724 33516
rect 10444 33348 10500 33358
rect 10444 33254 10500 33292
rect 10556 33236 10612 33246
rect 10556 33142 10612 33180
rect 10668 33234 10724 33246
rect 10668 33182 10670 33234
rect 10722 33182 10724 33234
rect 10220 32844 10500 32900
rect 9996 31892 10052 31902
rect 9884 31890 10052 31892
rect 9884 31838 9998 31890
rect 10050 31838 10052 31890
rect 9884 31836 10052 31838
rect 9996 31826 10052 31836
rect 9772 31780 9828 31790
rect 9772 31686 9828 31724
rect 10220 31778 10276 32844
rect 10444 32786 10500 32844
rect 10444 32734 10446 32786
rect 10498 32734 10500 32786
rect 10444 32722 10500 32734
rect 10668 32004 10724 33182
rect 10780 32116 10836 34078
rect 10892 32900 10948 38780
rect 11676 38724 11732 38734
rect 11676 38630 11732 38668
rect 11788 38612 11844 38892
rect 11788 38546 11844 38556
rect 11228 38500 11284 38510
rect 11116 38444 11228 38500
rect 11004 37380 11060 37390
rect 11004 37286 11060 37324
rect 11004 36932 11060 36942
rect 11004 35252 11060 36876
rect 11004 35186 11060 35196
rect 11004 34802 11060 34814
rect 11004 34750 11006 34802
rect 11058 34750 11060 34802
rect 11004 33012 11060 34750
rect 11116 34356 11172 38444
rect 11228 38434 11284 38444
rect 11418 38444 11682 38454
rect 11474 38388 11522 38444
rect 11578 38388 11626 38444
rect 11418 38378 11682 38388
rect 11788 38274 11844 38286
rect 11788 38222 11790 38274
rect 11842 38222 11844 38274
rect 11228 38164 11284 38174
rect 11284 38108 11396 38164
rect 11228 38098 11284 38108
rect 11228 37826 11284 37838
rect 11228 37774 11230 37826
rect 11282 37774 11284 37826
rect 11228 37604 11284 37774
rect 11228 37538 11284 37548
rect 11228 37380 11284 37390
rect 11340 37380 11396 38108
rect 11788 38162 11844 38222
rect 11788 38110 11790 38162
rect 11842 38110 11844 38162
rect 11452 37492 11508 37502
rect 11452 37490 11620 37492
rect 11452 37438 11454 37490
rect 11506 37438 11620 37490
rect 11452 37436 11620 37438
rect 11452 37426 11508 37436
rect 11228 37378 11396 37380
rect 11228 37326 11230 37378
rect 11282 37326 11396 37378
rect 11228 37324 11396 37326
rect 11228 35588 11284 37324
rect 11452 37266 11508 37278
rect 11452 37214 11454 37266
rect 11506 37214 11508 37266
rect 11452 37156 11508 37214
rect 11564 37268 11620 37436
rect 11564 37202 11620 37212
rect 11788 37378 11844 38110
rect 11788 37326 11790 37378
rect 11842 37326 11844 37378
rect 11452 37090 11508 37100
rect 11418 36876 11682 36886
rect 11474 36820 11522 36876
rect 11578 36820 11626 36876
rect 11418 36810 11682 36820
rect 11228 35522 11284 35532
rect 11676 35588 11732 35598
rect 11676 35494 11732 35532
rect 11418 35308 11682 35318
rect 11474 35252 11522 35308
rect 11578 35252 11626 35308
rect 11418 35242 11682 35252
rect 11676 35140 11732 35150
rect 11676 35046 11732 35084
rect 11340 34916 11396 34926
rect 11340 34822 11396 34860
rect 11116 34290 11172 34300
rect 11788 34804 11844 37326
rect 11788 34356 11844 34748
rect 11788 34290 11844 34300
rect 11116 34132 11172 34142
rect 11116 34038 11172 34076
rect 11564 34018 11620 34030
rect 11564 33966 11566 34018
rect 11618 33966 11620 34018
rect 11228 33908 11284 33918
rect 11564 33908 11620 33966
rect 11284 33852 11620 33908
rect 11116 33348 11172 33358
rect 11116 33254 11172 33292
rect 11004 32956 11172 33012
rect 10892 32834 10948 32844
rect 11004 32788 11060 32798
rect 11004 32694 11060 32732
rect 11116 32452 11172 32956
rect 10780 32050 10836 32060
rect 10892 32396 11172 32452
rect 10668 31938 10724 31948
rect 10220 31726 10222 31778
rect 10274 31726 10276 31778
rect 9996 31554 10052 31566
rect 9996 31502 9998 31554
rect 10050 31502 10052 31554
rect 9884 31444 9940 31454
rect 9884 31218 9940 31388
rect 9884 31166 9886 31218
rect 9938 31166 9940 31218
rect 9772 30324 9828 30334
rect 9660 30322 9828 30324
rect 9660 30270 9774 30322
rect 9826 30270 9828 30322
rect 9660 30268 9828 30270
rect 9548 30210 9604 30268
rect 9772 30258 9828 30268
rect 9548 30158 9550 30210
rect 9602 30158 9604 30210
rect 9548 30146 9604 30158
rect 9884 30210 9940 31166
rect 9884 30158 9886 30210
rect 9938 30158 9940 30210
rect 9884 30100 9940 30158
rect 9884 30034 9940 30044
rect 9660 29988 9716 29998
rect 9660 29316 9716 29932
rect 9660 29222 9716 29260
rect 9772 29986 9828 29998
rect 9772 29934 9774 29986
rect 9826 29934 9828 29986
rect 9660 27748 9716 27758
rect 9660 27654 9716 27692
rect 9548 27412 9604 27422
rect 9548 26516 9604 27356
rect 9660 27076 9716 27086
rect 9660 26982 9716 27020
rect 9660 26516 9716 26526
rect 9548 26514 9716 26516
rect 9548 26462 9662 26514
rect 9714 26462 9716 26514
rect 9548 26460 9716 26462
rect 9660 26450 9716 26460
rect 9548 26068 9604 26078
rect 9548 23940 9604 26012
rect 9660 25284 9716 25294
rect 9660 24722 9716 25228
rect 9660 24670 9662 24722
rect 9714 24670 9716 24722
rect 9660 24658 9716 24670
rect 9772 24724 9828 29934
rect 9884 28196 9940 28206
rect 9884 26292 9940 28140
rect 9996 26404 10052 31502
rect 10220 31444 10276 31726
rect 10220 31378 10276 31388
rect 10332 31892 10388 31902
rect 10220 31220 10276 31230
rect 10332 31220 10388 31836
rect 10220 31218 10612 31220
rect 10220 31166 10222 31218
rect 10274 31166 10612 31218
rect 10220 31164 10612 31166
rect 10220 31154 10276 31164
rect 10556 30324 10612 31164
rect 10332 30212 10388 30222
rect 10332 30118 10388 30156
rect 10556 30210 10612 30268
rect 10556 30158 10558 30210
rect 10610 30158 10612 30210
rect 10556 30146 10612 30158
rect 10668 30994 10724 31006
rect 10668 30942 10670 30994
rect 10722 30942 10724 30994
rect 10668 30212 10724 30942
rect 10892 30322 10948 32396
rect 11228 32340 11284 33852
rect 11418 33740 11682 33750
rect 11474 33684 11522 33740
rect 11578 33684 11626 33740
rect 11418 33674 11682 33684
rect 11900 33348 11956 44492
rect 12236 44324 12292 44334
rect 12236 44230 12292 44268
rect 12012 44212 12068 44222
rect 12012 44118 12068 44156
rect 12124 44098 12180 44110
rect 12124 44046 12126 44098
rect 12178 44046 12180 44098
rect 12124 43650 12180 44046
rect 12124 43598 12126 43650
rect 12178 43598 12180 43650
rect 12124 43586 12180 43598
rect 12124 42980 12180 42990
rect 12012 42924 12124 42980
rect 12012 42866 12068 42924
rect 12124 42914 12180 42924
rect 12012 42814 12014 42866
rect 12066 42814 12068 42866
rect 12012 42532 12068 42814
rect 12012 42466 12068 42476
rect 12348 42196 12404 44492
rect 12460 44100 12516 45612
rect 12572 45602 12628 45612
rect 12572 44436 12628 44446
rect 12572 44322 12628 44380
rect 12572 44270 12574 44322
rect 12626 44270 12628 44322
rect 12572 44258 12628 44270
rect 12460 44034 12516 44044
rect 12684 42868 12740 48412
rect 12908 47236 12964 47246
rect 12908 47142 12964 47180
rect 12796 46004 12852 46014
rect 12796 45330 12852 45948
rect 12796 45278 12798 45330
rect 12850 45278 12852 45330
rect 12796 45266 12852 45278
rect 12908 45108 12964 45118
rect 12908 44324 12964 45052
rect 13020 44436 13076 48412
rect 13132 48402 13188 48412
rect 13244 46788 13300 50876
rect 13244 46722 13300 46732
rect 13244 46562 13300 46574
rect 13244 46510 13246 46562
rect 13298 46510 13300 46562
rect 13244 45220 13300 46510
rect 13244 45154 13300 45164
rect 13244 44994 13300 45006
rect 13244 44942 13246 44994
rect 13298 44942 13300 44994
rect 13244 44882 13300 44942
rect 13244 44830 13246 44882
rect 13298 44830 13300 44882
rect 13244 44818 13300 44830
rect 13020 44380 13300 44436
rect 12460 42530 12516 42542
rect 12460 42478 12462 42530
rect 12514 42478 12516 42530
rect 12460 42420 12516 42478
rect 12460 42354 12516 42364
rect 12124 42140 12516 42196
rect 12124 41972 12180 42140
rect 12124 41906 12180 41916
rect 12348 41972 12404 41982
rect 12348 41878 12404 41916
rect 12236 41860 12292 41870
rect 12012 41300 12068 41310
rect 12236 41300 12292 41804
rect 12012 33572 12068 41244
rect 12124 41244 12236 41300
rect 12124 38274 12180 41244
rect 12236 41234 12292 41244
rect 12460 41188 12516 42140
rect 12348 41132 12516 41188
rect 12236 41076 12292 41086
rect 12348 41076 12404 41132
rect 12236 41074 12404 41076
rect 12236 41022 12238 41074
rect 12290 41022 12404 41074
rect 12236 41020 12404 41022
rect 12236 40852 12292 41020
rect 12236 40786 12292 40796
rect 12460 40404 12516 40414
rect 12236 40292 12292 40302
rect 12236 40198 12292 40236
rect 12348 40290 12404 40302
rect 12348 40238 12350 40290
rect 12402 40238 12404 40290
rect 12348 40068 12404 40238
rect 12348 40002 12404 40012
rect 12348 38836 12404 38846
rect 12460 38836 12516 40348
rect 12404 38780 12516 38836
rect 12572 40402 12628 40414
rect 12572 40350 12574 40402
rect 12626 40350 12628 40402
rect 12348 38742 12404 38780
rect 12124 38222 12126 38274
rect 12178 38222 12180 38274
rect 12124 38210 12180 38222
rect 12236 38276 12292 38286
rect 12236 38052 12292 38220
rect 12124 37996 12292 38052
rect 12124 37266 12180 37996
rect 12348 37940 12404 37950
rect 12236 37828 12292 37838
rect 12348 37828 12404 37884
rect 12236 37826 12404 37828
rect 12236 37774 12238 37826
rect 12290 37774 12404 37826
rect 12236 37772 12404 37774
rect 12572 37828 12628 40350
rect 12684 38052 12740 42812
rect 12796 44212 12852 44222
rect 12796 40964 12852 44156
rect 12908 42866 12964 44268
rect 12908 42814 12910 42866
rect 12962 42814 12964 42866
rect 12908 42802 12964 42814
rect 13020 41860 13076 41870
rect 13020 41766 13076 41804
rect 13244 41524 13300 44380
rect 13132 41468 13300 41524
rect 13020 41076 13076 41086
rect 12796 40962 12964 40964
rect 12796 40910 12798 40962
rect 12850 40910 12964 40962
rect 12796 40908 12964 40910
rect 12796 40898 12852 40908
rect 12908 40628 12964 40908
rect 12908 40562 12964 40572
rect 12796 40516 12852 40526
rect 12796 39058 12852 40460
rect 12796 39006 12798 39058
rect 12850 39006 12852 39058
rect 12796 38388 12852 39006
rect 12796 38322 12852 38332
rect 12908 39730 12964 39742
rect 12908 39678 12910 39730
rect 12962 39678 12964 39730
rect 12908 38052 12964 39678
rect 12684 37986 12740 37996
rect 12796 37996 12964 38052
rect 12796 37828 12852 37996
rect 12572 37772 12852 37828
rect 12908 37826 12964 37838
rect 12908 37774 12910 37826
rect 12962 37774 12964 37826
rect 12236 37762 12292 37772
rect 12572 37716 12628 37772
rect 12460 37660 12628 37716
rect 12124 37214 12126 37266
rect 12178 37214 12180 37266
rect 12124 37202 12180 37214
rect 12236 37604 12292 37614
rect 12124 36596 12180 36606
rect 12124 36502 12180 36540
rect 12124 36372 12180 36382
rect 12124 35698 12180 36316
rect 12124 35646 12126 35698
rect 12178 35646 12180 35698
rect 12124 35634 12180 35646
rect 12236 35698 12292 37548
rect 12460 35922 12516 37660
rect 12572 37266 12628 37278
rect 12572 37214 12574 37266
rect 12626 37214 12628 37266
rect 12572 36372 12628 37214
rect 12796 37268 12852 37278
rect 12908 37268 12964 37774
rect 12796 37266 12964 37268
rect 12796 37214 12798 37266
rect 12850 37214 12964 37266
rect 12796 37212 12964 37214
rect 12684 37154 12740 37166
rect 12684 37102 12686 37154
rect 12738 37102 12740 37154
rect 12684 36484 12740 37102
rect 12796 37044 12852 37212
rect 12796 36978 12852 36988
rect 12908 36932 12964 36942
rect 12684 36418 12740 36428
rect 12796 36820 12852 36830
rect 12572 36306 12628 36316
rect 12460 35870 12462 35922
rect 12514 35870 12516 35922
rect 12460 35858 12516 35870
rect 12572 36036 12628 36046
rect 12236 35646 12238 35698
rect 12290 35646 12292 35698
rect 12236 34692 12292 35646
rect 12572 35698 12628 35980
rect 12572 35646 12574 35698
rect 12626 35646 12628 35698
rect 12348 35586 12404 35598
rect 12348 35534 12350 35586
rect 12402 35534 12404 35586
rect 12348 34916 12404 35534
rect 12348 34850 12404 34860
rect 12572 35588 12628 35646
rect 12460 34692 12516 34702
rect 12236 34690 12516 34692
rect 12236 34638 12462 34690
rect 12514 34638 12516 34690
rect 12236 34636 12516 34638
rect 12124 34356 12180 34366
rect 12124 34262 12180 34300
rect 12348 33908 12404 34636
rect 12460 34626 12516 34636
rect 12460 34020 12516 34030
rect 12460 33926 12516 33964
rect 12348 33842 12404 33852
rect 12012 33506 12068 33516
rect 11788 33292 11956 33348
rect 12012 33348 12068 33358
rect 11676 33234 11732 33246
rect 11676 33182 11678 33234
rect 11730 33182 11732 33234
rect 11340 33124 11396 33134
rect 11340 33030 11396 33068
rect 11452 32788 11508 32798
rect 11452 32694 11508 32732
rect 11116 32284 11284 32340
rect 11676 32340 11732 33182
rect 10892 30270 10894 30322
rect 10946 30270 10948 30322
rect 10892 30258 10948 30270
rect 11004 31556 11060 31566
rect 10668 30146 10724 30156
rect 10444 30100 10500 30110
rect 10220 29988 10276 29998
rect 10108 29932 10220 29988
rect 10108 26740 10164 29932
rect 10220 29922 10276 29932
rect 10332 29538 10388 29550
rect 10332 29486 10334 29538
rect 10386 29486 10388 29538
rect 10332 28196 10388 29486
rect 10444 29426 10500 30044
rect 10892 30100 10948 30110
rect 10892 30006 10948 30044
rect 10780 29988 10836 29998
rect 10780 29894 10836 29932
rect 10556 29650 10612 29662
rect 11004 29652 11060 31500
rect 10556 29598 10558 29650
rect 10610 29598 10612 29650
rect 10556 29540 10612 29598
rect 10556 29474 10612 29484
rect 10780 29596 11060 29652
rect 10444 29374 10446 29426
rect 10498 29374 10500 29426
rect 10444 29362 10500 29374
rect 10332 28130 10388 28140
rect 10444 28756 10500 28766
rect 10220 27972 10276 27982
rect 10220 27878 10276 27916
rect 10444 27970 10500 28700
rect 10780 28196 10836 29596
rect 11116 29540 11172 32284
rect 11676 32274 11732 32284
rect 11418 32172 11682 32182
rect 11228 32116 11284 32126
rect 11474 32116 11522 32172
rect 11578 32116 11626 32172
rect 11418 32106 11682 32116
rect 11228 29764 11284 32060
rect 11564 31780 11620 31790
rect 11564 31686 11620 31724
rect 11340 31666 11396 31678
rect 11340 31614 11342 31666
rect 11394 31614 11396 31666
rect 11340 31556 11396 31614
rect 11340 31490 11396 31500
rect 11452 31554 11508 31566
rect 11452 31502 11454 31554
rect 11506 31502 11508 31554
rect 11340 31108 11396 31118
rect 11452 31108 11508 31502
rect 11340 31106 11508 31108
rect 11340 31054 11342 31106
rect 11394 31054 11508 31106
rect 11340 31052 11508 31054
rect 11340 31042 11396 31052
rect 11418 30604 11682 30614
rect 11474 30548 11522 30604
rect 11578 30548 11626 30604
rect 11418 30538 11682 30548
rect 11452 30324 11508 30334
rect 11452 30230 11508 30268
rect 11228 29708 11396 29764
rect 11228 29540 11284 29550
rect 11116 29538 11284 29540
rect 11116 29486 11230 29538
rect 11282 29486 11284 29538
rect 11116 29484 11284 29486
rect 10892 29428 10948 29438
rect 10892 29334 10948 29372
rect 11116 29204 11172 29484
rect 11228 29474 11284 29484
rect 11340 29204 11396 29708
rect 11788 29428 11844 33292
rect 12012 33254 12068 33292
rect 12348 33348 12404 33358
rect 12572 33348 12628 35532
rect 12796 35308 12852 36764
rect 12684 35252 12852 35308
rect 12908 36482 12964 36876
rect 12908 36430 12910 36482
rect 12962 36430 12964 36482
rect 12908 35812 12964 36430
rect 12684 35028 12740 35252
rect 12684 34962 12740 34972
rect 12908 35026 12964 35756
rect 12908 34974 12910 35026
rect 12962 34974 12964 35026
rect 12348 33346 12628 33348
rect 12348 33294 12350 33346
rect 12402 33294 12628 33346
rect 12348 33292 12628 33294
rect 12796 33908 12852 33918
rect 12796 33458 12852 33852
rect 12796 33406 12798 33458
rect 12850 33406 12852 33458
rect 11900 33122 11956 33134
rect 11900 33070 11902 33122
rect 11954 33070 11956 33122
rect 11900 32900 11956 33070
rect 12124 33122 12180 33134
rect 12124 33070 12126 33122
rect 12178 33070 12180 33122
rect 12012 32900 12068 32910
rect 11900 32844 12012 32900
rect 12012 32834 12068 32844
rect 12124 32676 12180 33070
rect 12348 33012 12404 33292
rect 12348 32946 12404 32956
rect 12684 33236 12740 33246
rect 12572 32788 12628 32798
rect 12684 32788 12740 33180
rect 12796 32900 12852 33406
rect 12796 32834 12852 32844
rect 12572 32786 12740 32788
rect 12572 32734 12574 32786
rect 12626 32734 12740 32786
rect 12572 32732 12740 32734
rect 12572 32722 12628 32732
rect 12124 32620 12516 32676
rect 12124 32450 12180 32462
rect 12124 32398 12126 32450
rect 12178 32398 12180 32450
rect 12124 32116 12180 32398
rect 12460 32228 12516 32620
rect 12460 32172 12628 32228
rect 12124 32050 12180 32060
rect 11900 32002 11956 32014
rect 11900 31950 11902 32002
rect 11954 31950 11956 32002
rect 11900 31948 11956 31950
rect 11900 31892 12516 31948
rect 12460 31890 12516 31892
rect 12460 31838 12462 31890
rect 12514 31838 12516 31890
rect 12460 31826 12516 31838
rect 12012 31778 12068 31790
rect 12012 31726 12014 31778
rect 12066 31726 12068 31778
rect 12012 31668 12068 31726
rect 12124 31668 12180 31678
rect 12012 31612 12124 31668
rect 12124 31602 12180 31612
rect 12572 31668 12628 32172
rect 12572 31574 12628 31612
rect 12684 32004 12740 32732
rect 12908 32562 12964 34974
rect 12908 32510 12910 32562
rect 12962 32510 12964 32562
rect 12908 32498 12964 32510
rect 12908 32116 12964 32126
rect 12796 32004 12852 32014
rect 12684 32002 12852 32004
rect 12684 31950 12798 32002
rect 12850 31950 12852 32002
rect 12684 31948 12852 31950
rect 12684 31444 12740 31948
rect 12796 31938 12852 31948
rect 12460 31388 12740 31444
rect 12012 30212 12068 30222
rect 12012 30118 12068 30156
rect 11900 30100 11956 30110
rect 11900 29652 11956 30044
rect 12460 29876 12516 31388
rect 12908 30996 12964 32060
rect 12908 30930 12964 30940
rect 12572 30324 12628 30334
rect 12572 30230 12628 30268
rect 12796 30212 12852 30222
rect 12684 29988 12740 29998
rect 12460 29820 12628 29876
rect 12348 29652 12404 29662
rect 11900 29650 12348 29652
rect 11900 29598 11902 29650
rect 11954 29598 12348 29650
rect 11900 29596 12348 29598
rect 11900 29586 11956 29596
rect 12348 29558 12404 29596
rect 11788 29372 12180 29428
rect 11116 29138 11172 29148
rect 11228 29148 11396 29204
rect 12012 29204 12068 29214
rect 11228 28868 11284 29148
rect 11418 29036 11682 29046
rect 11474 28980 11522 29036
rect 11578 28980 11626 29036
rect 11418 28970 11682 28980
rect 11228 28812 11620 28868
rect 11116 28756 11172 28766
rect 11116 28644 11172 28700
rect 11228 28644 11284 28654
rect 11116 28642 11284 28644
rect 11116 28590 11230 28642
rect 11282 28590 11284 28642
rect 11116 28588 11284 28590
rect 11228 28578 11284 28588
rect 10780 28130 10836 28140
rect 11452 28084 11508 28094
rect 11004 28082 11508 28084
rect 11004 28030 11454 28082
rect 11506 28030 11508 28082
rect 11004 28028 11508 28030
rect 10444 27918 10446 27970
rect 10498 27918 10500 27970
rect 10444 27906 10500 27918
rect 10780 27972 10836 27982
rect 10780 27878 10836 27916
rect 11004 27970 11060 28028
rect 11452 28018 11508 28028
rect 11564 28084 11620 28812
rect 11788 28756 11844 28766
rect 11788 28644 11844 28700
rect 11676 28588 11844 28644
rect 11676 28196 11732 28588
rect 11788 28420 11844 28430
rect 12012 28420 12068 29148
rect 11788 28418 12068 28420
rect 11788 28366 11790 28418
rect 11842 28366 12068 28418
rect 11788 28364 12068 28366
rect 11788 28354 11844 28364
rect 12124 28308 12180 29372
rect 12460 28868 12516 28878
rect 12460 28754 12516 28812
rect 12460 28702 12462 28754
rect 12514 28702 12516 28754
rect 12460 28690 12516 28702
rect 11900 28252 12180 28308
rect 11676 28140 11844 28196
rect 11564 27990 11620 28028
rect 11004 27918 11006 27970
rect 11058 27918 11060 27970
rect 11004 27906 11060 27918
rect 11340 27858 11396 27870
rect 11340 27806 11342 27858
rect 11394 27806 11396 27858
rect 10556 27748 10612 27758
rect 10332 27746 10612 27748
rect 10332 27694 10558 27746
rect 10610 27694 10612 27746
rect 10332 27692 10612 27694
rect 10332 27186 10388 27692
rect 10556 27682 10612 27692
rect 11004 27636 11060 27646
rect 10332 27134 10334 27186
rect 10386 27134 10388 27186
rect 10332 27122 10388 27134
rect 10556 27412 10612 27422
rect 10108 26684 10276 26740
rect 9996 26348 10164 26404
rect 9884 26290 10052 26292
rect 9884 26238 9886 26290
rect 9938 26238 10052 26290
rect 9884 26236 10052 26238
rect 9884 26226 9940 26236
rect 9996 25618 10052 26236
rect 9996 25566 9998 25618
rect 10050 25566 10052 25618
rect 9996 25554 10052 25566
rect 10108 25396 10164 26348
rect 9772 24658 9828 24668
rect 9996 25340 10164 25396
rect 9772 24388 9828 24398
rect 9772 24050 9828 24332
rect 9772 23998 9774 24050
rect 9826 23998 9828 24050
rect 9772 23986 9828 23998
rect 9548 23884 9716 23940
rect 9436 23772 9604 23828
rect 9324 23660 9492 23716
rect 8988 23436 9156 23492
rect 8876 23214 8878 23266
rect 8930 23214 8932 23266
rect 8876 23202 8932 23214
rect 8988 23042 9044 23054
rect 8988 22990 8990 23042
rect 9042 22990 9044 23042
rect 8876 22596 8932 22606
rect 8988 22596 9044 22990
rect 8932 22540 9044 22596
rect 8876 22482 8932 22540
rect 9100 22484 9156 23436
rect 8876 22430 8878 22482
rect 8930 22430 8932 22482
rect 8876 22418 8932 22430
rect 8988 22428 9156 22484
rect 8876 20244 8932 20254
rect 8876 20130 8932 20188
rect 8876 20078 8878 20130
rect 8930 20078 8932 20130
rect 8876 20066 8932 20078
rect 8988 19908 9044 22428
rect 9100 21028 9156 21038
rect 9100 20914 9156 20972
rect 9100 20862 9102 20914
rect 9154 20862 9156 20914
rect 9100 20850 9156 20862
rect 9100 19908 9156 19918
rect 8988 19852 9100 19908
rect 8652 19346 9044 19348
rect 8652 19294 8654 19346
rect 8706 19294 9044 19346
rect 8652 19292 9044 19294
rect 8652 19282 8708 19292
rect 7812 19180 7924 19236
rect 7756 19142 7812 19180
rect 6972 19122 7028 19134
rect 6972 19070 6974 19122
rect 7026 19070 7028 19122
rect 6972 19012 7028 19070
rect 6972 18946 7028 18956
rect 7532 19010 7588 19022
rect 7532 18958 7534 19010
rect 7586 18958 7588 19010
rect 7532 18452 7588 18958
rect 7644 19012 7700 19022
rect 7644 18918 7700 18956
rect 7868 18676 7924 19180
rect 8204 19234 8372 19236
rect 8204 19182 8206 19234
rect 8258 19182 8372 19234
rect 8204 19180 8372 19182
rect 8204 19170 8260 19180
rect 8316 19012 8372 19180
rect 8540 19170 8596 19180
rect 8988 19234 9044 19292
rect 8988 19182 8990 19234
rect 9042 19182 9044 19234
rect 8316 18956 8484 19012
rect 8016 18844 8280 18854
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8016 18778 8280 18788
rect 7868 18620 8148 18676
rect 7420 17108 7476 17118
rect 7532 17108 7588 18396
rect 8092 18338 8148 18620
rect 8092 18286 8094 18338
rect 8146 18286 8148 18338
rect 8092 18274 8148 18286
rect 7868 18116 7924 18126
rect 7644 17108 7700 17118
rect 7532 17106 7700 17108
rect 7532 17054 7646 17106
rect 7698 17054 7700 17106
rect 7532 17052 7700 17054
rect 6972 16996 7028 17006
rect 7196 16996 7252 17006
rect 6972 16994 7196 16996
rect 6972 16942 6974 16994
rect 7026 16942 7196 16994
rect 6972 16940 7196 16942
rect 7420 16996 7476 17052
rect 7420 16940 7588 16996
rect 6972 16930 7028 16940
rect 7196 16930 7252 16940
rect 6860 15484 7028 15540
rect 6860 15314 6916 15326
rect 6860 15262 6862 15314
rect 6914 15262 6916 15314
rect 6860 15204 6916 15262
rect 6860 15138 6916 15148
rect 6972 15092 7028 15484
rect 7084 15428 7140 15438
rect 7420 15428 7476 15438
rect 7140 15372 7364 15428
rect 7084 15362 7140 15372
rect 7308 15148 7364 15372
rect 7420 15334 7476 15372
rect 7420 15204 7476 15214
rect 7308 15092 7476 15148
rect 6972 15036 7252 15092
rect 6636 14478 6638 14530
rect 6690 14478 6692 14530
rect 6636 12738 6692 14478
rect 6972 13412 7028 13422
rect 6972 12962 7028 13356
rect 6972 12910 6974 12962
rect 7026 12910 7028 12962
rect 6972 12898 7028 12910
rect 7196 12962 7252 15036
rect 7308 14420 7364 14430
rect 7308 14326 7364 14364
rect 7420 13634 7476 15092
rect 7420 13582 7422 13634
rect 7474 13582 7476 13634
rect 7420 13570 7476 13582
rect 7196 12910 7198 12962
rect 7250 12910 7252 12962
rect 7084 12852 7140 12862
rect 7084 12758 7140 12796
rect 6636 12686 6638 12738
rect 6690 12686 6692 12738
rect 6636 11508 6692 12686
rect 7196 12068 7252 12910
rect 7420 12740 7476 12750
rect 7308 12068 7364 12078
rect 7196 12012 7308 12068
rect 7308 11974 7364 12012
rect 6076 11330 6132 11340
rect 6188 11452 6692 11508
rect 6748 11508 6804 11518
rect 5964 11172 6020 11182
rect 6188 11172 6244 11452
rect 6748 11396 6804 11452
rect 7196 11508 7252 11518
rect 7420 11508 7476 12684
rect 7196 11506 7476 11508
rect 7196 11454 7198 11506
rect 7250 11454 7476 11506
rect 7196 11452 7476 11454
rect 7196 11442 7252 11452
rect 7532 11396 7588 16940
rect 7644 15540 7700 17052
rect 7868 17106 7924 18060
rect 8428 17444 8484 18956
rect 8988 18674 9044 19182
rect 8988 18622 8990 18674
rect 9042 18622 9044 18674
rect 8540 18452 8596 18462
rect 8540 18358 8596 18396
rect 8540 18116 8596 18126
rect 8540 17778 8596 18060
rect 8988 17780 9044 18622
rect 9100 18340 9156 19852
rect 9100 18274 9156 18284
rect 9212 18116 9268 23660
rect 8540 17726 8542 17778
rect 8594 17726 8596 17778
rect 8540 17714 8596 17726
rect 8876 17724 8988 17780
rect 8016 17276 8280 17286
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8016 17210 8280 17220
rect 7868 17054 7870 17106
rect 7922 17054 7924 17106
rect 7868 17042 7924 17054
rect 8204 17108 8260 17118
rect 7756 16996 7812 17006
rect 7756 16902 7812 16940
rect 8204 16098 8260 17052
rect 8204 16046 8206 16098
rect 8258 16046 8260 16098
rect 8204 16034 8260 16046
rect 8316 16884 8372 16894
rect 8428 16884 8484 17388
rect 8316 16882 8484 16884
rect 8316 16830 8318 16882
rect 8370 16830 8484 16882
rect 8316 16828 8484 16830
rect 8316 15876 8372 16828
rect 8876 16210 8932 17724
rect 8988 17686 9044 17724
rect 9100 18060 9212 18116
rect 8988 17108 9044 17118
rect 9100 17108 9156 18060
rect 9212 18050 9268 18060
rect 9324 23492 9380 23502
rect 8988 17106 9156 17108
rect 8988 17054 8990 17106
rect 9042 17054 9156 17106
rect 8988 17052 9156 17054
rect 8988 17042 9044 17052
rect 8876 16158 8878 16210
rect 8930 16158 8932 16210
rect 8316 15820 8484 15876
rect 8016 15708 8280 15718
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8016 15642 8280 15652
rect 7756 15540 7812 15550
rect 8428 15540 8484 15820
rect 7644 15484 7756 15540
rect 7756 15446 7812 15484
rect 8316 15484 8484 15540
rect 8540 15540 8596 15550
rect 8876 15540 8932 16158
rect 8988 15540 9044 15550
rect 8876 15538 9044 15540
rect 8876 15486 8990 15538
rect 9042 15486 9044 15538
rect 8876 15484 9044 15486
rect 7868 15316 7924 15326
rect 7868 15202 7924 15260
rect 7868 15150 7870 15202
rect 7922 15150 7924 15202
rect 7868 15138 7924 15150
rect 7980 15314 8036 15326
rect 7980 15262 7982 15314
rect 8034 15262 8036 15314
rect 7980 15204 8036 15262
rect 8316 15314 8372 15484
rect 8316 15262 8318 15314
rect 8370 15262 8372 15314
rect 8316 15250 8372 15262
rect 7980 15138 8036 15148
rect 8540 15148 8596 15484
rect 8988 15474 9044 15484
rect 9324 15148 9380 23436
rect 9436 20916 9492 23660
rect 9436 20850 9492 20860
rect 9436 20692 9492 20702
rect 9436 20598 9492 20636
rect 9436 17444 9492 17454
rect 9436 17350 9492 17388
rect 9548 16884 9604 23772
rect 9660 22596 9716 23884
rect 9660 22530 9716 22540
rect 9996 22036 10052 25340
rect 10108 24164 10164 24174
rect 10108 23938 10164 24108
rect 10108 23886 10110 23938
rect 10162 23886 10164 23938
rect 10108 23874 10164 23886
rect 10220 22708 10276 26684
rect 10332 26178 10388 26190
rect 10332 26126 10334 26178
rect 10386 26126 10388 26178
rect 10332 26068 10388 26126
rect 10332 26002 10388 26012
rect 10444 25284 10500 25294
rect 10444 25190 10500 25228
rect 10332 24610 10388 24622
rect 10332 24558 10334 24610
rect 10386 24558 10388 24610
rect 10332 23714 10388 24558
rect 10444 24388 10500 24398
rect 10444 23938 10500 24332
rect 10444 23886 10446 23938
rect 10498 23886 10500 23938
rect 10444 23874 10500 23886
rect 10332 23662 10334 23714
rect 10386 23662 10388 23714
rect 10332 23650 10388 23662
rect 10220 22652 10500 22708
rect 10108 22596 10164 22606
rect 10164 22540 10276 22596
rect 10108 22530 10164 22540
rect 10220 22482 10276 22540
rect 10220 22430 10222 22482
rect 10274 22430 10276 22482
rect 10220 22418 10276 22430
rect 10444 22258 10500 22652
rect 10444 22206 10446 22258
rect 10498 22206 10500 22258
rect 9884 21980 10052 22036
rect 10332 22146 10388 22158
rect 10332 22094 10334 22146
rect 10386 22094 10388 22146
rect 9660 21812 9716 21822
rect 9660 21586 9716 21756
rect 9884 21700 9940 21980
rect 10332 21924 10388 22094
rect 9884 21634 9940 21644
rect 9996 21868 10388 21924
rect 9660 21534 9662 21586
rect 9714 21534 9716 21586
rect 9660 21522 9716 21534
rect 9996 21026 10052 21868
rect 9996 20974 9998 21026
rect 10050 20974 10052 21026
rect 9996 20962 10052 20974
rect 10332 21474 10388 21486
rect 10332 21422 10334 21474
rect 10386 21422 10388 21474
rect 10220 20916 10276 20926
rect 9772 20804 9828 20842
rect 10220 20804 10276 20860
rect 9828 20748 9940 20804
rect 9772 20738 9828 20748
rect 9772 20580 9828 20590
rect 9772 19346 9828 20524
rect 9772 19294 9774 19346
rect 9826 19294 9828 19346
rect 9772 19282 9828 19294
rect 9660 18452 9716 18462
rect 9660 17106 9716 18396
rect 9660 17054 9662 17106
rect 9714 17054 9716 17106
rect 9660 17042 9716 17054
rect 9884 16996 9940 20748
rect 9996 20802 10276 20804
rect 9996 20750 10222 20802
rect 10274 20750 10276 20802
rect 9996 20748 10276 20750
rect 9996 20244 10052 20748
rect 10220 20738 10276 20748
rect 10220 20580 10276 20590
rect 10332 20580 10388 21422
rect 10444 21476 10500 22206
rect 10444 21410 10500 21420
rect 10556 21140 10612 27356
rect 10780 26292 10836 26302
rect 10780 26198 10836 26236
rect 10780 25956 10836 25966
rect 10780 24164 10836 25900
rect 10668 23828 10724 23838
rect 10668 23734 10724 23772
rect 10780 23380 10836 24108
rect 10892 23380 10948 23390
rect 10780 23378 10948 23380
rect 10780 23326 10894 23378
rect 10946 23326 10948 23378
rect 10780 23324 10948 23326
rect 10892 23314 10948 23324
rect 11004 22820 11060 27580
rect 11340 27636 11396 27806
rect 11340 27570 11396 27580
rect 11418 27468 11682 27478
rect 11474 27412 11522 27468
rect 11578 27412 11626 27468
rect 11418 27402 11682 27412
rect 10556 21074 10612 21084
rect 10892 22764 11060 22820
rect 11116 26292 11172 26302
rect 10780 21028 10836 21038
rect 10780 20802 10836 20972
rect 10780 20750 10782 20802
rect 10834 20750 10836 20802
rect 10220 20578 10388 20580
rect 10220 20526 10222 20578
rect 10274 20526 10388 20578
rect 10220 20524 10388 20526
rect 10556 20692 10612 20702
rect 10220 20514 10276 20524
rect 9996 20130 10052 20188
rect 10444 20244 10500 20254
rect 10556 20244 10612 20636
rect 10668 20580 10724 20590
rect 10668 20486 10724 20524
rect 10780 20356 10836 20750
rect 10444 20242 10556 20244
rect 10444 20190 10446 20242
rect 10498 20190 10556 20242
rect 10444 20188 10556 20190
rect 10444 20178 10500 20188
rect 10556 20178 10612 20188
rect 10668 20300 10836 20356
rect 9996 20078 9998 20130
rect 10050 20078 10052 20130
rect 9996 20066 10052 20078
rect 10108 18564 10164 18574
rect 10108 17778 10164 18508
rect 10108 17726 10110 17778
rect 10162 17726 10164 17778
rect 10108 17714 10164 17726
rect 10332 18340 10388 18350
rect 10220 17444 10276 17454
rect 9884 16940 10164 16996
rect 9548 16828 9940 16884
rect 9772 16324 9828 16334
rect 9660 15316 9716 15326
rect 9772 15316 9828 16268
rect 9660 15314 9828 15316
rect 9660 15262 9662 15314
rect 9714 15262 9828 15314
rect 9660 15260 9828 15262
rect 9660 15250 9716 15260
rect 8540 15092 8708 15148
rect 9324 15092 9492 15148
rect 8540 14420 8596 14430
rect 8016 14140 8280 14150
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8016 14074 8280 14084
rect 8540 13970 8596 14364
rect 8540 13918 8542 13970
rect 8594 13918 8596 13970
rect 8540 13906 8596 13918
rect 8316 13860 8372 13870
rect 8092 13748 8148 13758
rect 8092 13654 8148 13692
rect 8316 13746 8372 13804
rect 8316 13694 8318 13746
rect 8370 13694 8372 13746
rect 7644 13412 7700 13422
rect 7644 11506 7700 13356
rect 8092 13076 8148 13086
rect 8316 13076 8372 13694
rect 8652 13412 8708 15092
rect 8652 13346 8708 13356
rect 8764 14644 8820 14654
rect 8764 13858 8820 14588
rect 9436 14642 9492 15092
rect 9436 14590 9438 14642
rect 9490 14590 9492 14642
rect 9436 14196 9492 14590
rect 9772 14532 9828 15260
rect 9884 14756 9940 16828
rect 10108 16548 10164 16940
rect 9884 14690 9940 14700
rect 9996 16492 10164 16548
rect 10220 16884 10276 17388
rect 10332 17108 10388 18284
rect 10444 17892 10500 17902
rect 10444 17666 10500 17836
rect 10444 17614 10446 17666
rect 10498 17614 10500 17666
rect 10444 17602 10500 17614
rect 10332 17014 10388 17052
rect 10556 17442 10612 17454
rect 10556 17390 10558 17442
rect 10610 17390 10612 17442
rect 9884 14532 9940 14542
rect 9772 14530 9940 14532
rect 9772 14478 9886 14530
rect 9938 14478 9940 14530
rect 9772 14476 9940 14478
rect 9436 14140 9828 14196
rect 9660 13972 9716 13982
rect 8764 13806 8766 13858
rect 8818 13806 8820 13858
rect 8148 13020 8372 13076
rect 8092 12982 8148 13020
rect 8540 12740 8596 12750
rect 8540 12646 8596 12684
rect 8016 12572 8280 12582
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8764 12516 8820 13806
rect 8988 13970 9716 13972
rect 8988 13918 9662 13970
rect 9714 13918 9716 13970
rect 8988 13916 9716 13918
rect 8988 13858 9044 13916
rect 9660 13906 9716 13916
rect 8988 13806 8990 13858
rect 9042 13806 9044 13858
rect 8988 13794 9044 13806
rect 9548 13746 9604 13758
rect 9548 13694 9550 13746
rect 9602 13694 9604 13746
rect 9548 13412 9604 13694
rect 9772 13746 9828 14140
rect 9884 13972 9940 14476
rect 9884 13906 9940 13916
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9772 13524 9828 13694
rect 9996 13636 10052 16492
rect 10220 16100 10276 16828
rect 9996 13570 10052 13580
rect 10108 13748 10164 13758
rect 10220 13748 10276 16044
rect 10332 15428 10388 15438
rect 10556 15428 10612 17390
rect 10332 15426 10612 15428
rect 10332 15374 10334 15426
rect 10386 15374 10612 15426
rect 10332 15372 10612 15374
rect 10332 15362 10388 15372
rect 10668 15148 10724 20300
rect 10780 20020 10836 20030
rect 10780 18564 10836 19964
rect 10780 17666 10836 18508
rect 10780 17614 10782 17666
rect 10834 17614 10836 17666
rect 10780 17602 10836 17614
rect 10892 17444 10948 22764
rect 11004 22596 11060 22606
rect 11004 22482 11060 22540
rect 11004 22430 11006 22482
rect 11058 22430 11060 22482
rect 11004 22418 11060 22430
rect 11004 21028 11060 21038
rect 11004 20934 11060 20972
rect 11116 19460 11172 26236
rect 11418 25900 11682 25910
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11418 25834 11682 25844
rect 11788 24948 11844 28140
rect 11900 26908 11956 28252
rect 12572 28196 12628 29820
rect 12572 28130 12628 28140
rect 12460 28084 12516 28094
rect 12012 27858 12068 27870
rect 12012 27806 12014 27858
rect 12066 27806 12068 27858
rect 12012 27748 12068 27806
rect 12348 27748 12404 27758
rect 12012 27746 12404 27748
rect 12012 27694 12350 27746
rect 12402 27694 12404 27746
rect 12012 27692 12404 27694
rect 12348 27636 12404 27692
rect 12348 27570 12404 27580
rect 12460 27186 12516 28028
rect 12460 27134 12462 27186
rect 12514 27134 12516 27186
rect 12460 27122 12516 27134
rect 12684 26908 12740 29932
rect 12796 29426 12852 30156
rect 12908 29988 12964 29998
rect 12908 29894 12964 29932
rect 12796 29374 12798 29426
rect 12850 29374 12852 29426
rect 12796 28196 12852 29374
rect 12908 28756 12964 28766
rect 12908 28662 12964 28700
rect 12796 28140 12964 28196
rect 12796 27746 12852 27758
rect 12796 27694 12798 27746
rect 12850 27694 12852 27746
rect 12796 27524 12852 27694
rect 12796 27458 12852 27468
rect 12908 27186 12964 28140
rect 12908 27134 12910 27186
rect 12962 27134 12964 27186
rect 12908 27076 12964 27134
rect 12908 27010 12964 27020
rect 11900 26852 12180 26908
rect 12124 26404 12180 26852
rect 12012 26348 12180 26404
rect 12348 26852 12740 26908
rect 11788 24882 11844 24892
rect 11900 25284 11956 25294
rect 11418 24332 11682 24342
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11418 24266 11682 24276
rect 11564 24052 11620 24062
rect 11228 23940 11284 23950
rect 11228 23846 11284 23884
rect 11564 23938 11620 23996
rect 11564 23886 11566 23938
rect 11618 23886 11620 23938
rect 11564 23716 11620 23886
rect 11788 23940 11844 23950
rect 11900 23940 11956 25228
rect 11788 23938 11956 23940
rect 11788 23886 11790 23938
rect 11842 23886 11956 23938
rect 11788 23884 11956 23886
rect 12012 23940 12068 26348
rect 11788 23874 11844 23884
rect 11676 23828 11732 23838
rect 12012 23828 12068 23884
rect 11676 23734 11732 23772
rect 11900 23826 12068 23828
rect 11900 23774 12014 23826
rect 12066 23774 12068 23826
rect 11900 23772 12068 23774
rect 11564 23650 11620 23660
rect 11900 23268 11956 23772
rect 12012 23762 12068 23772
rect 12124 26180 12180 26190
rect 11788 23212 11956 23268
rect 11418 22764 11682 22774
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11418 22698 11682 22708
rect 11788 22372 11844 23212
rect 11788 22306 11844 22316
rect 11900 23042 11956 23054
rect 11900 22990 11902 23042
rect 11954 22990 11956 23042
rect 11900 22932 11956 22990
rect 11418 21196 11682 21206
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11418 21130 11682 21140
rect 11676 21028 11732 21038
rect 11676 20934 11732 20972
rect 11340 20916 11396 20926
rect 11340 20802 11396 20860
rect 11340 20750 11342 20802
rect 11394 20750 11396 20802
rect 11340 20738 11396 20750
rect 11788 20804 11844 20814
rect 11788 20692 11844 20748
rect 11676 20690 11844 20692
rect 11676 20638 11790 20690
rect 11842 20638 11844 20690
rect 11676 20636 11844 20638
rect 11452 20244 11508 20254
rect 11452 20150 11508 20188
rect 11676 20242 11732 20636
rect 11788 20626 11844 20636
rect 11900 20356 11956 22876
rect 11676 20190 11678 20242
rect 11730 20190 11732 20242
rect 11676 20178 11732 20190
rect 11788 20300 11956 20356
rect 12012 22596 12068 22606
rect 12012 21026 12068 22540
rect 12012 20974 12014 21026
rect 12066 20974 12068 21026
rect 11418 19628 11682 19638
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11418 19562 11682 19572
rect 11116 19404 11620 19460
rect 11564 18452 11620 19404
rect 11564 18358 11620 18396
rect 11228 18338 11284 18350
rect 11228 18286 11230 18338
rect 11282 18286 11284 18338
rect 11228 17892 11284 18286
rect 11418 18060 11682 18070
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11418 17994 11682 18004
rect 11228 17826 11284 17836
rect 11004 17668 11060 17678
rect 11564 17668 11620 17678
rect 11004 17666 11620 17668
rect 11004 17614 11006 17666
rect 11058 17614 11566 17666
rect 11618 17614 11620 17666
rect 11004 17612 11620 17614
rect 11004 17602 11060 17612
rect 11564 17602 11620 17612
rect 11676 17668 11732 17678
rect 11676 17574 11732 17612
rect 10892 17388 11284 17444
rect 11228 17106 11284 17388
rect 11228 17054 11230 17106
rect 11282 17054 11284 17106
rect 10780 16884 10836 16894
rect 10780 16790 10836 16828
rect 11116 15876 11172 15886
rect 10668 15092 10836 15148
rect 10556 14418 10612 14430
rect 10556 14366 10558 14418
rect 10610 14366 10612 14418
rect 10556 13972 10612 14366
rect 10668 13972 10724 13982
rect 10556 13970 10724 13972
rect 10556 13918 10670 13970
rect 10722 13918 10724 13970
rect 10556 13916 10724 13918
rect 10668 13906 10724 13916
rect 10444 13860 10500 13870
rect 10444 13748 10500 13804
rect 10108 13746 10276 13748
rect 10108 13694 10110 13746
rect 10162 13694 10276 13746
rect 10108 13692 10276 13694
rect 10332 13746 10500 13748
rect 10332 13694 10446 13746
rect 10498 13694 10500 13746
rect 10332 13692 10500 13694
rect 9772 13458 9828 13468
rect 9324 12740 9380 12750
rect 9324 12646 9380 12684
rect 9548 12740 9604 13356
rect 9884 13412 9940 13422
rect 9660 12740 9716 12750
rect 9548 12738 9716 12740
rect 9548 12686 9662 12738
rect 9714 12686 9716 12738
rect 9548 12684 9716 12686
rect 8016 12506 8280 12516
rect 8428 12460 8820 12516
rect 8204 12404 8260 12414
rect 8428 12404 8484 12460
rect 8204 12402 8484 12404
rect 8204 12350 8206 12402
rect 8258 12350 8484 12402
rect 8204 12348 8484 12350
rect 7644 11454 7646 11506
rect 7698 11454 7700 11506
rect 7644 11442 7700 11454
rect 7868 11508 7924 11518
rect 7868 11414 7924 11452
rect 6524 11340 6804 11396
rect 6300 11284 6356 11294
rect 6300 11190 6356 11228
rect 6524 11282 6580 11340
rect 6524 11230 6526 11282
rect 6578 11230 6580 11282
rect 6524 11218 6580 11230
rect 5292 11170 6244 11172
rect 5292 11118 5966 11170
rect 6018 11118 6244 11170
rect 5292 11116 6244 11118
rect 6412 11170 6468 11182
rect 6412 11118 6414 11170
rect 6466 11118 6468 11170
rect 5964 9828 6020 11116
rect 6300 10388 6356 10398
rect 5964 9826 6244 9828
rect 5964 9774 5966 9826
rect 6018 9774 6244 9826
rect 5964 9772 6244 9774
rect 5964 9762 6020 9772
rect 5068 9602 5236 9604
rect 5068 9550 5070 9602
rect 5122 9550 5236 9602
rect 5068 9548 5236 9550
rect 5068 9538 5124 9548
rect 4508 9102 4510 9154
rect 4562 9102 4564 9154
rect 4508 9090 4564 9102
rect 4396 8990 4398 9042
rect 4450 8990 4452 9042
rect 4396 8978 4452 8990
rect 4614 8652 4878 8662
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4614 8586 4878 8596
rect 4732 8372 4788 8382
rect 4732 7474 4788 8316
rect 5068 8370 5124 8382
rect 5068 8318 5070 8370
rect 5122 8318 5124 8370
rect 5068 8036 5124 8318
rect 5068 7970 5124 7980
rect 5180 7924 5236 9548
rect 6076 9044 6132 9054
rect 5964 9042 6132 9044
rect 5964 8990 6078 9042
rect 6130 8990 6132 9042
rect 5964 8988 6132 8990
rect 5516 8930 5572 8942
rect 5516 8878 5518 8930
rect 5570 8878 5572 8930
rect 5516 8484 5572 8878
rect 5516 8418 5572 8428
rect 5180 7858 5236 7868
rect 5404 8036 5460 8046
rect 5068 7700 5124 7710
rect 5068 7606 5124 7644
rect 4732 7422 4734 7474
rect 4786 7422 4788 7474
rect 4732 7410 4788 7422
rect 5180 7474 5236 7486
rect 5180 7422 5182 7474
rect 5234 7422 5236 7474
rect 4956 7252 5012 7262
rect 4284 7250 5012 7252
rect 4284 7198 4958 7250
rect 5010 7198 5012 7250
rect 4284 7196 5012 7198
rect 4956 7186 5012 7196
rect 4614 7084 4878 7094
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4614 7018 4878 7028
rect 5180 6804 5236 7422
rect 4844 6748 5236 6804
rect 4732 6692 4788 6702
rect 4732 6598 4788 6636
rect 4844 6690 4900 6748
rect 5404 6692 5460 7980
rect 5516 7588 5572 7598
rect 5964 7588 6020 8988
rect 6076 8978 6132 8988
rect 6076 8034 6132 8046
rect 6076 7982 6078 8034
rect 6130 7982 6132 8034
rect 6076 7924 6132 7982
rect 6076 7858 6132 7868
rect 5572 7532 6020 7588
rect 6188 7700 6244 9772
rect 6300 9154 6356 10332
rect 6300 9102 6302 9154
rect 6354 9102 6356 9154
rect 6300 9090 6356 9102
rect 6412 9044 6468 11118
rect 6636 11172 6692 11182
rect 6636 9940 6692 11116
rect 6748 10612 6804 11340
rect 6748 10546 6804 10556
rect 7308 11340 7588 11396
rect 7308 10612 7364 11340
rect 8204 11172 8260 12348
rect 9548 12292 9604 12684
rect 9660 12674 9716 12684
rect 9772 12738 9828 12750
rect 9772 12686 9774 12738
rect 9826 12686 9828 12738
rect 9772 12404 9828 12686
rect 9548 12226 9604 12236
rect 9660 12348 9828 12404
rect 9884 12740 9940 13356
rect 10108 12852 10164 13692
rect 10108 12758 10164 12796
rect 10332 13076 10388 13692
rect 10444 13682 10500 13692
rect 10780 13748 10836 15092
rect 11116 13858 11172 15820
rect 11228 15764 11284 17054
rect 11452 17442 11508 17454
rect 11452 17390 11454 17442
rect 11506 17390 11508 17442
rect 11452 17108 11508 17390
rect 11676 17108 11732 17118
rect 11452 17052 11676 17108
rect 11676 17014 11732 17052
rect 11418 16492 11682 16502
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11418 16426 11682 16436
rect 11228 15698 11284 15708
rect 11418 14924 11682 14934
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11418 14858 11682 14868
rect 11564 13972 11620 13982
rect 11564 13878 11620 13916
rect 11116 13806 11118 13858
rect 11170 13806 11172 13858
rect 11116 13794 11172 13806
rect 8988 12180 9044 12190
rect 8652 12124 8988 12180
rect 8540 12068 8596 12078
rect 8540 11974 8596 12012
rect 7868 11116 8260 11172
rect 7756 10724 7812 10734
rect 7756 10630 7812 10668
rect 7308 10610 7588 10612
rect 7308 10558 7310 10610
rect 7362 10558 7588 10610
rect 7308 10556 7588 10558
rect 7308 10546 7364 10556
rect 6636 9874 6692 9884
rect 6636 9714 6692 9726
rect 6636 9662 6638 9714
rect 6690 9662 6692 9714
rect 6524 9268 6580 9278
rect 6636 9268 6692 9662
rect 6524 9266 6692 9268
rect 6524 9214 6526 9266
rect 6578 9214 6692 9266
rect 6524 9212 6692 9214
rect 7532 9266 7588 10556
rect 7644 10388 7700 10398
rect 7644 10294 7700 10332
rect 7532 9214 7534 9266
rect 7586 9214 7588 9266
rect 6524 9202 6580 9212
rect 7532 9202 7588 9214
rect 7868 9266 7924 11116
rect 8016 11004 8280 11014
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8016 10938 8280 10948
rect 8652 10834 8708 12124
rect 8988 12086 9044 12124
rect 9660 12178 9716 12348
rect 9660 12126 9662 12178
rect 9714 12126 9716 12178
rect 9660 12114 9716 12126
rect 9772 12180 9828 12190
rect 9772 12086 9828 12124
rect 8652 10782 8654 10834
rect 8706 10782 8708 10834
rect 8652 10770 8708 10782
rect 8764 11620 8820 11630
rect 8764 10724 8820 11564
rect 9884 11508 9940 12684
rect 10220 12180 10276 12190
rect 10332 12180 10388 13020
rect 10556 12292 10612 12302
rect 10556 12198 10612 12236
rect 10220 12178 10388 12180
rect 10220 12126 10222 12178
rect 10274 12126 10388 12178
rect 10220 12124 10388 12126
rect 10220 12114 10276 12124
rect 9884 11442 9940 11452
rect 9996 12066 10052 12078
rect 9996 12014 9998 12066
rect 10050 12014 10052 12066
rect 9996 11506 10052 12014
rect 9996 11454 9998 11506
rect 10050 11454 10052 11506
rect 9996 11442 10052 11454
rect 10108 11508 10164 11518
rect 8092 10612 8148 10622
rect 8092 10518 8148 10556
rect 8764 9940 8820 10668
rect 9212 11284 9268 11294
rect 8764 9938 8932 9940
rect 8764 9886 8766 9938
rect 8818 9886 8932 9938
rect 8764 9884 8932 9886
rect 8764 9874 8820 9884
rect 8016 9436 8280 9446
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8016 9370 8280 9380
rect 7868 9214 7870 9266
rect 7922 9214 7924 9266
rect 7868 9202 7924 9214
rect 8876 9266 8932 9884
rect 8876 9214 8878 9266
rect 8930 9214 8932 9266
rect 8876 9202 8932 9214
rect 9212 9602 9268 11228
rect 10108 11172 10164 11452
rect 10668 11394 10724 11406
rect 10668 11342 10670 11394
rect 10722 11342 10724 11394
rect 10668 11284 10724 11342
rect 10668 11218 10724 11228
rect 10108 11106 10164 11116
rect 10444 11060 10500 11070
rect 9884 10836 9940 10846
rect 9884 10742 9940 10780
rect 10220 10612 10276 10622
rect 10444 10612 10500 11004
rect 10220 10610 10500 10612
rect 10220 10558 10222 10610
rect 10274 10558 10446 10610
rect 10498 10558 10500 10610
rect 10220 10556 10500 10558
rect 10220 10546 10276 10556
rect 10444 10546 10500 10556
rect 10780 10836 10836 13692
rect 10892 13524 10948 13534
rect 10892 13074 10948 13468
rect 11418 13356 11682 13366
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11418 13290 11682 13300
rect 10892 13022 10894 13074
rect 10946 13022 10948 13074
rect 10892 13010 10948 13022
rect 11340 13076 11396 13086
rect 11340 12982 11396 13020
rect 11788 12964 11844 20300
rect 11900 20132 11956 20142
rect 12012 20132 12068 20974
rect 11900 20130 12068 20132
rect 11900 20078 11902 20130
rect 11954 20078 12068 20130
rect 11900 20076 12068 20078
rect 11900 20066 11956 20076
rect 11900 19794 11956 19806
rect 11900 19742 11902 19794
rect 11954 19742 11956 19794
rect 11900 19346 11956 19742
rect 11900 19294 11902 19346
rect 11954 19294 11956 19346
rect 11900 19282 11956 19294
rect 12124 19124 12180 26124
rect 12348 24836 12404 26852
rect 13020 26740 13076 41020
rect 13132 27412 13188 41468
rect 13244 41188 13300 41198
rect 13244 40626 13300 41132
rect 13244 40574 13246 40626
rect 13298 40574 13300 40626
rect 13244 40562 13300 40574
rect 13356 38668 13412 52332
rect 13468 51378 13524 51390
rect 13468 51326 13470 51378
rect 13522 51326 13524 51378
rect 13468 50708 13524 51326
rect 13468 50642 13524 50652
rect 13580 51156 13636 51166
rect 13580 50596 13636 51100
rect 13580 50530 13636 50540
rect 13468 50260 13524 50270
rect 13468 49700 13524 50204
rect 13580 49924 13636 49934
rect 13692 49924 13748 52668
rect 13916 51044 13972 53788
rect 13916 50978 13972 50988
rect 14028 52162 14084 55022
rect 14140 54404 14196 55468
rect 14140 54338 14196 54348
rect 14252 55410 14308 55422
rect 14252 55358 14254 55410
rect 14306 55358 14308 55410
rect 14140 52276 14196 52286
rect 14140 52182 14196 52220
rect 14028 52110 14030 52162
rect 14082 52110 14084 52162
rect 13580 49922 13748 49924
rect 13580 49870 13582 49922
rect 13634 49870 13748 49922
rect 13580 49868 13748 49870
rect 13580 49858 13636 49868
rect 13468 49644 13636 49700
rect 13468 49476 13524 49486
rect 13468 45332 13524 49420
rect 13580 49250 13636 49644
rect 13580 49198 13582 49250
rect 13634 49198 13636 49250
rect 13580 49186 13636 49198
rect 13468 45266 13524 45276
rect 13580 47234 13636 47246
rect 13580 47182 13582 47234
rect 13634 47182 13636 47234
rect 13468 45108 13524 45118
rect 13468 45014 13524 45052
rect 13468 44660 13524 44670
rect 13468 44322 13524 44604
rect 13580 44548 13636 47182
rect 13692 45668 13748 49868
rect 14028 49924 14084 52110
rect 14252 52052 14308 55358
rect 14364 55298 14420 55310
rect 14364 55246 14366 55298
rect 14418 55246 14420 55298
rect 14364 55076 14420 55246
rect 14476 55300 14532 55804
rect 14476 55234 14532 55244
rect 14364 55010 14420 55020
rect 14364 53508 14420 53546
rect 14364 53442 14420 53452
rect 14028 49858 14084 49868
rect 14140 51996 14308 52052
rect 14140 49476 14196 51996
rect 14140 49410 14196 49420
rect 14252 50596 14308 50606
rect 14252 49252 14308 50540
rect 14028 49196 14308 49252
rect 13916 49028 13972 49038
rect 13804 48916 13860 48926
rect 13804 48020 13860 48860
rect 13804 46900 13860 47964
rect 13916 47458 13972 48972
rect 14028 48804 14084 49196
rect 14588 49140 14644 56028
rect 14812 56018 14868 56028
rect 15372 55188 15428 56252
rect 15596 56196 15652 56206
rect 15708 56196 15764 58942
rect 15596 56194 15764 56196
rect 15596 56142 15598 56194
rect 15650 56142 15764 56194
rect 15596 56140 15764 56142
rect 15820 58996 15876 59006
rect 15596 56130 15652 56140
rect 15484 56084 15540 56094
rect 15820 56084 15876 58940
rect 15932 58772 15988 60060
rect 16380 60004 16436 60014
rect 15932 58706 15988 58716
rect 16044 60002 16436 60004
rect 16044 59950 16382 60002
rect 16434 59950 16436 60002
rect 16044 59948 16436 59950
rect 15484 55990 15540 56028
rect 15708 56028 15876 56084
rect 15932 56868 15988 56878
rect 15372 55122 15428 55132
rect 14820 54908 15084 54918
rect 14876 54852 14924 54908
rect 14980 54852 15028 54908
rect 14820 54842 15084 54852
rect 15372 54740 15428 54750
rect 15708 54740 15764 56028
rect 15932 55300 15988 56812
rect 15932 55234 15988 55244
rect 15372 54738 15764 54740
rect 15372 54686 15374 54738
rect 15426 54686 15764 54738
rect 15372 54684 15764 54686
rect 15372 54674 15428 54684
rect 15260 54514 15316 54526
rect 15260 54462 15262 54514
rect 15314 54462 15316 54514
rect 15036 54402 15092 54414
rect 15036 54350 15038 54402
rect 15090 54350 15092 54402
rect 14924 53732 14980 53742
rect 14700 53508 14756 53518
rect 14700 52948 14756 53452
rect 14924 53508 14980 53676
rect 15036 53620 15092 54350
rect 15036 53554 15092 53564
rect 15260 53618 15316 54462
rect 15260 53566 15262 53618
rect 15314 53566 15316 53618
rect 14924 53442 14980 53452
rect 14820 53340 15084 53350
rect 14876 53284 14924 53340
rect 14980 53284 15028 53340
rect 14820 53274 15084 53284
rect 15036 53060 15092 53070
rect 14812 52948 14868 52958
rect 14700 52946 14868 52948
rect 14700 52894 14814 52946
rect 14866 52894 14868 52946
rect 14700 52892 14868 52894
rect 14812 52612 14868 52892
rect 14812 52546 14868 52556
rect 15036 52052 15092 53004
rect 15260 53060 15316 53566
rect 15260 52994 15316 53004
rect 15372 53620 15428 53630
rect 14252 49084 14644 49140
rect 14700 52050 15092 52052
rect 14700 51998 15038 52050
rect 15090 51998 15092 52050
rect 14700 51996 15092 51998
rect 14140 49028 14196 49038
rect 14140 48934 14196 48972
rect 14028 48738 14084 48748
rect 14140 48356 14196 48366
rect 14140 48262 14196 48300
rect 14140 48132 14196 48142
rect 13916 47406 13918 47458
rect 13970 47406 13972 47458
rect 13916 47394 13972 47406
rect 14028 48076 14140 48132
rect 14028 47124 14084 48076
rect 14140 48066 14196 48076
rect 14140 47460 14196 47470
rect 14140 47366 14196 47404
rect 14028 47058 14084 47068
rect 13916 46900 13972 46910
rect 13804 46898 13972 46900
rect 13804 46846 13918 46898
rect 13970 46846 13972 46898
rect 13804 46844 13972 46846
rect 13804 45892 13860 46844
rect 13916 46834 13972 46844
rect 13804 45826 13860 45836
rect 13804 45668 13860 45678
rect 13692 45666 13860 45668
rect 13692 45614 13806 45666
rect 13858 45614 13860 45666
rect 13692 45612 13860 45614
rect 13692 45332 13748 45612
rect 13804 45602 13860 45612
rect 14252 45444 14308 49084
rect 14364 48914 14420 48926
rect 14364 48862 14366 48914
rect 14418 48862 14420 48914
rect 14364 48692 14420 48862
rect 14364 48626 14420 48636
rect 14476 48916 14532 48926
rect 14364 47348 14420 47358
rect 14364 47254 14420 47292
rect 14364 47124 14420 47134
rect 14364 45890 14420 47068
rect 14364 45838 14366 45890
rect 14418 45838 14420 45890
rect 14364 45826 14420 45838
rect 13692 45266 13748 45276
rect 13804 45388 14308 45444
rect 13692 45106 13748 45118
rect 13692 45054 13694 45106
rect 13746 45054 13748 45106
rect 13692 44996 13748 45054
rect 13692 44930 13748 44940
rect 13580 44482 13636 44492
rect 13692 44436 13748 44446
rect 13468 44270 13470 44322
rect 13522 44270 13524 44322
rect 13468 44212 13524 44270
rect 13580 44324 13636 44334
rect 13692 44324 13748 44380
rect 13580 44322 13748 44324
rect 13580 44270 13582 44322
rect 13634 44270 13748 44322
rect 13580 44268 13748 44270
rect 13580 44258 13636 44268
rect 13468 44146 13524 44156
rect 13692 44098 13748 44110
rect 13692 44046 13694 44098
rect 13746 44046 13748 44098
rect 13692 43988 13748 44046
rect 13692 43922 13748 43932
rect 13804 43428 13860 45388
rect 13916 45218 13972 45230
rect 13916 45166 13918 45218
rect 13970 45166 13972 45218
rect 13916 44436 13972 45166
rect 14028 45220 14084 45230
rect 14364 45220 14420 45230
rect 14028 45218 14420 45220
rect 14028 45166 14030 45218
rect 14082 45166 14366 45218
rect 14418 45166 14420 45218
rect 14028 45164 14420 45166
rect 14028 45154 14084 45164
rect 14364 45154 14420 45164
rect 14476 44436 14532 48860
rect 14588 48914 14644 48926
rect 14588 48862 14590 48914
rect 14642 48862 14644 48914
rect 14588 48692 14644 48862
rect 14700 48804 14756 51996
rect 15036 51986 15092 51996
rect 15148 52946 15204 52958
rect 15148 52894 15150 52946
rect 15202 52894 15204 52946
rect 15148 52164 15204 52894
rect 15372 52948 15428 53564
rect 15372 52882 15428 52892
rect 14820 51772 15084 51782
rect 14876 51716 14924 51772
rect 14980 51716 15028 51772
rect 14820 51706 15084 51716
rect 14812 50820 14868 50830
rect 14812 50482 14868 50764
rect 15148 50820 15204 52108
rect 15372 51268 15428 51278
rect 15148 50754 15204 50764
rect 15260 51266 15428 51268
rect 15260 51214 15374 51266
rect 15426 51214 15428 51266
rect 15260 51212 15428 51214
rect 14812 50430 14814 50482
rect 14866 50430 14868 50482
rect 14812 50418 14868 50430
rect 15036 50484 15092 50494
rect 15036 50390 15092 50428
rect 14820 50204 15084 50214
rect 14876 50148 14924 50204
rect 14980 50148 15028 50204
rect 14820 50138 15084 50148
rect 15260 50148 15316 51212
rect 15372 51202 15428 51212
rect 15260 50082 15316 50092
rect 15372 51044 15428 51054
rect 15372 50594 15428 50988
rect 15372 50542 15374 50594
rect 15426 50542 15428 50594
rect 15148 49812 15204 49822
rect 15372 49812 15428 50542
rect 15148 49810 15428 49812
rect 15148 49758 15150 49810
rect 15202 49758 15428 49810
rect 15148 49756 15428 49758
rect 15148 49028 15204 49756
rect 15484 49588 15540 54684
rect 15820 54628 15876 54638
rect 15820 54626 15988 54628
rect 15820 54574 15822 54626
rect 15874 54574 15988 54626
rect 15820 54572 15988 54574
rect 15820 54562 15876 54572
rect 15596 53284 15652 53294
rect 15596 52162 15652 53228
rect 15708 53060 15764 53070
rect 15708 52966 15764 53004
rect 15932 53060 15988 54572
rect 15932 52994 15988 53004
rect 15596 52110 15598 52162
rect 15650 52110 15652 52162
rect 15596 51380 15652 52110
rect 15596 51314 15652 51324
rect 15932 51154 15988 51166
rect 15932 51102 15934 51154
rect 15986 51102 15988 51154
rect 15932 50820 15988 51102
rect 15932 50754 15988 50764
rect 15596 50370 15652 50382
rect 15596 50318 15598 50370
rect 15650 50318 15652 50370
rect 15596 50036 15652 50318
rect 15932 50148 15988 50158
rect 15652 49980 15764 50036
rect 15596 49970 15652 49980
rect 15484 49522 15540 49532
rect 15372 49140 15428 49150
rect 15204 48972 15316 49028
rect 15148 48962 15204 48972
rect 14924 48914 14980 48926
rect 14924 48862 14926 48914
rect 14978 48862 14980 48914
rect 14924 48804 14980 48862
rect 14700 48748 15204 48804
rect 14588 48636 14756 48692
rect 14588 48242 14644 48254
rect 14588 48190 14590 48242
rect 14642 48190 14644 48242
rect 14588 45332 14644 48190
rect 14700 48020 14756 48636
rect 14820 48636 15084 48646
rect 14876 48580 14924 48636
rect 14980 48580 15028 48636
rect 14820 48570 15084 48580
rect 15036 48468 15092 48478
rect 15036 48242 15092 48412
rect 15036 48190 15038 48242
rect 15090 48190 15092 48242
rect 15036 48178 15092 48190
rect 15148 48244 15204 48748
rect 14700 47458 14756 47964
rect 14700 47406 14702 47458
rect 14754 47406 14756 47458
rect 14700 47394 14756 47406
rect 14700 47236 14756 47246
rect 14700 45892 14756 47180
rect 14820 47068 15084 47078
rect 14876 47012 14924 47068
rect 14980 47012 15028 47068
rect 14820 47002 15084 47012
rect 15036 46788 15092 46798
rect 15036 46674 15092 46732
rect 15036 46622 15038 46674
rect 15090 46622 15092 46674
rect 15036 46610 15092 46622
rect 15148 46676 15204 48188
rect 15260 47684 15316 48972
rect 15260 47458 15316 47628
rect 15260 47406 15262 47458
rect 15314 47406 15316 47458
rect 15260 47394 15316 47406
rect 15372 47012 15428 49084
rect 15372 46956 15652 47012
rect 15260 46900 15316 46910
rect 15260 46898 15428 46900
rect 15260 46846 15262 46898
rect 15314 46846 15428 46898
rect 15260 46844 15428 46846
rect 15260 46834 15316 46844
rect 15260 46676 15316 46686
rect 15148 46674 15316 46676
rect 15148 46622 15262 46674
rect 15314 46622 15316 46674
rect 15148 46620 15316 46622
rect 15260 46610 15316 46620
rect 14700 45826 14756 45836
rect 14700 45668 14756 45678
rect 14700 45574 14756 45612
rect 14820 45500 15084 45510
rect 14876 45444 14924 45500
rect 14980 45444 15028 45500
rect 14820 45434 15084 45444
rect 14588 44548 14644 45276
rect 14924 45332 14980 45342
rect 14812 45218 14868 45230
rect 14812 45166 14814 45218
rect 14866 45166 14868 45218
rect 14812 44772 14868 45166
rect 14812 44706 14868 44716
rect 14588 44482 14644 44492
rect 13916 44370 13972 44380
rect 14028 44380 14532 44436
rect 13916 44100 13972 44110
rect 13916 44006 13972 44044
rect 13804 43362 13860 43372
rect 13916 43764 13972 43774
rect 13804 42868 13860 42878
rect 13692 42812 13804 42868
rect 13580 41860 13636 41870
rect 13580 41186 13636 41804
rect 13580 41134 13582 41186
rect 13634 41134 13636 41186
rect 13580 41122 13636 41134
rect 13468 41074 13524 41086
rect 13468 41022 13470 41074
rect 13522 41022 13524 41074
rect 13468 40628 13524 41022
rect 13468 40562 13524 40572
rect 13580 40628 13636 40638
rect 13692 40628 13748 42812
rect 13804 42802 13860 42812
rect 13916 42866 13972 43708
rect 13916 42814 13918 42866
rect 13970 42814 13972 42866
rect 13916 42802 13972 42814
rect 14028 41412 14084 44380
rect 14700 44324 14756 44334
rect 14252 44322 14756 44324
rect 14252 44270 14702 44322
rect 14754 44270 14756 44322
rect 14252 44268 14756 44270
rect 14252 43988 14308 44268
rect 14700 44258 14756 44268
rect 14924 44322 14980 45276
rect 15260 45106 15316 45118
rect 15260 45054 15262 45106
rect 15314 45054 15316 45106
rect 15260 44434 15316 45054
rect 15372 44884 15428 46844
rect 15484 46676 15540 46686
rect 15484 45218 15540 46620
rect 15484 45166 15486 45218
rect 15538 45166 15540 45218
rect 15484 45154 15540 45166
rect 15596 44996 15652 46956
rect 15708 45332 15764 49980
rect 15932 49026 15988 50092
rect 15932 48974 15934 49026
rect 15986 48974 15988 49026
rect 15932 48468 15988 48974
rect 15932 48402 15988 48412
rect 16044 47684 16100 59948
rect 16380 59938 16436 59948
rect 16156 59780 16212 59790
rect 16156 59444 16212 59724
rect 16156 58546 16212 59388
rect 16492 58660 16548 63532
rect 16604 63026 16660 64428
rect 16604 62974 16606 63026
rect 16658 62974 16660 63026
rect 16604 62962 16660 62974
rect 16604 61572 16660 61582
rect 16604 60564 16660 61516
rect 16604 60498 16660 60508
rect 16156 58494 16158 58546
rect 16210 58494 16212 58546
rect 16156 58482 16212 58494
rect 16268 58604 16548 58660
rect 16604 59220 16660 59230
rect 16716 59220 16772 66892
rect 16828 66164 16884 66174
rect 16828 66070 16884 66108
rect 16940 65604 16996 68348
rect 16828 65548 16996 65604
rect 16828 65266 16884 65548
rect 16828 65214 16830 65266
rect 16882 65214 16884 65266
rect 16828 64708 16884 65214
rect 16940 65378 16996 65390
rect 16940 65326 16942 65378
rect 16994 65326 16996 65378
rect 16940 64930 16996 65326
rect 16940 64878 16942 64930
rect 16994 64878 16996 64930
rect 16940 64866 16996 64878
rect 16940 64708 16996 64718
rect 16828 64706 16996 64708
rect 16828 64654 16942 64706
rect 16994 64654 16996 64706
rect 16828 64652 16996 64654
rect 16940 64642 16996 64652
rect 17052 64260 17108 77980
rect 17164 77364 17220 77374
rect 17276 77364 17332 82292
rect 17724 82068 17780 83468
rect 17500 82066 17780 82068
rect 17500 82014 17726 82066
rect 17778 82014 17780 82066
rect 17500 82012 17780 82014
rect 17500 81394 17556 82012
rect 17724 82002 17780 82012
rect 17836 83410 17892 84924
rect 17836 83358 17838 83410
rect 17890 83358 17892 83410
rect 17724 81732 17780 81742
rect 17836 81732 17892 83358
rect 17780 81676 17892 81732
rect 17948 85090 18004 85102
rect 17948 85038 17950 85090
rect 18002 85038 18004 85090
rect 17948 83524 18004 85038
rect 18620 85092 18676 85102
rect 18620 84998 18676 85036
rect 18620 84194 18676 84206
rect 18620 84142 18622 84194
rect 18674 84142 18676 84194
rect 18620 83972 18676 84142
rect 18732 84084 18788 85820
rect 18732 84018 18788 84028
rect 18222 83916 18486 83926
rect 18278 83860 18326 83916
rect 18382 83860 18430 83916
rect 18222 83850 18486 83860
rect 18396 83634 18452 83646
rect 18396 83582 18398 83634
rect 18450 83582 18452 83634
rect 18060 83524 18116 83534
rect 17948 83522 18116 83524
rect 17948 83470 18062 83522
rect 18114 83470 18116 83522
rect 17948 83468 18116 83470
rect 17724 81666 17780 81676
rect 17500 81342 17502 81394
rect 17554 81342 17556 81394
rect 17500 81330 17556 81342
rect 17836 81396 17892 81406
rect 17948 81396 18004 83468
rect 18060 83458 18116 83468
rect 18396 83524 18452 83582
rect 18396 83458 18452 83468
rect 17836 81394 18004 81396
rect 17836 81342 17838 81394
rect 17890 81342 18004 81394
rect 17836 81340 18004 81342
rect 18060 82626 18116 82638
rect 18060 82574 18062 82626
rect 18114 82574 18116 82626
rect 18060 82514 18116 82574
rect 18508 82628 18564 82638
rect 18620 82628 18676 83916
rect 18844 83636 18900 86156
rect 19404 85876 19460 87612
rect 19740 88338 19796 88350
rect 19740 88286 19742 88338
rect 19794 88286 19796 88338
rect 19516 87332 19572 87342
rect 19516 87330 19684 87332
rect 19516 87278 19518 87330
rect 19570 87278 19684 87330
rect 19516 87276 19684 87278
rect 19516 87266 19572 87276
rect 19404 85810 19460 85820
rect 19516 86546 19572 86558
rect 19516 86494 19518 86546
rect 19570 86494 19572 86546
rect 19068 85764 19124 85774
rect 19516 85708 19572 86494
rect 19068 83972 19124 85708
rect 19404 85652 19572 85708
rect 19628 85764 19684 87276
rect 19740 86882 19796 88286
rect 19852 88114 19908 89292
rect 19852 88062 19854 88114
rect 19906 88062 19908 88114
rect 19852 88050 19908 88062
rect 19964 88900 20020 88910
rect 19964 87666 20020 88844
rect 20076 88340 20132 88350
rect 20076 88246 20132 88284
rect 19964 87614 19966 87666
rect 20018 87614 20020 87666
rect 19964 87602 20020 87614
rect 20300 87556 20356 90524
rect 20412 90578 20468 90590
rect 20412 90526 20414 90578
rect 20466 90526 20468 90578
rect 20412 90468 20468 90526
rect 20636 90578 20692 90860
rect 20860 90692 20916 92988
rect 21196 92260 21252 94446
rect 21644 94500 21700 94510
rect 21756 94500 21812 94556
rect 21644 94498 21812 94500
rect 21644 94446 21646 94498
rect 21698 94446 21812 94498
rect 21644 94444 21812 94446
rect 21644 94434 21700 94444
rect 21868 94388 21924 94398
rect 21420 94274 21476 94286
rect 21420 94222 21422 94274
rect 21474 94222 21476 94274
rect 21308 93828 21364 93838
rect 21308 92370 21364 93772
rect 21420 92930 21476 94222
rect 21756 94276 21812 94286
rect 21868 94276 21924 94332
rect 21812 94220 21924 94276
rect 21756 94210 21812 94220
rect 21624 94108 21888 94118
rect 21680 94052 21728 94108
rect 21784 94052 21832 94108
rect 21980 94108 22036 94556
rect 22428 94274 22484 94286
rect 22428 94222 22430 94274
rect 22482 94222 22484 94274
rect 21980 94052 22372 94108
rect 21624 94042 21888 94052
rect 21644 93940 21700 93950
rect 21644 93042 21700 93884
rect 21980 93940 22036 93950
rect 21644 92990 21646 93042
rect 21698 92990 21700 93042
rect 21644 92978 21700 92990
rect 21756 93828 21812 93838
rect 21420 92878 21422 92930
rect 21474 92878 21476 92930
rect 21420 92866 21476 92878
rect 21756 92930 21812 93772
rect 21756 92878 21758 92930
rect 21810 92878 21812 92930
rect 21756 92866 21812 92878
rect 21980 92930 22036 93884
rect 22316 93938 22372 94052
rect 22316 93886 22318 93938
rect 22370 93886 22372 93938
rect 22316 93874 22372 93886
rect 22428 93940 22484 94222
rect 22428 93874 22484 93884
rect 22540 93716 22596 93726
rect 22428 93714 22596 93716
rect 22428 93662 22542 93714
rect 22594 93662 22596 93714
rect 22428 93660 22596 93662
rect 22316 93156 22372 93166
rect 22428 93156 22484 93660
rect 22540 93650 22596 93660
rect 22316 93154 22484 93156
rect 22316 93102 22318 93154
rect 22370 93102 22484 93154
rect 22316 93100 22484 93102
rect 22540 93100 22820 93156
rect 22316 93090 22372 93100
rect 22540 93044 22596 93100
rect 22428 92988 22596 93044
rect 22764 93044 22820 93100
rect 22876 93044 22932 93054
rect 22764 93042 22932 93044
rect 22764 92990 22878 93042
rect 22930 92990 22932 93042
rect 22764 92988 22932 92990
rect 22428 92932 22484 92988
rect 22876 92978 22932 92988
rect 21980 92878 21982 92930
rect 22034 92878 22036 92930
rect 21980 92866 22036 92878
rect 22204 92876 22484 92932
rect 22652 92930 22708 92942
rect 22652 92878 22654 92930
rect 22706 92878 22708 92930
rect 21532 92820 21588 92830
rect 21532 92706 21588 92764
rect 21532 92654 21534 92706
rect 21586 92654 21588 92706
rect 21532 92642 21588 92654
rect 21624 92540 21888 92550
rect 21680 92484 21728 92540
rect 21784 92484 21832 92540
rect 21624 92474 21888 92484
rect 21308 92318 21310 92370
rect 21362 92318 21364 92370
rect 21308 92306 21364 92318
rect 21196 92194 21252 92204
rect 22092 92260 22148 92270
rect 21980 92146 22036 92158
rect 21980 92094 21982 92146
rect 22034 92094 22036 92146
rect 21980 91364 22036 92094
rect 21980 91298 22036 91308
rect 22092 91250 22148 92204
rect 22204 91362 22260 92876
rect 22540 92820 22596 92830
rect 22428 92764 22540 92820
rect 22428 92370 22484 92764
rect 22540 92754 22596 92764
rect 22428 92318 22430 92370
rect 22482 92318 22484 92370
rect 22428 92306 22484 92318
rect 22316 92260 22372 92270
rect 22316 92166 22372 92204
rect 22428 92148 22484 92158
rect 22204 91310 22206 91362
rect 22258 91310 22260 91362
rect 22204 91298 22260 91310
rect 22316 91364 22372 91374
rect 22316 91270 22372 91308
rect 22092 91198 22094 91250
rect 22146 91198 22148 91250
rect 21624 90972 21888 90982
rect 21680 90916 21728 90972
rect 21784 90916 21832 90972
rect 21624 90906 21888 90916
rect 22092 90804 22148 91198
rect 22428 91140 22484 92092
rect 22540 92146 22596 92158
rect 22540 92094 22542 92146
rect 22594 92094 22596 92146
rect 22540 91252 22596 92094
rect 22652 92036 22708 92878
rect 22876 92148 22932 92158
rect 22876 92054 22932 92092
rect 22652 91970 22708 91980
rect 22988 91700 23044 102396
rect 23660 102450 23716 102956
rect 23660 102398 23662 102450
rect 23714 102398 23716 102450
rect 23660 102386 23716 102398
rect 23212 102340 23268 102350
rect 23212 102246 23268 102284
rect 23772 102228 23828 104188
rect 23996 104132 24052 105982
rect 23996 104066 24052 104076
rect 24108 103682 24164 103694
rect 24108 103630 24110 103682
rect 24162 103630 24164 103682
rect 24108 103572 24164 103630
rect 23884 103516 24164 103572
rect 23884 102452 23940 103516
rect 23996 103348 24052 103358
rect 24220 103348 24276 114212
rect 24668 109228 24724 117070
rect 25026 116844 25290 116854
rect 25082 116788 25130 116844
rect 25186 116788 25234 116844
rect 25026 116778 25290 116788
rect 25026 115276 25290 115286
rect 25082 115220 25130 115276
rect 25186 115220 25234 115276
rect 25026 115210 25290 115220
rect 24780 114660 24836 114670
rect 24780 112532 24836 114604
rect 28252 114268 28308 119600
rect 28428 117628 28692 117638
rect 28484 117572 28532 117628
rect 28588 117572 28636 117628
rect 28428 117562 28692 117572
rect 28428 116060 28692 116070
rect 28484 116004 28532 116060
rect 28588 116004 28636 116060
rect 28428 115994 28692 116004
rect 28428 114492 28692 114502
rect 28484 114436 28532 114492
rect 28588 114436 28636 114492
rect 28428 114426 28692 114436
rect 28140 114212 28308 114268
rect 25026 113708 25290 113718
rect 25082 113652 25130 113708
rect 25186 113652 25234 113708
rect 25026 113642 25290 113652
rect 25900 113316 25956 113326
rect 24780 112530 24948 112532
rect 24780 112478 24782 112530
rect 24834 112478 24948 112530
rect 24780 112476 24948 112478
rect 24780 112466 24836 112476
rect 24892 111972 24948 112476
rect 25900 112530 25956 113260
rect 25900 112478 25902 112530
rect 25954 112478 25956 112530
rect 25026 112140 25290 112150
rect 25082 112084 25130 112140
rect 25186 112084 25234 112140
rect 25026 112074 25290 112084
rect 25228 111972 25284 111982
rect 24892 111970 25284 111972
rect 24892 111918 25230 111970
rect 25282 111918 25284 111970
rect 24892 111916 25284 111918
rect 25228 111906 25284 111916
rect 25788 111748 25844 111758
rect 25900 111748 25956 112478
rect 25788 111746 25956 111748
rect 25788 111694 25790 111746
rect 25842 111694 25956 111746
rect 25788 111692 25956 111694
rect 26684 113314 26740 113326
rect 26684 113262 26686 113314
rect 26738 113262 26740 113314
rect 26684 112530 26740 113262
rect 26684 112478 26686 112530
rect 26738 112478 26740 112530
rect 26684 111748 26740 112478
rect 28028 111972 28084 111982
rect 28028 111858 28084 111916
rect 28028 111806 28030 111858
rect 28082 111806 28084 111858
rect 28028 111794 28084 111806
rect 25788 110964 25844 111692
rect 25900 110964 25956 110974
rect 25788 110962 25956 110964
rect 25788 110910 25902 110962
rect 25954 110910 25956 110962
rect 25788 110908 25956 110910
rect 25026 110572 25290 110582
rect 25082 110516 25130 110572
rect 25186 110516 25234 110572
rect 25026 110506 25290 110516
rect 24444 109172 24724 109228
rect 25900 110178 25956 110908
rect 25900 110126 25902 110178
rect 25954 110126 25956 110178
rect 25900 109394 25956 110126
rect 25900 109342 25902 109394
rect 25954 109342 25956 109394
rect 24332 107604 24388 107614
rect 24332 107510 24388 107548
rect 24332 106036 24388 106046
rect 24332 105942 24388 105980
rect 24444 105700 24500 109172
rect 25026 109004 25290 109014
rect 25082 108948 25130 109004
rect 25186 108948 25234 109004
rect 25026 108938 25290 108948
rect 24892 108724 24948 108734
rect 24892 108610 24948 108668
rect 25900 108724 25956 109342
rect 24892 108558 24894 108610
rect 24946 108558 24948 108610
rect 24892 108546 24948 108558
rect 25676 108612 25732 108622
rect 25676 108518 25732 108556
rect 24668 108388 24724 108398
rect 24668 107604 24724 108332
rect 24668 106820 24724 107548
rect 25900 107826 25956 108668
rect 25900 107774 25902 107826
rect 25954 107774 25956 107826
rect 24780 107492 24836 107502
rect 24836 107436 24948 107492
rect 24780 107426 24836 107436
rect 24892 107156 24948 107436
rect 25026 107436 25290 107446
rect 25082 107380 25130 107436
rect 25186 107380 25234 107436
rect 25026 107370 25290 107380
rect 25004 107156 25060 107166
rect 24892 107154 25060 107156
rect 24892 107102 25006 107154
rect 25058 107102 25060 107154
rect 24892 107100 25060 107102
rect 25004 107090 25060 107100
rect 25900 107042 25956 107774
rect 25900 106990 25902 107042
rect 25954 106990 25956 107042
rect 24668 106818 24836 106820
rect 24668 106766 24670 106818
rect 24722 106766 24836 106818
rect 24668 106764 24836 106766
rect 24668 106754 24724 106764
rect 24444 105634 24500 105644
rect 24444 105476 24500 105486
rect 23996 103346 24276 103348
rect 23996 103294 23998 103346
rect 24050 103294 24276 103346
rect 23996 103292 24276 103294
rect 24332 105474 24500 105476
rect 24332 105422 24446 105474
rect 24498 105422 24500 105474
rect 24332 105420 24500 105422
rect 23996 103282 24052 103292
rect 24220 103124 24276 103134
rect 24220 103030 24276 103068
rect 23884 102386 23940 102396
rect 24220 102452 24276 102462
rect 24332 102452 24388 105420
rect 24444 105410 24500 105420
rect 24780 105364 24836 106764
rect 25340 106260 25396 106270
rect 25340 106166 25396 106204
rect 25900 106258 25956 106990
rect 25900 106206 25902 106258
rect 25954 106206 25956 106258
rect 25900 106194 25956 106206
rect 26684 110962 26740 111692
rect 26684 110910 26686 110962
rect 26738 110910 26740 110962
rect 26684 110178 26740 110910
rect 26684 110126 26686 110178
rect 26738 110126 26740 110178
rect 26684 109394 26740 110126
rect 26684 109342 26686 109394
rect 26738 109342 26740 109394
rect 26684 108612 26740 109342
rect 26684 107826 26740 108556
rect 27244 108388 27300 108398
rect 27244 108294 27300 108332
rect 26684 107774 26686 107826
rect 26738 107774 26740 107826
rect 26684 107042 26740 107774
rect 26684 106990 26686 107042
rect 26738 106990 26740 107042
rect 26684 106258 26740 106990
rect 26684 106206 26686 106258
rect 26738 106206 26740 106258
rect 26684 106194 26740 106206
rect 24892 106036 24948 106046
rect 24892 105476 24948 105980
rect 25026 105868 25290 105878
rect 25082 105812 25130 105868
rect 25186 105812 25234 105868
rect 25026 105802 25290 105812
rect 26236 105588 26292 105598
rect 26236 105494 26292 105532
rect 28028 105588 28084 105598
rect 25004 105476 25060 105486
rect 24892 105474 25060 105476
rect 24892 105422 25006 105474
rect 25058 105422 25060 105474
rect 24892 105420 25060 105422
rect 25004 105410 25060 105420
rect 24780 105298 24836 105308
rect 24668 105252 24724 105262
rect 24220 102450 24388 102452
rect 24220 102398 24222 102450
rect 24274 102398 24388 102450
rect 24220 102396 24388 102398
rect 24444 104132 24500 104142
rect 24444 103906 24500 104076
rect 24668 104018 24724 105196
rect 25340 105250 25396 105262
rect 25340 105198 25342 105250
rect 25394 105198 25396 105250
rect 25228 104804 25284 104814
rect 24668 103966 24670 104018
rect 24722 103966 24724 104018
rect 24668 103954 24724 103966
rect 24892 104802 25284 104804
rect 24892 104750 25230 104802
rect 25282 104750 25284 104802
rect 24892 104748 25284 104750
rect 24444 103854 24446 103906
rect 24498 103854 24500 103906
rect 24220 102386 24276 102396
rect 23996 102338 24052 102350
rect 23996 102286 23998 102338
rect 24050 102286 24052 102338
rect 23996 102228 24052 102286
rect 23772 102172 24052 102228
rect 24332 102228 24388 102238
rect 24444 102228 24500 103854
rect 24892 103906 24948 104748
rect 25228 104738 25284 104748
rect 25340 104692 25396 105198
rect 25676 105252 25732 105262
rect 25676 105158 25732 105196
rect 26012 105252 26068 105262
rect 25676 104692 25732 104702
rect 25340 104690 25732 104692
rect 25340 104638 25678 104690
rect 25730 104638 25732 104690
rect 25340 104636 25732 104638
rect 25676 104626 25732 104636
rect 25026 104300 25290 104310
rect 25082 104244 25130 104300
rect 25186 104244 25234 104300
rect 25026 104234 25290 104244
rect 26012 104018 26068 105196
rect 26684 105252 26740 105262
rect 26684 105158 26740 105196
rect 28028 104914 28084 105532
rect 28028 104862 28030 104914
rect 28082 104862 28084 104914
rect 28028 104850 28084 104862
rect 26684 104690 26740 104702
rect 26684 104638 26686 104690
rect 26738 104638 26740 104690
rect 26684 104132 26740 104638
rect 26684 104066 26740 104076
rect 27580 104132 27636 104142
rect 27580 104038 27636 104076
rect 26012 103966 26014 104018
rect 26066 103966 26068 104018
rect 26012 103954 26068 103966
rect 27692 103908 27748 103918
rect 24892 103854 24894 103906
rect 24946 103854 24948 103906
rect 24892 103842 24948 103854
rect 26908 103906 27748 103908
rect 26908 103854 27694 103906
rect 27746 103854 27748 103906
rect 26908 103852 27748 103854
rect 26908 103794 26964 103852
rect 27692 103842 27748 103852
rect 26908 103742 26910 103794
rect 26962 103742 26964 103794
rect 26908 103730 26964 103742
rect 24332 102226 24500 102228
rect 24332 102174 24334 102226
rect 24386 102174 24500 102226
rect 24332 102172 24500 102174
rect 24556 103012 24612 103022
rect 24332 102162 24388 102172
rect 24556 101892 24612 102956
rect 25340 103012 25396 103022
rect 25340 102918 25396 102956
rect 25026 102732 25290 102742
rect 25082 102676 25130 102732
rect 25186 102676 25234 102732
rect 25026 102666 25290 102676
rect 24780 102452 24836 102462
rect 24780 102358 24836 102396
rect 24444 101836 24612 101892
rect 23324 101554 23380 101566
rect 23324 101502 23326 101554
rect 23378 101502 23380 101554
rect 23324 100772 23380 101502
rect 23660 101554 23716 101566
rect 23660 101502 23662 101554
rect 23714 101502 23716 101554
rect 23324 100706 23380 100716
rect 23548 101442 23604 101454
rect 23548 101390 23550 101442
rect 23602 101390 23604 101442
rect 23436 100658 23492 100670
rect 23436 100606 23438 100658
rect 23490 100606 23492 100658
rect 23436 100210 23492 100606
rect 23436 100158 23438 100210
rect 23490 100158 23492 100210
rect 23436 100146 23492 100158
rect 23548 100210 23604 101390
rect 23548 100158 23550 100210
rect 23602 100158 23604 100210
rect 23548 100146 23604 100158
rect 23324 99988 23380 99998
rect 23324 99894 23380 99932
rect 23660 99204 23716 101502
rect 23884 101556 23940 101566
rect 23884 101462 23940 101500
rect 24332 101332 24388 101342
rect 24108 101330 24388 101332
rect 24108 101278 24334 101330
rect 24386 101278 24388 101330
rect 24108 101276 24388 101278
rect 24108 99988 24164 101276
rect 24332 101266 24388 101276
rect 24220 100772 24276 100782
rect 24220 100678 24276 100716
rect 24444 99988 24500 101836
rect 24556 101666 24612 101678
rect 24556 101614 24558 101666
rect 24610 101614 24612 101666
rect 24556 100884 24612 101614
rect 25340 101442 25396 101454
rect 25340 101390 25342 101442
rect 25394 101390 25396 101442
rect 24668 101332 24724 101342
rect 25340 101332 25396 101390
rect 24668 101330 24948 101332
rect 24668 101278 24670 101330
rect 24722 101278 24948 101330
rect 24668 101276 24948 101278
rect 25340 101276 25620 101332
rect 24668 101266 24724 101276
rect 24892 100996 24948 101276
rect 25026 101164 25290 101174
rect 25082 101108 25130 101164
rect 25186 101108 25234 101164
rect 25026 101098 25290 101108
rect 24892 100940 25172 100996
rect 24556 100882 24724 100884
rect 24556 100830 24558 100882
rect 24610 100830 24724 100882
rect 24556 100828 24724 100830
rect 24556 100818 24612 100828
rect 24108 99894 24164 99932
rect 24332 99932 24500 99988
rect 23660 99138 23716 99148
rect 23884 99874 23940 99886
rect 23884 99822 23886 99874
rect 23938 99822 23940 99874
rect 23884 99092 23940 99822
rect 23884 99026 23940 99036
rect 23772 98980 23828 98990
rect 23772 98644 23828 98924
rect 23884 98644 23940 98654
rect 23772 98642 23940 98644
rect 23772 98590 23886 98642
rect 23938 98590 23940 98642
rect 23772 98588 23940 98590
rect 23884 98578 23940 98588
rect 23996 98418 24052 98430
rect 23996 98366 23998 98418
rect 24050 98366 24052 98418
rect 23548 98308 23604 98318
rect 23548 98306 23828 98308
rect 23548 98254 23550 98306
rect 23602 98254 23828 98306
rect 23548 98252 23828 98254
rect 23548 98242 23604 98252
rect 23436 97858 23492 97870
rect 23436 97806 23438 97858
rect 23490 97806 23492 97858
rect 23100 97636 23156 97646
rect 23100 97542 23156 97580
rect 23324 97636 23380 97646
rect 23324 97412 23380 97580
rect 23436 97468 23492 97806
rect 23660 97748 23716 97758
rect 23548 97692 23660 97748
rect 23548 97634 23604 97692
rect 23660 97682 23716 97692
rect 23548 97582 23550 97634
rect 23602 97582 23604 97634
rect 23548 97570 23604 97582
rect 23772 97524 23828 98252
rect 23884 98196 23940 98206
rect 23884 98102 23940 98140
rect 23996 97972 24052 98366
rect 23996 97906 24052 97916
rect 24220 97634 24276 97646
rect 24220 97582 24222 97634
rect 24274 97582 24276 97634
rect 24220 97524 24276 97582
rect 23436 97412 23716 97468
rect 23772 97412 23940 97468
rect 24220 97458 24276 97468
rect 23212 97410 23380 97412
rect 23212 97358 23326 97410
rect 23378 97358 23380 97410
rect 23212 97356 23380 97358
rect 23212 95956 23268 97356
rect 23324 97318 23380 97356
rect 23548 97076 23604 97086
rect 23212 95862 23268 95900
rect 23436 97074 23604 97076
rect 23436 97022 23550 97074
rect 23602 97022 23604 97074
rect 23436 97020 23604 97022
rect 23324 95844 23380 95854
rect 23324 95750 23380 95788
rect 23436 95508 23492 97020
rect 23548 97010 23604 97020
rect 23660 96066 23716 97412
rect 23884 96740 23940 97412
rect 23884 96646 23940 96684
rect 24332 96180 24388 99932
rect 24444 99764 24500 99774
rect 24444 99762 24612 99764
rect 24444 99710 24446 99762
rect 24498 99710 24612 99762
rect 24444 99708 24612 99710
rect 24444 99698 24500 99708
rect 24444 98532 24500 98542
rect 24444 98438 24500 98476
rect 24556 98420 24612 99708
rect 24668 99092 24724 100828
rect 24892 100772 24948 100782
rect 24892 99988 24948 100716
rect 25116 100212 25172 100940
rect 25452 100660 25508 100670
rect 25340 100604 25452 100660
rect 25228 100212 25284 100222
rect 25116 100210 25284 100212
rect 25116 100158 25230 100210
rect 25282 100158 25284 100210
rect 25116 100156 25284 100158
rect 25228 100146 25284 100156
rect 25340 100210 25396 100604
rect 25452 100594 25508 100604
rect 25340 100158 25342 100210
rect 25394 100158 25396 100210
rect 25340 100146 25396 100158
rect 25564 100100 25620 101276
rect 27356 100770 27412 100782
rect 27356 100718 27358 100770
rect 27410 100718 27412 100770
rect 26684 100660 26740 100670
rect 26684 100566 26740 100604
rect 25676 100100 25732 100110
rect 25564 100098 25732 100100
rect 25564 100046 25678 100098
rect 25730 100046 25732 100098
rect 25564 100044 25732 100046
rect 24892 99316 24948 99932
rect 25452 99986 25508 99998
rect 25452 99934 25454 99986
rect 25506 99934 25508 99986
rect 25026 99596 25290 99606
rect 25082 99540 25130 99596
rect 25186 99540 25234 99596
rect 25026 99530 25290 99540
rect 24668 99026 24724 99036
rect 24780 99314 24948 99316
rect 24780 99262 24894 99314
rect 24946 99262 24948 99314
rect 24780 99260 24948 99262
rect 24556 98418 24724 98420
rect 24556 98366 24558 98418
rect 24610 98366 24724 98418
rect 24556 98364 24724 98366
rect 24556 98354 24612 98364
rect 23660 96014 23662 96066
rect 23714 96014 23716 96066
rect 23660 96002 23716 96014
rect 24108 96178 24388 96180
rect 24108 96126 24334 96178
rect 24386 96126 24388 96178
rect 24108 96124 24388 96126
rect 23436 95442 23492 95452
rect 24108 95506 24164 96124
rect 24108 95454 24110 95506
rect 24162 95454 24164 95506
rect 24108 95442 24164 95454
rect 24332 95508 24388 96124
rect 24444 98194 24500 98206
rect 24444 98142 24446 98194
rect 24498 98142 24500 98194
rect 24444 97746 24500 98142
rect 24444 97694 24446 97746
rect 24498 97694 24500 97746
rect 24444 96068 24500 97694
rect 24668 97748 24724 98364
rect 24668 97682 24724 97692
rect 24780 96180 24836 99260
rect 24892 99250 24948 99260
rect 25228 98532 25284 98542
rect 25228 98306 25284 98476
rect 25228 98254 25230 98306
rect 25282 98254 25284 98306
rect 25228 98242 25284 98254
rect 25026 98028 25290 98038
rect 25082 97972 25130 98028
rect 25186 97972 25234 98028
rect 25026 97962 25290 97972
rect 25340 97860 25396 97870
rect 25340 97766 25396 97804
rect 25452 97748 25508 99934
rect 25676 99876 25732 100044
rect 27356 99988 27412 100718
rect 27356 99922 27412 99932
rect 28028 99988 28084 99998
rect 26236 99876 26292 99886
rect 26684 99876 26740 99886
rect 25676 99874 26740 99876
rect 25676 99822 26238 99874
rect 26290 99822 26686 99874
rect 26738 99822 26740 99874
rect 25676 99820 26740 99822
rect 25676 98980 25732 99820
rect 26236 99810 26292 99820
rect 26684 99810 26740 99820
rect 25452 97654 25508 97692
rect 25564 98924 25676 98980
rect 25116 97636 25172 97646
rect 24892 97524 24948 97562
rect 24892 97458 24948 97468
rect 25116 97468 25172 97580
rect 25564 97636 25620 98924
rect 25676 98914 25732 98924
rect 25116 97412 25284 97468
rect 25228 96738 25284 97412
rect 25228 96686 25230 96738
rect 25282 96686 25284 96738
rect 25228 96674 25284 96686
rect 25026 96460 25290 96470
rect 25082 96404 25130 96460
rect 25186 96404 25234 96460
rect 25026 96394 25290 96404
rect 24780 96124 24948 96180
rect 24444 96002 24500 96012
rect 24556 95956 24612 95966
rect 24444 95508 24500 95518
rect 24332 95506 24500 95508
rect 24332 95454 24446 95506
rect 24498 95454 24500 95506
rect 24332 95452 24500 95454
rect 24444 95442 24500 95452
rect 24556 95394 24612 95900
rect 24556 95342 24558 95394
rect 24610 95342 24612 95394
rect 24556 95330 24612 95342
rect 24220 95284 24276 95294
rect 24220 95190 24276 95228
rect 24892 94500 24948 96124
rect 25228 96068 25284 96078
rect 25228 95974 25284 96012
rect 25340 95956 25396 95966
rect 25340 95862 25396 95900
rect 25452 95844 25508 95854
rect 25452 95750 25508 95788
rect 25452 95396 25508 95406
rect 25564 95396 25620 97580
rect 25676 98532 25732 98542
rect 25676 97634 25732 98476
rect 28028 98418 28084 99932
rect 28028 98366 28030 98418
rect 28082 98366 28084 98418
rect 27356 98306 27412 98318
rect 27356 98254 27358 98306
rect 27410 98254 27412 98306
rect 27356 98196 27412 98254
rect 27356 98130 27412 98140
rect 25676 97582 25678 97634
rect 25730 97582 25732 97634
rect 25676 97570 25732 97582
rect 26796 97636 26852 97646
rect 26684 97524 26740 97562
rect 26684 97458 26740 97468
rect 26796 97522 26852 97580
rect 27356 97636 27412 97646
rect 27356 97542 27412 97580
rect 26796 97470 26798 97522
rect 26850 97470 26852 97522
rect 26796 97458 26852 97470
rect 27020 97412 27076 97422
rect 27020 97410 27300 97412
rect 27020 97358 27022 97410
rect 27074 97358 27300 97410
rect 27020 97356 27300 97358
rect 27020 97346 27076 97356
rect 27244 96964 27300 97356
rect 27356 96964 27412 96974
rect 27244 96962 27412 96964
rect 27244 96910 27358 96962
rect 27410 96910 27412 96962
rect 27244 96908 27412 96910
rect 27356 96898 27412 96908
rect 28028 96850 28084 98366
rect 28028 96798 28030 96850
rect 28082 96798 28084 96850
rect 28028 96786 28084 96798
rect 26236 96740 26292 96750
rect 25452 95394 25620 95396
rect 25452 95342 25454 95394
rect 25506 95342 25620 95394
rect 25452 95340 25620 95342
rect 25452 95330 25508 95340
rect 25340 95284 25396 95294
rect 25340 95190 25396 95228
rect 25564 95284 25620 95340
rect 25900 96066 25956 96078
rect 25900 96014 25902 96066
rect 25954 96014 25956 96066
rect 25026 94892 25290 94902
rect 25082 94836 25130 94892
rect 25186 94836 25234 94892
rect 25026 94826 25290 94836
rect 25004 94500 25060 94510
rect 24892 94498 25060 94500
rect 24892 94446 25006 94498
rect 25058 94446 25060 94498
rect 24892 94444 25060 94446
rect 25004 94434 25060 94444
rect 23100 93604 23156 93614
rect 23100 93510 23156 93548
rect 25026 93324 25290 93334
rect 25082 93268 25130 93324
rect 25186 93268 25234 93324
rect 25026 93258 25290 93268
rect 25228 93044 25284 93054
rect 23660 92932 23716 92942
rect 23660 92930 24052 92932
rect 23660 92878 23662 92930
rect 23714 92878 24052 92930
rect 23660 92876 24052 92878
rect 23660 92866 23716 92876
rect 23324 92820 23380 92830
rect 23324 92726 23380 92764
rect 23996 92818 24052 92876
rect 23996 92766 23998 92818
rect 24050 92766 24052 92818
rect 23996 92754 24052 92766
rect 24108 92818 24164 92830
rect 24108 92766 24110 92818
rect 24162 92766 24164 92818
rect 23436 92706 23492 92718
rect 23436 92654 23438 92706
rect 23490 92654 23492 92706
rect 23436 92372 23492 92654
rect 23772 92708 23828 92718
rect 23772 92614 23828 92652
rect 24108 92484 24164 92766
rect 23996 92428 24164 92484
rect 23212 92316 23492 92372
rect 23548 92372 23604 92382
rect 23100 92260 23156 92270
rect 23100 92166 23156 92204
rect 23212 91700 23268 92316
rect 23548 92258 23604 92316
rect 23996 92370 24052 92428
rect 24332 92372 24388 92382
rect 23996 92318 23998 92370
rect 24050 92318 24052 92370
rect 23996 92306 24052 92318
rect 24108 92316 24332 92372
rect 23548 92206 23550 92258
rect 23602 92206 23604 92258
rect 23548 92194 23604 92206
rect 24108 92258 24164 92316
rect 24108 92206 24110 92258
rect 24162 92206 24164 92258
rect 24108 92194 24164 92206
rect 22988 91634 23044 91644
rect 23100 91644 23268 91700
rect 23324 92146 23380 92158
rect 23324 92094 23326 92146
rect 23378 92094 23380 92146
rect 22876 91588 22932 91598
rect 22876 91494 22932 91532
rect 22540 91158 22596 91196
rect 22988 91476 23044 91486
rect 23100 91476 23156 91644
rect 22988 91474 23156 91476
rect 22988 91422 22990 91474
rect 23042 91422 23156 91474
rect 22988 91420 23156 91422
rect 22428 91074 22484 91084
rect 22764 91140 22820 91150
rect 22092 90738 22148 90748
rect 22764 90802 22820 91084
rect 22764 90750 22766 90802
rect 22818 90750 22820 90802
rect 22764 90738 22820 90750
rect 22876 90916 22932 90926
rect 20860 90626 20916 90636
rect 21868 90690 21924 90702
rect 21868 90638 21870 90690
rect 21922 90638 21924 90690
rect 20636 90526 20638 90578
rect 20690 90526 20692 90578
rect 20636 90514 20692 90526
rect 21084 90580 21140 90590
rect 21308 90580 21364 90590
rect 21084 90578 21252 90580
rect 21084 90526 21086 90578
rect 21138 90526 21252 90578
rect 21084 90524 21252 90526
rect 21084 90514 21140 90524
rect 20412 90402 20468 90412
rect 20860 90468 20916 90478
rect 20860 90374 20916 90412
rect 21196 90356 21252 90524
rect 21308 90486 21364 90524
rect 21644 90578 21700 90590
rect 21644 90526 21646 90578
rect 21698 90526 21700 90578
rect 21644 90356 21700 90526
rect 21196 90300 21700 90356
rect 21756 89908 21812 89918
rect 21868 89908 21924 90638
rect 22876 90690 22932 90860
rect 22876 90638 22878 90690
rect 22930 90638 22932 90690
rect 22876 90626 22932 90638
rect 21980 90580 22036 90590
rect 22540 90580 22596 90590
rect 21980 90578 22596 90580
rect 21980 90526 21982 90578
rect 22034 90526 22542 90578
rect 22594 90526 22596 90578
rect 21980 90524 22596 90526
rect 21980 90514 22036 90524
rect 22540 90514 22596 90524
rect 22652 90356 22708 90366
rect 22988 90356 23044 91420
rect 23324 91364 23380 92094
rect 23884 92146 23940 92158
rect 23884 92094 23886 92146
rect 23938 92094 23940 92146
rect 23436 92036 23492 92046
rect 23436 91922 23492 91980
rect 23436 91870 23438 91922
rect 23490 91870 23492 91922
rect 23436 91858 23492 91870
rect 23884 91588 23940 92094
rect 23884 91522 23940 91532
rect 23548 91364 23604 91374
rect 23324 91308 23492 91364
rect 23212 91138 23268 91150
rect 23212 91086 23214 91138
rect 23266 91086 23268 91138
rect 23212 90916 23268 91086
rect 23212 90850 23268 90860
rect 23324 91138 23380 91150
rect 23324 91086 23326 91138
rect 23378 91086 23380 91138
rect 23324 90692 23380 91086
rect 23436 91140 23492 91308
rect 23436 91074 23492 91084
rect 23548 90916 23604 91308
rect 23772 91252 23828 91262
rect 23996 91252 24052 91262
rect 23548 90850 23604 90860
rect 23660 91196 23772 91252
rect 23828 91250 24052 91252
rect 23828 91198 23998 91250
rect 24050 91198 24052 91250
rect 23828 91196 24052 91198
rect 23436 90692 23492 90702
rect 23324 90636 23436 90692
rect 21868 89852 22148 89908
rect 21756 89796 21812 89852
rect 21420 89794 21812 89796
rect 21420 89742 21758 89794
rect 21810 89742 21812 89794
rect 21420 89740 21812 89742
rect 21420 89236 21476 89740
rect 21756 89730 21812 89740
rect 22092 89796 22148 89852
rect 22540 89796 22596 89806
rect 22092 89794 22596 89796
rect 22092 89742 22542 89794
rect 22594 89742 22596 89794
rect 22092 89740 22596 89742
rect 21868 89684 21924 89694
rect 21868 89590 21924 89628
rect 21980 89570 22036 89582
rect 21980 89518 21982 89570
rect 22034 89518 22036 89570
rect 21980 89460 22036 89518
rect 21624 89404 21888 89414
rect 21680 89348 21728 89404
rect 21784 89348 21832 89404
rect 21980 89394 22036 89404
rect 21624 89338 21888 89348
rect 21644 89236 21700 89246
rect 21420 89234 21700 89236
rect 21420 89182 21646 89234
rect 21698 89182 21700 89234
rect 21420 89180 21700 89182
rect 21644 89170 21700 89180
rect 21420 89012 21476 89022
rect 21420 88918 21476 88956
rect 22092 89010 22148 89740
rect 22540 89730 22596 89740
rect 22204 89572 22260 89582
rect 22260 89516 22484 89572
rect 22204 89478 22260 89516
rect 22428 89234 22484 89516
rect 22652 89460 22708 90300
rect 22764 90300 23044 90356
rect 23212 90356 23268 90366
rect 23324 90356 23380 90636
rect 23436 90598 23492 90636
rect 23548 90692 23604 90702
rect 23660 90692 23716 91196
rect 23772 91158 23828 91196
rect 23996 91186 24052 91196
rect 24220 91250 24276 92316
rect 24332 92306 24388 92316
rect 25228 92260 25284 92988
rect 25452 92820 25508 92830
rect 25228 92166 25284 92204
rect 25340 92818 25508 92820
rect 25340 92766 25454 92818
rect 25506 92766 25508 92818
rect 25340 92764 25508 92766
rect 24332 92146 24388 92158
rect 24332 92094 24334 92146
rect 24386 92094 24388 92146
rect 24332 92036 24388 92094
rect 24668 92148 24724 92158
rect 24668 92054 24724 92092
rect 25340 92036 25396 92764
rect 25452 92754 25508 92764
rect 25452 92372 25508 92382
rect 25452 92258 25508 92316
rect 25452 92206 25454 92258
rect 25506 92206 25508 92258
rect 25452 92194 25508 92206
rect 25340 91980 25508 92036
rect 24332 91970 24388 91980
rect 25026 91756 25290 91766
rect 25082 91700 25130 91756
rect 25186 91700 25234 91756
rect 25026 91690 25290 91700
rect 25228 91588 25284 91598
rect 24220 91198 24222 91250
rect 24274 91198 24276 91250
rect 24220 91028 24276 91198
rect 24220 90962 24276 90972
rect 24332 91250 24388 91262
rect 24332 91198 24334 91250
rect 24386 91198 24388 91250
rect 24332 91140 24388 91198
rect 23548 90690 23716 90692
rect 23548 90638 23550 90690
rect 23602 90638 23716 90690
rect 23548 90636 23716 90638
rect 23884 90916 23940 90926
rect 23548 90626 23604 90636
rect 23268 90300 23380 90356
rect 23436 90354 23492 90366
rect 23436 90302 23438 90354
rect 23490 90302 23492 90354
rect 22764 89908 22820 90300
rect 23212 90290 23268 90300
rect 22764 89684 22820 89852
rect 22876 90020 22932 90030
rect 23212 90020 23268 90030
rect 22932 90018 23268 90020
rect 22932 89966 23214 90018
rect 23266 89966 23268 90018
rect 22932 89964 23268 89966
rect 22876 89794 22932 89964
rect 23212 89954 23268 89964
rect 22876 89742 22878 89794
rect 22930 89742 22932 89794
rect 22876 89730 22932 89742
rect 22764 89590 22820 89628
rect 23324 89682 23380 89694
rect 23324 89630 23326 89682
rect 23378 89630 23380 89682
rect 23324 89572 23380 89630
rect 23324 89506 23380 89516
rect 22652 89404 22820 89460
rect 22428 89182 22430 89234
rect 22482 89182 22484 89234
rect 22428 89170 22484 89182
rect 22092 88958 22094 89010
rect 22146 88958 22148 89010
rect 22092 88946 22148 88958
rect 22652 89012 22708 89022
rect 20748 88900 20804 88910
rect 20524 88340 20580 88350
rect 20524 88246 20580 88284
rect 20748 88226 20804 88844
rect 21532 88900 21588 88910
rect 21532 88806 21588 88844
rect 22652 88450 22708 88956
rect 22652 88398 22654 88450
rect 22706 88398 22708 88450
rect 22652 88386 22708 88398
rect 22764 88786 22820 89404
rect 22988 89348 23044 89358
rect 22764 88734 22766 88786
rect 22818 88734 22820 88786
rect 20748 88174 20750 88226
rect 20802 88174 20804 88226
rect 20748 88162 20804 88174
rect 20412 88114 20468 88126
rect 20412 88062 20414 88114
rect 20466 88062 20468 88114
rect 20412 87892 20468 88062
rect 20412 87826 20468 87836
rect 21624 87836 21888 87846
rect 21680 87780 21728 87836
rect 21784 87780 21832 87836
rect 21624 87770 21888 87780
rect 20188 87500 20356 87556
rect 20188 86884 20244 87500
rect 20300 87330 20356 87342
rect 20300 87278 20302 87330
rect 20354 87278 20356 87330
rect 20300 87108 20356 87278
rect 20300 87042 20356 87052
rect 20860 87330 20916 87342
rect 21308 87332 21364 87342
rect 20860 87278 20862 87330
rect 20914 87278 20916 87330
rect 20860 87218 20916 87278
rect 20860 87166 20862 87218
rect 20914 87166 20916 87218
rect 19740 86830 19742 86882
rect 19794 86830 19796 86882
rect 19740 86818 19796 86830
rect 19852 86828 20244 86884
rect 19628 85698 19684 85708
rect 19180 85316 19236 85326
rect 19180 85222 19236 85260
rect 19068 83906 19124 83916
rect 19404 84196 19460 85652
rect 18508 82626 18676 82628
rect 18508 82574 18510 82626
rect 18562 82574 18676 82626
rect 18508 82572 18676 82574
rect 18508 82562 18564 82572
rect 18060 82462 18062 82514
rect 18114 82462 18116 82514
rect 18060 81396 18116 82462
rect 18222 82348 18486 82358
rect 18278 82292 18326 82348
rect 18382 82292 18430 82348
rect 18222 82282 18486 82292
rect 18620 82348 18676 82572
rect 18396 82068 18452 82078
rect 18396 81974 18452 82012
rect 18060 81340 18340 81396
rect 17836 81330 17892 81340
rect 17724 81172 17780 81182
rect 17948 81172 18004 81182
rect 18172 81172 18228 81182
rect 17724 81078 17780 81116
rect 17836 81170 18004 81172
rect 17836 81118 17950 81170
rect 18002 81118 18004 81170
rect 17836 81116 18004 81118
rect 17612 80948 17668 80958
rect 17836 80948 17892 81116
rect 17948 81106 18004 81116
rect 18060 81170 18228 81172
rect 18060 81118 18174 81170
rect 18226 81118 18228 81170
rect 18060 81116 18228 81118
rect 17668 80892 17892 80948
rect 17948 80948 18004 80958
rect 17612 80882 17668 80892
rect 17836 80612 17892 80622
rect 17500 80498 17556 80510
rect 17500 80446 17502 80498
rect 17554 80446 17556 80498
rect 17388 80386 17444 80398
rect 17388 80334 17390 80386
rect 17442 80334 17444 80386
rect 17388 79716 17444 80334
rect 17500 80276 17556 80446
rect 17836 80386 17892 80556
rect 17836 80334 17838 80386
rect 17890 80334 17892 80386
rect 17836 80322 17892 80334
rect 17500 80210 17556 80220
rect 17836 79940 17892 79950
rect 17724 79828 17780 79838
rect 17724 79734 17780 79772
rect 17612 79716 17668 79726
rect 17388 79660 17612 79716
rect 17612 79622 17668 79660
rect 17724 78930 17780 78942
rect 17724 78878 17726 78930
rect 17778 78878 17780 78930
rect 17500 78260 17556 78270
rect 17500 78166 17556 78204
rect 17724 78260 17780 78878
rect 17836 78820 17892 79884
rect 17948 79604 18004 80892
rect 18060 80386 18116 81116
rect 18172 81106 18228 81116
rect 18172 80948 18228 80958
rect 18284 80948 18340 81340
rect 18396 81282 18452 81294
rect 18396 81230 18398 81282
rect 18450 81230 18452 81282
rect 18396 80948 18452 81230
rect 18508 81284 18564 81294
rect 18620 81284 18676 82292
rect 18508 81282 18676 81284
rect 18508 81230 18510 81282
rect 18562 81230 18676 81282
rect 18508 81228 18676 81230
rect 18732 83580 18900 83636
rect 18956 83636 19012 83646
rect 18508 81218 18564 81228
rect 18228 80892 18452 80948
rect 18172 80882 18228 80892
rect 18222 80780 18486 80790
rect 18278 80724 18326 80780
rect 18382 80724 18430 80780
rect 18222 80714 18486 80724
rect 18284 80500 18340 80510
rect 18732 80500 18788 83580
rect 18956 83542 19012 83580
rect 19292 83524 19348 83534
rect 19292 83430 19348 83468
rect 18844 83412 18900 83422
rect 19404 83412 19460 84140
rect 19516 84868 19572 84878
rect 19516 83634 19572 84812
rect 19852 84530 19908 86828
rect 20076 86548 20132 86558
rect 19852 84478 19854 84530
rect 19906 84478 19908 84530
rect 19852 84466 19908 84478
rect 19964 86546 20132 86548
rect 19964 86494 20078 86546
rect 20130 86494 20132 86546
rect 19964 86492 20132 86494
rect 19964 86324 20020 86492
rect 20076 86482 20132 86492
rect 20188 86436 20244 86446
rect 20188 86342 20244 86380
rect 20412 86434 20468 86446
rect 20412 86382 20414 86434
rect 20466 86382 20468 86434
rect 19964 85764 20020 86268
rect 19964 84530 20020 85708
rect 20412 85652 20468 86382
rect 20748 86436 20804 86446
rect 20860 86436 20916 87166
rect 21196 87330 21364 87332
rect 21196 87278 21310 87330
rect 21362 87278 21364 87330
rect 21196 87276 21364 87278
rect 20748 86434 20916 86436
rect 20748 86382 20750 86434
rect 20802 86382 20916 86434
rect 20748 86380 20916 86382
rect 21084 86660 21140 86670
rect 20748 86324 20804 86380
rect 20748 86258 20804 86268
rect 20300 85596 20468 85652
rect 20300 84532 20356 85596
rect 20636 85316 20692 85326
rect 20636 85314 21028 85316
rect 20636 85262 20638 85314
rect 20690 85262 21028 85314
rect 20636 85260 21028 85262
rect 20636 85250 20692 85260
rect 19964 84478 19966 84530
rect 20018 84478 20020 84530
rect 19964 84466 20020 84478
rect 20188 84476 20356 84532
rect 20524 84980 20580 84990
rect 20076 84420 20132 84430
rect 20076 84326 20132 84364
rect 20188 84418 20244 84476
rect 20188 84366 20190 84418
rect 20242 84366 20244 84418
rect 20188 84354 20244 84366
rect 19740 84308 19796 84318
rect 20524 84308 20580 84924
rect 20748 84980 20804 84990
rect 20748 84978 20916 84980
rect 20748 84926 20750 84978
rect 20802 84926 20916 84978
rect 20748 84924 20916 84926
rect 20748 84914 20804 84924
rect 20636 84868 20692 84878
rect 20636 84774 20692 84812
rect 20860 84532 20916 84924
rect 19516 83582 19518 83634
rect 19570 83582 19572 83634
rect 19516 83570 19572 83582
rect 19628 84306 19796 84308
rect 19628 84254 19742 84306
rect 19794 84254 19796 84306
rect 19628 84252 19796 84254
rect 19404 83356 19572 83412
rect 18844 83318 18900 83356
rect 18956 82626 19012 82638
rect 19404 82628 19460 82638
rect 18956 82574 18958 82626
rect 19010 82574 19012 82626
rect 18956 82514 19012 82574
rect 18956 82462 18958 82514
rect 19010 82462 19012 82514
rect 18956 82450 19012 82462
rect 19292 82626 19460 82628
rect 19292 82574 19406 82626
rect 19458 82574 19460 82626
rect 19292 82572 19460 82574
rect 19292 82292 19348 82572
rect 19404 82562 19460 82572
rect 18844 81732 18900 81742
rect 19292 81732 19348 82236
rect 18844 81730 19460 81732
rect 18844 81678 18846 81730
rect 18898 81678 19294 81730
rect 19346 81678 19460 81730
rect 18844 81676 19460 81678
rect 18844 81666 18900 81676
rect 19292 81666 19348 81676
rect 19068 81396 19124 81406
rect 19068 81060 19124 81340
rect 19292 81396 19348 81406
rect 19292 81302 19348 81340
rect 19404 81172 19460 81676
rect 19404 81078 19460 81116
rect 19068 80994 19124 81004
rect 19292 80946 19348 80958
rect 19516 80948 19572 83356
rect 19292 80894 19294 80946
rect 19346 80894 19348 80946
rect 18284 80498 18788 80500
rect 18284 80446 18286 80498
rect 18338 80446 18788 80498
rect 18284 80444 18788 80446
rect 18844 80612 18900 80622
rect 18284 80434 18340 80444
rect 18060 80334 18062 80386
rect 18114 80334 18116 80386
rect 18060 80322 18116 80334
rect 18844 80386 18900 80556
rect 18844 80334 18846 80386
rect 18898 80334 18900 80386
rect 18844 80322 18900 80334
rect 19292 80386 19348 80894
rect 19292 80334 19294 80386
rect 19346 80334 19348 80386
rect 19292 80322 19348 80334
rect 19404 80892 19572 80948
rect 19628 83300 19684 84252
rect 19740 84242 19796 84252
rect 20300 84252 20580 84308
rect 20188 83972 20244 83982
rect 20076 83916 20188 83972
rect 18732 80276 18788 80286
rect 17948 79510 18004 79548
rect 18172 79602 18228 79614
rect 18172 79550 18174 79602
rect 18226 79550 18228 79602
rect 18172 79380 18228 79550
rect 18172 79314 18228 79324
rect 18222 79212 18486 79222
rect 18278 79156 18326 79212
rect 18382 79156 18430 79212
rect 18222 79146 18486 79156
rect 18732 79156 18788 80220
rect 19068 79716 19124 79726
rect 19124 79660 19348 79716
rect 19068 79602 19124 79660
rect 19068 79550 19070 79602
rect 19122 79550 19124 79602
rect 19068 79538 19124 79550
rect 19180 79490 19236 79502
rect 19180 79438 19182 79490
rect 19234 79438 19236 79490
rect 19068 79380 19124 79390
rect 18732 79100 19012 79156
rect 18060 78820 18116 78830
rect 17836 78818 18116 78820
rect 17836 78766 18062 78818
rect 18114 78766 18116 78818
rect 17836 78764 18116 78766
rect 18060 78754 18116 78764
rect 18620 78594 18676 78606
rect 18620 78542 18622 78594
rect 18674 78542 18676 78594
rect 18172 78260 18228 78270
rect 17724 78194 17780 78204
rect 18060 78204 18172 78260
rect 17220 77308 17332 77364
rect 17388 78034 17444 78046
rect 17388 77982 17390 78034
rect 17442 77982 17444 78034
rect 17388 77924 17444 77982
rect 17388 77476 17444 77868
rect 17164 65156 17220 77308
rect 17388 75572 17444 77420
rect 17500 78036 17556 78046
rect 17500 76690 17556 77980
rect 17612 78034 17668 78046
rect 17612 77982 17614 78034
rect 17666 77982 17668 78034
rect 17612 77924 17668 77982
rect 17948 78036 18004 78046
rect 17948 77942 18004 77980
rect 17612 77364 17668 77868
rect 17836 77812 17892 77822
rect 17836 77718 17892 77756
rect 17612 77298 17668 77308
rect 17500 76638 17502 76690
rect 17554 76638 17556 76690
rect 17500 75684 17556 76638
rect 18060 76580 18116 78204
rect 18172 78194 18228 78204
rect 18508 78260 18564 78270
rect 18508 78034 18564 78204
rect 18508 77982 18510 78034
rect 18562 77982 18564 78034
rect 18508 77970 18564 77982
rect 18508 77812 18564 77850
rect 18508 77746 18564 77756
rect 18222 77644 18486 77654
rect 18278 77588 18326 77644
rect 18382 77588 18430 77644
rect 18222 77578 18486 77588
rect 18396 77140 18452 77150
rect 18396 77046 18452 77084
rect 18172 76580 18228 76590
rect 18060 76578 18228 76580
rect 18060 76526 18174 76578
rect 18226 76526 18228 76578
rect 18060 76524 18228 76526
rect 18172 76514 18228 76524
rect 17500 75618 17556 75628
rect 17612 76356 17668 76366
rect 17388 75506 17444 75516
rect 17276 75460 17332 75470
rect 17276 75366 17332 75404
rect 17500 74900 17556 74910
rect 17612 74900 17668 76300
rect 18060 76242 18116 76254
rect 18060 76190 18062 76242
rect 18114 76190 18116 76242
rect 17724 75572 17780 75582
rect 17724 75478 17780 75516
rect 17948 75570 18004 75582
rect 17948 75518 17950 75570
rect 18002 75518 18004 75570
rect 17948 75460 18004 75518
rect 17500 74898 17668 74900
rect 17500 74846 17502 74898
rect 17554 74846 17668 74898
rect 17500 74844 17668 74846
rect 17724 75124 17780 75134
rect 17276 74676 17332 74686
rect 17276 74226 17332 74620
rect 17276 74174 17278 74226
rect 17330 74174 17332 74226
rect 17276 74162 17332 74174
rect 17500 73948 17556 74844
rect 17388 73892 17556 73948
rect 17276 73106 17332 73118
rect 17276 73054 17278 73106
rect 17330 73054 17332 73106
rect 17276 72548 17332 73054
rect 17276 72482 17332 72492
rect 17276 71540 17332 71550
rect 17276 71446 17332 71484
rect 17276 71316 17332 71326
rect 17276 70978 17332 71260
rect 17276 70926 17278 70978
rect 17330 70926 17332 70978
rect 17276 70914 17332 70926
rect 17388 70194 17444 73892
rect 17724 73444 17780 75068
rect 17948 73556 18004 75404
rect 18060 75124 18116 76190
rect 18222 76076 18486 76086
rect 18278 76020 18326 76076
rect 18382 76020 18430 76076
rect 18222 76010 18486 76020
rect 18284 75908 18340 75918
rect 18284 75906 18452 75908
rect 18284 75854 18286 75906
rect 18338 75854 18452 75906
rect 18284 75852 18452 75854
rect 18284 75842 18340 75852
rect 18284 75684 18340 75694
rect 18284 75590 18340 75628
rect 18060 75058 18116 75068
rect 18172 75458 18228 75470
rect 18172 75406 18174 75458
rect 18226 75406 18228 75458
rect 18172 75010 18228 75406
rect 18172 74958 18174 75010
rect 18226 74958 18228 75010
rect 18172 74946 18228 74958
rect 18396 74788 18452 75852
rect 18620 75124 18676 78542
rect 18732 77588 18788 79100
rect 18956 79042 19012 79100
rect 18956 78990 18958 79042
rect 19010 78990 19012 79042
rect 18956 78978 19012 78990
rect 19068 78930 19124 79324
rect 19068 78878 19070 78930
rect 19122 78878 19124 78930
rect 19068 78866 19124 78878
rect 19180 78484 19236 79438
rect 19292 78818 19348 79660
rect 19292 78766 19294 78818
rect 19346 78766 19348 78818
rect 19292 78596 19348 78766
rect 19292 78530 19348 78540
rect 18844 78372 18900 78382
rect 18844 78146 18900 78316
rect 18844 78094 18846 78146
rect 18898 78094 18900 78146
rect 18844 77812 18900 78094
rect 19180 78036 19236 78428
rect 18844 77746 18900 77756
rect 19068 77980 19236 78036
rect 18732 77532 18900 77588
rect 18620 75058 18676 75068
rect 18396 74732 18788 74788
rect 18620 74564 18676 74574
rect 18222 74508 18486 74518
rect 18278 74452 18326 74508
rect 18382 74452 18430 74508
rect 18222 74442 18486 74452
rect 18620 74338 18676 74508
rect 18620 74286 18622 74338
rect 18674 74286 18676 74338
rect 18620 74274 18676 74286
rect 17612 73388 17780 73444
rect 17836 73500 18004 73556
rect 18508 74228 18564 74238
rect 17500 73330 17556 73342
rect 17500 73278 17502 73330
rect 17554 73278 17556 73330
rect 17500 73220 17556 73278
rect 17500 73154 17556 73164
rect 17500 71988 17556 71998
rect 17500 71762 17556 71932
rect 17500 71710 17502 71762
rect 17554 71710 17556 71762
rect 17500 70644 17556 71710
rect 17500 70578 17556 70588
rect 17388 70142 17390 70194
rect 17442 70142 17444 70194
rect 17388 70130 17444 70142
rect 17612 69972 17668 73388
rect 17836 73332 17892 73500
rect 18060 73444 18116 73454
rect 18060 73350 18116 73388
rect 17276 69916 17668 69972
rect 17724 73276 17892 73332
rect 17948 73332 18004 73342
rect 17276 66836 17332 69916
rect 17388 69188 17444 69198
rect 17388 69094 17444 69132
rect 17388 68626 17444 68638
rect 17388 68574 17390 68626
rect 17442 68574 17444 68626
rect 17388 68516 17444 68574
rect 17612 68628 17668 68638
rect 17612 68534 17668 68572
rect 17388 68450 17444 68460
rect 17500 68514 17556 68526
rect 17500 68462 17502 68514
rect 17554 68462 17556 68514
rect 17500 67058 17556 68462
rect 17500 67006 17502 67058
rect 17554 67006 17556 67058
rect 17500 66994 17556 67006
rect 17612 67060 17668 67070
rect 17612 66966 17668 67004
rect 17276 66780 17668 66836
rect 17500 66274 17556 66286
rect 17500 66222 17502 66274
rect 17554 66222 17556 66274
rect 17500 66052 17556 66222
rect 17612 66162 17668 66780
rect 17612 66110 17614 66162
rect 17666 66110 17668 66162
rect 17612 66098 17668 66110
rect 17500 65986 17556 65996
rect 17276 65492 17332 65502
rect 17276 65398 17332 65436
rect 17500 65490 17556 65502
rect 17500 65438 17502 65490
rect 17554 65438 17556 65490
rect 17164 65100 17332 65156
rect 16940 64204 17108 64260
rect 17164 64930 17220 64942
rect 17164 64878 17166 64930
rect 17218 64878 17220 64930
rect 16828 63810 16884 63822
rect 16828 63758 16830 63810
rect 16882 63758 16884 63810
rect 16828 63364 16884 63758
rect 16828 62804 16884 63308
rect 16828 62738 16884 62748
rect 16828 62356 16884 62366
rect 16828 61908 16884 62300
rect 16828 61842 16884 61852
rect 16828 61570 16884 61582
rect 16828 61518 16830 61570
rect 16882 61518 16884 61570
rect 16828 61460 16884 61518
rect 16828 61394 16884 61404
rect 16940 61124 16996 64204
rect 17164 64148 17220 64878
rect 17276 64708 17332 65100
rect 17500 64930 17556 65438
rect 17724 65268 17780 73276
rect 17948 73238 18004 73276
rect 18284 73332 18340 73342
rect 18284 73238 18340 73276
rect 18508 73220 18564 74172
rect 18732 74226 18788 74732
rect 18732 74174 18734 74226
rect 18786 74174 18788 74226
rect 18732 74162 18788 74174
rect 18844 73948 18900 77532
rect 18956 76466 19012 76478
rect 18956 76414 18958 76466
rect 19010 76414 19012 76466
rect 18956 76356 19012 76414
rect 18956 76132 19012 76300
rect 18956 76066 19012 76076
rect 18956 74228 19012 74238
rect 18956 74114 19012 74172
rect 18956 74062 18958 74114
rect 19010 74062 19012 74114
rect 18956 74050 19012 74062
rect 19068 73948 19124 77980
rect 19292 77924 19348 77934
rect 19292 77830 19348 77868
rect 19180 77812 19236 77822
rect 19180 75794 19236 77756
rect 19180 75742 19182 75794
rect 19234 75742 19236 75794
rect 19180 74564 19236 75742
rect 19180 74498 19236 74508
rect 19292 74338 19348 74350
rect 19292 74286 19294 74338
rect 19346 74286 19348 74338
rect 19292 74228 19348 74286
rect 18844 73892 19012 73948
rect 19068 73892 19236 73948
rect 18732 73780 18788 73790
rect 18508 73164 18676 73220
rect 18222 72940 18486 72950
rect 18278 72884 18326 72940
rect 18382 72884 18430 72940
rect 18222 72874 18486 72884
rect 18620 72772 18676 73164
rect 18508 72716 18676 72772
rect 18732 73218 18788 73724
rect 18732 73166 18734 73218
rect 18786 73166 18788 73218
rect 17836 72660 17892 72670
rect 17836 71204 17892 72604
rect 18508 72434 18564 72716
rect 18508 72382 18510 72434
rect 18562 72382 18564 72434
rect 18508 72370 18564 72382
rect 18620 72548 18676 72558
rect 18732 72548 18788 73166
rect 18620 72546 18788 72548
rect 18620 72494 18622 72546
rect 18674 72494 18788 72546
rect 18620 72492 18788 72494
rect 18844 73668 18900 73678
rect 18620 71988 18676 72492
rect 18844 72212 18900 73612
rect 18956 72658 19012 73892
rect 19180 72772 19236 73892
rect 19292 73442 19348 74172
rect 19292 73390 19294 73442
rect 19346 73390 19348 73442
rect 19292 73378 19348 73390
rect 19404 73444 19460 80892
rect 19516 80612 19572 80622
rect 19516 79714 19572 80556
rect 19516 79662 19518 79714
rect 19570 79662 19572 79714
rect 19516 79650 19572 79662
rect 19628 79492 19684 83244
rect 19964 83524 20020 83534
rect 19964 82962 20020 83468
rect 19964 82910 19966 82962
rect 20018 82910 20020 82962
rect 19964 82898 20020 82910
rect 19852 82626 19908 82638
rect 19852 82574 19854 82626
rect 19906 82574 19908 82626
rect 19740 81730 19796 81742
rect 19740 81678 19742 81730
rect 19794 81678 19796 81730
rect 19740 81172 19796 81678
rect 19740 81106 19796 81116
rect 19852 80612 19908 82574
rect 20076 81732 20132 83916
rect 20188 83906 20244 83916
rect 20300 83636 20356 84252
rect 20188 83634 20356 83636
rect 20188 83582 20302 83634
rect 20354 83582 20356 83634
rect 20188 83580 20356 83582
rect 20188 81956 20244 83580
rect 20300 83570 20356 83580
rect 20412 84084 20468 84094
rect 20188 81862 20244 81900
rect 20300 83412 20356 83422
rect 20300 82738 20356 83356
rect 20300 82686 20302 82738
rect 20354 82686 20356 82738
rect 20300 81844 20356 82686
rect 20300 81778 20356 81788
rect 20076 81676 20244 81732
rect 19852 80546 19908 80556
rect 19964 81282 20020 81294
rect 19964 81230 19966 81282
rect 20018 81230 20020 81282
rect 19964 81172 20020 81230
rect 19964 80388 20020 81116
rect 20188 80610 20244 81676
rect 20188 80558 20190 80610
rect 20242 80558 20244 80610
rect 20188 80546 20244 80558
rect 19852 80386 20020 80388
rect 19852 80334 19966 80386
rect 20018 80334 20020 80386
rect 19852 80332 20020 80334
rect 19516 79436 19684 79492
rect 19740 79602 19796 79614
rect 19740 79550 19742 79602
rect 19794 79550 19796 79602
rect 19516 75348 19572 79436
rect 19740 79042 19796 79550
rect 19740 78990 19742 79042
rect 19794 78990 19796 79042
rect 19740 78978 19796 78990
rect 19628 78706 19684 78718
rect 19628 78654 19630 78706
rect 19682 78654 19684 78706
rect 19628 78596 19684 78654
rect 19740 78708 19796 78718
rect 19740 78614 19796 78652
rect 19628 78484 19684 78540
rect 19852 78484 19908 80332
rect 19964 80322 20020 80332
rect 19964 79716 20020 79726
rect 19964 79490 20020 79660
rect 19964 79438 19966 79490
rect 20018 79438 20020 79490
rect 19964 79426 20020 79438
rect 20188 78820 20244 78830
rect 20188 78726 20244 78764
rect 19628 78428 19908 78484
rect 19740 78036 19796 78046
rect 19740 77942 19796 77980
rect 19628 76354 19684 76366
rect 19628 76302 19630 76354
rect 19682 76302 19684 76354
rect 19628 75796 19684 76302
rect 19740 75796 19796 75806
rect 19628 75794 19796 75796
rect 19628 75742 19742 75794
rect 19794 75742 19796 75794
rect 19628 75740 19796 75742
rect 19740 75730 19796 75740
rect 19628 75572 19684 75582
rect 19628 75478 19684 75516
rect 19516 75292 19684 75348
rect 19516 74004 19572 74042
rect 19516 73938 19572 73948
rect 19404 73388 19572 73444
rect 18956 72606 18958 72658
rect 19010 72606 19012 72658
rect 18956 72594 19012 72606
rect 19068 72716 19236 72772
rect 19404 73106 19460 73118
rect 19404 73054 19406 73106
rect 19458 73054 19460 73106
rect 18620 71922 18676 71932
rect 18732 72156 18900 72212
rect 18956 72436 19012 72446
rect 18060 71876 18116 71886
rect 17948 71762 18004 71774
rect 17948 71710 17950 71762
rect 18002 71710 18004 71762
rect 17948 71428 18004 71710
rect 17948 71362 18004 71372
rect 18060 71762 18116 71820
rect 18060 71710 18062 71762
rect 18114 71710 18116 71762
rect 17948 71204 18004 71214
rect 17836 71148 17948 71204
rect 17948 71138 18004 71148
rect 17948 70866 18004 70878
rect 17948 70814 17950 70866
rect 18002 70814 18004 70866
rect 17836 70754 17892 70766
rect 17836 70702 17838 70754
rect 17890 70702 17892 70754
rect 17836 69412 17892 70702
rect 17836 69346 17892 69356
rect 17836 69186 17892 69198
rect 17836 69134 17838 69186
rect 17890 69134 17892 69186
rect 17836 68964 17892 69134
rect 17836 68898 17892 68908
rect 17948 68852 18004 70814
rect 18060 70644 18116 71710
rect 18284 71652 18340 71662
rect 18284 71558 18340 71596
rect 18222 71372 18486 71382
rect 18278 71316 18326 71372
rect 18382 71316 18430 71372
rect 18222 71306 18486 71316
rect 18396 70866 18452 70878
rect 18396 70814 18398 70866
rect 18450 70814 18452 70866
rect 18284 70756 18340 70766
rect 18284 70662 18340 70700
rect 18172 70644 18228 70654
rect 18060 70588 18172 70644
rect 18172 70578 18228 70588
rect 18396 70308 18452 70814
rect 18732 70588 18788 72156
rect 18844 71988 18900 71998
rect 18956 71988 19012 72380
rect 19068 72324 19124 72716
rect 19180 72548 19236 72558
rect 19180 72454 19236 72492
rect 19068 72268 19236 72324
rect 18844 71986 19012 71988
rect 18844 71934 18846 71986
rect 18898 71934 19012 71986
rect 18844 71932 19012 71934
rect 19068 71988 19124 71998
rect 18844 71922 18900 71932
rect 19068 71762 19124 71932
rect 19068 71710 19070 71762
rect 19122 71710 19124 71762
rect 18844 71204 18900 71214
rect 18844 71090 18900 71148
rect 18844 71038 18846 71090
rect 18898 71038 18900 71090
rect 18844 71026 18900 71038
rect 19068 70980 19124 71710
rect 19068 70914 19124 70924
rect 19068 70644 19124 70654
rect 18732 70532 18900 70588
rect 18396 70242 18452 70252
rect 18172 70084 18228 70094
rect 18172 70082 18676 70084
rect 18172 70030 18174 70082
rect 18226 70030 18676 70082
rect 18172 70028 18676 70030
rect 18172 70018 18228 70028
rect 18222 69804 18486 69814
rect 18278 69748 18326 69804
rect 18382 69748 18430 69804
rect 18222 69738 18486 69748
rect 18284 69410 18340 69422
rect 18284 69358 18286 69410
rect 18338 69358 18340 69410
rect 18284 69076 18340 69358
rect 18620 69186 18676 70028
rect 18732 69300 18788 69310
rect 18732 69206 18788 69244
rect 18620 69134 18622 69186
rect 18674 69134 18676 69186
rect 18620 69122 18676 69134
rect 18284 69010 18340 69020
rect 17948 68786 18004 68796
rect 17836 68740 17892 68750
rect 17836 68646 17892 68684
rect 18508 68516 18564 68526
rect 18508 68514 18676 68516
rect 18508 68462 18510 68514
rect 18562 68462 18676 68514
rect 18508 68460 18676 68462
rect 18508 68450 18564 68460
rect 18222 68236 18486 68246
rect 18278 68180 18326 68236
rect 18382 68180 18430 68236
rect 18222 68170 18486 68180
rect 18172 67732 18228 67742
rect 17836 67730 18228 67732
rect 17836 67678 18174 67730
rect 18226 67678 18228 67730
rect 17836 67676 18228 67678
rect 17836 67282 17892 67676
rect 18172 67666 18228 67676
rect 17836 67230 17838 67282
rect 17890 67230 17892 67282
rect 17836 67218 17892 67230
rect 18060 67396 18116 67406
rect 17948 67172 18004 67182
rect 17948 67078 18004 67116
rect 17836 66948 17892 66958
rect 18060 66948 18116 67340
rect 18620 67172 18676 68460
rect 18732 67956 18788 67966
rect 18732 67282 18788 67900
rect 18732 67230 18734 67282
rect 18786 67230 18788 67282
rect 18732 67218 18788 67230
rect 18620 67106 18676 67116
rect 18396 67060 18452 67070
rect 18844 67060 18900 70532
rect 18956 69524 19012 69534
rect 18956 69410 19012 69468
rect 18956 69358 18958 69410
rect 19010 69358 19012 69410
rect 18956 69346 19012 69358
rect 19068 68852 19124 70588
rect 19180 70532 19236 72268
rect 19404 71874 19460 73054
rect 19516 72548 19572 73388
rect 19516 72482 19572 72492
rect 19516 72324 19572 72334
rect 19516 72230 19572 72268
rect 19404 71822 19406 71874
rect 19458 71822 19460 71874
rect 19404 71810 19460 71822
rect 19292 71540 19348 71550
rect 19292 70978 19348 71484
rect 19292 70926 19294 70978
rect 19346 70926 19348 70978
rect 19292 70914 19348 70926
rect 19516 70756 19572 70766
rect 19516 70662 19572 70700
rect 19628 70754 19684 75292
rect 19852 74564 19908 78428
rect 20188 78148 20244 78158
rect 20412 78148 20468 84028
rect 20524 82738 20580 84252
rect 20636 84476 20916 84532
rect 20636 83300 20692 84476
rect 20860 84306 20916 84318
rect 20860 84254 20862 84306
rect 20914 84254 20916 84306
rect 20748 84196 20804 84206
rect 20860 84196 20916 84254
rect 20972 84308 21028 85260
rect 20972 84242 21028 84252
rect 21084 84306 21140 86604
rect 21196 86548 21252 87276
rect 21308 87266 21364 87276
rect 21756 87330 21812 87342
rect 21756 87278 21758 87330
rect 21810 87278 21812 87330
rect 21756 87220 21812 87278
rect 21756 87218 21924 87220
rect 21756 87166 21758 87218
rect 21810 87166 21924 87218
rect 21756 87164 21924 87166
rect 21756 87154 21812 87164
rect 21196 86482 21252 86492
rect 21308 86658 21364 86670
rect 21308 86606 21310 86658
rect 21362 86606 21364 86658
rect 21308 85204 21364 86606
rect 21868 86658 21924 87164
rect 22764 86884 22820 88734
rect 22764 86818 22820 86828
rect 22876 89236 22932 89246
rect 22876 86772 22932 89180
rect 22988 88450 23044 89292
rect 23324 89348 23380 89358
rect 23436 89348 23492 90302
rect 23380 89292 23492 89348
rect 23324 89282 23380 89292
rect 23212 89236 23268 89246
rect 23212 89124 23268 89180
rect 23324 89124 23380 89134
rect 23212 89122 23380 89124
rect 23212 89070 23326 89122
rect 23378 89070 23380 89122
rect 23212 89068 23380 89070
rect 23324 89058 23380 89068
rect 23548 89012 23604 89022
rect 23548 88918 23604 88956
rect 23884 88788 23940 90860
rect 24220 89794 24276 89806
rect 24220 89742 24222 89794
rect 24274 89742 24276 89794
rect 23996 89682 24052 89694
rect 23996 89630 23998 89682
rect 24050 89630 24052 89682
rect 23996 89012 24052 89630
rect 24108 89570 24164 89582
rect 24108 89518 24110 89570
rect 24162 89518 24164 89570
rect 24108 89124 24164 89518
rect 24220 89348 24276 89742
rect 24220 89282 24276 89292
rect 24108 89058 24164 89068
rect 23996 88946 24052 88956
rect 24332 88900 24388 91084
rect 24556 91252 24612 91262
rect 24556 89794 24612 91196
rect 25116 91250 25172 91262
rect 25116 91198 25118 91250
rect 25170 91198 25172 91250
rect 25116 90804 25172 91198
rect 25228 91138 25284 91532
rect 25228 91086 25230 91138
rect 25282 91086 25284 91138
rect 25228 90916 25284 91086
rect 25452 90916 25508 91980
rect 25564 91700 25620 95228
rect 25676 95282 25732 95294
rect 25676 95230 25678 95282
rect 25730 95230 25732 95282
rect 25676 94612 25732 95230
rect 25788 94612 25844 94622
rect 25676 94610 25844 94612
rect 25676 94558 25790 94610
rect 25842 94558 25844 94610
rect 25676 94556 25844 94558
rect 25788 94546 25844 94556
rect 25900 94164 25956 96014
rect 26236 95844 26292 96684
rect 26236 95750 26292 95788
rect 27132 95844 27188 95854
rect 26012 95284 26068 95294
rect 26012 95190 26068 95228
rect 25900 94098 25956 94108
rect 26908 94164 26964 94174
rect 26908 93938 26964 94108
rect 26908 93886 26910 93938
rect 26962 93886 26964 93938
rect 25788 93042 25844 93054
rect 25788 92990 25790 93042
rect 25842 92990 25844 93042
rect 25788 92932 25844 92990
rect 26124 93044 26180 93054
rect 26124 92932 26180 92988
rect 26236 92932 26292 92942
rect 26124 92930 26292 92932
rect 26124 92878 26238 92930
rect 26290 92878 26292 92930
rect 26124 92876 26292 92878
rect 25788 92866 25844 92876
rect 26236 92866 26292 92876
rect 26348 92932 26404 92942
rect 26348 92838 26404 92876
rect 26572 92930 26628 92942
rect 26572 92878 26574 92930
rect 26626 92878 26628 92930
rect 25676 92708 25732 92718
rect 26012 92708 26068 92718
rect 26236 92708 26292 92718
rect 26572 92708 26628 92878
rect 25676 92706 25956 92708
rect 25676 92654 25678 92706
rect 25730 92654 25956 92706
rect 25676 92652 25956 92654
rect 25676 92642 25732 92652
rect 25788 92484 25844 92494
rect 25788 92148 25844 92428
rect 25564 91634 25620 91644
rect 25676 92034 25732 92046
rect 25676 91982 25678 92034
rect 25730 91982 25732 92034
rect 25676 91588 25732 91982
rect 25676 91522 25732 91532
rect 25564 91364 25620 91374
rect 25564 91270 25620 91308
rect 25788 91364 25844 92092
rect 25788 91298 25844 91308
rect 25676 91250 25732 91262
rect 25676 91198 25678 91250
rect 25730 91198 25732 91250
rect 25676 91140 25732 91198
rect 25900 91140 25956 92652
rect 26068 92652 26180 92708
rect 26012 92642 26068 92652
rect 26124 92148 26180 92652
rect 26236 92706 26516 92708
rect 26236 92654 26238 92706
rect 26290 92654 26516 92706
rect 26236 92652 26516 92654
rect 26236 92642 26292 92652
rect 26236 92148 26292 92158
rect 26124 92146 26404 92148
rect 26124 92094 26238 92146
rect 26290 92094 26404 92146
rect 26124 92092 26404 92094
rect 26236 92082 26292 92092
rect 26012 92036 26068 92046
rect 26012 91588 26068 91980
rect 26124 91588 26180 91598
rect 26012 91586 26180 91588
rect 26012 91534 26126 91586
rect 26178 91534 26180 91586
rect 26012 91532 26180 91534
rect 26124 91522 26180 91532
rect 26348 91586 26404 92092
rect 26460 92146 26516 92652
rect 26572 92642 26628 92652
rect 26908 92484 26964 93886
rect 27132 93714 27188 95788
rect 28140 95396 28196 114212
rect 28252 113090 28308 113102
rect 28252 113038 28254 113090
rect 28306 113038 28308 113090
rect 28252 112754 28308 113038
rect 28428 112924 28692 112934
rect 28484 112868 28532 112924
rect 28588 112868 28636 112924
rect 28428 112858 28692 112868
rect 28252 112702 28254 112754
rect 28306 112702 28308 112754
rect 28252 111972 28308 112702
rect 28252 111186 28308 111916
rect 28428 111356 28692 111366
rect 28484 111300 28532 111356
rect 28588 111300 28636 111356
rect 28428 111290 28692 111300
rect 28252 111134 28254 111186
rect 28306 111134 28308 111186
rect 28252 110290 28308 111134
rect 28252 110238 28254 110290
rect 28306 110238 28308 110290
rect 28252 109618 28308 110238
rect 28428 109788 28692 109798
rect 28484 109732 28532 109788
rect 28588 109732 28636 109788
rect 28428 109722 28692 109732
rect 28252 109566 28254 109618
rect 28306 109566 28308 109618
rect 28252 108388 28308 109566
rect 28252 108050 28308 108332
rect 28428 108220 28692 108230
rect 28484 108164 28532 108220
rect 28588 108164 28636 108220
rect 28428 108154 28692 108164
rect 28252 107998 28254 108050
rect 28306 107998 28308 108050
rect 28252 107154 28308 107998
rect 28252 107102 28254 107154
rect 28306 107102 28308 107154
rect 28252 106482 28308 107102
rect 28428 106652 28692 106662
rect 28484 106596 28532 106652
rect 28588 106596 28636 106652
rect 28428 106586 28692 106596
rect 28252 106430 28254 106482
rect 28306 106430 28308 106482
rect 28252 105588 28308 106430
rect 28252 105522 28308 105532
rect 28428 105084 28692 105094
rect 28484 105028 28532 105084
rect 28588 105028 28636 105084
rect 28428 105018 28692 105028
rect 28428 103516 28692 103526
rect 28484 103460 28532 103516
rect 28588 103460 28636 103516
rect 28428 103450 28692 103460
rect 28428 101948 28692 101958
rect 28484 101892 28532 101948
rect 28588 101892 28636 101948
rect 28428 101882 28692 101892
rect 28428 100380 28692 100390
rect 28484 100324 28532 100380
rect 28588 100324 28636 100380
rect 28428 100314 28692 100324
rect 28428 98812 28692 98822
rect 28484 98756 28532 98812
rect 28588 98756 28636 98812
rect 28428 98746 28692 98756
rect 28428 97244 28692 97254
rect 28484 97188 28532 97244
rect 28588 97188 28636 97244
rect 28428 97178 28692 97188
rect 28428 95676 28692 95686
rect 28484 95620 28532 95676
rect 28588 95620 28636 95676
rect 28428 95610 28692 95620
rect 28140 95330 28196 95340
rect 27132 93662 27134 93714
rect 27186 93662 27188 93714
rect 27132 93604 27188 93662
rect 28028 94274 28084 94286
rect 28028 94222 28030 94274
rect 28082 94222 28084 94274
rect 27804 93604 27860 93614
rect 28028 93604 28084 94222
rect 28428 94108 28692 94118
rect 28484 94052 28532 94108
rect 28588 94052 28636 94108
rect 28428 94042 28692 94052
rect 27132 93602 28196 93604
rect 27132 93550 27806 93602
rect 27858 93550 28196 93602
rect 27132 93548 28196 93550
rect 27804 93538 27860 93548
rect 27132 92818 27188 92830
rect 27132 92766 27134 92818
rect 27186 92766 27188 92818
rect 26460 92094 26462 92146
rect 26514 92094 26516 92146
rect 26460 92082 26516 92094
rect 26572 92428 26964 92484
rect 27020 92706 27076 92718
rect 27020 92654 27022 92706
rect 27074 92654 27076 92706
rect 27020 92484 27076 92654
rect 26348 91534 26350 91586
rect 26402 91534 26404 91586
rect 26348 91522 26404 91534
rect 26460 91588 26516 91598
rect 26572 91588 26628 92428
rect 27020 92418 27076 92428
rect 27132 92484 27188 92766
rect 27132 92428 28084 92484
rect 26796 92260 26852 92270
rect 27132 92260 27188 92428
rect 26796 92258 27188 92260
rect 26796 92206 26798 92258
rect 26850 92206 27188 92258
rect 26796 92204 27188 92206
rect 26796 92194 26852 92204
rect 27356 92148 27412 92158
rect 26908 92146 27412 92148
rect 26908 92094 27358 92146
rect 27410 92094 27412 92146
rect 26908 92092 27412 92094
rect 26684 92034 26740 92046
rect 26684 91982 26686 92034
rect 26738 91982 26740 92034
rect 26684 91924 26740 91982
rect 26684 91858 26740 91868
rect 26908 91812 26964 92092
rect 27356 92082 27412 92092
rect 27580 92146 27636 92158
rect 27580 92094 27582 92146
rect 27634 92094 27636 92146
rect 27468 92034 27524 92046
rect 27468 91982 27470 92034
rect 27522 91982 27524 92034
rect 27020 91924 27076 91934
rect 27468 91924 27524 91982
rect 27020 91922 27524 91924
rect 27020 91870 27022 91922
rect 27074 91870 27524 91922
rect 27020 91868 27524 91870
rect 27020 91858 27076 91868
rect 26908 91746 26964 91756
rect 27244 91588 27300 91598
rect 27580 91588 27636 92094
rect 26572 91532 27076 91588
rect 26460 91494 26516 91532
rect 26908 91364 26964 91374
rect 26908 91270 26964 91308
rect 26012 91252 26068 91262
rect 26012 91158 26068 91196
rect 25732 91084 25956 91140
rect 25676 91074 25732 91084
rect 25228 90860 25508 90916
rect 25116 90738 25172 90748
rect 25026 90188 25290 90198
rect 25082 90132 25130 90188
rect 25186 90132 25234 90188
rect 25026 90122 25290 90132
rect 24556 89742 24558 89794
rect 24610 89742 24612 89794
rect 24556 89730 24612 89742
rect 24892 89684 24948 89694
rect 24668 89682 24948 89684
rect 24668 89630 24894 89682
rect 24946 89630 24948 89682
rect 24668 89628 24948 89630
rect 23996 88788 24052 88798
rect 22988 88398 22990 88450
rect 23042 88398 23044 88450
rect 22988 88386 23044 88398
rect 23212 88786 24052 88788
rect 23212 88734 23998 88786
rect 24050 88734 24052 88786
rect 23212 88732 24052 88734
rect 23212 88338 23268 88732
rect 23996 88722 24052 88732
rect 24332 88786 24388 88844
rect 24556 89236 24612 89246
rect 24556 88900 24612 89180
rect 24556 88806 24612 88844
rect 24332 88734 24334 88786
rect 24386 88734 24388 88786
rect 24332 88452 24388 88734
rect 24332 88386 24388 88396
rect 23212 88286 23214 88338
rect 23266 88286 23268 88338
rect 23212 88274 23268 88286
rect 24556 88228 24612 88238
rect 24556 88134 24612 88172
rect 24108 88116 24164 88126
rect 24108 87442 24164 88060
rect 24668 87554 24724 89628
rect 24892 89618 24948 89628
rect 25116 89460 25172 89470
rect 25452 89460 25508 90860
rect 26012 91028 26068 91038
rect 25788 90468 25844 90478
rect 25788 89684 25844 90412
rect 25172 89404 25508 89460
rect 25564 89572 25620 89582
rect 25116 89010 25172 89404
rect 25564 89122 25620 89516
rect 25564 89070 25566 89122
rect 25618 89070 25620 89122
rect 25116 88958 25118 89010
rect 25170 88958 25172 89010
rect 25116 88946 25172 88958
rect 25340 89012 25396 89022
rect 25340 88918 25396 88956
rect 25564 88900 25620 89070
rect 25788 89010 25844 89628
rect 26012 89572 26068 90972
rect 26348 90580 26404 90590
rect 26012 89478 26068 89516
rect 26124 89794 26180 89806
rect 26124 89742 26126 89794
rect 26178 89742 26180 89794
rect 25788 88958 25790 89010
rect 25842 88958 25844 89010
rect 25788 88946 25844 88958
rect 25564 88834 25620 88844
rect 25026 88620 25290 88630
rect 25082 88564 25130 88620
rect 25186 88564 25234 88620
rect 25026 88554 25290 88564
rect 24780 88452 24836 88462
rect 24780 88358 24836 88396
rect 25004 88226 25060 88238
rect 25004 88174 25006 88226
rect 25058 88174 25060 88226
rect 25004 88116 25060 88174
rect 25004 88050 25060 88060
rect 26124 87668 26180 89742
rect 26348 89010 26404 90524
rect 27020 90578 27076 91532
rect 27244 91586 27636 91588
rect 27244 91534 27246 91586
rect 27298 91534 27636 91586
rect 27244 91532 27636 91534
rect 28028 92146 28084 92428
rect 28028 92094 28030 92146
rect 28082 92094 28084 92146
rect 27244 91522 27300 91532
rect 27132 91140 27188 91150
rect 27132 91046 27188 91084
rect 27020 90526 27022 90578
rect 27074 90526 27076 90578
rect 27020 89794 27076 90526
rect 27580 90580 27636 90590
rect 27580 90486 27636 90524
rect 28028 90468 28084 92094
rect 28140 91588 28196 93548
rect 28428 92540 28692 92550
rect 28484 92484 28532 92540
rect 28588 92484 28636 92540
rect 28428 92474 28692 92484
rect 28140 91474 28196 91532
rect 28140 91422 28142 91474
rect 28194 91422 28196 91474
rect 28140 90748 28196 91422
rect 28428 90972 28692 90982
rect 28484 90916 28532 90972
rect 28588 90916 28636 90972
rect 28428 90906 28692 90916
rect 28140 90692 28308 90748
rect 28028 90374 28084 90412
rect 27020 89742 27022 89794
rect 27074 89742 27076 89794
rect 27020 89684 27076 89742
rect 27020 89618 27076 89628
rect 27132 90354 27188 90366
rect 27132 90302 27134 90354
rect 27186 90302 27188 90354
rect 27132 89124 27188 90302
rect 26348 88958 26350 89010
rect 26402 88958 26404 89010
rect 26348 88946 26404 88958
rect 26796 89122 27188 89124
rect 26796 89070 27134 89122
rect 27186 89070 27188 89122
rect 26796 89068 27188 89070
rect 26236 88898 26292 88910
rect 26236 88846 26238 88898
rect 26290 88846 26292 88898
rect 26236 88340 26292 88846
rect 26236 88284 26404 88340
rect 24668 87502 24670 87554
rect 24722 87502 24724 87554
rect 24668 87490 24724 87502
rect 25676 87666 26180 87668
rect 25676 87614 26126 87666
rect 26178 87614 26180 87666
rect 25676 87612 26180 87614
rect 24108 87390 24110 87442
rect 24162 87390 24164 87442
rect 23996 86884 24052 86894
rect 23996 86790 24052 86828
rect 22876 86716 23044 86772
rect 21868 86606 21870 86658
rect 21922 86606 21924 86658
rect 21868 86594 21924 86606
rect 21980 86548 22036 86558
rect 21532 86436 21588 86474
rect 21980 86454 22036 86492
rect 22876 86548 22932 86558
rect 22876 86454 22932 86492
rect 21532 86370 21588 86380
rect 21624 86268 21888 86278
rect 21680 86212 21728 86268
rect 21784 86212 21832 86268
rect 21624 86202 21888 86212
rect 22988 85986 23044 86716
rect 24108 86770 24164 87390
rect 24108 86718 24110 86770
rect 24162 86718 24164 86770
rect 24108 86706 24164 86718
rect 24332 87330 24388 87342
rect 24332 87278 24334 87330
rect 24386 87278 24388 87330
rect 24332 86772 24388 87278
rect 24332 86706 24388 86716
rect 24444 87332 24500 87342
rect 22988 85934 22990 85986
rect 23042 85934 23044 85986
rect 22988 85708 23044 85934
rect 23548 86660 23604 86670
rect 22988 85652 23156 85708
rect 22988 85314 23044 85326
rect 22988 85262 22990 85314
rect 23042 85262 23044 85314
rect 21084 84254 21086 84306
rect 21138 84254 21140 84306
rect 21084 84242 21140 84254
rect 21196 85148 21364 85204
rect 21980 85204 22036 85214
rect 21980 85202 22148 85204
rect 21980 85150 21982 85202
rect 22034 85150 22148 85202
rect 21980 85148 22148 85150
rect 20804 84140 20916 84196
rect 20748 84130 20804 84140
rect 21196 84084 21252 85148
rect 21980 85138 22036 85148
rect 21308 84980 21364 84990
rect 21308 84886 21364 84924
rect 21420 84866 21476 84878
rect 21420 84814 21422 84866
rect 21474 84814 21476 84866
rect 21420 84532 21476 84814
rect 21624 84700 21888 84710
rect 21680 84644 21728 84700
rect 21784 84644 21832 84700
rect 21624 84634 21888 84644
rect 21420 84476 21812 84532
rect 21308 84420 21364 84430
rect 21308 84196 21364 84364
rect 21756 84306 21812 84476
rect 21756 84254 21758 84306
rect 21810 84254 21812 84306
rect 21756 84242 21812 84254
rect 21420 84196 21476 84206
rect 21308 84194 21476 84196
rect 21308 84142 21422 84194
rect 21474 84142 21476 84194
rect 21308 84140 21476 84142
rect 21420 84130 21476 84140
rect 21196 84018 21252 84028
rect 21532 84084 21588 84094
rect 20748 83748 20804 83758
rect 20748 83522 20804 83692
rect 21532 83634 21588 84028
rect 21532 83582 21534 83634
rect 21586 83582 21588 83634
rect 21532 83570 21588 83582
rect 21644 83972 21700 83982
rect 20748 83470 20750 83522
rect 20802 83470 20804 83522
rect 20748 83458 20804 83470
rect 21308 83410 21364 83422
rect 21308 83358 21310 83410
rect 21362 83358 21364 83410
rect 21308 83300 21364 83358
rect 21532 83300 21588 83310
rect 21644 83300 21700 83916
rect 21980 83524 22036 83534
rect 21980 83430 22036 83468
rect 20636 83244 21140 83300
rect 20524 82686 20526 82738
rect 20578 82686 20580 82738
rect 20524 82674 20580 82686
rect 20860 83076 20916 83086
rect 20524 81844 20580 81854
rect 20524 81058 20580 81788
rect 20636 81730 20692 81742
rect 20636 81678 20638 81730
rect 20690 81678 20692 81730
rect 20636 81284 20692 81678
rect 20748 81732 20804 81742
rect 20748 81638 20804 81676
rect 20636 81218 20692 81228
rect 20748 81396 20804 81406
rect 20748 81170 20804 81340
rect 20748 81118 20750 81170
rect 20802 81118 20804 81170
rect 20748 81106 20804 81118
rect 20524 81006 20526 81058
rect 20578 81006 20580 81058
rect 20524 80994 20580 81006
rect 20524 80276 20580 80286
rect 20524 80182 20580 80220
rect 20860 79716 20916 83020
rect 21084 82852 21140 83244
rect 21308 83234 21364 83244
rect 21420 83298 21700 83300
rect 21420 83246 21534 83298
rect 21586 83246 21700 83298
rect 21420 83244 21700 83246
rect 21084 82758 21140 82796
rect 21308 81954 21364 81966
rect 21308 81902 21310 81954
rect 21362 81902 21364 81954
rect 21308 81844 21364 81902
rect 21308 81778 21364 81788
rect 21308 80386 21364 80398
rect 21308 80334 21310 80386
rect 21362 80334 21364 80386
rect 21196 80276 21252 80286
rect 21308 80276 21364 80334
rect 21252 80220 21364 80276
rect 21196 80210 21252 80220
rect 20860 79650 20916 79660
rect 21420 80164 21476 83244
rect 21532 83234 21588 83244
rect 21624 83132 21888 83142
rect 21680 83076 21728 83132
rect 21784 83076 21832 83132
rect 22092 83076 22148 85148
rect 22316 85090 22372 85102
rect 22316 85038 22318 85090
rect 22370 85038 22372 85090
rect 22316 84644 22372 85038
rect 22764 84978 22820 84990
rect 22764 84926 22766 84978
rect 22818 84926 22820 84978
rect 22316 84588 22596 84644
rect 22540 84306 22596 84588
rect 22540 84254 22542 84306
rect 22594 84254 22596 84306
rect 22540 83636 22596 84254
rect 22652 84194 22708 84206
rect 22652 84142 22654 84194
rect 22706 84142 22708 84194
rect 22652 83860 22708 84142
rect 22764 83972 22820 84926
rect 22764 83906 22820 83916
rect 22876 84868 22932 84878
rect 22876 84418 22932 84812
rect 22876 84366 22878 84418
rect 22930 84366 22932 84418
rect 22652 83794 22708 83804
rect 22652 83636 22708 83646
rect 22540 83580 22652 83636
rect 22652 83542 22708 83580
rect 21624 83066 21888 83076
rect 21980 83020 22148 83076
rect 22428 83524 22484 83534
rect 21980 82178 22036 83020
rect 22092 82852 22148 82862
rect 22092 82758 22148 82796
rect 21980 82126 21982 82178
rect 22034 82126 22036 82178
rect 21532 81956 21588 81966
rect 21532 81862 21588 81900
rect 21980 81732 22036 82126
rect 21624 81564 21888 81574
rect 21680 81508 21728 81564
rect 21784 81508 21832 81564
rect 21624 81498 21888 81508
rect 21644 81170 21700 81182
rect 21644 81118 21646 81170
rect 21698 81118 21700 81170
rect 21644 80610 21700 81118
rect 21980 81172 22036 81676
rect 22428 81172 22484 83468
rect 22764 83524 22820 83534
rect 22876 83524 22932 84366
rect 22764 83522 22932 83524
rect 22764 83470 22766 83522
rect 22818 83470 22932 83522
rect 22764 83468 22932 83470
rect 22540 82740 22596 82750
rect 22764 82740 22820 83468
rect 22988 82740 23044 85262
rect 22540 82738 22820 82740
rect 22540 82686 22542 82738
rect 22594 82686 22820 82738
rect 22540 82684 22820 82686
rect 22876 82684 23044 82740
rect 22540 81956 22596 82684
rect 22540 81890 22596 81900
rect 22652 81844 22708 81854
rect 22652 81282 22708 81788
rect 22876 81620 22932 82684
rect 22764 81564 22932 81620
rect 22988 82516 23044 82526
rect 22764 81396 22820 81564
rect 22764 81330 22820 81340
rect 22876 81396 22932 81406
rect 22988 81396 23044 82460
rect 22876 81394 23044 81396
rect 22876 81342 22878 81394
rect 22930 81342 23044 81394
rect 22876 81340 23044 81342
rect 22876 81330 22932 81340
rect 22652 81230 22654 81282
rect 22706 81230 22708 81282
rect 22652 81218 22708 81230
rect 22540 81172 22596 81182
rect 22428 81170 22596 81172
rect 22428 81118 22542 81170
rect 22594 81118 22596 81170
rect 22428 81116 22596 81118
rect 21980 81106 22036 81116
rect 21644 80558 21646 80610
rect 21698 80558 21700 80610
rect 21644 80546 21700 80558
rect 22540 80612 22596 81116
rect 22988 81172 23044 81182
rect 22988 81078 23044 81116
rect 22092 80500 22148 80510
rect 22092 80386 22148 80444
rect 22092 80334 22094 80386
rect 22146 80334 22148 80386
rect 21532 80164 21588 80174
rect 21420 80162 21588 80164
rect 21420 80110 21534 80162
rect 21586 80110 21588 80162
rect 21420 80108 21588 80110
rect 21084 79604 21140 79614
rect 21420 79604 21476 80108
rect 21532 80098 21588 80108
rect 22092 80052 22148 80334
rect 22428 80276 22484 80286
rect 21624 79996 21888 80006
rect 21680 79940 21728 79996
rect 21784 79940 21832 79996
rect 22092 79986 22148 79996
rect 22316 80274 22484 80276
rect 22316 80222 22430 80274
rect 22482 80222 22484 80274
rect 22316 80220 22484 80222
rect 21624 79930 21888 79940
rect 21532 79604 21588 79614
rect 21084 79602 21252 79604
rect 21084 79550 21086 79602
rect 21138 79550 21252 79602
rect 21084 79548 21252 79550
rect 21420 79548 21532 79604
rect 21084 79538 21140 79548
rect 21196 78932 21252 79548
rect 21420 78932 21476 78942
rect 21196 78930 21476 78932
rect 21196 78878 21422 78930
rect 21474 78878 21476 78930
rect 21196 78876 21476 78878
rect 21420 78866 21476 78876
rect 20188 78146 20468 78148
rect 20188 78094 20190 78146
rect 20242 78094 20468 78146
rect 20188 78092 20468 78094
rect 20524 78706 20580 78718
rect 20524 78654 20526 78706
rect 20578 78654 20580 78706
rect 20188 77140 20244 78092
rect 20412 77812 20468 77822
rect 20412 77474 20468 77756
rect 20412 77422 20414 77474
rect 20466 77422 20468 77474
rect 20412 77410 20468 77422
rect 20524 77364 20580 78654
rect 21308 78706 21364 78718
rect 21308 78654 21310 78706
rect 21362 78654 21364 78706
rect 21308 78484 21364 78654
rect 21532 78596 21588 79548
rect 21868 79602 21924 79614
rect 21868 79550 21870 79602
rect 21922 79550 21924 79602
rect 21868 78708 21924 79550
rect 21868 78642 21924 78652
rect 21532 78530 21588 78540
rect 22092 78596 22148 78606
rect 21308 78418 21364 78428
rect 21624 78428 21888 78438
rect 21680 78372 21728 78428
rect 21784 78372 21832 78428
rect 21624 78362 21888 78372
rect 21868 78034 21924 78046
rect 21868 77982 21870 78034
rect 21922 77982 21924 78034
rect 20636 77922 20692 77934
rect 20636 77870 20638 77922
rect 20690 77870 20692 77922
rect 20636 77810 20692 77870
rect 20636 77758 20638 77810
rect 20690 77758 20692 77810
rect 20636 77476 20692 77758
rect 20636 77410 20692 77420
rect 21084 77922 21140 77934
rect 21084 77870 21086 77922
rect 21138 77870 21140 77922
rect 20524 77298 20580 77308
rect 21084 77252 21140 77870
rect 21084 77186 21140 77196
rect 21420 77810 21476 77822
rect 21420 77758 21422 77810
rect 21474 77758 21476 77810
rect 21420 77362 21476 77758
rect 21420 77310 21422 77362
rect 21474 77310 21476 77362
rect 21420 77252 21476 77310
rect 20188 77074 20244 77084
rect 19964 77028 20020 77038
rect 19964 75682 20020 76972
rect 20524 77026 20580 77038
rect 20524 76974 20526 77026
rect 20578 76974 20580 77026
rect 20524 76916 20580 76974
rect 20188 76860 20580 76916
rect 20636 77026 20692 77038
rect 20636 76974 20638 77026
rect 20690 76974 20692 77026
rect 20188 75906 20244 76860
rect 20636 76356 20692 76974
rect 21420 76580 21476 77196
rect 21868 77028 21924 77982
rect 22092 77812 22148 78540
rect 21980 77252 22036 77262
rect 21980 77158 22036 77196
rect 21868 76972 22036 77028
rect 21624 76860 21888 76870
rect 21680 76804 21728 76860
rect 21784 76804 21832 76860
rect 21624 76794 21888 76804
rect 21420 76524 21924 76580
rect 20636 76290 20692 76300
rect 21420 76356 21476 76366
rect 20188 75854 20190 75906
rect 20242 75854 20244 75906
rect 20188 75842 20244 75854
rect 20748 75796 20804 75806
rect 19964 75630 19966 75682
rect 20018 75630 20020 75682
rect 19964 74788 20020 75630
rect 20188 75684 20244 75694
rect 20188 75590 20244 75628
rect 20412 75460 20468 75470
rect 19964 74722 20020 74732
rect 20300 74786 20356 74798
rect 20300 74734 20302 74786
rect 20354 74734 20356 74786
rect 19852 74508 20020 74564
rect 19852 74116 19908 74126
rect 19852 74022 19908 74060
rect 19852 73218 19908 73230
rect 19852 73166 19854 73218
rect 19906 73166 19908 73218
rect 19852 73108 19908 73166
rect 19964 73108 20020 74508
rect 20300 74338 20356 74734
rect 20300 74286 20302 74338
rect 20354 74286 20356 74338
rect 20300 74274 20356 74286
rect 20300 74116 20356 74126
rect 20300 74022 20356 74060
rect 20300 73556 20356 73566
rect 20300 73462 20356 73500
rect 19852 73052 20356 73108
rect 20188 72322 20244 72334
rect 20188 72270 20190 72322
rect 20242 72270 20244 72322
rect 19628 70702 19630 70754
rect 19682 70702 19684 70754
rect 19628 70690 19684 70702
rect 19740 70980 19796 70990
rect 19180 70476 19684 70532
rect 19516 70308 19572 70318
rect 19404 69524 19460 69534
rect 19404 69430 19460 69468
rect 19516 69410 19572 70252
rect 19516 69358 19518 69410
rect 19570 69358 19572 69410
rect 19516 69346 19572 69358
rect 19068 68786 19124 68796
rect 19292 69186 19348 69198
rect 19292 69134 19294 69186
rect 19346 69134 19348 69186
rect 18956 68516 19012 68526
rect 19292 68516 19348 69134
rect 19516 69188 19572 69198
rect 19404 68852 19460 68862
rect 19404 68758 19460 68796
rect 18956 68514 19124 68516
rect 18956 68462 18958 68514
rect 19010 68462 19124 68514
rect 18956 68460 19124 68462
rect 18956 68450 19012 68460
rect 18956 67844 19012 67854
rect 18956 67750 19012 67788
rect 19068 67732 19124 68460
rect 19292 68402 19348 68460
rect 19292 68350 19294 68402
rect 19346 68350 19348 68402
rect 19292 68338 19348 68350
rect 19292 67956 19348 67966
rect 19292 67842 19348 67900
rect 19292 67790 19294 67842
rect 19346 67790 19348 67842
rect 19292 67778 19348 67790
rect 19068 67620 19124 67676
rect 18396 66966 18452 67004
rect 18732 67004 18900 67060
rect 18956 67564 19124 67620
rect 19404 67620 19460 67630
rect 17836 66386 17892 66892
rect 17836 66334 17838 66386
rect 17890 66334 17892 66386
rect 17836 66322 17892 66334
rect 17948 66892 18116 66948
rect 17948 65602 18004 66892
rect 18222 66668 18486 66678
rect 18278 66612 18326 66668
rect 18382 66612 18430 66668
rect 18222 66602 18486 66612
rect 18508 66274 18564 66286
rect 18508 66222 18510 66274
rect 18562 66222 18564 66274
rect 17948 65550 17950 65602
rect 18002 65550 18004 65602
rect 17948 65538 18004 65550
rect 18060 65604 18116 65614
rect 18060 65510 18116 65548
rect 18508 65492 18564 66222
rect 18732 65828 18788 67004
rect 18956 66164 19012 67564
rect 19404 67526 19460 67564
rect 19516 67396 19572 69132
rect 19628 67618 19684 70476
rect 19740 68292 19796 70924
rect 20188 70980 20244 72270
rect 20300 71764 20356 73052
rect 20412 71988 20468 75404
rect 20748 75122 20804 75740
rect 21420 75794 21476 76300
rect 21756 76356 21812 76366
rect 21756 76262 21812 76300
rect 21420 75742 21422 75794
rect 21474 75742 21476 75794
rect 21420 75730 21476 75742
rect 21532 76132 21588 76142
rect 21308 75460 21364 75470
rect 21532 75460 21588 76076
rect 21868 75906 21924 76524
rect 21868 75854 21870 75906
rect 21922 75854 21924 75906
rect 21868 75794 21924 75854
rect 21868 75742 21870 75794
rect 21922 75742 21924 75794
rect 21868 75730 21924 75742
rect 21980 76242 22036 76972
rect 22092 76692 22148 77756
rect 22204 77140 22260 77150
rect 22204 77046 22260 77084
rect 22204 76692 22260 76702
rect 22092 76690 22260 76692
rect 22092 76638 22206 76690
rect 22258 76638 22260 76690
rect 22092 76636 22260 76638
rect 22204 76626 22260 76636
rect 21980 76190 21982 76242
rect 22034 76190 22036 76242
rect 20748 75070 20750 75122
rect 20802 75070 20804 75122
rect 20748 75058 20804 75070
rect 20860 75458 21364 75460
rect 20860 75406 21310 75458
rect 21362 75406 21364 75458
rect 20860 75404 21364 75406
rect 20748 74002 20804 74014
rect 20748 73950 20750 74002
rect 20802 73950 20804 74002
rect 20748 73948 20804 73950
rect 20636 73892 20804 73948
rect 20636 72548 20692 73892
rect 20748 73444 20804 73454
rect 20748 73350 20804 73388
rect 20524 72492 20692 72548
rect 20524 72324 20580 72492
rect 20524 72258 20580 72268
rect 20636 72324 20692 72334
rect 20636 72322 20804 72324
rect 20636 72270 20638 72322
rect 20690 72270 20804 72322
rect 20636 72268 20804 72270
rect 20636 72258 20692 72268
rect 20412 71932 20692 71988
rect 20412 71764 20468 71774
rect 20300 71762 20468 71764
rect 20300 71710 20414 71762
rect 20466 71710 20468 71762
rect 20300 71708 20468 71710
rect 20412 71698 20468 71708
rect 20188 70886 20244 70924
rect 20524 70980 20580 70990
rect 20188 70756 20244 70766
rect 19852 69410 19908 69422
rect 19852 69358 19854 69410
rect 19906 69358 19908 69410
rect 19852 68852 19908 69358
rect 19852 68786 19908 68796
rect 20076 69188 20132 69198
rect 19852 68514 19908 68526
rect 19852 68462 19854 68514
rect 19906 68462 19908 68514
rect 19852 68404 19908 68462
rect 19964 68404 20020 68414
rect 19852 68402 20020 68404
rect 19852 68350 19966 68402
rect 20018 68350 20020 68402
rect 19852 68348 20020 68350
rect 19964 68338 20020 68348
rect 19740 68236 19908 68292
rect 19852 67732 19908 68236
rect 19852 67666 19908 67676
rect 19628 67566 19630 67618
rect 19682 67566 19684 67618
rect 19628 67554 19684 67566
rect 19740 67620 19796 67630
rect 19404 67340 19572 67396
rect 19404 67170 19460 67340
rect 19404 67118 19406 67170
rect 19458 67118 19460 67170
rect 19404 67106 19460 67118
rect 18956 66098 19012 66108
rect 19068 67058 19124 67070
rect 19068 67006 19070 67058
rect 19122 67006 19124 67058
rect 18508 65426 18564 65436
rect 18620 65772 18788 65828
rect 18844 66050 18900 66062
rect 18844 65998 18846 66050
rect 18898 65998 18900 66050
rect 18284 65380 18340 65390
rect 18284 65286 18340 65324
rect 17724 65212 18116 65268
rect 17500 64878 17502 64930
rect 17554 64878 17556 64930
rect 17500 64866 17556 64878
rect 17276 64642 17332 64652
rect 16940 61058 16996 61068
rect 17052 64092 17220 64148
rect 17388 64484 17444 64494
rect 17052 60564 17108 64092
rect 17388 63924 17444 64428
rect 17388 63858 17444 63868
rect 17724 64036 17780 64046
rect 17612 63810 17668 63822
rect 17612 63758 17614 63810
rect 17666 63758 17668 63810
rect 17612 63362 17668 63758
rect 17612 63310 17614 63362
rect 17666 63310 17668 63362
rect 17612 63298 17668 63310
rect 17724 63250 17780 63980
rect 17724 63198 17726 63250
rect 17778 63198 17780 63250
rect 17164 63140 17220 63150
rect 17164 63046 17220 63084
rect 17500 62804 17556 62814
rect 17164 62692 17220 62702
rect 17164 61572 17220 62636
rect 17500 62466 17556 62748
rect 17724 62692 17780 63198
rect 17724 62626 17780 62636
rect 17500 62414 17502 62466
rect 17554 62414 17556 62466
rect 17500 62402 17556 62414
rect 17612 62354 17668 62366
rect 17612 62302 17614 62354
rect 17666 62302 17668 62354
rect 17500 62244 17556 62254
rect 17500 62150 17556 62188
rect 17612 62132 17668 62302
rect 17612 62066 17668 62076
rect 17724 61796 17780 61806
rect 17276 61572 17332 61582
rect 17164 61570 17332 61572
rect 17164 61518 17278 61570
rect 17330 61518 17332 61570
rect 17164 61516 17332 61518
rect 17164 61012 17220 61516
rect 17276 61506 17332 61516
rect 17388 61348 17444 61358
rect 17164 60946 17220 60956
rect 17276 61346 17444 61348
rect 17276 61294 17390 61346
rect 17442 61294 17444 61346
rect 17276 61292 17444 61294
rect 17276 60788 17332 61292
rect 17388 61282 17444 61292
rect 17612 60900 17668 60910
rect 17500 60898 17668 60900
rect 17500 60846 17614 60898
rect 17666 60846 17668 60898
rect 17500 60844 17668 60846
rect 17388 60788 17444 60798
rect 17276 60786 17444 60788
rect 17276 60734 17390 60786
rect 17442 60734 17444 60786
rect 17276 60732 17444 60734
rect 17388 60722 17444 60732
rect 16828 60508 17108 60564
rect 17276 60562 17332 60574
rect 17276 60510 17278 60562
rect 17330 60510 17332 60562
rect 16828 59444 16884 60508
rect 17276 60452 17332 60510
rect 16940 60396 17332 60452
rect 17388 60452 17444 60462
rect 16940 60002 16996 60396
rect 16940 59950 16942 60002
rect 16994 59950 16996 60002
rect 16940 59938 16996 59950
rect 17276 60228 17332 60238
rect 16828 59388 16996 59444
rect 16604 59218 16772 59220
rect 16604 59166 16606 59218
rect 16658 59166 16772 59218
rect 16604 59164 16772 59166
rect 16828 59220 16884 59230
rect 16156 56082 16212 56094
rect 16156 56030 16158 56082
rect 16210 56030 16212 56082
rect 16156 53508 16212 56030
rect 16268 54068 16324 58604
rect 16380 58436 16436 58446
rect 16380 58342 16436 58380
rect 16492 58322 16548 58334
rect 16492 58270 16494 58322
rect 16546 58270 16548 58322
rect 16492 57652 16548 58270
rect 16492 57586 16548 57596
rect 16492 57092 16548 57102
rect 16268 54012 16436 54068
rect 16268 53732 16324 53770
rect 16268 53666 16324 53676
rect 16268 53508 16324 53518
rect 16156 53452 16268 53508
rect 16268 53442 16324 53452
rect 16268 52948 16324 52958
rect 16268 51716 16324 52892
rect 16156 51380 16212 51390
rect 16156 51286 16212 51324
rect 16268 51378 16324 51660
rect 16268 51326 16270 51378
rect 16322 51326 16324 51378
rect 16268 51314 16324 51326
rect 15932 47628 16100 47684
rect 16156 50820 16212 50830
rect 15932 46676 15988 47628
rect 16156 47068 16212 50764
rect 16380 50428 16436 54012
rect 16492 53842 16548 57036
rect 16604 56980 16660 59164
rect 16828 59126 16884 59164
rect 16604 56866 16660 56924
rect 16604 56814 16606 56866
rect 16658 56814 16660 56866
rect 16604 56802 16660 56814
rect 16828 57652 16884 57662
rect 16828 57538 16884 57596
rect 16828 57486 16830 57538
rect 16882 57486 16884 57538
rect 16604 56308 16660 56318
rect 16604 56082 16660 56252
rect 16604 56030 16606 56082
rect 16658 56030 16660 56082
rect 16604 55524 16660 56030
rect 16604 55458 16660 55468
rect 16492 53790 16494 53842
rect 16546 53790 16548 53842
rect 16492 53778 16548 53790
rect 16716 53732 16772 53742
rect 16268 50372 16436 50428
rect 16492 53060 16548 53070
rect 16492 50484 16548 53004
rect 16716 52724 16772 53676
rect 16828 52948 16884 57486
rect 16940 56420 16996 59388
rect 17052 58324 17108 58334
rect 17052 56868 17108 58268
rect 17052 56774 17108 56812
rect 16940 56354 16996 56364
rect 16940 55972 16996 55982
rect 16940 55878 16996 55916
rect 17164 55188 17220 55198
rect 17164 55094 17220 55132
rect 17276 53508 17332 60172
rect 17388 59890 17444 60396
rect 17388 59838 17390 59890
rect 17442 59838 17444 59890
rect 17388 59826 17444 59838
rect 17500 59892 17556 60844
rect 17612 60834 17668 60844
rect 17500 59826 17556 59836
rect 17612 60452 17668 60462
rect 17500 59108 17556 59118
rect 17388 59106 17556 59108
rect 17388 59054 17502 59106
rect 17554 59054 17556 59106
rect 17388 59052 17556 59054
rect 17388 57650 17444 59052
rect 17500 58994 17556 59052
rect 17500 58942 17502 58994
rect 17554 58942 17556 58994
rect 17500 58930 17556 58942
rect 17500 57874 17556 57886
rect 17500 57822 17502 57874
rect 17554 57822 17556 57874
rect 17500 57764 17556 57822
rect 17500 57698 17556 57708
rect 17388 57598 17390 57650
rect 17442 57598 17444 57650
rect 17388 56420 17444 57598
rect 17388 56354 17444 56364
rect 17612 56196 17668 60396
rect 17724 56308 17780 61740
rect 17836 61682 17892 61694
rect 17836 61630 17838 61682
rect 17890 61630 17892 61682
rect 17836 61236 17892 61630
rect 17836 61170 17892 61180
rect 17948 60788 18004 60798
rect 17948 60694 18004 60732
rect 17836 60564 17892 60574
rect 17836 58994 17892 60508
rect 17836 58942 17838 58994
rect 17890 58942 17892 58994
rect 17836 58930 17892 58942
rect 17948 57764 18004 57774
rect 17836 57762 18004 57764
rect 17836 57710 17950 57762
rect 18002 57710 18004 57762
rect 17836 57708 18004 57710
rect 17836 57652 17892 57708
rect 17948 57698 18004 57708
rect 17836 57586 17892 57596
rect 18060 56868 18116 65212
rect 18222 65100 18486 65110
rect 18278 65044 18326 65100
rect 18382 65044 18430 65100
rect 18222 65034 18486 65044
rect 18222 63532 18486 63542
rect 18278 63476 18326 63532
rect 18382 63476 18430 63532
rect 18222 63466 18486 63476
rect 18172 63364 18228 63374
rect 18620 63364 18676 65772
rect 18732 65604 18788 65614
rect 18732 65510 18788 65548
rect 18844 65044 18900 65998
rect 19068 66052 19124 67006
rect 19516 67058 19572 67070
rect 19516 67006 19518 67058
rect 19570 67006 19572 67058
rect 19068 65986 19124 65996
rect 19404 66052 19460 66062
rect 19404 65958 19460 65996
rect 19516 65604 19572 67006
rect 19628 67060 19684 67070
rect 19740 67060 19796 67564
rect 19628 67058 19796 67060
rect 19628 67006 19630 67058
rect 19682 67006 19796 67058
rect 19628 67004 19796 67006
rect 19628 66994 19684 67004
rect 20076 66836 20132 69132
rect 20188 68180 20244 70700
rect 20300 70308 20356 70318
rect 20300 70082 20356 70252
rect 20300 70030 20302 70082
rect 20354 70030 20356 70082
rect 20300 70018 20356 70030
rect 20412 69188 20468 69198
rect 20412 69094 20468 69132
rect 20524 68964 20580 70924
rect 20188 68114 20244 68124
rect 20300 68908 20580 68964
rect 20300 68850 20356 68908
rect 20300 68798 20302 68850
rect 20354 68798 20356 68850
rect 20188 67842 20244 67854
rect 20188 67790 20190 67842
rect 20242 67790 20244 67842
rect 20188 67732 20244 67790
rect 20188 67666 20244 67676
rect 20300 67844 20356 68798
rect 20188 67060 20244 67070
rect 20300 67060 20356 67788
rect 20524 67732 20580 67742
rect 20636 67732 20692 71932
rect 20748 71876 20804 72268
rect 20748 71810 20804 71820
rect 20860 71652 20916 75404
rect 21308 75394 21364 75404
rect 21420 75404 21588 75460
rect 21420 75236 21476 75404
rect 21196 75180 21476 75236
rect 21624 75292 21888 75302
rect 21680 75236 21728 75292
rect 21784 75236 21832 75292
rect 21624 75226 21888 75236
rect 21084 73330 21140 73342
rect 21084 73278 21086 73330
rect 21138 73278 21140 73330
rect 21084 72996 21140 73278
rect 21084 72930 21140 72940
rect 21196 72772 21252 75180
rect 21980 75124 22036 76190
rect 22316 76020 22372 80220
rect 22428 80210 22484 80220
rect 22540 80164 22596 80556
rect 23100 80500 23156 85652
rect 23324 85314 23380 85326
rect 23324 85262 23326 85314
rect 23378 85262 23380 85314
rect 23324 85202 23380 85262
rect 23324 85150 23326 85202
rect 23378 85150 23380 85202
rect 23324 85138 23380 85150
rect 23548 84194 23604 86604
rect 23884 86436 23940 86446
rect 23884 86100 23940 86380
rect 24444 86100 24500 87276
rect 25564 87332 25620 87342
rect 25564 87238 25620 87276
rect 23884 86098 24500 86100
rect 23884 86046 24446 86098
rect 24498 86046 24500 86098
rect 23884 86044 24500 86046
rect 23884 85986 23940 86044
rect 24444 86034 24500 86044
rect 24892 87220 24948 87230
rect 23884 85934 23886 85986
rect 23938 85934 23940 85986
rect 23884 85922 23940 85934
rect 24668 85876 24724 85886
rect 24556 85764 24612 85802
rect 24556 85698 24612 85708
rect 24668 85762 24724 85820
rect 24668 85710 24670 85762
rect 24722 85710 24724 85762
rect 23996 85652 24052 85662
rect 23996 85558 24052 85596
rect 24668 85314 24724 85710
rect 24668 85262 24670 85314
rect 24722 85262 24724 85314
rect 24668 85250 24724 85262
rect 24892 85316 24948 87164
rect 25026 87052 25290 87062
rect 25082 86996 25130 87052
rect 25186 86996 25234 87052
rect 25026 86986 25290 86996
rect 25004 86658 25060 86670
rect 25004 86606 25006 86658
rect 25058 86606 25060 86658
rect 25004 86100 25060 86606
rect 25004 86034 25060 86044
rect 25676 86098 25732 87612
rect 26124 87602 26180 87612
rect 25788 87444 25844 87454
rect 25788 87350 25844 87388
rect 26348 87332 26404 88284
rect 26348 87266 26404 87276
rect 26460 88226 26516 88238
rect 26460 88174 26462 88226
rect 26514 88174 26516 88226
rect 26460 87444 26516 88174
rect 26012 87108 26068 87118
rect 26012 86658 26068 87052
rect 26012 86606 26014 86658
rect 26066 86606 26068 86658
rect 26012 86594 26068 86606
rect 26460 86324 26516 87388
rect 26796 88228 26852 89068
rect 27132 89058 27188 89068
rect 27244 89682 27300 89694
rect 27244 89630 27246 89682
rect 27298 89630 27300 89682
rect 26684 87218 26740 87230
rect 26684 87166 26686 87218
rect 26738 87166 26740 87218
rect 26460 86268 26628 86324
rect 25676 86046 25678 86098
rect 25730 86046 25732 86098
rect 25676 86034 25732 86046
rect 25788 86100 25844 86110
rect 25788 86006 25844 86044
rect 26460 85986 26516 85998
rect 26460 85934 26462 85986
rect 26514 85934 26516 85986
rect 25452 85876 25508 85886
rect 25452 85782 25508 85820
rect 26348 85874 26404 85886
rect 26348 85822 26350 85874
rect 26402 85822 26404 85874
rect 26348 85764 26404 85822
rect 26348 85698 26404 85708
rect 26460 85652 26516 85934
rect 25026 85484 25290 85494
rect 25082 85428 25130 85484
rect 25186 85428 25234 85484
rect 25026 85418 25290 85428
rect 25116 85316 25172 85326
rect 24892 85314 25172 85316
rect 24892 85262 25118 85314
rect 25170 85262 25172 85314
rect 24892 85260 25172 85262
rect 25116 85250 25172 85260
rect 25452 85316 25508 85326
rect 25452 85222 25508 85260
rect 24220 85204 24276 85214
rect 24220 85110 24276 85148
rect 25564 85204 25620 85214
rect 24780 84978 24836 84990
rect 24780 84926 24782 84978
rect 24834 84926 24836 84978
rect 23548 84142 23550 84194
rect 23602 84142 23604 84194
rect 23212 83748 23268 83758
rect 23268 83692 23380 83748
rect 23212 83682 23268 83692
rect 23324 82292 23380 83692
rect 23548 83636 23604 84142
rect 23660 84866 23716 84878
rect 23660 84814 23662 84866
rect 23714 84814 23716 84866
rect 23660 84196 23716 84814
rect 24668 84868 24724 84878
rect 24668 84774 24724 84812
rect 23660 84130 23716 84140
rect 23772 84306 23828 84318
rect 23772 84254 23774 84306
rect 23826 84254 23828 84306
rect 23436 83410 23492 83422
rect 23436 83358 23438 83410
rect 23490 83358 23492 83410
rect 23436 82740 23492 83358
rect 23548 82962 23604 83580
rect 23660 83972 23716 83982
rect 23660 83522 23716 83916
rect 23660 83470 23662 83522
rect 23714 83470 23716 83522
rect 23660 83458 23716 83470
rect 23772 83524 23828 84254
rect 24444 84308 24500 84318
rect 24444 84214 24500 84252
rect 24780 84084 24836 84926
rect 25564 84532 25620 85148
rect 25676 85092 25732 85102
rect 25676 84998 25732 85036
rect 26124 85092 26180 85102
rect 26124 84532 26180 85036
rect 26236 85092 26292 85102
rect 26460 85092 26516 85596
rect 26572 85316 26628 86268
rect 26572 85202 26628 85260
rect 26572 85150 26574 85202
rect 26626 85150 26628 85202
rect 26572 85138 26628 85150
rect 26236 85090 26516 85092
rect 26236 85038 26238 85090
rect 26290 85038 26516 85090
rect 26236 85036 26516 85038
rect 26236 85026 26292 85036
rect 25564 84476 25732 84532
rect 26124 84476 26292 84532
rect 25564 84308 25620 84318
rect 24780 84018 24836 84028
rect 25452 84252 25564 84308
rect 25026 83916 25290 83926
rect 23772 83458 23828 83468
rect 24220 83860 24276 83870
rect 25082 83860 25130 83916
rect 25186 83860 25234 83916
rect 25026 83850 25290 83860
rect 23548 82910 23550 82962
rect 23602 82910 23604 82962
rect 23548 82898 23604 82910
rect 24220 82850 24276 83804
rect 24332 83636 24388 83646
rect 24332 83542 24388 83580
rect 24444 83524 24500 83534
rect 24444 83430 24500 83468
rect 24220 82798 24222 82850
rect 24274 82798 24276 82850
rect 24220 82786 24276 82798
rect 24556 83410 24612 83422
rect 24556 83358 24558 83410
rect 24610 83358 24612 83410
rect 24556 82852 24612 83358
rect 25452 82962 25508 84252
rect 25564 84214 25620 84252
rect 25452 82910 25454 82962
rect 25506 82910 25508 82962
rect 25452 82898 25508 82910
rect 23436 82738 23716 82740
rect 23436 82686 23438 82738
rect 23490 82686 23716 82738
rect 23436 82684 23716 82686
rect 23436 82674 23492 82684
rect 23324 82236 23492 82292
rect 23212 81956 23268 81966
rect 23212 81862 23268 81900
rect 23436 81396 23492 82236
rect 22876 80444 23156 80500
rect 23212 81394 23492 81396
rect 23212 81342 23438 81394
rect 23490 81342 23492 81394
rect 23212 81340 23492 81342
rect 22652 80164 22708 80174
rect 22540 80108 22652 80164
rect 22652 79490 22708 80108
rect 22652 79438 22654 79490
rect 22706 79438 22708 79490
rect 22652 79426 22708 79438
rect 22540 78706 22596 78718
rect 22540 78654 22542 78706
rect 22594 78654 22596 78706
rect 22540 78596 22596 78654
rect 22540 78530 22596 78540
rect 22652 78594 22708 78606
rect 22652 78542 22654 78594
rect 22706 78542 22708 78594
rect 22540 77924 22596 77934
rect 22428 77922 22596 77924
rect 22428 77870 22542 77922
rect 22594 77870 22596 77922
rect 22428 77868 22596 77870
rect 22428 77026 22484 77868
rect 22540 77858 22596 77868
rect 22540 77476 22596 77486
rect 22652 77476 22708 78542
rect 22764 78596 22820 78606
rect 22764 78502 22820 78540
rect 22540 77474 22708 77476
rect 22540 77422 22542 77474
rect 22594 77422 22708 77474
rect 22540 77420 22708 77422
rect 22540 77410 22596 77420
rect 22428 76974 22430 77026
rect 22482 76974 22484 77026
rect 22428 76962 22484 76974
rect 22540 77250 22596 77262
rect 22540 77198 22542 77250
rect 22594 77198 22596 77250
rect 22540 76356 22596 77198
rect 22316 75964 22484 76020
rect 21420 75068 22036 75124
rect 22092 75906 22148 75918
rect 22092 75854 22094 75906
rect 22146 75854 22148 75906
rect 21308 74786 21364 74798
rect 21308 74734 21310 74786
rect 21362 74734 21364 74786
rect 21308 73330 21364 74734
rect 21308 73278 21310 73330
rect 21362 73278 21364 73330
rect 21308 73108 21364 73278
rect 21308 73042 21364 73052
rect 21420 74114 21476 75068
rect 21980 74900 22036 74910
rect 22092 74900 22148 75854
rect 22316 75796 22372 75806
rect 21980 74898 22260 74900
rect 21980 74846 21982 74898
rect 22034 74846 22260 74898
rect 21980 74844 22260 74846
rect 21980 74834 22036 74844
rect 21420 74062 21422 74114
rect 21474 74062 21476 74114
rect 21420 72884 21476 74062
rect 22204 74674 22260 74844
rect 22204 74622 22206 74674
rect 22258 74622 22260 74674
rect 22092 74002 22148 74014
rect 22092 73950 22094 74002
rect 22146 73950 22148 74002
rect 22092 73948 22148 73950
rect 21980 73892 22148 73948
rect 21624 73724 21888 73734
rect 21680 73668 21728 73724
rect 21784 73668 21832 73724
rect 21624 73658 21888 73668
rect 21868 73556 21924 73566
rect 21980 73556 22036 73892
rect 21868 73554 22036 73556
rect 21868 73502 21870 73554
rect 21922 73502 22036 73554
rect 21868 73500 22036 73502
rect 21868 73490 21924 73500
rect 21868 73330 21924 73342
rect 22204 73332 22260 74622
rect 22316 73444 22372 75740
rect 22428 74452 22484 75964
rect 22540 75796 22596 76300
rect 22652 76692 22708 76702
rect 22876 76692 22932 80444
rect 23100 80276 23156 80286
rect 23212 80276 23268 81340
rect 23436 81330 23492 81340
rect 23660 81394 23716 82684
rect 24556 82348 24612 82796
rect 24444 82292 24612 82348
rect 24668 82740 24724 82750
rect 23660 81342 23662 81394
rect 23714 81342 23716 81394
rect 23660 81330 23716 81342
rect 23772 82068 23828 82078
rect 23772 81394 23828 82012
rect 24444 81956 24500 82292
rect 24668 82068 24724 82684
rect 25452 82738 25508 82750
rect 25452 82686 25454 82738
rect 25506 82686 25508 82738
rect 25026 82348 25290 82358
rect 25082 82292 25130 82348
rect 25186 82292 25234 82348
rect 25026 82282 25290 82292
rect 25228 82180 25284 82190
rect 25228 82086 25284 82124
rect 24332 81954 24500 81956
rect 24332 81902 24446 81954
rect 24498 81902 24500 81954
rect 24332 81900 24500 81902
rect 23772 81342 23774 81394
rect 23826 81342 23828 81394
rect 23772 81330 23828 81342
rect 24220 81844 24276 81854
rect 23884 81284 23940 81294
rect 24220 81284 24276 81788
rect 24332 81620 24388 81900
rect 24444 81890 24500 81900
rect 24556 82012 24724 82068
rect 24780 82068 24836 82078
rect 24556 81844 24612 82012
rect 24780 82010 24836 82012
rect 24780 81958 24782 82010
rect 24834 81958 24836 82010
rect 24780 81946 24836 81958
rect 25452 81956 25508 82686
rect 25676 82348 25732 84476
rect 26236 84420 26292 84476
rect 26236 84326 26292 84364
rect 26124 84308 26180 84318
rect 26012 83524 26068 83534
rect 25900 83522 26068 83524
rect 25900 83470 26014 83522
rect 26066 83470 26068 83522
rect 25900 83468 26068 83470
rect 25340 81954 25508 81956
rect 25340 81902 25454 81954
rect 25506 81902 25508 81954
rect 25340 81900 25508 81902
rect 24668 81844 24724 81854
rect 24612 81842 24724 81844
rect 24612 81790 24670 81842
rect 24722 81790 24724 81842
rect 24612 81788 24724 81790
rect 24556 81778 24612 81788
rect 24668 81778 24724 81788
rect 24332 81564 24836 81620
rect 24556 81394 24612 81564
rect 24556 81342 24558 81394
rect 24610 81342 24612 81394
rect 24556 81330 24612 81342
rect 24668 81396 24724 81406
rect 24444 81284 24500 81294
rect 24220 81282 24500 81284
rect 24220 81230 24446 81282
rect 24498 81230 24500 81282
rect 24220 81228 24500 81230
rect 23884 81190 23940 81228
rect 24108 81060 24164 81070
rect 24108 80610 24164 81004
rect 24444 80724 24500 81228
rect 24556 80948 24612 80958
rect 24556 80854 24612 80892
rect 24444 80668 24612 80724
rect 24108 80558 24110 80610
rect 24162 80558 24164 80610
rect 24108 80546 24164 80558
rect 24556 80612 24612 80668
rect 24556 80518 24612 80556
rect 23436 80500 23492 80510
rect 23436 80406 23492 80444
rect 24444 80500 24500 80510
rect 24444 80386 24500 80444
rect 24444 80334 24446 80386
rect 24498 80334 24500 80386
rect 24444 80322 24500 80334
rect 23100 80274 23268 80276
rect 23100 80222 23102 80274
rect 23154 80222 23268 80274
rect 23100 80220 23268 80222
rect 23996 80274 24052 80286
rect 23996 80222 23998 80274
rect 24050 80222 24052 80274
rect 23100 80210 23156 80220
rect 23324 80164 23380 80174
rect 23324 80070 23380 80108
rect 23996 79828 24052 80222
rect 23996 79762 24052 79772
rect 24556 79828 24612 79838
rect 23772 79604 23828 79614
rect 23772 79510 23828 79548
rect 24220 79604 24276 79614
rect 23324 79490 23380 79502
rect 23324 79438 23326 79490
rect 23378 79438 23380 79490
rect 23324 78708 23380 79438
rect 24220 78930 24276 79548
rect 24220 78878 24222 78930
rect 24274 78878 24276 78930
rect 24220 78866 24276 78878
rect 23772 78820 23828 78830
rect 23772 78726 23828 78764
rect 23324 78614 23380 78652
rect 23212 78596 23268 78606
rect 23212 77812 23268 78540
rect 23212 77362 23268 77756
rect 23212 77310 23214 77362
rect 23266 77310 23268 77362
rect 23212 77298 23268 77310
rect 24220 78596 24276 78606
rect 23660 77140 23716 77150
rect 23660 77046 23716 77084
rect 22652 76690 22876 76692
rect 22652 76638 22654 76690
rect 22706 76638 22876 76690
rect 22652 76636 22876 76638
rect 22652 76132 22708 76636
rect 22876 76598 22932 76636
rect 23100 77026 23156 77038
rect 23100 76974 23102 77026
rect 23154 76974 23156 77026
rect 22652 76066 22708 76076
rect 22876 76242 22932 76254
rect 22876 76190 22878 76242
rect 22930 76190 22932 76242
rect 22540 75730 22596 75740
rect 22876 75682 22932 76190
rect 22876 75630 22878 75682
rect 22930 75630 22932 75682
rect 22876 75618 22932 75630
rect 23100 75684 23156 76974
rect 23772 76692 23828 76702
rect 23100 75618 23156 75628
rect 23212 76354 23268 76366
rect 23212 76302 23214 76354
rect 23266 76302 23268 76354
rect 22540 74788 22596 74798
rect 22540 74694 22596 74732
rect 22988 74786 23044 74798
rect 22988 74734 22990 74786
rect 23042 74734 23044 74786
rect 22428 74396 22708 74452
rect 22540 74228 22596 74238
rect 22316 73388 22484 73444
rect 21868 73278 21870 73330
rect 21922 73278 21924 73330
rect 21868 73220 21924 73278
rect 21868 73154 21924 73164
rect 22092 73276 22260 73332
rect 21644 73108 21700 73118
rect 21644 73014 21700 73052
rect 21868 72996 21924 73006
rect 22092 72996 22148 73276
rect 22316 73218 22372 73230
rect 22316 73166 22318 73218
rect 22370 73166 22372 73218
rect 21924 72940 22148 72996
rect 22204 73106 22260 73118
rect 22204 73054 22206 73106
rect 22258 73054 22260 73106
rect 22204 72996 22260 73054
rect 22316 73108 22372 73166
rect 22316 73042 22372 73052
rect 22428 73220 22484 73388
rect 21420 72828 21588 72884
rect 21196 72716 21476 72772
rect 21420 72658 21476 72716
rect 21420 72606 21422 72658
rect 21474 72606 21476 72658
rect 21420 72594 21476 72606
rect 21196 72548 21252 72558
rect 20748 71596 20916 71652
rect 21084 72324 21140 72334
rect 20748 70866 20804 71596
rect 21084 71204 21140 72268
rect 20748 70814 20750 70866
rect 20802 70814 20804 70866
rect 20748 70802 20804 70814
rect 20972 71148 21140 71204
rect 20860 70644 20916 70654
rect 20748 70084 20804 70094
rect 20748 69990 20804 70028
rect 20748 69186 20804 69198
rect 20748 69134 20750 69186
rect 20802 69134 20804 69186
rect 20748 69076 20804 69134
rect 20748 69010 20804 69020
rect 20748 68852 20804 68862
rect 20748 68758 20804 68796
rect 20524 67730 20692 67732
rect 20524 67678 20526 67730
rect 20578 67678 20692 67730
rect 20524 67676 20692 67678
rect 20524 67666 20580 67676
rect 20860 67172 20916 70588
rect 20188 67058 20356 67060
rect 20188 67006 20190 67058
rect 20242 67006 20356 67058
rect 20188 67004 20356 67006
rect 20188 66994 20244 67004
rect 19516 65538 19572 65548
rect 19852 66780 20132 66836
rect 18732 64988 18900 65044
rect 19404 65378 19460 65390
rect 19404 65326 19406 65378
rect 19458 65326 19460 65378
rect 18732 63588 18788 64988
rect 18732 63522 18788 63532
rect 18844 64818 18900 64830
rect 18844 64766 18846 64818
rect 18898 64766 18900 64818
rect 18620 63308 18788 63364
rect 18172 62356 18228 63308
rect 18732 63140 18788 63308
rect 18844 63362 18900 64766
rect 19180 64594 19236 64606
rect 19180 64542 19182 64594
rect 19234 64542 19236 64594
rect 18844 63310 18846 63362
rect 18898 63310 18900 63362
rect 18844 63298 18900 63310
rect 18956 64482 19012 64494
rect 18956 64430 18958 64482
rect 19010 64430 19012 64482
rect 18956 63364 19012 64430
rect 19180 64372 19236 64542
rect 19180 64306 19236 64316
rect 19404 64260 19460 65326
rect 19404 64194 19460 64204
rect 19628 64708 19684 64718
rect 19628 64482 19684 64652
rect 19628 64430 19630 64482
rect 19682 64430 19684 64482
rect 19292 63588 19348 63598
rect 19348 63532 19572 63588
rect 19292 63522 19348 63532
rect 18956 63298 19012 63308
rect 19292 63362 19348 63374
rect 19292 63310 19294 63362
rect 19346 63310 19348 63362
rect 19180 63140 19236 63178
rect 18732 63084 18900 63140
rect 18396 63026 18452 63038
rect 18396 62974 18398 63026
rect 18450 62974 18452 63026
rect 18396 62468 18452 62974
rect 18620 63028 18676 63038
rect 18620 62934 18676 62972
rect 18396 62402 18452 62412
rect 18620 62466 18676 62478
rect 18620 62414 18622 62466
rect 18674 62414 18676 62466
rect 18284 62356 18340 62366
rect 18172 62354 18340 62356
rect 18172 62302 18286 62354
rect 18338 62302 18340 62354
rect 18172 62300 18340 62302
rect 18284 62290 18340 62300
rect 18620 62356 18676 62414
rect 18620 62290 18676 62300
rect 18222 61964 18486 61974
rect 18278 61908 18326 61964
rect 18382 61908 18430 61964
rect 18222 61898 18486 61908
rect 18172 61124 18228 61134
rect 18228 61068 18340 61124
rect 18172 61058 18228 61068
rect 18284 60676 18340 61068
rect 18620 60788 18676 60798
rect 18508 60786 18676 60788
rect 18508 60734 18622 60786
rect 18674 60734 18676 60786
rect 18508 60732 18676 60734
rect 18508 60676 18564 60732
rect 18620 60722 18676 60732
rect 18732 60788 18788 60798
rect 18284 60620 18564 60676
rect 18620 60564 18676 60574
rect 18222 60396 18486 60406
rect 18278 60340 18326 60396
rect 18382 60340 18430 60396
rect 18222 60330 18486 60340
rect 18172 60004 18228 60014
rect 18172 59220 18228 59948
rect 18508 59780 18564 59790
rect 18508 59686 18564 59724
rect 18172 59106 18228 59164
rect 18172 59054 18174 59106
rect 18226 59054 18228 59106
rect 18172 59042 18228 59054
rect 18222 58828 18486 58838
rect 18278 58772 18326 58828
rect 18382 58772 18430 58828
rect 18222 58762 18486 58772
rect 18396 58434 18452 58446
rect 18396 58382 18398 58434
rect 18450 58382 18452 58434
rect 18396 58324 18452 58382
rect 18396 58258 18452 58268
rect 18222 57260 18486 57270
rect 18278 57204 18326 57260
rect 18382 57204 18430 57260
rect 18222 57194 18486 57204
rect 17948 56812 18116 56868
rect 17836 56308 17892 56318
rect 17724 56306 17892 56308
rect 17724 56254 17838 56306
rect 17890 56254 17892 56306
rect 17724 56252 17892 56254
rect 17948 56308 18004 56812
rect 18172 56754 18228 56766
rect 18172 56702 18174 56754
rect 18226 56702 18228 56754
rect 17948 56252 18116 56308
rect 17836 56242 17892 56252
rect 17612 56140 17780 56196
rect 17724 56084 17780 56140
rect 17948 56084 18004 56094
rect 17724 56028 17892 56084
rect 17612 55972 17668 55982
rect 17612 55878 17668 55916
rect 16828 52882 16884 52892
rect 17164 53452 17332 53508
rect 17388 55524 17444 55534
rect 17388 54402 17444 55468
rect 17388 54350 17390 54402
rect 17442 54350 17444 54402
rect 16716 52050 16772 52668
rect 16716 51998 16718 52050
rect 16770 51998 16772 52050
rect 16716 51604 16772 51998
rect 17052 52724 17108 52734
rect 16716 51538 16772 51548
rect 16828 51716 16884 51726
rect 16828 51602 16884 51660
rect 16828 51550 16830 51602
rect 16882 51550 16884 51602
rect 16828 51538 16884 51550
rect 16492 50390 16548 50428
rect 16268 49140 16324 50372
rect 16716 50034 16772 50046
rect 16716 49982 16718 50034
rect 16770 49982 16772 50034
rect 16268 49074 16324 49084
rect 16380 49588 16436 49598
rect 15932 46610 15988 46620
rect 16044 47012 16212 47068
rect 16268 48356 16324 48366
rect 16268 47348 16324 48300
rect 16380 48244 16436 49532
rect 16716 48692 16772 49982
rect 16828 49924 16884 49934
rect 16828 49830 16884 49868
rect 17052 49252 17108 52668
rect 16828 49196 17108 49252
rect 16828 48804 16884 49196
rect 17052 48916 17108 48926
rect 16828 48748 16996 48804
rect 16716 48626 16772 48636
rect 16604 48468 16660 48478
rect 16604 48466 16772 48468
rect 16604 48414 16606 48466
rect 16658 48414 16772 48466
rect 16604 48412 16772 48414
rect 16604 48402 16660 48412
rect 16380 48188 16660 48244
rect 16380 47348 16436 47358
rect 16268 47346 16436 47348
rect 16268 47294 16382 47346
rect 16434 47294 16436 47346
rect 16268 47292 16436 47294
rect 15708 45266 15764 45276
rect 15820 45892 15876 45902
rect 15372 44818 15428 44828
rect 15484 44940 15652 44996
rect 15260 44382 15262 44434
rect 15314 44382 15316 44434
rect 15260 44370 15316 44382
rect 14924 44270 14926 44322
rect 14978 44270 14980 44322
rect 14924 44258 14980 44270
rect 15372 44322 15428 44334
rect 15372 44270 15374 44322
rect 15426 44270 15428 44322
rect 15148 44100 15204 44110
rect 15148 44098 15316 44100
rect 15148 44046 15150 44098
rect 15202 44046 15316 44098
rect 15148 44044 15316 44046
rect 15148 44034 15204 44044
rect 14252 43426 14308 43932
rect 14820 43932 15084 43942
rect 14252 43374 14254 43426
rect 14306 43374 14308 43426
rect 14252 43362 14308 43374
rect 14364 43876 14420 43886
rect 14364 43316 14420 43820
rect 14364 43250 14420 43260
rect 14588 43876 14644 43886
rect 14876 43876 14924 43932
rect 14980 43876 15028 43932
rect 14820 43866 15084 43876
rect 15260 43876 15316 44044
rect 14588 42642 14644 43820
rect 15260 43810 15316 43820
rect 14588 42590 14590 42642
rect 14642 42590 14644 42642
rect 14140 42532 14196 42542
rect 14140 42438 14196 42476
rect 14252 42530 14308 42542
rect 14252 42478 14254 42530
rect 14306 42478 14308 42530
rect 13916 41356 14084 41412
rect 13804 41076 13860 41086
rect 13804 40982 13860 41020
rect 13916 40964 13972 41356
rect 14028 41188 14084 41198
rect 14252 41188 14308 42478
rect 14364 42532 14420 42542
rect 14364 42438 14420 42476
rect 14588 41636 14644 42590
rect 14588 41570 14644 41580
rect 14700 43540 14756 43550
rect 14588 41300 14644 41310
rect 14700 41300 14756 43484
rect 15036 43540 15092 43550
rect 15036 43446 15092 43484
rect 15148 42754 15204 42766
rect 15148 42702 15150 42754
rect 15202 42702 15204 42754
rect 14820 42364 15084 42374
rect 14876 42308 14924 42364
rect 14980 42308 15028 42364
rect 14820 42298 15084 42308
rect 15148 42084 15204 42702
rect 15036 42028 15204 42084
rect 15260 42532 15316 42542
rect 14588 41298 14756 41300
rect 14588 41246 14590 41298
rect 14642 41246 14756 41298
rect 14588 41244 14756 41246
rect 14812 41972 14868 41982
rect 15036 41972 15092 42028
rect 14868 41916 15092 41972
rect 14588 41234 14644 41244
rect 14812 41188 14868 41916
rect 15148 41860 15204 41870
rect 15260 41860 15316 42476
rect 15148 41858 15316 41860
rect 15148 41806 15150 41858
rect 15202 41806 15316 41858
rect 15148 41804 15316 41806
rect 15372 41860 15428 44270
rect 15148 41794 15204 41804
rect 14924 41636 14980 41646
rect 14980 41580 15204 41636
rect 14924 41570 14980 41580
rect 14028 41186 14308 41188
rect 14028 41134 14030 41186
rect 14082 41134 14308 41186
rect 14028 41132 14308 41134
rect 14700 41186 14868 41188
rect 14700 41134 14814 41186
rect 14866 41134 14868 41186
rect 14700 41132 14868 41134
rect 14028 41122 14084 41132
rect 13916 40908 14308 40964
rect 14028 40628 14084 40638
rect 13580 40626 13972 40628
rect 13580 40574 13582 40626
rect 13634 40574 13972 40626
rect 13580 40572 13972 40574
rect 13580 40292 13636 40572
rect 13580 40226 13636 40236
rect 13580 39842 13636 39854
rect 13580 39790 13582 39842
rect 13634 39790 13636 39842
rect 13580 39394 13636 39790
rect 13580 39342 13582 39394
rect 13634 39342 13636 39394
rect 13580 39172 13636 39342
rect 13580 39106 13636 39116
rect 13244 38612 13412 38668
rect 13244 34020 13300 38612
rect 13580 38276 13636 38286
rect 13580 38162 13636 38220
rect 13580 38110 13582 38162
rect 13634 38110 13636 38162
rect 13580 38098 13636 38110
rect 13692 38274 13748 38286
rect 13692 38222 13694 38274
rect 13746 38222 13748 38274
rect 13580 37492 13636 37502
rect 13580 37044 13636 37436
rect 13580 36978 13636 36988
rect 13692 36932 13748 38222
rect 13916 37492 13972 40572
rect 14028 40534 14084 40572
rect 14028 39844 14084 39854
rect 14028 38834 14084 39788
rect 14140 39620 14196 39630
rect 14140 39526 14196 39564
rect 14028 38782 14030 38834
rect 14082 38782 14084 38834
rect 14028 38274 14084 38782
rect 14028 38222 14030 38274
rect 14082 38222 14084 38274
rect 14028 38210 14084 38222
rect 13916 37398 13972 37436
rect 14140 37826 14196 37838
rect 14140 37774 14142 37826
rect 14194 37774 14196 37826
rect 14140 37268 14196 37774
rect 13692 36866 13748 36876
rect 13804 37212 14196 37268
rect 14252 37266 14308 40908
rect 14476 40290 14532 40302
rect 14476 40238 14478 40290
rect 14530 40238 14532 40290
rect 14476 39842 14532 40238
rect 14476 39790 14478 39842
rect 14530 39790 14532 39842
rect 14476 39778 14532 39790
rect 14700 39844 14756 41132
rect 14812 41122 14868 41132
rect 15148 40964 15204 41580
rect 15372 41524 15428 41804
rect 15260 41468 15428 41524
rect 15260 41076 15316 41468
rect 15372 41300 15428 41310
rect 15484 41300 15540 44940
rect 15820 44210 15876 45836
rect 15932 45332 15988 45342
rect 16044 45332 16100 47012
rect 16268 46786 16324 47292
rect 16380 47282 16436 47292
rect 16268 46734 16270 46786
rect 16322 46734 16324 46786
rect 16268 45778 16324 46734
rect 16268 45726 16270 45778
rect 16322 45726 16324 45778
rect 16268 45714 16324 45726
rect 15932 45330 16100 45332
rect 15932 45278 15934 45330
rect 15986 45278 16100 45330
rect 15932 45276 16100 45278
rect 16156 45332 16212 45342
rect 15932 45266 15988 45276
rect 15820 44158 15822 44210
rect 15874 44158 15876 44210
rect 15820 44146 15876 44158
rect 16156 45106 16212 45276
rect 16156 45054 16158 45106
rect 16210 45054 16212 45106
rect 16044 44098 16100 44110
rect 16044 44046 16046 44098
rect 16098 44046 16100 44098
rect 15596 43538 15652 43550
rect 15596 43486 15598 43538
rect 15650 43486 15652 43538
rect 15596 41524 15652 43486
rect 15932 43538 15988 43550
rect 15932 43486 15934 43538
rect 15986 43486 15988 43538
rect 15708 43428 15764 43438
rect 15708 43426 15876 43428
rect 15708 43374 15710 43426
rect 15762 43374 15876 43426
rect 15708 43372 15876 43374
rect 15708 43362 15764 43372
rect 15820 42866 15876 43372
rect 15820 42814 15822 42866
rect 15874 42814 15876 42866
rect 15820 42802 15876 42814
rect 15932 42196 15988 43486
rect 16044 43316 16100 44046
rect 16156 44100 16212 45054
rect 16380 45106 16436 45118
rect 16380 45054 16382 45106
rect 16434 45054 16436 45106
rect 16156 44034 16212 44044
rect 16268 44994 16324 45006
rect 16268 44942 16270 44994
rect 16322 44942 16324 44994
rect 16156 43540 16212 43550
rect 16156 43446 16212 43484
rect 16044 43250 16100 43260
rect 15932 42140 16100 42196
rect 15708 42084 15764 42094
rect 15708 41990 15764 42028
rect 15932 41970 15988 41982
rect 15932 41918 15934 41970
rect 15986 41918 15988 41970
rect 15820 41860 15876 41870
rect 15596 41458 15652 41468
rect 15708 41858 15876 41860
rect 15708 41806 15822 41858
rect 15874 41806 15876 41858
rect 15708 41804 15876 41806
rect 15428 41244 15540 41300
rect 15596 41300 15652 41310
rect 15708 41300 15764 41804
rect 15820 41794 15876 41804
rect 15596 41298 15764 41300
rect 15596 41246 15598 41298
rect 15650 41246 15764 41298
rect 15596 41244 15764 41246
rect 15932 41748 15988 41918
rect 15372 41234 15428 41244
rect 15596 41234 15652 41244
rect 15260 41020 15652 41076
rect 14820 40796 15084 40806
rect 14876 40740 14924 40796
rect 14980 40740 15028 40796
rect 14820 40730 15084 40740
rect 15148 40626 15204 40908
rect 15148 40574 15150 40626
rect 15202 40574 15204 40626
rect 15148 40562 15204 40574
rect 15596 40626 15652 41020
rect 15596 40574 15598 40626
rect 15650 40574 15652 40626
rect 15596 40562 15652 40574
rect 14700 39778 14756 39788
rect 15932 39732 15988 41692
rect 16044 41188 16100 42140
rect 16268 41972 16324 44942
rect 16380 43652 16436 45054
rect 16604 45106 16660 48188
rect 16604 45054 16606 45106
rect 16658 45054 16660 45106
rect 16604 43764 16660 45054
rect 16604 43698 16660 43708
rect 16380 43586 16436 43596
rect 16604 43426 16660 43438
rect 16604 43374 16606 43426
rect 16658 43374 16660 43426
rect 16492 43314 16548 43326
rect 16492 43262 16494 43314
rect 16546 43262 16548 43314
rect 16492 42868 16548 43262
rect 16492 42802 16548 42812
rect 16604 42196 16660 43374
rect 16044 40626 16100 41132
rect 16044 40574 16046 40626
rect 16098 40574 16100 40626
rect 16044 40562 16100 40574
rect 16156 41916 16324 41972
rect 16380 42140 16660 42196
rect 16156 40292 16212 41916
rect 16268 41748 16324 41758
rect 16380 41748 16436 42140
rect 16268 41746 16436 41748
rect 16268 41694 16270 41746
rect 16322 41694 16436 41746
rect 16268 41692 16436 41694
rect 16492 41970 16548 41982
rect 16492 41918 16494 41970
rect 16546 41918 16548 41970
rect 16268 41682 16324 41692
rect 16492 41636 16548 41918
rect 16156 40226 16212 40236
rect 16380 41580 16548 41636
rect 16380 40180 16436 41580
rect 16716 41076 16772 48412
rect 16828 48354 16884 48366
rect 16828 48302 16830 48354
rect 16882 48302 16884 48354
rect 16828 48020 16884 48302
rect 16828 47954 16884 47964
rect 16828 47796 16884 47806
rect 16828 45218 16884 47740
rect 16828 45166 16830 45218
rect 16882 45166 16884 45218
rect 16828 45154 16884 45166
rect 16940 44436 16996 48748
rect 17052 47572 17108 48860
rect 17164 48020 17220 53452
rect 17388 53396 17444 54350
rect 17164 47954 17220 47964
rect 17276 53340 17444 53396
rect 17612 55300 17668 55310
rect 17276 47796 17332 53340
rect 17388 52948 17444 52958
rect 17388 51380 17444 52892
rect 17612 52724 17668 55244
rect 17612 52658 17668 52668
rect 17724 54516 17780 54526
rect 17724 52500 17780 54460
rect 17612 52276 17668 52286
rect 17612 52162 17668 52220
rect 17612 52110 17614 52162
rect 17666 52110 17668 52162
rect 17612 52098 17668 52110
rect 17724 51938 17780 52444
rect 17724 51886 17726 51938
rect 17778 51886 17780 51938
rect 17500 51716 17556 51726
rect 17500 51602 17556 51660
rect 17500 51550 17502 51602
rect 17554 51550 17556 51602
rect 17500 51538 17556 51550
rect 17388 51324 17556 51380
rect 17388 50594 17444 50606
rect 17388 50542 17390 50594
rect 17442 50542 17444 50594
rect 17388 49924 17444 50542
rect 17388 49858 17444 49868
rect 17388 48916 17444 48926
rect 17500 48916 17556 51324
rect 17724 50484 17780 51886
rect 17724 50418 17780 50428
rect 17444 48860 17556 48916
rect 17612 50372 17668 50382
rect 17388 48850 17444 48860
rect 17500 48580 17556 48590
rect 17388 48524 17500 48580
rect 17388 48242 17444 48524
rect 17500 48514 17556 48524
rect 17500 48356 17556 48366
rect 17612 48356 17668 50316
rect 17724 49924 17780 49934
rect 17724 48804 17780 49868
rect 17724 48738 17780 48748
rect 17556 48300 17668 48356
rect 17500 48262 17556 48300
rect 17388 48190 17390 48242
rect 17442 48190 17444 48242
rect 17388 48178 17444 48190
rect 17276 47730 17332 47740
rect 17612 48020 17668 48030
rect 17052 47516 17332 47572
rect 17052 47346 17108 47358
rect 17052 47294 17054 47346
rect 17106 47294 17108 47346
rect 17052 46004 17108 47294
rect 17276 47236 17332 47516
rect 17276 47180 17444 47236
rect 17052 45938 17108 45948
rect 17276 47068 17332 47078
rect 17164 45668 17220 45678
rect 16940 44370 16996 44380
rect 17052 45666 17220 45668
rect 17052 45614 17166 45666
rect 17218 45614 17220 45666
rect 17052 45612 17220 45614
rect 16828 43538 16884 43550
rect 16828 43486 16830 43538
rect 16882 43486 16884 43538
rect 16828 42308 16884 43486
rect 16828 42242 16884 42252
rect 16716 41010 16772 41020
rect 16828 42084 16884 42094
rect 16716 40740 16772 40750
rect 16828 40740 16884 42028
rect 16772 40684 16884 40740
rect 16716 40626 16772 40684
rect 16716 40574 16718 40626
rect 16770 40574 16772 40626
rect 16716 40562 16772 40574
rect 16380 40114 16436 40124
rect 16380 39844 16436 39854
rect 16044 39732 16100 39742
rect 15932 39730 16100 39732
rect 15932 39678 16046 39730
rect 16098 39678 16100 39730
rect 15932 39676 16100 39678
rect 16044 39666 16100 39676
rect 16380 39730 16436 39788
rect 16380 39678 16382 39730
rect 16434 39678 16436 39730
rect 15148 39620 15204 39630
rect 15148 39526 15204 39564
rect 14588 39508 14644 39518
rect 14924 39508 14980 39518
rect 14588 39506 14924 39508
rect 14588 39454 14590 39506
rect 14642 39454 14924 39506
rect 14588 39452 14924 39454
rect 14588 39442 14644 39452
rect 14924 39414 14980 39452
rect 15484 39508 15540 39518
rect 15484 39414 15540 39452
rect 15148 39394 15204 39406
rect 15148 39342 15150 39394
rect 15202 39342 15204 39394
rect 14820 39228 15084 39238
rect 14876 39172 14924 39228
rect 14980 39172 15028 39228
rect 14820 39162 15084 39172
rect 15148 39060 15204 39342
rect 16044 39284 16100 39294
rect 14700 39004 15204 39060
rect 15372 39060 15428 39070
rect 14700 38946 14756 39004
rect 14700 38894 14702 38946
rect 14754 38894 14756 38946
rect 14700 38882 14756 38894
rect 14820 37660 15084 37670
rect 14876 37604 14924 37660
rect 14980 37604 15028 37660
rect 14820 37594 15084 37604
rect 14252 37214 14254 37266
rect 14306 37214 14308 37266
rect 13804 36708 13860 37212
rect 14252 37202 14308 37214
rect 14364 37492 14420 37502
rect 14028 36708 14084 36718
rect 13804 36652 14028 36708
rect 13692 36484 13748 36494
rect 13468 36372 13524 36382
rect 13468 36278 13524 36316
rect 13356 35812 13412 35822
rect 13356 35698 13412 35756
rect 13356 35646 13358 35698
rect 13410 35646 13412 35698
rect 13356 35634 13412 35646
rect 13692 35308 13748 36428
rect 13916 36484 13972 36494
rect 13916 36390 13972 36428
rect 14028 36482 14084 36652
rect 14364 36708 14420 37436
rect 15260 37492 15316 37502
rect 15260 37398 15316 37436
rect 14364 36614 14420 36652
rect 14476 37266 14532 37278
rect 14476 37214 14478 37266
rect 14530 37214 14532 37266
rect 14028 36430 14030 36482
rect 14082 36430 14084 36482
rect 14028 36418 14084 36430
rect 13580 35252 13748 35308
rect 13804 36372 13860 36382
rect 14476 36372 14532 37214
rect 14588 37268 14644 37278
rect 14588 37174 14644 37212
rect 15036 37268 15092 37278
rect 15036 37174 15092 37212
rect 15148 36820 15204 36830
rect 13580 35138 13636 35252
rect 13580 35086 13582 35138
rect 13634 35086 13636 35138
rect 13580 35026 13636 35086
rect 13580 34974 13582 35026
rect 13634 34974 13636 35026
rect 13580 34962 13636 34974
rect 13244 33964 13412 34020
rect 13132 27346 13188 27356
rect 13244 33572 13300 33582
rect 12684 26684 13076 26740
rect 12572 26514 12628 26526
rect 12572 26462 12574 26514
rect 12626 26462 12628 26514
rect 12460 26404 12516 26414
rect 12572 26404 12628 26462
rect 12516 26348 12628 26404
rect 12460 26338 12516 26348
rect 12348 24770 12404 24780
rect 12460 25284 12516 25294
rect 12460 24610 12516 25228
rect 12460 24558 12462 24610
rect 12514 24558 12516 24610
rect 12460 24546 12516 24558
rect 12684 24052 12740 26684
rect 12796 26290 12852 26302
rect 12796 26238 12798 26290
rect 12850 26238 12852 26290
rect 12796 25620 12852 26238
rect 13132 26290 13188 26302
rect 13132 26238 13134 26290
rect 13186 26238 13188 26290
rect 13132 26180 13188 26238
rect 13132 26114 13188 26124
rect 12796 25554 12852 25564
rect 12908 26068 12964 26078
rect 12908 25618 12964 26012
rect 13244 25956 13300 33516
rect 13356 29092 13412 33964
rect 13580 33124 13636 33134
rect 13468 33122 13636 33124
rect 13468 33070 13582 33122
rect 13634 33070 13636 33122
rect 13468 33068 13636 33070
rect 13468 33012 13524 33068
rect 13580 33058 13636 33068
rect 13468 32004 13524 32956
rect 13804 32788 13860 36316
rect 14140 36316 14532 36372
rect 14588 36594 14644 36606
rect 14588 36542 14590 36594
rect 14642 36542 14644 36594
rect 14140 35924 14196 36316
rect 14140 35868 14308 35924
rect 14140 35588 14196 35598
rect 14140 35494 14196 35532
rect 13916 35138 13972 35150
rect 13916 35086 13918 35138
rect 13970 35086 13972 35138
rect 13916 34916 13972 35086
rect 13916 34354 13972 34860
rect 13916 34302 13918 34354
rect 13970 34302 13972 34354
rect 13916 34290 13972 34302
rect 14140 34914 14196 34926
rect 14140 34862 14142 34914
rect 14194 34862 14196 34914
rect 14140 34020 14196 34862
rect 14140 33954 14196 33964
rect 13468 31938 13524 31948
rect 13580 32732 13860 32788
rect 13468 31668 13524 31678
rect 13468 30882 13524 31612
rect 13468 30830 13470 30882
rect 13522 30830 13524 30882
rect 13468 30818 13524 30830
rect 13580 30660 13636 32732
rect 13692 32450 13748 32462
rect 13692 32398 13694 32450
rect 13746 32398 13748 32450
rect 13692 31220 13748 32398
rect 14140 31220 14196 31230
rect 13692 31218 14196 31220
rect 13692 31166 14142 31218
rect 14194 31166 14196 31218
rect 13692 31164 14196 31166
rect 14252 31220 14308 35868
rect 14588 35812 14644 36542
rect 14700 36484 14756 36494
rect 14700 36390 14756 36428
rect 15148 36482 15204 36764
rect 15148 36430 15150 36482
rect 15202 36430 15204 36482
rect 15148 36418 15204 36430
rect 15260 36484 15316 36494
rect 15372 36484 15428 39004
rect 15932 38052 15988 38062
rect 15932 37604 15988 37996
rect 15932 37538 15988 37548
rect 16044 37940 16100 39228
rect 16380 38164 16436 39678
rect 17052 39620 17108 45612
rect 17164 45602 17220 45612
rect 16716 39564 17108 39620
rect 17164 45332 17220 45342
rect 16492 38164 16548 38174
rect 16380 38108 16492 38164
rect 16492 38070 16548 38108
rect 16044 37490 16100 37884
rect 16044 37438 16046 37490
rect 16098 37438 16100 37490
rect 15596 37156 15652 37166
rect 15260 36482 15428 36484
rect 15260 36430 15262 36482
rect 15314 36430 15428 36482
rect 15260 36428 15428 36430
rect 15484 37044 15540 37054
rect 15484 36482 15540 36988
rect 15484 36430 15486 36482
rect 15538 36430 15540 36482
rect 15260 36418 15316 36428
rect 15372 36260 15428 36270
rect 15372 36166 15428 36204
rect 14820 36092 15084 36102
rect 14876 36036 14924 36092
rect 14980 36036 15028 36092
rect 14820 36026 15084 36036
rect 15260 35924 15316 35934
rect 14476 35756 14644 35812
rect 15148 35868 15260 35924
rect 14364 35364 14420 35374
rect 14364 33236 14420 35308
rect 14476 35138 14532 35756
rect 14812 35588 14868 35598
rect 14476 35086 14478 35138
rect 14530 35086 14532 35138
rect 14476 35074 14532 35086
rect 14588 35308 14644 35318
rect 14588 34916 14644 35252
rect 14812 35026 14868 35532
rect 14812 34974 14814 35026
rect 14866 34974 14868 35026
rect 14812 34962 14868 34974
rect 14924 35028 14980 35038
rect 14364 33170 14420 33180
rect 14476 34860 14644 34916
rect 14700 34916 14756 34926
rect 14252 31164 14420 31220
rect 14140 31154 14196 31164
rect 13356 28756 13412 29036
rect 13356 28690 13412 28700
rect 13468 30604 13636 30660
rect 14028 30994 14084 31006
rect 14028 30942 14030 30994
rect 14082 30942 14084 30994
rect 13356 28420 13412 28430
rect 13356 27524 13412 28364
rect 13468 28308 13524 30604
rect 13804 29988 13860 29998
rect 14028 29988 14084 30942
rect 13804 29986 14084 29988
rect 13804 29934 13806 29986
rect 13858 29934 14084 29986
rect 13804 29932 14084 29934
rect 14140 30996 14196 31006
rect 14140 29986 14196 30940
rect 14252 30994 14308 31006
rect 14252 30942 14254 30994
rect 14306 30942 14308 30994
rect 14252 30884 14308 30942
rect 14252 30324 14308 30828
rect 14252 30258 14308 30268
rect 14140 29934 14142 29986
rect 14194 29934 14196 29986
rect 13804 29922 13860 29932
rect 13580 29314 13636 29326
rect 13580 29262 13582 29314
rect 13634 29262 13636 29314
rect 13580 28756 13636 29262
rect 13804 28756 13860 28766
rect 13580 28754 13860 28756
rect 13580 28702 13806 28754
rect 13858 28702 13860 28754
rect 13580 28700 13860 28702
rect 13804 28690 13860 28700
rect 13916 28756 13972 29932
rect 13916 28690 13972 28700
rect 14028 29092 14084 29102
rect 14028 28642 14084 29036
rect 14140 28868 14196 29934
rect 14140 28802 14196 28812
rect 14252 28980 14308 28990
rect 14028 28590 14030 28642
rect 14082 28590 14084 28642
rect 14028 28578 14084 28590
rect 14140 28644 14196 28654
rect 14140 28550 14196 28588
rect 14252 28642 14308 28924
rect 14252 28590 14254 28642
rect 14306 28590 14308 28642
rect 13692 28532 13748 28542
rect 13692 28438 13748 28476
rect 14252 28420 14308 28590
rect 14140 28364 14308 28420
rect 13468 28252 13860 28308
rect 13692 27524 13748 27534
rect 13356 27458 13412 27468
rect 13468 27468 13692 27524
rect 13468 26514 13524 27468
rect 13692 27458 13748 27468
rect 13580 27076 13636 27086
rect 13580 26982 13636 27020
rect 13692 26852 13748 26862
rect 13468 26462 13470 26514
rect 13522 26462 13524 26514
rect 13468 26450 13524 26462
rect 13580 26796 13692 26852
rect 13356 26402 13412 26414
rect 13356 26350 13358 26402
rect 13410 26350 13412 26402
rect 13356 26068 13412 26350
rect 13356 26002 13412 26012
rect 12908 25566 12910 25618
rect 12962 25566 12964 25618
rect 12908 25554 12964 25566
rect 13132 25900 13300 25956
rect 12908 24610 12964 24622
rect 12908 24558 12910 24610
rect 12962 24558 12964 24610
rect 12460 23996 12740 24052
rect 12796 24276 12852 24286
rect 12796 24050 12852 24220
rect 12796 23998 12798 24050
rect 12850 23998 12852 24050
rect 12348 23938 12404 23950
rect 12348 23886 12350 23938
rect 12402 23886 12404 23938
rect 12348 23548 12404 23886
rect 12236 23492 12404 23548
rect 12236 23154 12292 23492
rect 12460 23380 12516 23996
rect 12796 23986 12852 23998
rect 12908 23940 12964 24558
rect 12908 23884 13076 23940
rect 12684 23828 12740 23838
rect 12236 23102 12238 23154
rect 12290 23102 12292 23154
rect 12236 23044 12292 23102
rect 12236 22978 12292 22988
rect 12348 23324 12516 23380
rect 12572 23826 12740 23828
rect 12572 23774 12686 23826
rect 12738 23774 12740 23826
rect 12572 23772 12740 23774
rect 12348 22036 12404 23324
rect 12460 23154 12516 23166
rect 12460 23102 12462 23154
rect 12514 23102 12516 23154
rect 12460 22932 12516 23102
rect 12460 22866 12516 22876
rect 12236 21980 12404 22036
rect 12236 21026 12292 21980
rect 12236 20974 12238 21026
rect 12290 20974 12292 21026
rect 12236 20962 12292 20974
rect 12348 21812 12404 21822
rect 11900 19068 12180 19124
rect 12348 20018 12404 21756
rect 12460 21476 12516 21486
rect 12460 21382 12516 21420
rect 12348 19966 12350 20018
rect 12402 19966 12404 20018
rect 11900 17220 11956 19068
rect 12348 18452 12404 19966
rect 12460 21026 12516 21038
rect 12460 20974 12462 21026
rect 12514 20974 12516 21026
rect 12460 20914 12516 20974
rect 12460 20862 12462 20914
rect 12514 20862 12516 20914
rect 12460 20692 12516 20862
rect 12460 20020 12516 20636
rect 12460 19954 12516 19964
rect 12460 19796 12516 19806
rect 12460 19346 12516 19740
rect 12460 19294 12462 19346
rect 12514 19294 12516 19346
rect 12460 19236 12516 19294
rect 12460 19170 12516 19180
rect 12124 18396 12348 18452
rect 12012 17666 12068 17678
rect 12012 17614 12014 17666
rect 12066 17614 12068 17666
rect 12012 17444 12068 17614
rect 12012 17378 12068 17388
rect 11900 17164 12068 17220
rect 12012 15148 12068 17164
rect 12124 16882 12180 18396
rect 12348 18386 12404 18396
rect 12572 17668 12628 23772
rect 12684 23762 12740 23772
rect 12796 23828 12852 23838
rect 12684 23604 12740 23614
rect 12684 23378 12740 23548
rect 12684 23326 12686 23378
rect 12738 23326 12740 23378
rect 12684 23156 12740 23326
rect 12796 23378 12852 23772
rect 12908 23714 12964 23726
rect 12908 23662 12910 23714
rect 12962 23662 12964 23714
rect 12908 23604 12964 23662
rect 12908 23538 12964 23548
rect 13020 23716 13076 23884
rect 12796 23326 12798 23378
rect 12850 23326 12852 23378
rect 12796 23314 12852 23326
rect 13020 23380 13076 23660
rect 13020 23314 13076 23324
rect 12684 23100 13076 23156
rect 13020 22482 13076 23100
rect 13020 22430 13022 22482
rect 13074 22430 13076 22482
rect 13020 22418 13076 22430
rect 12684 22372 12740 22382
rect 12684 17890 12740 22316
rect 12908 21812 12964 21822
rect 12908 21718 12964 21756
rect 13132 21812 13188 25900
rect 13356 25620 13412 25630
rect 13412 25564 13524 25620
rect 13356 25554 13412 25564
rect 13356 24724 13412 24734
rect 13468 24724 13524 25564
rect 13356 24722 13524 24724
rect 13356 24670 13358 24722
rect 13410 24670 13524 24722
rect 13356 24668 13524 24670
rect 13244 23716 13300 23726
rect 13244 23378 13300 23660
rect 13244 23326 13246 23378
rect 13298 23326 13300 23378
rect 13244 23314 13300 23326
rect 13356 23044 13412 24668
rect 13468 24276 13524 24286
rect 13468 24050 13524 24220
rect 13468 23998 13470 24050
rect 13522 23998 13524 24050
rect 13468 23986 13524 23998
rect 13356 22978 13412 22988
rect 13580 23154 13636 26796
rect 13692 26786 13748 26796
rect 13804 26068 13860 28252
rect 14028 27860 14084 27870
rect 14028 26402 14084 27804
rect 14140 26852 14196 28364
rect 14252 28196 14308 28206
rect 14252 28082 14308 28140
rect 14252 28030 14254 28082
rect 14306 28030 14308 28082
rect 14252 28018 14308 28030
rect 14364 27524 14420 31164
rect 14364 27458 14420 27468
rect 14140 26786 14196 26796
rect 14252 26962 14308 26974
rect 14252 26910 14254 26962
rect 14306 26910 14308 26962
rect 14252 26514 14308 26910
rect 14252 26462 14254 26514
rect 14306 26462 14308 26514
rect 14252 26450 14308 26462
rect 14364 26516 14420 26526
rect 14028 26350 14030 26402
rect 14082 26350 14084 26402
rect 14028 26338 14084 26350
rect 14364 26292 14420 26460
rect 14252 26290 14420 26292
rect 14252 26238 14366 26290
rect 14418 26238 14420 26290
rect 14252 26236 14420 26238
rect 13804 26012 14196 26068
rect 13804 25620 13860 25630
rect 13804 25526 13860 25564
rect 14140 25506 14196 26012
rect 14140 25454 14142 25506
rect 14194 25454 14196 25506
rect 14140 25442 14196 25454
rect 14252 24946 14308 26236
rect 14364 26226 14420 26236
rect 14476 25394 14532 34860
rect 14700 34822 14756 34860
rect 14924 34914 14980 34972
rect 14924 34862 14926 34914
rect 14978 34862 14980 34914
rect 14924 34850 14980 34862
rect 14820 34524 15084 34534
rect 14876 34468 14924 34524
rect 14980 34468 15028 34524
rect 14820 34458 15084 34468
rect 14924 33460 14980 33470
rect 14700 33458 14980 33460
rect 14700 33406 14926 33458
rect 14978 33406 14980 33458
rect 14700 33404 14980 33406
rect 14588 33348 14644 33358
rect 14588 31220 14644 33292
rect 14588 31154 14644 31164
rect 14588 30996 14644 31006
rect 14588 30902 14644 30940
rect 14588 30772 14644 30782
rect 14700 30772 14756 33404
rect 14924 33394 14980 33404
rect 15148 33346 15204 35868
rect 15260 35858 15316 35868
rect 15484 35812 15540 36430
rect 15484 35746 15540 35756
rect 15596 35140 15652 37100
rect 16044 36820 16100 37438
rect 16044 36754 16100 36764
rect 15708 36708 15764 36718
rect 15708 36482 15764 36652
rect 15708 36430 15710 36482
rect 15762 36430 15764 36482
rect 15708 36418 15764 36430
rect 16156 36484 16212 36494
rect 16044 36370 16100 36382
rect 16044 36318 16046 36370
rect 16098 36318 16100 36370
rect 15708 36260 15764 36270
rect 15764 36204 15876 36260
rect 15708 36194 15764 36204
rect 15148 33294 15150 33346
rect 15202 33294 15204 33346
rect 14812 33236 14868 33246
rect 14812 33142 14868 33180
rect 14820 32956 15084 32966
rect 14876 32900 14924 32956
rect 14980 32900 15028 32956
rect 14820 32890 15084 32900
rect 15148 32452 15204 33294
rect 15148 32386 15204 32396
rect 15260 35084 15652 35140
rect 15708 35476 15764 35486
rect 15820 35476 15876 36204
rect 16044 35924 16100 36318
rect 16044 35858 16100 35868
rect 16044 35700 16100 35710
rect 15820 35420 15988 35476
rect 14820 31388 15084 31398
rect 14876 31332 14924 31388
rect 14980 31332 15028 31388
rect 14820 31322 15084 31332
rect 14588 30770 14756 30772
rect 14588 30718 14590 30770
rect 14642 30718 14756 30770
rect 14588 30716 14756 30718
rect 14812 31220 14868 31230
rect 14588 30706 14644 30716
rect 14812 30322 14868 31164
rect 15260 30884 15316 35084
rect 15596 34916 15652 34926
rect 15596 34356 15652 34860
rect 15708 34802 15764 35420
rect 15932 34914 15988 35420
rect 15932 34862 15934 34914
rect 15986 34862 15988 34914
rect 15932 34850 15988 34862
rect 15708 34750 15710 34802
rect 15762 34750 15764 34802
rect 15708 34738 15764 34750
rect 15820 34802 15876 34814
rect 15820 34750 15822 34802
rect 15874 34750 15876 34802
rect 15820 34580 15876 34750
rect 15820 34524 15988 34580
rect 15820 34356 15876 34366
rect 15596 34354 15876 34356
rect 15596 34302 15822 34354
rect 15874 34302 15876 34354
rect 15596 34300 15876 34302
rect 15820 34290 15876 34300
rect 15372 34020 15428 34030
rect 15372 31108 15428 33964
rect 15932 33348 15988 34524
rect 15932 33282 15988 33292
rect 15596 33236 15652 33246
rect 15596 33142 15652 33180
rect 15820 32452 15876 32462
rect 15820 32358 15876 32396
rect 16044 32116 16100 35644
rect 16156 35588 16212 36428
rect 16492 36484 16548 36494
rect 16492 36390 16548 36428
rect 16604 36372 16660 36382
rect 16604 36278 16660 36316
rect 16268 36260 16324 36270
rect 16268 36166 16324 36204
rect 16380 36258 16436 36270
rect 16380 36206 16382 36258
rect 16434 36206 16436 36258
rect 16268 35588 16324 35598
rect 16156 35586 16324 35588
rect 16156 35534 16270 35586
rect 16322 35534 16324 35586
rect 16156 35532 16324 35534
rect 16268 35522 16324 35532
rect 16380 35476 16436 36206
rect 16716 36148 16772 39564
rect 16940 39394 16996 39406
rect 16940 39342 16942 39394
rect 16994 39342 16996 39394
rect 16940 39060 16996 39342
rect 16940 38994 16996 39004
rect 16828 38724 16884 38734
rect 16828 38630 16884 38668
rect 16380 35410 16436 35420
rect 16492 36092 16772 36148
rect 16828 38164 16884 38174
rect 16828 37490 16884 38108
rect 16828 37438 16830 37490
rect 16882 37438 16884 37490
rect 16380 35140 16436 35150
rect 16380 35046 16436 35084
rect 16492 32788 16548 36092
rect 16716 35924 16772 35934
rect 16828 35924 16884 37438
rect 17164 36484 17220 45276
rect 17276 36596 17332 47012
rect 17388 46674 17444 47180
rect 17388 46622 17390 46674
rect 17442 46622 17444 46674
rect 17388 45892 17444 46622
rect 17388 45826 17444 45836
rect 17500 45780 17556 45790
rect 17500 45330 17556 45724
rect 17500 45278 17502 45330
rect 17554 45278 17556 45330
rect 17500 45266 17556 45278
rect 17612 45332 17668 47964
rect 17836 47236 17892 56028
rect 17948 55990 18004 56028
rect 17948 53060 18004 53070
rect 17948 52966 18004 53004
rect 17948 52612 18004 52622
rect 17948 51266 18004 52556
rect 17948 51214 17950 51266
rect 18002 51214 18004 51266
rect 17948 49812 18004 51214
rect 17948 49746 18004 49756
rect 18060 47348 18116 56252
rect 18172 55972 18228 56702
rect 18284 56084 18340 56094
rect 18284 55990 18340 56028
rect 18172 55906 18228 55916
rect 18222 55692 18486 55702
rect 18278 55636 18326 55692
rect 18382 55636 18430 55692
rect 18222 55626 18486 55636
rect 18222 54124 18486 54134
rect 18278 54068 18326 54124
rect 18382 54068 18430 54124
rect 18222 54058 18486 54068
rect 18396 53732 18452 53742
rect 18396 53284 18452 53676
rect 18508 53620 18564 53630
rect 18508 53526 18564 53564
rect 18396 53218 18452 53228
rect 18620 52948 18676 60508
rect 18732 53954 18788 60732
rect 18732 53902 18734 53954
rect 18786 53902 18788 53954
rect 18732 53890 18788 53902
rect 18620 52882 18676 52892
rect 18620 52724 18676 52734
rect 18222 52556 18486 52566
rect 18278 52500 18326 52556
rect 18382 52500 18430 52556
rect 18222 52490 18486 52500
rect 18172 52052 18228 52062
rect 18172 51156 18228 51996
rect 18396 51940 18452 51950
rect 18396 51378 18452 51884
rect 18620 51490 18676 52668
rect 18620 51438 18622 51490
rect 18674 51438 18676 51490
rect 18620 51426 18676 51438
rect 18732 51940 18788 51950
rect 18732 51492 18788 51884
rect 18732 51398 18788 51436
rect 18396 51326 18398 51378
rect 18450 51326 18452 51378
rect 18396 51314 18452 51326
rect 18172 51090 18228 51100
rect 18222 50988 18486 50998
rect 18278 50932 18326 50988
rect 18382 50932 18430 50988
rect 18222 50922 18486 50932
rect 18508 50820 18564 50830
rect 18508 49924 18564 50764
rect 18844 50148 18900 63084
rect 19180 63074 19236 63084
rect 19180 62916 19236 62926
rect 19292 62916 19348 63310
rect 19180 62914 19348 62916
rect 19180 62862 19182 62914
rect 19234 62862 19348 62914
rect 19180 62860 19348 62862
rect 19180 62850 19236 62860
rect 19292 62580 19348 62590
rect 19292 62486 19348 62524
rect 19180 62468 19236 62478
rect 19180 60900 19236 62412
rect 19516 62188 19572 63532
rect 19628 63140 19684 64430
rect 19740 63810 19796 63822
rect 19740 63758 19742 63810
rect 19794 63758 19796 63810
rect 19740 63362 19796 63758
rect 19740 63310 19742 63362
rect 19794 63310 19796 63362
rect 19740 63298 19796 63310
rect 19628 63046 19684 63084
rect 19852 62916 19908 66780
rect 19964 66050 20020 66062
rect 19964 65998 19966 66050
rect 20018 65998 20020 66050
rect 19964 65604 20020 65998
rect 19964 65538 20020 65548
rect 19964 65380 20020 65390
rect 19964 65378 20132 65380
rect 19964 65326 19966 65378
rect 20018 65326 20132 65378
rect 19964 65324 20132 65326
rect 19964 65314 20020 65324
rect 19964 64596 20020 64606
rect 20076 64596 20132 65324
rect 20300 64932 20356 67004
rect 20636 67116 20916 67172
rect 20188 64596 20244 64606
rect 20076 64594 20244 64596
rect 20076 64542 20190 64594
rect 20242 64542 20244 64594
rect 20076 64540 20244 64542
rect 19964 64502 20020 64540
rect 20188 64036 20244 64540
rect 18956 60898 19236 60900
rect 18956 60846 19182 60898
rect 19234 60846 19236 60898
rect 18956 60844 19236 60846
rect 18956 60002 19012 60844
rect 19180 60834 19236 60844
rect 19292 62132 19572 62188
rect 19628 62860 19908 62916
rect 19964 63980 20244 64036
rect 18956 59950 18958 60002
rect 19010 59950 19012 60002
rect 18956 59938 19012 59950
rect 19180 59892 19236 59930
rect 19180 59826 19236 59836
rect 19068 59780 19124 59790
rect 18956 59778 19124 59780
rect 18956 59726 19070 59778
rect 19122 59726 19124 59778
rect 18956 59724 19124 59726
rect 18956 59332 19012 59724
rect 19068 59714 19124 59724
rect 18956 59266 19012 59276
rect 19180 59668 19236 59678
rect 19180 57204 19236 59612
rect 19180 57138 19236 57148
rect 19292 56868 19348 62132
rect 19516 62020 19572 62030
rect 19516 61460 19572 61964
rect 19404 60900 19460 60910
rect 19404 60806 19460 60844
rect 19516 60564 19572 61404
rect 19628 60788 19684 62860
rect 19628 60722 19684 60732
rect 19740 62692 19796 62702
rect 19740 62578 19796 62636
rect 19740 62526 19742 62578
rect 19794 62526 19796 62578
rect 19740 60786 19796 62526
rect 19964 62188 20020 63980
rect 20300 63924 20356 64876
rect 20524 66052 20580 66062
rect 20412 64706 20468 64718
rect 20412 64654 20414 64706
rect 20466 64654 20468 64706
rect 20412 64148 20468 64654
rect 20524 64708 20580 65996
rect 20524 64614 20580 64652
rect 20412 64092 20580 64148
rect 20412 63924 20468 63934
rect 20300 63922 20468 63924
rect 20300 63870 20414 63922
rect 20466 63870 20468 63922
rect 20300 63868 20468 63870
rect 20412 63858 20468 63868
rect 20524 63812 20580 64092
rect 20524 63746 20580 63756
rect 20636 63588 20692 67116
rect 20860 66948 20916 66958
rect 20748 66946 20916 66948
rect 20748 66894 20862 66946
rect 20914 66894 20916 66946
rect 20748 66892 20916 66894
rect 20748 66612 20804 66892
rect 20860 66882 20916 66892
rect 20748 66546 20804 66556
rect 20748 66052 20804 66062
rect 20748 65958 20804 65996
rect 20972 65604 21028 71148
rect 21196 68740 21252 72492
rect 21532 72436 21588 72828
rect 21420 72380 21588 72436
rect 21868 72436 21924 72940
rect 22204 72930 22260 72940
rect 22316 72546 22372 72558
rect 22316 72494 22318 72546
rect 22370 72494 22372 72546
rect 21420 71988 21476 72380
rect 21868 72342 21924 72380
rect 22092 72434 22148 72446
rect 22092 72382 22094 72434
rect 22146 72382 22148 72434
rect 22092 72324 22148 72382
rect 21980 72212 22036 72222
rect 21624 72156 21888 72166
rect 21680 72100 21728 72156
rect 21784 72100 21832 72156
rect 21624 72090 21888 72100
rect 21532 71988 21588 71998
rect 21420 71932 21532 71988
rect 21420 71540 21476 71550
rect 21308 70420 21364 70430
rect 21308 70326 21364 70364
rect 21084 68684 21252 68740
rect 21084 66948 21140 68684
rect 21084 66882 21140 66892
rect 21196 68514 21252 68526
rect 21196 68462 21198 68514
rect 21250 68462 21252 68514
rect 21196 68402 21252 68462
rect 21196 68350 21198 68402
rect 21250 68350 21252 68402
rect 21196 66836 21252 68350
rect 21420 68180 21476 71484
rect 21532 70980 21588 71932
rect 21532 70886 21588 70924
rect 21980 71874 22036 72156
rect 21980 71822 21982 71874
rect 22034 71822 22036 71874
rect 21980 70644 22036 71822
rect 22092 70868 22148 72268
rect 22204 72322 22260 72334
rect 22204 72270 22206 72322
rect 22258 72270 22260 72322
rect 22204 71090 22260 72270
rect 22316 72100 22372 72494
rect 22428 72546 22484 73164
rect 22428 72494 22430 72546
rect 22482 72494 22484 72546
rect 22428 72482 22484 72494
rect 22540 73330 22596 74172
rect 22540 73278 22542 73330
rect 22594 73278 22596 73330
rect 22540 72548 22596 73278
rect 22540 72482 22596 72492
rect 22316 72034 22372 72044
rect 22652 71988 22708 74396
rect 22764 73780 22820 73790
rect 22764 72996 22820 73724
rect 22988 73444 23044 74734
rect 23212 73892 23268 76302
rect 23548 76356 23604 76366
rect 23548 76262 23604 76300
rect 23548 75570 23604 75582
rect 23548 75518 23550 75570
rect 23602 75518 23604 75570
rect 23324 74786 23380 74798
rect 23324 74734 23326 74786
rect 23378 74734 23380 74786
rect 23324 74674 23380 74734
rect 23324 74622 23326 74674
rect 23378 74622 23380 74674
rect 23324 74610 23380 74622
rect 23548 74452 23604 75518
rect 23548 74386 23604 74396
rect 23660 75572 23716 75582
rect 23660 74116 23716 75516
rect 23772 75122 23828 76636
rect 24108 76354 24164 76366
rect 24108 76302 24110 76354
rect 24162 76302 24164 76354
rect 23884 75908 23940 75918
rect 23940 75852 24052 75908
rect 23884 75842 23940 75852
rect 23772 75070 23774 75122
rect 23826 75070 23828 75122
rect 23772 75058 23828 75070
rect 23548 74060 23716 74116
rect 23996 74116 24052 75852
rect 24108 75012 24164 76302
rect 24108 74946 24164 74956
rect 24220 75124 24276 78540
rect 24444 77924 24500 77934
rect 24444 77250 24500 77868
rect 24444 77198 24446 77250
rect 24498 77198 24500 77250
rect 24444 77186 24500 77198
rect 24332 77140 24388 77150
rect 24332 77046 24388 77084
rect 24444 76692 24500 76702
rect 24556 76692 24612 79772
rect 24668 79826 24724 81340
rect 24780 80388 24836 81564
rect 25228 81060 25284 81070
rect 25340 81060 25396 81900
rect 25452 81890 25508 81900
rect 25564 82292 25732 82348
rect 25788 83410 25844 83422
rect 25788 83358 25790 83410
rect 25842 83358 25844 83410
rect 25284 81004 25396 81060
rect 25228 80966 25284 81004
rect 25452 80948 25508 80958
rect 25452 80854 25508 80892
rect 25026 80780 25290 80790
rect 25082 80724 25130 80780
rect 25186 80724 25234 80780
rect 25026 80714 25290 80724
rect 24780 80322 24836 80332
rect 25228 80612 25284 80622
rect 25564 80612 25620 82292
rect 25788 82180 25844 83358
rect 25788 81060 25844 82124
rect 25676 80948 25732 80958
rect 25788 80948 25844 81004
rect 25676 80946 25844 80948
rect 25676 80894 25678 80946
rect 25730 80894 25844 80946
rect 25676 80892 25844 80894
rect 25676 80882 25732 80892
rect 25900 80724 25956 83468
rect 26012 83458 26068 83468
rect 26124 83300 26180 84252
rect 26348 84308 26404 85036
rect 26572 84980 26628 84990
rect 26348 83746 26404 84252
rect 26348 83694 26350 83746
rect 26402 83694 26404 83746
rect 26348 83682 26404 83694
rect 26460 84924 26572 84980
rect 26460 84084 26516 84924
rect 26572 84914 26628 84924
rect 26572 84420 26628 84430
rect 26684 84420 26740 87166
rect 26796 87108 26852 88172
rect 27132 88898 27188 88910
rect 27132 88846 27134 88898
rect 27186 88846 27188 88898
rect 27132 88116 27188 88846
rect 27132 87442 27188 88060
rect 27132 87390 27134 87442
rect 27186 87390 27188 87442
rect 27132 87378 27188 87390
rect 26908 87220 26964 87230
rect 26908 87126 26964 87164
rect 26796 87042 26852 87052
rect 27244 86884 27300 89630
rect 28140 89012 28196 89022
rect 28252 89012 28308 90692
rect 28428 89404 28692 89414
rect 28484 89348 28532 89404
rect 28588 89348 28636 89404
rect 28428 89338 28692 89348
rect 28140 89010 28308 89012
rect 28140 88958 28142 89010
rect 28194 88958 28308 89010
rect 28140 88956 28308 88958
rect 28140 88946 28196 88956
rect 27580 88228 27636 88238
rect 27580 87666 27636 88172
rect 28428 87836 28692 87846
rect 28484 87780 28532 87836
rect 28588 87780 28636 87836
rect 28428 87770 28692 87780
rect 27580 87614 27582 87666
rect 27634 87614 27636 87666
rect 27580 87602 27636 87614
rect 27132 86828 27300 86884
rect 27356 87442 27412 87454
rect 27356 87390 27358 87442
rect 27410 87390 27412 87442
rect 27132 85988 27188 86828
rect 27244 86660 27300 86670
rect 27244 86566 27300 86604
rect 26908 85932 27188 85988
rect 26572 84418 26740 84420
rect 26572 84366 26574 84418
rect 26626 84366 26740 84418
rect 26572 84364 26740 84366
rect 26796 85540 26852 85550
rect 26572 84354 26628 84364
rect 26684 84196 26740 84206
rect 26796 84196 26852 85484
rect 26908 84644 26964 85932
rect 27244 85876 27300 85886
rect 27020 85874 27300 85876
rect 27020 85822 27246 85874
rect 27298 85822 27300 85874
rect 27020 85820 27300 85822
rect 27356 85876 27412 87390
rect 27468 87332 27524 87342
rect 27468 87238 27524 87276
rect 28140 87330 28196 87342
rect 28140 87278 28142 87330
rect 28194 87278 28196 87330
rect 27692 86772 27748 86782
rect 27748 86716 27860 86772
rect 27692 86706 27748 86716
rect 27804 85986 27860 86716
rect 27804 85934 27806 85986
rect 27858 85934 27860 85986
rect 27804 85922 27860 85934
rect 27916 86658 27972 86670
rect 27916 86606 27918 86658
rect 27970 86606 27972 86658
rect 27356 85820 27636 85876
rect 27020 85090 27076 85820
rect 27244 85810 27300 85820
rect 27468 85652 27524 85662
rect 27468 85558 27524 85596
rect 27356 85540 27412 85550
rect 27356 85316 27412 85484
rect 27356 85260 27524 85316
rect 27020 85038 27022 85090
rect 27074 85038 27076 85090
rect 27020 84756 27076 85038
rect 27132 84980 27188 84990
rect 27356 84980 27412 84990
rect 27132 84978 27412 84980
rect 27132 84926 27134 84978
rect 27186 84926 27358 84978
rect 27410 84926 27412 84978
rect 27132 84924 27412 84926
rect 27132 84914 27188 84924
rect 27356 84914 27412 84924
rect 27468 84978 27524 85260
rect 27468 84926 27470 84978
rect 27522 84926 27524 84978
rect 27468 84914 27524 84926
rect 27020 84700 27188 84756
rect 26908 84578 26964 84588
rect 27132 84420 27188 84700
rect 27580 84532 27636 85820
rect 27916 85708 27972 86606
rect 27692 85650 27748 85662
rect 27692 85598 27694 85650
rect 27746 85598 27748 85650
rect 27692 85540 27748 85598
rect 27692 85474 27748 85484
rect 27804 85652 27972 85708
rect 27692 84868 27748 84878
rect 27692 84774 27748 84812
rect 27580 84476 27748 84532
rect 27132 84306 27188 84364
rect 27468 84308 27524 84318
rect 27132 84254 27134 84306
rect 27186 84254 27188 84306
rect 27132 84242 27188 84254
rect 27244 84306 27524 84308
rect 27244 84254 27470 84306
rect 27522 84254 27524 84306
rect 27244 84252 27524 84254
rect 26684 84194 26852 84196
rect 26684 84142 26686 84194
rect 26738 84142 26852 84194
rect 26684 84140 26852 84142
rect 26684 84130 26740 84140
rect 26012 83244 26180 83300
rect 26012 82178 26068 83244
rect 26236 82852 26292 82862
rect 26236 82758 26292 82796
rect 26124 82740 26180 82750
rect 26124 82646 26180 82684
rect 26348 82626 26404 82638
rect 26348 82574 26350 82626
rect 26402 82574 26404 82626
rect 26012 82126 26014 82178
rect 26066 82126 26068 82178
rect 26012 82114 26068 82126
rect 26236 82180 26292 82190
rect 26236 81954 26292 82124
rect 26236 81902 26238 81954
rect 26290 81902 26292 81954
rect 26236 81890 26292 81902
rect 26348 81956 26404 82574
rect 26348 81890 26404 81900
rect 26460 81620 26516 84028
rect 26908 84084 26964 84094
rect 27244 84084 27300 84252
rect 27468 84242 27524 84252
rect 27580 84308 27636 84318
rect 27580 84214 27636 84252
rect 27692 84084 27748 84476
rect 26908 84082 27300 84084
rect 26908 84030 26910 84082
rect 26962 84030 27300 84082
rect 26908 84028 27300 84030
rect 27468 84028 27748 84084
rect 26908 84018 26964 84028
rect 26684 83972 26740 83982
rect 26236 81564 26516 81620
rect 26572 82066 26628 82078
rect 26572 82014 26574 82066
rect 26626 82014 26628 82066
rect 26572 81956 26628 82014
rect 26124 81396 26180 81406
rect 26236 81396 26292 81564
rect 26124 81394 26292 81396
rect 26124 81342 26126 81394
rect 26178 81342 26292 81394
rect 26124 81340 26292 81342
rect 26124 81330 26180 81340
rect 26348 81284 26404 81294
rect 26348 81282 26516 81284
rect 26348 81230 26350 81282
rect 26402 81230 26516 81282
rect 26348 81228 26516 81230
rect 26348 81218 26404 81228
rect 26460 81172 26516 81228
rect 26460 81106 26516 81116
rect 26348 81060 26404 81070
rect 25228 80386 25284 80556
rect 25228 80334 25230 80386
rect 25282 80334 25284 80386
rect 25228 80322 25284 80334
rect 25452 80556 25620 80612
rect 25788 80668 25956 80724
rect 26236 80948 26292 80958
rect 24668 79774 24670 79826
rect 24722 79774 24724 79826
rect 24668 79762 24724 79774
rect 25004 80162 25060 80174
rect 25004 80110 25006 80162
rect 25058 80110 25060 80162
rect 25004 79604 25060 80110
rect 25452 79716 25508 80556
rect 25564 80388 25620 80426
rect 25564 80322 25620 80332
rect 25564 80164 25620 80174
rect 25788 80164 25844 80668
rect 26236 80612 26292 80892
rect 25900 80610 26292 80612
rect 25900 80558 26238 80610
rect 26290 80558 26292 80610
rect 25900 80556 26292 80558
rect 25900 80386 25956 80556
rect 26236 80546 26292 80556
rect 25900 80334 25902 80386
rect 25954 80334 25956 80386
rect 25900 80322 25956 80334
rect 26348 80276 26404 81004
rect 26460 80946 26516 80958
rect 26460 80894 26462 80946
rect 26514 80894 26516 80946
rect 26460 80612 26516 80894
rect 26572 80948 26628 81900
rect 26572 80882 26628 80892
rect 26460 80546 26516 80556
rect 26572 80724 26628 80734
rect 26572 80610 26628 80668
rect 26572 80558 26574 80610
rect 26626 80558 26628 80610
rect 26572 80546 26628 80558
rect 26460 80276 26516 80286
rect 26348 80274 26516 80276
rect 26348 80222 26462 80274
rect 26514 80222 26516 80274
rect 26348 80220 26516 80222
rect 26460 80210 26516 80220
rect 25564 80162 25844 80164
rect 25564 80110 25566 80162
rect 25618 80110 25844 80162
rect 25564 80108 25844 80110
rect 26684 80164 26740 83916
rect 27468 83746 27524 84028
rect 27468 83694 27470 83746
rect 27522 83694 27524 83746
rect 27468 83682 27524 83694
rect 27132 83410 27188 83422
rect 27132 83358 27134 83410
rect 27186 83358 27188 83410
rect 25564 80098 25620 80108
rect 26684 80098 26740 80108
rect 26796 83298 26852 83310
rect 26796 83246 26798 83298
rect 26850 83246 26852 83298
rect 26236 79828 26292 79838
rect 26684 79828 26740 79838
rect 26796 79828 26852 83246
rect 27020 82738 27076 82750
rect 27020 82686 27022 82738
rect 27074 82686 27076 82738
rect 26908 82292 26964 82302
rect 26908 81170 26964 82236
rect 27020 81284 27076 82686
rect 27132 82626 27188 83358
rect 27356 83298 27412 83310
rect 27356 83246 27358 83298
rect 27410 83246 27412 83298
rect 27244 82740 27300 82750
rect 27244 82646 27300 82684
rect 27132 82574 27134 82626
rect 27186 82574 27188 82626
rect 27132 81844 27188 82574
rect 27244 82180 27300 82190
rect 27244 82066 27300 82124
rect 27244 82014 27246 82066
rect 27298 82014 27300 82066
rect 27244 82002 27300 82014
rect 27132 81788 27300 81844
rect 27020 81218 27076 81228
rect 26908 81118 26910 81170
rect 26962 81118 26964 81170
rect 26908 80724 26964 81118
rect 27132 81172 27188 81182
rect 27132 81078 27188 81116
rect 26908 80658 26964 80668
rect 27244 80610 27300 81788
rect 27356 81172 27412 83246
rect 27468 82850 27524 82862
rect 27468 82798 27470 82850
rect 27522 82798 27524 82850
rect 27468 82292 27524 82798
rect 27468 82226 27524 82236
rect 27692 82180 27748 82190
rect 27804 82180 27860 85652
rect 28140 85204 28196 87278
rect 28428 86268 28692 86278
rect 28484 86212 28532 86268
rect 28588 86212 28636 86268
rect 28428 86202 28692 86212
rect 28140 85138 28196 85148
rect 27916 84980 27972 84990
rect 27916 84886 27972 84924
rect 28428 84700 28692 84710
rect 28140 84644 28196 84654
rect 28484 84644 28532 84700
rect 28588 84644 28636 84700
rect 28428 84634 28692 84644
rect 28028 84194 28084 84206
rect 28028 84142 28030 84194
rect 28082 84142 28084 84194
rect 28028 84082 28084 84142
rect 28028 84030 28030 84082
rect 28082 84030 28084 84082
rect 28028 84018 28084 84030
rect 28028 83298 28084 83310
rect 28028 83246 28030 83298
rect 28082 83246 28084 83298
rect 28028 82852 28084 83246
rect 28028 82786 28084 82796
rect 28028 82628 28084 82638
rect 27580 82178 27860 82180
rect 27580 82126 27694 82178
rect 27746 82126 27860 82178
rect 27580 82124 27860 82126
rect 27916 82626 28084 82628
rect 27916 82574 28030 82626
rect 28082 82574 28084 82626
rect 27916 82572 28084 82574
rect 27468 81956 27524 81966
rect 27468 81862 27524 81900
rect 27356 81106 27412 81116
rect 27468 80836 27524 80846
rect 27244 80558 27246 80610
rect 27298 80558 27300 80610
rect 27244 80546 27300 80558
rect 27356 80780 27468 80836
rect 27020 80500 27076 80510
rect 27020 80406 27076 80444
rect 26236 79734 26292 79772
rect 26460 79826 26852 79828
rect 26460 79774 26686 79826
rect 26738 79774 26852 79826
rect 26460 79772 26852 79774
rect 27132 80052 27188 80062
rect 27132 79826 27188 79996
rect 27132 79774 27134 79826
rect 27186 79774 27188 79826
rect 25452 79660 25620 79716
rect 25004 79538 25060 79548
rect 25452 79490 25508 79502
rect 25452 79438 25454 79490
rect 25506 79438 25508 79490
rect 25026 79212 25290 79222
rect 25082 79156 25130 79212
rect 25186 79156 25234 79212
rect 25026 79146 25290 79156
rect 25340 79042 25396 79054
rect 25340 78990 25342 79042
rect 25394 78990 25396 79042
rect 24668 78596 24724 78606
rect 25116 78596 25172 78606
rect 24668 78594 24836 78596
rect 24668 78542 24670 78594
rect 24722 78542 24836 78594
rect 24668 78540 24836 78542
rect 24668 78530 24724 78540
rect 24668 77922 24724 77934
rect 24668 77870 24670 77922
rect 24722 77870 24724 77922
rect 24668 77812 24724 77870
rect 24668 77746 24724 77756
rect 24780 77252 24836 78540
rect 25116 78502 25172 78540
rect 25340 78034 25396 78990
rect 25340 77982 25342 78034
rect 25394 77982 25396 78034
rect 25340 77970 25396 77982
rect 25026 77644 25290 77654
rect 25082 77588 25130 77644
rect 25186 77588 25234 77644
rect 25026 77578 25290 77588
rect 25452 77476 25508 79438
rect 25564 79042 25620 79660
rect 25788 79604 25844 79614
rect 25788 79510 25844 79548
rect 25564 78990 25566 79042
rect 25618 78990 25620 79042
rect 25564 78932 25620 78990
rect 25564 78866 25620 78876
rect 26460 78930 26516 79772
rect 26684 79762 26740 79772
rect 27132 79762 27188 79774
rect 27356 79604 27412 80780
rect 27468 80770 27524 80780
rect 27580 80610 27636 82124
rect 27692 82114 27748 82124
rect 27580 80558 27582 80610
rect 27634 80558 27636 80610
rect 27580 80546 27636 80558
rect 27916 79828 27972 82572
rect 28028 82562 28084 82572
rect 28140 82404 28196 84588
rect 28028 82348 28196 82404
rect 28252 84082 28308 84094
rect 28252 84030 28254 84082
rect 28306 84030 28308 84082
rect 28028 81058 28084 82348
rect 28140 81730 28196 81742
rect 28140 81678 28142 81730
rect 28194 81678 28196 81730
rect 28140 81170 28196 81678
rect 28140 81118 28142 81170
rect 28194 81118 28196 81170
rect 28140 81106 28196 81118
rect 28028 81006 28030 81058
rect 28082 81006 28084 81058
rect 28028 80994 28084 81006
rect 28028 80836 28084 80846
rect 28028 80498 28084 80780
rect 28028 80446 28030 80498
rect 28082 80446 28084 80498
rect 28028 80434 28084 80446
rect 28252 79940 28308 84030
rect 28428 83132 28692 83142
rect 28484 83076 28532 83132
rect 28588 83076 28636 83132
rect 28428 83066 28692 83076
rect 28428 81564 28692 81574
rect 28484 81508 28532 81564
rect 28588 81508 28636 81564
rect 28428 81498 28692 81508
rect 27916 79762 27972 79772
rect 28028 79884 28308 79940
rect 28428 79996 28692 80006
rect 28484 79940 28532 79996
rect 28588 79940 28636 79996
rect 28428 79930 28692 79940
rect 28028 79826 28084 79884
rect 28028 79774 28030 79826
rect 28082 79774 28084 79826
rect 26460 78878 26462 78930
rect 26514 78878 26516 78930
rect 25676 78594 25732 78606
rect 25676 78542 25678 78594
rect 25730 78542 25732 78594
rect 25452 77420 25620 77476
rect 25228 77364 25284 77374
rect 25228 77362 25508 77364
rect 25228 77310 25230 77362
rect 25282 77310 25508 77362
rect 25228 77308 25508 77310
rect 25228 77298 25284 77308
rect 24780 77186 24836 77196
rect 24444 76690 24612 76692
rect 24444 76638 24446 76690
rect 24498 76638 24612 76690
rect 24444 76636 24612 76638
rect 24668 77138 24724 77150
rect 24668 77086 24670 77138
rect 24722 77086 24724 77138
rect 24668 77028 24724 77086
rect 24444 76242 24500 76636
rect 24444 76190 24446 76242
rect 24498 76190 24500 76242
rect 24444 76178 24500 76190
rect 24556 75908 24612 75918
rect 24668 75908 24724 76972
rect 24892 77138 24948 77150
rect 24892 77086 24894 77138
rect 24946 77086 24948 77138
rect 24892 76692 24948 77086
rect 24892 76626 24948 76636
rect 25340 76804 25396 76814
rect 25340 76690 25396 76748
rect 25340 76638 25342 76690
rect 25394 76638 25396 76690
rect 25340 76626 25396 76638
rect 25026 76076 25290 76086
rect 25082 76020 25130 76076
rect 25186 76020 25234 76076
rect 25026 76010 25290 76020
rect 24612 75852 24724 75908
rect 24556 75842 24612 75852
rect 24780 75796 24836 75806
rect 24668 75124 24724 75134
rect 24220 75122 24724 75124
rect 24220 75070 24670 75122
rect 24722 75070 24724 75122
rect 24220 75068 24724 75070
rect 24220 74788 24276 75068
rect 24668 75058 24724 75068
rect 24220 74786 24388 74788
rect 24220 74734 24222 74786
rect 24274 74734 24388 74786
rect 24220 74732 24388 74734
rect 24220 74722 24276 74732
rect 24220 74228 24276 74238
rect 24220 74134 24276 74172
rect 23996 74060 24164 74116
rect 23548 74004 23604 74060
rect 23212 73826 23268 73836
rect 23324 73948 23604 74004
rect 24108 73948 24164 74060
rect 22988 73378 23044 73388
rect 22988 73220 23044 73230
rect 22988 73126 23044 73164
rect 23212 73108 23268 73118
rect 22764 72100 22820 72940
rect 23100 73052 23212 73108
rect 22988 72548 23044 72558
rect 22988 72454 23044 72492
rect 23100 72324 23156 73052
rect 23212 73042 23268 73052
rect 23212 72548 23268 72558
rect 23324 72548 23380 73948
rect 23660 73892 23716 73902
rect 23660 73780 23716 73836
rect 23884 73892 23940 73902
rect 24108 73892 24276 73948
rect 23660 73724 23828 73780
rect 23548 73668 23604 73678
rect 23548 73554 23604 73612
rect 23548 73502 23550 73554
rect 23602 73502 23604 73554
rect 23548 73490 23604 73502
rect 23660 73556 23716 73566
rect 23436 73330 23492 73342
rect 23436 73278 23438 73330
rect 23490 73278 23492 73330
rect 23436 72772 23492 73278
rect 23436 72706 23492 72716
rect 23548 73332 23604 73342
rect 23436 72548 23492 72558
rect 23324 72546 23492 72548
rect 23324 72494 23438 72546
rect 23490 72494 23492 72546
rect 23324 72492 23492 72494
rect 23212 72454 23268 72492
rect 23436 72482 23492 72492
rect 23324 72324 23380 72334
rect 23548 72324 23604 73276
rect 23100 72322 23380 72324
rect 23100 72270 23326 72322
rect 23378 72270 23380 72322
rect 23100 72268 23380 72270
rect 23324 72258 23380 72268
rect 23436 72322 23604 72324
rect 23436 72270 23550 72322
rect 23602 72270 23604 72322
rect 23436 72268 23604 72270
rect 22764 72044 22932 72100
rect 22652 71932 22820 71988
rect 22652 71762 22708 71774
rect 22652 71710 22654 71762
rect 22706 71710 22708 71762
rect 22204 71038 22206 71090
rect 22258 71038 22260 71090
rect 22204 71026 22260 71038
rect 22540 71540 22596 71550
rect 22092 70812 22484 70868
rect 21624 70588 21888 70598
rect 21680 70532 21728 70588
rect 21784 70532 21832 70588
rect 21980 70578 22036 70588
rect 21624 70522 21888 70532
rect 21644 70420 21700 70430
rect 21644 69522 21700 70364
rect 22092 70194 22148 70206
rect 22092 70142 22094 70194
rect 22146 70142 22148 70194
rect 21756 70084 21812 70094
rect 21756 69990 21812 70028
rect 21644 69470 21646 69522
rect 21698 69470 21700 69522
rect 21644 69458 21700 69470
rect 21980 69524 22036 69534
rect 22092 69524 22148 70142
rect 21980 69522 22372 69524
rect 21980 69470 21982 69522
rect 22034 69470 22372 69522
rect 21980 69468 22372 69470
rect 21980 69458 22036 69468
rect 22316 69410 22372 69468
rect 22316 69358 22318 69410
rect 22370 69358 22372 69410
rect 21624 69020 21888 69030
rect 21680 68964 21728 69020
rect 21784 68964 21832 69020
rect 21624 68954 21888 68964
rect 22316 68626 22372 69358
rect 22316 68574 22318 68626
rect 22370 68574 22372 68626
rect 22316 68562 22372 68574
rect 21756 68516 21812 68526
rect 21756 68422 21812 68460
rect 21420 68114 21476 68124
rect 21644 67956 21700 67966
rect 21420 67954 21700 67956
rect 21420 67902 21646 67954
rect 21698 67902 21700 67954
rect 21420 67900 21700 67902
rect 21420 66948 21476 67900
rect 21644 67890 21700 67900
rect 21868 67844 21924 67854
rect 21868 67750 21924 67788
rect 21532 67732 21588 67742
rect 21532 67638 21588 67676
rect 22204 67732 22260 67742
rect 22204 67620 22260 67676
rect 22316 67620 22372 67630
rect 22204 67618 22372 67620
rect 22204 67566 22318 67618
rect 22370 67566 22372 67618
rect 22204 67564 22372 67566
rect 21624 67452 21888 67462
rect 21680 67396 21728 67452
rect 21784 67396 21832 67452
rect 21624 67386 21888 67396
rect 21420 66892 21588 66948
rect 21196 66780 21476 66836
rect 21196 66612 21252 66622
rect 20860 65548 21028 65604
rect 21084 66276 21140 66286
rect 20748 64596 20804 64606
rect 20748 64482 20804 64540
rect 20748 64430 20750 64482
rect 20802 64430 20804 64482
rect 20748 64418 20804 64430
rect 20748 64260 20804 64270
rect 20748 63700 20804 64204
rect 20748 63634 20804 63644
rect 20188 63532 20692 63588
rect 20076 63140 20132 63150
rect 20076 63046 20132 63084
rect 19740 60734 19742 60786
rect 19794 60734 19796 60786
rect 19404 60508 19572 60564
rect 19628 60564 19684 60574
rect 19404 58546 19460 60508
rect 19628 60470 19684 60508
rect 19516 60340 19572 60350
rect 19516 60226 19572 60284
rect 19516 60174 19518 60226
rect 19570 60174 19572 60226
rect 19516 60162 19572 60174
rect 19740 60116 19796 60734
rect 19628 60060 19796 60116
rect 19852 62132 20020 62188
rect 20188 62578 20244 63532
rect 20188 62526 20190 62578
rect 20242 62526 20244 62578
rect 19516 60004 19572 60014
rect 19628 60004 19684 60060
rect 19852 60004 19908 62132
rect 19964 61458 20020 61470
rect 19964 61406 19966 61458
rect 20018 61406 20020 61458
rect 19964 61010 20020 61406
rect 19964 60958 19966 61010
rect 20018 60958 20020 61010
rect 19964 60946 20020 60958
rect 20188 60900 20244 62526
rect 20524 62914 20580 62926
rect 20524 62862 20526 62914
rect 20578 62862 20580 62914
rect 20524 62580 20580 62862
rect 20636 62580 20692 62590
rect 20524 62524 20636 62580
rect 20636 62486 20692 62524
rect 20860 62356 20916 65548
rect 20972 65378 21028 65390
rect 20972 65326 20974 65378
rect 21026 65326 21028 65378
rect 20972 65266 21028 65326
rect 20972 65214 20974 65266
rect 21026 65214 21028 65266
rect 20972 64484 21028 65214
rect 20972 64418 21028 64428
rect 20972 64148 21028 64158
rect 21084 64148 21140 66220
rect 21196 66052 21252 66556
rect 21308 66052 21364 66062
rect 21196 66050 21364 66052
rect 21196 65998 21310 66050
rect 21362 65998 21364 66050
rect 21196 65996 21364 65998
rect 21308 65986 21364 65996
rect 21308 65716 21364 65726
rect 21420 65716 21476 66780
rect 21532 66498 21588 66892
rect 21532 66446 21534 66498
rect 21586 66446 21588 66498
rect 21532 66434 21588 66446
rect 21532 66274 21588 66286
rect 21532 66222 21534 66274
rect 21586 66222 21588 66274
rect 21532 66052 21588 66222
rect 21868 66164 21924 66174
rect 22092 66164 22148 66174
rect 21868 66162 22036 66164
rect 21868 66110 21870 66162
rect 21922 66110 22036 66162
rect 21868 66108 22036 66110
rect 21868 66098 21924 66108
rect 21532 65986 21588 65996
rect 21624 65884 21888 65894
rect 21680 65828 21728 65884
rect 21784 65828 21832 65884
rect 21624 65818 21888 65828
rect 21980 65716 22036 66108
rect 21420 65660 21588 65716
rect 21308 65604 21364 65660
rect 21308 65548 21476 65604
rect 21420 65490 21476 65548
rect 21420 65438 21422 65490
rect 21474 65438 21476 65490
rect 21420 65426 21476 65438
rect 20972 64146 21140 64148
rect 20972 64094 20974 64146
rect 21026 64094 21140 64146
rect 20972 64092 21140 64094
rect 20972 64082 21028 64092
rect 20524 62300 20916 62356
rect 20972 63700 21028 63710
rect 20412 61236 20468 61246
rect 20412 61010 20468 61180
rect 20412 60958 20414 61010
rect 20466 60958 20468 61010
rect 20412 60946 20468 60958
rect 20188 60834 20244 60844
rect 19516 60002 19684 60004
rect 19516 59950 19518 60002
rect 19570 59950 19684 60002
rect 19516 59948 19684 59950
rect 19740 59948 19908 60004
rect 19964 60788 20020 60798
rect 19516 58884 19572 59948
rect 19740 59892 19796 59948
rect 19516 58818 19572 58828
rect 19628 59836 19796 59892
rect 19404 58494 19406 58546
rect 19458 58494 19460 58546
rect 19404 58482 19460 58494
rect 19516 58324 19572 58334
rect 19180 56812 19348 56868
rect 19404 58322 19572 58324
rect 19404 58270 19518 58322
rect 19570 58270 19572 58322
rect 19404 58268 19572 58270
rect 19404 57764 19460 58268
rect 19516 58258 19572 58268
rect 18956 56642 19012 56654
rect 18956 56590 18958 56642
rect 19010 56590 19012 56642
rect 18956 56084 19012 56590
rect 19068 56644 19124 56654
rect 19068 56550 19124 56588
rect 18956 56018 19012 56028
rect 19068 56420 19124 56430
rect 19068 55970 19124 56364
rect 19068 55918 19070 55970
rect 19122 55918 19124 55970
rect 19068 54180 19124 55918
rect 19180 54852 19236 56812
rect 19292 56642 19348 56654
rect 19292 56590 19294 56642
rect 19346 56590 19348 56642
rect 19292 56084 19348 56590
rect 19292 56018 19348 56028
rect 19180 54786 19236 54796
rect 19068 54124 19348 54180
rect 19068 53954 19124 53966
rect 19068 53902 19070 53954
rect 19122 53902 19124 53954
rect 18956 53508 19012 53518
rect 18956 53414 19012 53452
rect 19068 51828 19124 53902
rect 19180 53508 19236 53518
rect 19180 52834 19236 53452
rect 19180 52782 19182 52834
rect 19234 52782 19236 52834
rect 19180 52052 19236 52782
rect 19180 51986 19236 51996
rect 19068 51762 19124 51772
rect 19180 51604 19236 51614
rect 19292 51604 19348 54124
rect 19404 53508 19460 57708
rect 19516 56756 19572 56766
rect 19516 56662 19572 56700
rect 19516 56082 19572 56094
rect 19516 56030 19518 56082
rect 19570 56030 19572 56082
rect 19516 55748 19572 56030
rect 19628 55972 19684 59836
rect 19964 58660 20020 60732
rect 20300 60564 20356 60574
rect 20300 60470 20356 60508
rect 20412 60452 20468 60462
rect 20076 60340 20132 60350
rect 20076 60226 20132 60284
rect 20076 60174 20078 60226
rect 20130 60174 20132 60226
rect 20076 60162 20132 60174
rect 20412 60226 20468 60396
rect 20412 60174 20414 60226
rect 20466 60174 20468 60226
rect 20412 60162 20468 60174
rect 20076 60004 20132 60014
rect 20076 59910 20132 59948
rect 20300 59332 20356 59342
rect 20300 59238 20356 59276
rect 19852 58604 20020 58660
rect 19852 57540 19908 58604
rect 20188 58212 20244 58222
rect 19964 57764 20020 57774
rect 19964 57670 20020 57708
rect 20188 57764 20244 58156
rect 19852 57474 19908 57484
rect 19628 55906 19684 55916
rect 19852 57204 19908 57214
rect 19516 55682 19572 55692
rect 19852 55300 19908 57148
rect 20188 57090 20244 57708
rect 20188 57038 20190 57090
rect 20242 57038 20244 57090
rect 20188 57026 20244 57038
rect 19964 56642 20020 56654
rect 19964 56590 19966 56642
rect 20018 56590 20020 56642
rect 19964 55524 20020 56590
rect 20076 56642 20132 56654
rect 20076 56590 20078 56642
rect 20130 56590 20132 56642
rect 20076 56196 20132 56590
rect 20076 56140 20356 56196
rect 20188 55972 20244 56010
rect 20188 55906 20244 55916
rect 19964 55458 20020 55468
rect 20188 55748 20244 55758
rect 20076 55300 20132 55310
rect 19852 55298 20132 55300
rect 19852 55246 20078 55298
rect 20130 55246 20132 55298
rect 19852 55244 20132 55246
rect 19964 55076 20020 55086
rect 19516 55074 20020 55076
rect 19516 55022 19966 55074
rect 20018 55022 20020 55074
rect 19516 55020 20020 55022
rect 19516 54626 19572 55020
rect 19964 55010 20020 55020
rect 19516 54574 19518 54626
rect 19570 54574 19572 54626
rect 19516 54562 19572 54574
rect 19628 54852 19684 54862
rect 19628 53730 19684 54796
rect 19628 53678 19630 53730
rect 19682 53678 19684 53730
rect 19628 53666 19684 53678
rect 19740 54740 19796 54750
rect 19404 53414 19460 53452
rect 19740 53170 19796 54684
rect 20076 54180 20132 55244
rect 20076 54114 20132 54124
rect 20188 54514 20244 55692
rect 20300 55522 20356 56140
rect 20300 55470 20302 55522
rect 20354 55470 20356 55522
rect 20300 55458 20356 55470
rect 20524 55412 20580 62300
rect 20972 61796 21028 63644
rect 21084 63698 21140 64092
rect 21084 63646 21086 63698
rect 21138 63646 21140 63698
rect 21084 63634 21140 63646
rect 21308 64932 21364 64942
rect 21308 64706 21364 64876
rect 21532 64932 21588 65660
rect 21980 65650 22036 65660
rect 21868 65378 21924 65390
rect 21868 65326 21870 65378
rect 21922 65326 21924 65378
rect 21868 65156 21924 65326
rect 22092 65266 22148 66108
rect 22092 65214 22094 65266
rect 22146 65214 22148 65266
rect 22092 65202 22148 65214
rect 21868 65090 21924 65100
rect 21532 64866 21588 64876
rect 21308 64654 21310 64706
rect 21362 64654 21364 64706
rect 21308 64036 21364 64654
rect 22092 64596 22148 64606
rect 22092 64502 22148 64540
rect 22204 64372 22260 67564
rect 22316 67554 22372 67564
rect 22428 65828 22484 70812
rect 22540 66164 22596 71484
rect 22540 66070 22596 66108
rect 22428 65762 22484 65772
rect 22316 65604 22372 65614
rect 22316 65378 22372 65548
rect 22316 65326 22318 65378
rect 22370 65326 22372 65378
rect 22316 64820 22372 65326
rect 22316 64754 22372 64764
rect 22428 65492 22484 65502
rect 21624 64316 21888 64326
rect 21680 64260 21728 64316
rect 21784 64260 21832 64316
rect 21624 64250 21888 64260
rect 22092 64316 22260 64372
rect 21868 64148 21924 64158
rect 21868 64054 21924 64092
rect 21308 62356 21364 63980
rect 21756 63922 21812 63934
rect 21756 63870 21758 63922
rect 21810 63870 21812 63922
rect 21756 63812 21812 63870
rect 21756 63746 21812 63756
rect 21420 63698 21476 63710
rect 21420 63646 21422 63698
rect 21474 63646 21476 63698
rect 21420 63138 21476 63646
rect 21644 63700 21700 63710
rect 21644 63606 21700 63644
rect 22092 63700 22148 64316
rect 22316 64260 22372 64270
rect 22092 63634 22148 63644
rect 22204 64204 22316 64260
rect 21420 63086 21422 63138
rect 21474 63086 21476 63138
rect 21420 63074 21476 63086
rect 21624 62748 21888 62758
rect 21680 62692 21728 62748
rect 21784 62692 21832 62748
rect 21624 62682 21888 62692
rect 21308 62354 21476 62356
rect 21308 62302 21310 62354
rect 21362 62302 21476 62354
rect 21308 62300 21476 62302
rect 21308 62290 21364 62300
rect 20636 61740 21028 61796
rect 20636 61348 20692 61740
rect 21420 61684 21476 62300
rect 22092 62244 22148 62282
rect 22092 62178 22148 62188
rect 20748 61682 21476 61684
rect 20748 61630 21422 61682
rect 21474 61630 21476 61682
rect 20748 61628 21476 61630
rect 20748 61570 20804 61628
rect 20748 61518 20750 61570
rect 20802 61518 20804 61570
rect 20748 61506 20804 61518
rect 20636 61292 20804 61348
rect 20636 60564 20692 60574
rect 20636 60470 20692 60508
rect 20636 59892 20692 59902
rect 20636 58660 20692 59836
rect 20636 58546 20692 58604
rect 20636 58494 20638 58546
rect 20690 58494 20692 58546
rect 20636 58482 20692 58494
rect 20748 57764 20804 61292
rect 20748 57698 20804 57708
rect 20972 60900 21028 60910
rect 20636 56642 20692 56654
rect 20636 56590 20638 56642
rect 20690 56590 20692 56642
rect 20636 56308 20692 56590
rect 20636 56242 20692 56252
rect 20748 55412 20804 55422
rect 20524 55356 20692 55412
rect 20188 54462 20190 54514
rect 20242 54462 20244 54514
rect 20076 53730 20132 53742
rect 20076 53678 20078 53730
rect 20130 53678 20132 53730
rect 20076 53620 20132 53678
rect 20076 53554 20132 53564
rect 19740 53118 19742 53170
rect 19794 53118 19796 53170
rect 19740 53106 19796 53118
rect 19740 52836 19796 52846
rect 19740 52274 19796 52780
rect 20076 52388 20132 52398
rect 19740 52222 19742 52274
rect 19794 52222 19796 52274
rect 19740 52210 19796 52222
rect 19964 52276 20020 52286
rect 19964 52162 20020 52220
rect 19964 52110 19966 52162
rect 20018 52110 20020 52162
rect 19964 52098 20020 52110
rect 20076 52162 20132 52332
rect 20076 52110 20078 52162
rect 20130 52110 20132 52162
rect 20076 52098 20132 52110
rect 19236 51548 19348 51604
rect 19404 51828 19460 51838
rect 19404 51602 19460 51772
rect 19404 51550 19406 51602
rect 19458 51550 19460 51602
rect 19180 51538 19236 51548
rect 19404 51538 19460 51550
rect 19740 51604 19796 51614
rect 19740 51510 19796 51548
rect 19180 51378 19236 51390
rect 19180 51326 19182 51378
rect 19234 51326 19236 51378
rect 19180 50708 19236 51326
rect 19180 50642 19236 50652
rect 19628 51380 19684 51390
rect 19628 50820 19684 51324
rect 20188 51378 20244 54462
rect 20524 55186 20580 55198
rect 20524 55134 20526 55186
rect 20578 55134 20580 55186
rect 20524 54628 20580 55134
rect 20524 54292 20580 54572
rect 20524 54226 20580 54236
rect 20300 54068 20356 54078
rect 20636 54068 20692 55356
rect 20748 55186 20804 55356
rect 20972 55300 21028 60844
rect 21084 59218 21140 61628
rect 21420 61618 21476 61628
rect 21980 61346 22036 61358
rect 21980 61294 21982 61346
rect 22034 61294 22036 61346
rect 21624 61180 21888 61190
rect 21680 61124 21728 61180
rect 21784 61124 21832 61180
rect 21624 61114 21888 61124
rect 21308 60788 21364 60798
rect 21084 59166 21086 59218
rect 21138 59166 21140 59218
rect 21084 58212 21140 59166
rect 21084 58146 21140 58156
rect 21196 60676 21252 60686
rect 21196 57650 21252 60620
rect 21196 57598 21198 57650
rect 21250 57598 21252 57650
rect 21196 56196 21252 57598
rect 21196 56130 21252 56140
rect 21308 55748 21364 60732
rect 21868 60788 21924 60798
rect 21980 60788 22036 61294
rect 21868 60786 22036 60788
rect 21868 60734 21870 60786
rect 21922 60734 22036 60786
rect 21868 60732 22036 60734
rect 21420 60564 21476 60574
rect 21420 58212 21476 60508
rect 21868 60564 21924 60732
rect 21868 60498 21924 60508
rect 22092 60676 22148 60686
rect 21644 60116 21700 60126
rect 21644 60022 21700 60060
rect 21624 59612 21888 59622
rect 21680 59556 21728 59612
rect 21784 59556 21832 59612
rect 21624 59546 21888 59556
rect 21532 59106 21588 59118
rect 21532 59054 21534 59106
rect 21586 59054 21588 59106
rect 21532 58884 21588 59054
rect 21980 59108 22036 59118
rect 22092 59108 22148 60620
rect 21980 59106 22148 59108
rect 21980 59054 21982 59106
rect 22034 59054 22148 59106
rect 21980 59052 22148 59054
rect 21980 59042 22036 59052
rect 21532 58818 21588 58828
rect 21868 58212 21924 58222
rect 21420 58210 22036 58212
rect 21420 58158 21422 58210
rect 21474 58158 21870 58210
rect 21922 58158 22036 58210
rect 21420 58156 22036 58158
rect 21420 58146 21476 58156
rect 21868 58146 21924 58156
rect 21624 58044 21888 58054
rect 21680 57988 21728 58044
rect 21784 57988 21832 58044
rect 21624 57978 21888 57988
rect 21644 57764 21700 57774
rect 21644 57670 21700 57708
rect 21980 57204 22036 58156
rect 21980 57138 22036 57148
rect 21980 56868 22036 56878
rect 21420 56756 21476 56766
rect 21420 56662 21476 56700
rect 21624 56476 21888 56486
rect 21680 56420 21728 56476
rect 21784 56420 21832 56476
rect 21624 56410 21888 56420
rect 21532 56308 21588 56318
rect 20972 55234 21028 55244
rect 21196 55692 21364 55748
rect 21420 55972 21476 55982
rect 20748 55134 20750 55186
rect 20802 55134 20804 55186
rect 20748 54292 20804 55134
rect 20860 55076 20916 55086
rect 21196 55076 21252 55692
rect 21308 55524 21364 55534
rect 21308 55298 21364 55468
rect 21420 55410 21476 55916
rect 21420 55358 21422 55410
rect 21474 55358 21476 55410
rect 21420 55346 21476 55358
rect 21308 55246 21310 55298
rect 21362 55246 21364 55298
rect 21308 55234 21364 55246
rect 21532 55188 21588 56252
rect 21868 55748 21924 55758
rect 21980 55748 22036 56812
rect 21924 55692 22036 55748
rect 21868 55682 21924 55692
rect 22092 55636 22148 59052
rect 22204 58546 22260 64204
rect 22316 64194 22372 64204
rect 22428 64036 22484 65436
rect 22652 65156 22708 71710
rect 22428 63942 22484 63980
rect 22540 65100 22708 65156
rect 22204 58494 22206 58546
rect 22258 58494 22260 58546
rect 22204 56308 22260 58494
rect 22316 63588 22372 63598
rect 22316 61458 22372 63532
rect 22428 62244 22484 62254
rect 22428 61682 22484 62188
rect 22428 61630 22430 61682
rect 22482 61630 22484 61682
rect 22428 61618 22484 61630
rect 22316 61406 22318 61458
rect 22370 61406 22372 61458
rect 22316 61236 22372 61406
rect 22316 58548 22372 61180
rect 22428 60676 22484 60686
rect 22428 60582 22484 60620
rect 22428 59780 22484 59790
rect 22540 59780 22596 65100
rect 22764 64708 22820 71932
rect 22876 68068 22932 72044
rect 23436 71762 23492 72268
rect 23548 72258 23604 72268
rect 23548 71988 23604 71998
rect 23660 71988 23716 73500
rect 23772 73330 23828 73724
rect 23772 73278 23774 73330
rect 23826 73278 23828 73330
rect 23772 72324 23828 73278
rect 23772 72258 23828 72268
rect 23548 71986 23716 71988
rect 23548 71934 23550 71986
rect 23602 71934 23716 71986
rect 23548 71932 23716 71934
rect 23548 71922 23604 71932
rect 23436 71710 23438 71762
rect 23490 71710 23492 71762
rect 23436 71540 23492 71710
rect 23772 71762 23828 71774
rect 23772 71710 23774 71762
rect 23826 71710 23828 71762
rect 23660 71652 23716 71662
rect 23660 71558 23716 71596
rect 23436 71474 23492 71484
rect 23436 71316 23492 71326
rect 23772 71316 23828 71710
rect 23492 71260 23828 71316
rect 23324 70980 23380 70990
rect 23100 70868 23156 70878
rect 22876 68002 22932 68012
rect 22988 68516 23044 68526
rect 22876 67844 22932 67854
rect 22876 66948 22932 67788
rect 22988 67618 23044 68460
rect 23100 68292 23156 70812
rect 23324 70084 23380 70924
rect 23324 70018 23380 70028
rect 23436 68516 23492 71260
rect 23884 70082 23940 73836
rect 23996 73444 24052 73454
rect 23996 73350 24052 73388
rect 24108 72324 24164 72334
rect 24108 72230 24164 72268
rect 24220 71988 24276 73892
rect 24332 73780 24388 74732
rect 24780 74114 24836 75740
rect 25228 75684 25284 75694
rect 25228 75460 25284 75628
rect 25228 75394 25284 75404
rect 24892 74676 24948 74686
rect 24892 74340 24948 74620
rect 25026 74508 25290 74518
rect 25082 74452 25130 74508
rect 25186 74452 25234 74508
rect 25026 74442 25290 74452
rect 24892 74284 25060 74340
rect 24780 74062 24782 74114
rect 24834 74062 24836 74114
rect 24556 73892 24612 73902
rect 24556 73798 24612 73836
rect 24668 73890 24724 73902
rect 24668 73838 24670 73890
rect 24722 73838 24724 73890
rect 24332 73714 24388 73724
rect 24332 73444 24388 73454
rect 24668 73444 24724 73838
rect 24388 73388 24724 73444
rect 24332 73378 24388 73388
rect 24780 73332 24836 74062
rect 25004 74228 25060 74284
rect 25004 74002 25060 74172
rect 25004 73950 25006 74002
rect 25058 73950 25060 74002
rect 25004 73938 25060 73950
rect 24444 73276 24836 73332
rect 24892 73892 24948 73902
rect 24444 73218 24500 73276
rect 24444 73166 24446 73218
rect 24498 73166 24500 73218
rect 24444 73154 24500 73166
rect 24332 73106 24388 73118
rect 24332 73054 24334 73106
rect 24386 73054 24388 73106
rect 24332 72548 24388 73054
rect 24668 72996 24724 73006
rect 24724 72940 24836 72996
rect 24668 72930 24724 72940
rect 24332 72492 24724 72548
rect 24556 72324 24612 72362
rect 24556 72258 24612 72268
rect 24556 72100 24612 72110
rect 24220 71932 24500 71988
rect 23996 71764 24052 71774
rect 24332 71764 24388 71774
rect 23996 71762 24388 71764
rect 23996 71710 23998 71762
rect 24050 71710 24334 71762
rect 24386 71710 24388 71762
rect 23996 71708 24388 71710
rect 23996 71698 24052 71708
rect 24220 71092 24276 71708
rect 24332 71698 24388 71708
rect 24332 71092 24388 71102
rect 24220 71090 24388 71092
rect 24220 71038 24334 71090
rect 24386 71038 24388 71090
rect 24220 71036 24388 71038
rect 24332 71026 24388 71036
rect 24444 70868 24500 71932
rect 24556 71986 24612 72044
rect 24556 71934 24558 71986
rect 24610 71934 24612 71986
rect 24556 71922 24612 71934
rect 24668 71764 24724 72492
rect 24668 71698 24724 71708
rect 24668 71540 24724 71550
rect 24780 71540 24836 72940
rect 24668 71538 24836 71540
rect 24668 71486 24670 71538
rect 24722 71486 24836 71538
rect 24668 71484 24836 71486
rect 24668 71474 24724 71484
rect 23884 70030 23886 70082
rect 23938 70030 23940 70082
rect 23548 69522 23604 69534
rect 23548 69470 23550 69522
rect 23602 69470 23604 69522
rect 23548 68852 23604 69470
rect 23548 68786 23604 68796
rect 23436 68450 23492 68460
rect 23100 68236 23492 68292
rect 23212 67732 23268 67742
rect 23212 67638 23268 67676
rect 22988 67566 22990 67618
rect 23042 67566 23044 67618
rect 22988 67172 23044 67566
rect 23100 67620 23156 67630
rect 23100 67526 23156 67564
rect 23324 67620 23380 67630
rect 23324 67526 23380 67564
rect 23436 67172 23492 68236
rect 22988 67116 23156 67172
rect 23436 67116 23604 67172
rect 22988 66948 23044 66958
rect 22876 66946 23044 66948
rect 22876 66894 22990 66946
rect 23042 66894 23044 66946
rect 22876 66892 23044 66894
rect 22988 66882 23044 66892
rect 22876 66276 22932 66286
rect 22876 66182 22932 66220
rect 23100 65604 23156 67116
rect 23436 66946 23492 66958
rect 23436 66894 23438 66946
rect 23490 66894 23492 66946
rect 23324 66836 23380 66846
rect 23324 65714 23380 66780
rect 23436 66276 23492 66894
rect 23436 66210 23492 66220
rect 23548 66052 23604 67116
rect 23324 65662 23326 65714
rect 23378 65662 23380 65714
rect 23324 65650 23380 65662
rect 23436 65996 23604 66052
rect 23100 65510 23156 65548
rect 22764 64642 22820 64652
rect 22876 65490 22932 65502
rect 22876 65438 22878 65490
rect 22930 65438 22932 65490
rect 22876 64820 22932 65438
rect 23212 65378 23268 65390
rect 23212 65326 23214 65378
rect 23266 65326 23268 65378
rect 23212 65268 23268 65326
rect 23212 65202 23268 65212
rect 22876 64148 22932 64764
rect 23436 64260 23492 65996
rect 23548 65490 23604 65502
rect 23548 65438 23550 65490
rect 23602 65438 23604 65490
rect 23548 65268 23604 65438
rect 23548 65202 23604 65212
rect 23436 64194 23492 64204
rect 22876 64082 22932 64092
rect 23100 63924 23156 63934
rect 23100 63830 23156 63868
rect 23548 63922 23604 63934
rect 23548 63870 23550 63922
rect 23602 63870 23604 63922
rect 22876 63810 22932 63822
rect 22876 63758 22878 63810
rect 22930 63758 22932 63810
rect 22876 63700 22932 63758
rect 22876 63634 22932 63644
rect 23436 63812 23492 63822
rect 23100 63476 23156 63486
rect 22876 63028 22932 63038
rect 22652 61572 22708 61582
rect 22652 61478 22708 61516
rect 22876 61570 22932 62972
rect 22876 61518 22878 61570
rect 22930 61518 22932 61570
rect 22876 61506 22932 61518
rect 23100 62580 23156 63420
rect 23100 60676 23156 62524
rect 23436 62916 23492 63756
rect 23100 60610 23156 60620
rect 23212 62244 23268 62254
rect 23100 60452 23156 60462
rect 22764 60340 22820 60350
rect 22764 60228 22820 60284
rect 22764 60172 22932 60228
rect 22484 59724 22596 59780
rect 22764 59892 22820 59902
rect 22428 59714 22484 59724
rect 22652 59444 22708 59454
rect 22316 58482 22372 58492
rect 22428 59388 22652 59444
rect 22316 58212 22372 58222
rect 22316 56868 22372 58156
rect 22316 56802 22372 56812
rect 22204 56242 22260 56252
rect 22428 56084 22484 59388
rect 22652 59378 22708 59388
rect 22764 59442 22820 59836
rect 22764 59390 22766 59442
rect 22818 59390 22820 59442
rect 22764 59378 22820 59390
rect 22876 59330 22932 60172
rect 22876 59278 22878 59330
rect 22930 59278 22932 59330
rect 22540 59218 22596 59230
rect 22540 59166 22542 59218
rect 22594 59166 22596 59218
rect 22540 58658 22596 59166
rect 22876 58828 22932 59278
rect 22988 59220 23044 59230
rect 22988 59126 23044 59164
rect 22540 58606 22542 58658
rect 22594 58606 22596 58658
rect 22540 58594 22596 58606
rect 22764 58772 22932 58828
rect 22764 58210 22820 58772
rect 22764 58158 22766 58210
rect 22818 58158 22820 58210
rect 22540 57540 22596 57550
rect 22540 57446 22596 57484
rect 22764 57316 22820 58158
rect 22876 58548 22932 58558
rect 22876 57762 22932 58492
rect 22876 57710 22878 57762
rect 22930 57710 22932 57762
rect 22876 57698 22932 57710
rect 22540 57260 22820 57316
rect 22988 57538 23044 57550
rect 22988 57486 22990 57538
rect 23042 57486 23044 57538
rect 22540 56308 22596 57260
rect 22988 57204 23044 57486
rect 22652 57148 23044 57204
rect 22652 56978 22708 57148
rect 22652 56926 22654 56978
rect 22706 56926 22708 56978
rect 22652 56914 22708 56926
rect 22540 56242 22596 56252
rect 22652 56196 22708 56206
rect 22428 56028 22596 56084
rect 22316 55972 22372 55982
rect 22316 55970 22484 55972
rect 22316 55918 22318 55970
rect 22370 55918 22484 55970
rect 22316 55916 22484 55918
rect 22316 55906 22372 55916
rect 22092 55570 22148 55580
rect 22316 55524 22372 55534
rect 21756 55412 22372 55468
rect 21420 55132 21588 55188
rect 21644 55188 21700 55198
rect 21756 55188 21812 55412
rect 21868 55300 21924 55310
rect 22316 55300 22372 55310
rect 21868 55298 22372 55300
rect 21868 55246 21870 55298
rect 21922 55246 22318 55298
rect 22370 55246 22372 55298
rect 21868 55244 22372 55246
rect 21868 55234 21924 55244
rect 22316 55234 22372 55244
rect 21700 55132 21812 55188
rect 21196 55020 21364 55076
rect 20860 54404 20916 55020
rect 21084 54628 21140 54638
rect 20972 54514 21028 54526
rect 20972 54462 20974 54514
rect 21026 54462 21028 54514
rect 20972 54404 21028 54462
rect 20916 54348 21028 54404
rect 21084 54404 21140 54572
rect 21196 54516 21252 54526
rect 21196 54422 21252 54460
rect 20860 54338 20916 54348
rect 21084 54338 21140 54348
rect 20748 54226 20804 54236
rect 21196 54292 21252 54302
rect 20636 54012 20804 54068
rect 20300 53732 20356 54012
rect 20300 53638 20356 53676
rect 20636 53732 20692 53742
rect 20636 53638 20692 53676
rect 20524 53618 20580 53630
rect 20524 53566 20526 53618
rect 20578 53566 20580 53618
rect 20300 53508 20356 53518
rect 20524 53508 20580 53566
rect 20356 53452 20580 53508
rect 20300 53442 20356 53452
rect 20300 53172 20356 53182
rect 20300 52946 20356 53116
rect 20524 53060 20580 53070
rect 20524 52966 20580 53004
rect 20636 53058 20692 53070
rect 20636 53006 20638 53058
rect 20690 53006 20692 53058
rect 20300 52894 20302 52946
rect 20354 52894 20356 52946
rect 20300 52882 20356 52894
rect 20636 52948 20692 53006
rect 20636 52882 20692 52892
rect 20188 51326 20190 51378
rect 20242 51326 20244 51378
rect 19628 50706 19684 50764
rect 19628 50654 19630 50706
rect 19682 50654 19684 50706
rect 19628 50642 19684 50654
rect 19964 51156 20020 51166
rect 19180 50482 19236 50494
rect 19180 50430 19182 50482
rect 19234 50430 19236 50482
rect 19180 50372 19236 50430
rect 19180 50306 19236 50316
rect 18844 50092 19460 50148
rect 18564 49868 18676 49924
rect 18508 49830 18564 49868
rect 18222 49420 18486 49430
rect 18278 49364 18326 49420
rect 18382 49364 18430 49420
rect 18222 49354 18486 49364
rect 18620 49026 18676 49868
rect 18620 48974 18622 49026
rect 18674 48974 18676 49026
rect 18620 48962 18676 48974
rect 18956 49812 19012 49822
rect 18956 49028 19012 49756
rect 18956 48934 19012 48972
rect 19068 49700 19124 49710
rect 18844 48914 18900 48926
rect 18844 48862 18846 48914
rect 18898 48862 18900 48914
rect 18222 47852 18486 47862
rect 18278 47796 18326 47852
rect 18382 47796 18430 47852
rect 18222 47786 18486 47796
rect 18396 47684 18452 47694
rect 18060 47292 18228 47348
rect 17612 45266 17668 45276
rect 17724 47180 17892 47236
rect 17948 47236 18004 47246
rect 17500 44548 17556 44558
rect 17500 44322 17556 44492
rect 17500 44270 17502 44322
rect 17554 44270 17556 44322
rect 17500 44258 17556 44270
rect 17500 44100 17556 44110
rect 17556 44044 17668 44100
rect 17500 44034 17556 44044
rect 17612 43650 17668 44044
rect 17612 43598 17614 43650
rect 17666 43598 17668 43650
rect 17612 43586 17668 43598
rect 17612 42308 17668 42318
rect 17724 42308 17780 47180
rect 17836 47012 17892 47022
rect 17836 45890 17892 46956
rect 17948 46786 18004 47180
rect 18172 47068 18228 47292
rect 18396 47346 18452 47628
rect 18396 47294 18398 47346
rect 18450 47294 18452 47346
rect 18396 47282 18452 47294
rect 18620 47460 18676 47470
rect 17948 46734 17950 46786
rect 18002 46734 18004 46786
rect 17948 46722 18004 46734
rect 18060 47012 18228 47068
rect 17836 45838 17838 45890
rect 17890 45838 17892 45890
rect 17836 45780 17892 45838
rect 17836 45714 17892 45724
rect 17948 44994 18004 45006
rect 17948 44942 17950 44994
rect 18002 44942 18004 44994
rect 17948 44884 18004 44942
rect 17836 44828 18004 44884
rect 17836 44548 17892 44828
rect 17836 44482 17892 44492
rect 17948 44660 18004 44670
rect 17948 44100 18004 44604
rect 17836 44044 18004 44100
rect 17836 43538 17892 44044
rect 17836 43486 17838 43538
rect 17890 43486 17892 43538
rect 17836 43474 17892 43486
rect 17948 43652 18004 43662
rect 17948 42866 18004 43596
rect 17948 42814 17950 42866
rect 18002 42814 18004 42866
rect 17948 42802 18004 42814
rect 17724 42252 18004 42308
rect 17612 42196 17668 42252
rect 17612 42140 17892 42196
rect 17500 41970 17556 41982
rect 17500 41918 17502 41970
rect 17554 41918 17556 41970
rect 17500 39620 17556 41918
rect 17612 41972 17668 41982
rect 17612 41878 17668 41916
rect 17724 41970 17780 41982
rect 17724 41918 17726 41970
rect 17778 41918 17780 41970
rect 17724 41524 17780 41918
rect 17724 41458 17780 41468
rect 17724 41300 17780 41310
rect 17836 41300 17892 42140
rect 17724 41298 17892 41300
rect 17724 41246 17726 41298
rect 17778 41246 17892 41298
rect 17724 41244 17892 41246
rect 17724 41234 17780 41244
rect 17500 39554 17556 39564
rect 17724 40402 17780 40414
rect 17724 40350 17726 40402
rect 17778 40350 17780 40402
rect 17388 39508 17444 39518
rect 17388 37492 17444 39452
rect 17724 39396 17780 40350
rect 17724 38948 17780 39340
rect 17500 38892 17780 38948
rect 17836 39842 17892 39854
rect 17836 39790 17838 39842
rect 17890 39790 17892 39842
rect 17836 39394 17892 39790
rect 17836 39342 17838 39394
rect 17890 39342 17892 39394
rect 17836 38948 17892 39342
rect 17948 38948 18004 42252
rect 18060 39172 18116 47012
rect 18222 46284 18486 46294
rect 18278 46228 18326 46284
rect 18382 46228 18430 46284
rect 18222 46218 18486 46228
rect 18284 45892 18340 45902
rect 18620 45892 18676 47404
rect 18284 45890 18676 45892
rect 18284 45838 18286 45890
rect 18338 45838 18676 45890
rect 18284 45836 18676 45838
rect 18284 45826 18340 45836
rect 18844 45444 18900 48862
rect 18956 48804 19012 48814
rect 18956 47458 19012 48748
rect 18956 47406 18958 47458
rect 19010 47406 19012 47458
rect 18956 47394 19012 47406
rect 18732 45388 18900 45444
rect 18956 46898 19012 46910
rect 18956 46846 18958 46898
rect 19010 46846 19012 46898
rect 18396 45220 18452 45230
rect 18396 44994 18452 45164
rect 18396 44942 18398 44994
rect 18450 44942 18452 44994
rect 18396 44930 18452 44942
rect 18222 44716 18486 44726
rect 18278 44660 18326 44716
rect 18382 44660 18430 44716
rect 18222 44650 18486 44660
rect 18508 43538 18564 43550
rect 18508 43486 18510 43538
rect 18562 43486 18564 43538
rect 18172 43428 18228 43438
rect 18172 43334 18228 43372
rect 18508 43428 18564 43486
rect 18508 43362 18564 43372
rect 18222 43148 18486 43158
rect 18278 43092 18326 43148
rect 18382 43092 18430 43148
rect 18222 43082 18486 43092
rect 18172 42924 18676 42980
rect 18172 41970 18228 42924
rect 18620 42866 18676 42924
rect 18620 42814 18622 42866
rect 18674 42814 18676 42866
rect 18620 42802 18676 42814
rect 18732 42756 18788 45388
rect 18844 45220 18900 45230
rect 18844 43650 18900 45164
rect 18844 43598 18846 43650
rect 18898 43598 18900 43650
rect 18844 43586 18900 43598
rect 18732 42700 18900 42756
rect 18284 42642 18340 42654
rect 18284 42590 18286 42642
rect 18338 42590 18340 42642
rect 18284 42532 18340 42590
rect 18844 42642 18900 42700
rect 18844 42590 18846 42642
rect 18898 42590 18900 42642
rect 18284 42466 18340 42476
rect 18508 42530 18564 42542
rect 18508 42478 18510 42530
rect 18562 42478 18564 42530
rect 18508 42084 18564 42478
rect 18732 42530 18788 42542
rect 18732 42478 18734 42530
rect 18786 42478 18788 42530
rect 18732 42308 18788 42478
rect 18732 42242 18788 42252
rect 18508 42018 18564 42028
rect 18172 41918 18174 41970
rect 18226 41918 18228 41970
rect 18172 41906 18228 41918
rect 18396 41972 18452 41982
rect 18396 41878 18452 41916
rect 18844 41972 18900 42590
rect 18844 41906 18900 41916
rect 18222 41580 18486 41590
rect 18278 41524 18326 41580
rect 18382 41524 18430 41580
rect 18222 41514 18486 41524
rect 18284 41412 18340 41422
rect 18284 41074 18340 41356
rect 18844 41300 18900 41310
rect 18844 41186 18900 41244
rect 18844 41134 18846 41186
rect 18898 41134 18900 41186
rect 18844 41122 18900 41134
rect 18284 41022 18286 41074
rect 18338 41022 18340 41074
rect 18284 40404 18340 41022
rect 18620 41074 18676 41086
rect 18620 41022 18622 41074
rect 18674 41022 18676 41074
rect 18508 40962 18564 40974
rect 18508 40910 18510 40962
rect 18562 40910 18564 40962
rect 18508 40514 18564 40910
rect 18620 40628 18676 41022
rect 18620 40572 18788 40628
rect 18508 40462 18510 40514
rect 18562 40462 18564 40514
rect 18508 40450 18564 40462
rect 18284 40338 18340 40348
rect 18222 40012 18486 40022
rect 18278 39956 18326 40012
rect 18382 39956 18430 40012
rect 18222 39946 18486 39956
rect 18732 39842 18788 40572
rect 18732 39790 18734 39842
rect 18786 39790 18788 39842
rect 18732 39778 18788 39790
rect 18844 40292 18900 40302
rect 18620 39620 18676 39630
rect 18172 39396 18228 39406
rect 18172 39302 18228 39340
rect 18620 39394 18676 39564
rect 18620 39342 18622 39394
rect 18674 39342 18676 39394
rect 18060 39116 18228 39172
rect 18060 38948 18116 38958
rect 17948 38946 18116 38948
rect 17948 38894 18062 38946
rect 18114 38894 18116 38946
rect 17948 38892 18116 38894
rect 17500 38722 17556 38892
rect 17836 38882 17892 38892
rect 18060 38882 18116 38892
rect 17500 38670 17502 38722
rect 17554 38670 17556 38722
rect 17500 38164 17556 38670
rect 17500 38098 17556 38108
rect 17612 38724 17668 38734
rect 17500 37492 17556 37502
rect 17388 37490 17556 37492
rect 17388 37438 17502 37490
rect 17554 37438 17556 37490
rect 17388 37436 17556 37438
rect 17500 37426 17556 37436
rect 17612 37490 17668 38668
rect 17612 37438 17614 37490
rect 17666 37438 17668 37490
rect 17612 37426 17668 37438
rect 17948 38612 18004 38622
rect 18172 38612 18228 39116
rect 18508 38836 18564 38846
rect 18508 38742 18564 38780
rect 17388 37266 17444 37278
rect 17388 37214 17390 37266
rect 17442 37214 17444 37266
rect 17388 37156 17444 37214
rect 17388 37090 17444 37100
rect 17948 37266 18004 38556
rect 17948 37214 17950 37266
rect 18002 37214 18004 37266
rect 17948 37044 18004 37214
rect 17948 36978 18004 36988
rect 18060 38556 18228 38612
rect 18060 36820 18116 38556
rect 18222 38444 18486 38454
rect 18278 38388 18326 38444
rect 18382 38388 18430 38444
rect 18222 38378 18486 38388
rect 18396 37492 18452 37502
rect 18396 37156 18452 37436
rect 18396 37090 18452 37100
rect 17724 36764 18116 36820
rect 18222 36876 18486 36886
rect 18278 36820 18326 36876
rect 18382 36820 18430 36876
rect 18222 36810 18486 36820
rect 17276 36540 17444 36596
rect 16716 35922 16884 35924
rect 16716 35870 16718 35922
rect 16770 35870 16884 35922
rect 16716 35868 16884 35870
rect 17052 36428 17220 36484
rect 16604 35812 16660 35822
rect 16604 33572 16660 35756
rect 16604 33506 16660 33516
rect 16716 35700 16772 35868
rect 16716 34580 16772 35644
rect 17052 35308 17108 36428
rect 17164 36260 17220 36270
rect 17164 36166 17220 36204
rect 17388 35924 17444 36540
rect 17612 36372 17668 36382
rect 17612 36278 17668 36316
rect 17276 35868 17444 35924
rect 17500 36148 17556 36158
rect 17052 35252 17220 35308
rect 17052 34690 17108 34702
rect 17052 34638 17054 34690
rect 17106 34638 17108 34690
rect 17052 34580 17108 34638
rect 16716 34524 17108 34580
rect 16604 32788 16660 32798
rect 16492 32732 16604 32788
rect 16604 32722 16660 32732
rect 16268 32452 16324 32462
rect 16716 32452 16772 34524
rect 17052 33684 17108 33694
rect 16940 33572 16996 33582
rect 16268 32450 16772 32452
rect 16268 32398 16270 32450
rect 16322 32398 16772 32450
rect 16268 32396 16772 32398
rect 16828 32452 16884 32462
rect 16268 32386 16324 32396
rect 15932 32060 16100 32116
rect 15372 31042 15428 31052
rect 15484 31220 15540 31230
rect 15484 31106 15540 31164
rect 15484 31054 15486 31106
rect 15538 31054 15540 31106
rect 15484 31042 15540 31054
rect 15932 31218 15988 32060
rect 15932 31166 15934 31218
rect 15986 31166 15988 31218
rect 15708 30994 15764 31006
rect 15708 30942 15710 30994
rect 15762 30942 15764 30994
rect 15260 30828 15540 30884
rect 14812 30270 14814 30322
rect 14866 30270 14868 30322
rect 14812 30258 14868 30270
rect 15148 30098 15204 30110
rect 15148 30046 15150 30098
rect 15202 30046 15204 30098
rect 14588 29986 14644 29998
rect 14588 29934 14590 29986
rect 14642 29934 14644 29986
rect 14588 29652 14644 29934
rect 14588 28196 14644 29596
rect 14588 28130 14644 28140
rect 14700 29986 14756 29998
rect 14700 29934 14702 29986
rect 14754 29934 14756 29986
rect 14700 27860 14756 29934
rect 14924 29988 14980 30026
rect 14924 29922 14980 29932
rect 14820 29820 15084 29830
rect 14876 29764 14924 29820
rect 14980 29764 15028 29820
rect 14820 29754 15084 29764
rect 14812 29652 14868 29662
rect 14812 29316 14868 29596
rect 14812 29250 14868 29260
rect 15148 29204 15204 30046
rect 15372 30100 15428 30110
rect 15036 28868 15092 28878
rect 14812 28756 14868 28766
rect 14812 28662 14868 28700
rect 14924 28644 14980 28654
rect 14924 28550 14980 28588
rect 15036 28420 15092 28812
rect 15148 28642 15204 29148
rect 15260 29988 15316 29998
rect 15260 28756 15316 29932
rect 15260 28690 15316 28700
rect 15148 28590 15150 28642
rect 15202 28590 15204 28642
rect 15148 28578 15204 28590
rect 15036 28364 15204 28420
rect 14820 28252 15084 28262
rect 14876 28196 14924 28252
rect 14980 28196 15028 28252
rect 14820 28186 15084 28196
rect 14924 27860 14980 27898
rect 14700 27804 14924 27860
rect 14924 27794 14980 27804
rect 15036 27748 15092 27758
rect 15148 27748 15204 28364
rect 15092 27692 15204 27748
rect 15036 27682 15092 27692
rect 14924 27634 14980 27646
rect 14924 27582 14926 27634
rect 14978 27582 14980 27634
rect 14924 26908 14980 27582
rect 15148 27076 15204 27692
rect 15260 28084 15316 28094
rect 15260 27748 15316 28028
rect 15260 27654 15316 27692
rect 15260 27076 15316 27086
rect 15148 27020 15260 27076
rect 14700 26852 14980 26908
rect 14588 26068 14644 26078
rect 14700 26068 14756 26852
rect 14820 26684 15084 26694
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 14820 26618 15084 26628
rect 15260 26516 15316 27020
rect 14812 26514 15316 26516
rect 14812 26462 15262 26514
rect 15314 26462 15316 26514
rect 14812 26460 15316 26462
rect 14812 26290 14868 26460
rect 15260 26450 15316 26460
rect 14812 26238 14814 26290
rect 14866 26238 14868 26290
rect 14812 26226 14868 26238
rect 15372 26292 15428 30044
rect 15372 26226 15428 26236
rect 14588 26066 14756 26068
rect 14588 26014 14590 26066
rect 14642 26014 14756 26066
rect 14588 26012 14756 26014
rect 15148 26068 15204 26078
rect 14588 26002 14644 26012
rect 14476 25342 14478 25394
rect 14530 25342 14532 25394
rect 14364 25284 14420 25294
rect 14476 25284 14532 25342
rect 14924 25284 14980 25294
rect 14476 25282 14980 25284
rect 14476 25230 14926 25282
rect 14978 25230 14980 25282
rect 14476 25228 14980 25230
rect 14364 25190 14420 25228
rect 14252 24894 14254 24946
rect 14306 24894 14308 24946
rect 14252 24498 14308 24894
rect 14700 24612 14756 25228
rect 14924 25218 14980 25228
rect 14820 25116 15084 25126
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 14820 25050 15084 25060
rect 15148 24946 15204 26012
rect 15148 24894 15150 24946
rect 15202 24894 15204 24946
rect 15148 24612 15204 24894
rect 14700 24610 14868 24612
rect 14700 24558 14702 24610
rect 14754 24558 14868 24610
rect 14700 24556 14868 24558
rect 14700 24546 14756 24556
rect 14252 24446 14254 24498
rect 14306 24446 14308 24498
rect 14252 24434 14308 24446
rect 13916 24164 13972 24174
rect 13692 23938 13748 23950
rect 13692 23886 13694 23938
rect 13746 23886 13748 23938
rect 13692 23828 13748 23886
rect 13692 23762 13748 23772
rect 13580 23102 13582 23154
rect 13634 23102 13636 23154
rect 13580 22484 13636 23102
rect 13356 21812 13412 21822
rect 13132 21810 13412 21812
rect 13132 21758 13358 21810
rect 13410 21758 13412 21810
rect 13132 21756 13412 21758
rect 12908 20916 12964 20926
rect 12908 20822 12964 20860
rect 13132 20804 13188 21756
rect 13356 21746 13412 21756
rect 13580 21812 13636 22428
rect 13692 23044 13748 23054
rect 13692 22482 13748 22988
rect 13692 22430 13694 22482
rect 13746 22430 13748 22482
rect 13692 22418 13748 22430
rect 13580 21746 13636 21756
rect 13132 20738 13188 20748
rect 13468 20690 13524 20702
rect 13468 20638 13470 20690
rect 13522 20638 13524 20690
rect 13468 20580 13524 20638
rect 13692 20692 13748 20702
rect 13692 20598 13748 20636
rect 13468 20514 13524 20524
rect 13580 20578 13636 20590
rect 13580 20526 13582 20578
rect 13634 20526 13636 20578
rect 13580 20356 13636 20526
rect 13020 20300 13636 20356
rect 12908 20132 12964 20142
rect 12908 19348 12964 20076
rect 13020 20130 13076 20300
rect 13020 20078 13022 20130
rect 13074 20078 13076 20130
rect 13020 20066 13076 20078
rect 13916 20132 13972 24108
rect 14476 24164 14532 24174
rect 14028 24052 14084 24062
rect 14028 23958 14084 23996
rect 14476 23938 14532 24108
rect 14476 23886 14478 23938
rect 14530 23886 14532 23938
rect 14476 23874 14532 23886
rect 14812 23828 14868 24556
rect 15148 24546 15204 24556
rect 15372 25732 15428 25742
rect 15372 25282 15428 25676
rect 15372 25230 15374 25282
rect 15426 25230 15428 25282
rect 14924 24498 14980 24510
rect 14924 24446 14926 24498
rect 14978 24446 14980 24498
rect 14924 23938 14980 24446
rect 15372 24164 15428 25230
rect 15372 24098 15428 24108
rect 14924 23886 14926 23938
rect 14978 23886 14980 23938
rect 14924 23874 14980 23886
rect 14812 23762 14868 23772
rect 15148 23828 15204 23838
rect 15148 23826 15316 23828
rect 15148 23774 15150 23826
rect 15202 23774 15316 23826
rect 15148 23772 15316 23774
rect 15148 23762 15204 23772
rect 14700 23714 14756 23726
rect 14700 23662 14702 23714
rect 14754 23662 14756 23714
rect 14700 23380 14756 23662
rect 14820 23548 15084 23558
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 14820 23482 15084 23492
rect 14252 23324 14756 23380
rect 15148 23380 15204 23390
rect 14252 23266 14308 23324
rect 14252 23214 14254 23266
rect 14306 23214 14308 23266
rect 14252 23202 14308 23214
rect 14476 23156 14532 23166
rect 14532 23100 14644 23156
rect 14476 23090 14532 23100
rect 14476 21700 14532 21710
rect 14476 21606 14532 21644
rect 14252 21476 14308 21486
rect 14252 21382 14308 21420
rect 14364 21474 14420 21486
rect 14364 21422 14366 21474
rect 14418 21422 14420 21474
rect 14364 21140 14420 21422
rect 14028 21084 14420 21140
rect 14028 21026 14084 21084
rect 14028 20974 14030 21026
rect 14082 20974 14084 21026
rect 14028 20962 14084 20974
rect 14252 20916 14308 20926
rect 14252 20802 14308 20860
rect 14252 20750 14254 20802
rect 14306 20750 14308 20802
rect 14252 20738 14308 20750
rect 14588 20132 14644 23100
rect 14700 22484 14756 22494
rect 14700 21028 14756 22428
rect 15148 22148 15204 23324
rect 15260 22820 15316 23772
rect 15484 22932 15540 30828
rect 15708 30324 15764 30942
rect 15708 30258 15764 30268
rect 15596 30212 15652 30222
rect 15596 30118 15652 30156
rect 15932 29764 15988 31166
rect 16044 31556 16100 31566
rect 16044 31218 16100 31500
rect 16044 31166 16046 31218
rect 16098 31166 16100 31218
rect 16044 31154 16100 31166
rect 16268 31444 16324 31454
rect 16268 30210 16324 31388
rect 16268 30158 16270 30210
rect 16322 30158 16324 30210
rect 16268 30146 16324 30158
rect 16380 30212 16436 32396
rect 16716 31666 16772 31678
rect 16716 31614 16718 31666
rect 16770 31614 16772 31666
rect 16492 31220 16548 31230
rect 16492 31126 16548 31164
rect 16380 30146 16436 30156
rect 16716 30100 16772 31614
rect 16828 30884 16884 32396
rect 16940 31218 16996 33516
rect 16940 31166 16942 31218
rect 16994 31166 16996 31218
rect 16940 30996 16996 31166
rect 16940 30930 16996 30940
rect 16828 30818 16884 30828
rect 16716 30034 16772 30044
rect 15820 29708 16212 29764
rect 15708 29316 15764 29326
rect 15596 29314 15764 29316
rect 15596 29262 15710 29314
rect 15762 29262 15764 29314
rect 15596 29260 15764 29262
rect 15596 29204 15652 29260
rect 15708 29250 15764 29260
rect 15596 29138 15652 29148
rect 15708 28756 15764 28766
rect 15708 28662 15764 28700
rect 15708 28532 15764 28542
rect 15708 28082 15764 28476
rect 15708 28030 15710 28082
rect 15762 28030 15764 28082
rect 15596 27412 15652 27422
rect 15596 24948 15652 27356
rect 15708 26514 15764 28030
rect 15708 26462 15710 26514
rect 15762 26462 15764 26514
rect 15708 26404 15764 26462
rect 15708 26338 15764 26348
rect 15820 26066 15876 29708
rect 16156 29650 16212 29708
rect 16156 29598 16158 29650
rect 16210 29598 16212 29650
rect 16156 29586 16212 29598
rect 16604 29316 16660 29326
rect 16604 29314 16772 29316
rect 16604 29262 16606 29314
rect 16658 29262 16772 29314
rect 16604 29260 16772 29262
rect 16604 29250 16660 29260
rect 16044 28644 16100 28654
rect 16044 28550 16100 28588
rect 16380 27860 16436 27870
rect 16156 27748 16212 27758
rect 16156 27654 16212 27692
rect 16380 27186 16436 27804
rect 16380 27134 16382 27186
rect 16434 27134 16436 27186
rect 16380 27122 16436 27134
rect 16716 27188 16772 29260
rect 16940 28642 16996 28654
rect 16940 28590 16942 28642
rect 16994 28590 16996 28642
rect 16940 27972 16996 28590
rect 16940 27906 16996 27916
rect 17052 28084 17108 33628
rect 16940 27748 16996 27758
rect 17052 27748 17108 28028
rect 16940 27746 17108 27748
rect 16940 27694 16942 27746
rect 16994 27694 17108 27746
rect 16940 27692 17108 27694
rect 16940 27682 16996 27692
rect 16828 27188 16884 27198
rect 16772 27186 16884 27188
rect 16772 27134 16830 27186
rect 16882 27134 16884 27186
rect 16772 27132 16884 27134
rect 16716 27094 16772 27132
rect 16828 27122 16884 27132
rect 17164 26908 17220 35252
rect 17276 31778 17332 35868
rect 17388 35700 17444 35710
rect 17388 35606 17444 35644
rect 17500 32788 17556 36092
rect 17612 34804 17668 34814
rect 17612 33684 17668 34748
rect 17612 33618 17668 33628
rect 17500 32722 17556 32732
rect 17724 32788 17780 36764
rect 18620 36706 18676 39342
rect 18844 38946 18900 40236
rect 18844 38894 18846 38946
rect 18898 38894 18900 38946
rect 18844 38882 18900 38894
rect 18620 36654 18622 36706
rect 18674 36654 18676 36706
rect 18620 36642 18676 36654
rect 18732 38834 18788 38846
rect 18732 38782 18734 38834
rect 18786 38782 18788 38834
rect 18396 36596 18452 36606
rect 18396 36502 18452 36540
rect 18732 36484 18788 38782
rect 18844 37716 18900 37726
rect 18956 37716 19012 46846
rect 19068 42980 19124 49644
rect 19292 48916 19348 48926
rect 19292 48132 19348 48860
rect 19180 47684 19236 47694
rect 19180 46564 19236 47628
rect 19180 46470 19236 46508
rect 19292 45778 19348 48076
rect 19292 45726 19294 45778
rect 19346 45726 19348 45778
rect 19292 45714 19348 45726
rect 19180 44212 19236 44222
rect 19180 43762 19236 44156
rect 19404 43876 19460 50092
rect 19516 50036 19572 50046
rect 19516 49812 19572 49980
rect 19964 49924 20020 51100
rect 20188 50818 20244 51326
rect 20188 50766 20190 50818
rect 20242 50766 20244 50818
rect 20188 50754 20244 50766
rect 20412 52836 20468 52846
rect 20076 50372 20132 50382
rect 20132 50316 20244 50372
rect 20076 50278 20132 50316
rect 19516 49718 19572 49756
rect 19628 49922 20020 49924
rect 19628 49870 19966 49922
rect 20018 49870 20020 49922
rect 19628 49868 20020 49870
rect 19516 48244 19572 48254
rect 19628 48244 19684 49868
rect 19964 49858 20020 49868
rect 19740 49700 19796 49710
rect 19740 49698 19908 49700
rect 19740 49646 19742 49698
rect 19794 49646 19908 49698
rect 19740 49644 19908 49646
rect 19740 49634 19796 49644
rect 19516 48242 19684 48244
rect 19516 48190 19518 48242
rect 19570 48190 19684 48242
rect 19516 48188 19684 48190
rect 19740 48692 19796 48702
rect 19516 47570 19572 48188
rect 19516 47518 19518 47570
rect 19570 47518 19572 47570
rect 19516 47460 19572 47518
rect 19516 47394 19572 47404
rect 19740 47908 19796 48636
rect 19740 47124 19796 47852
rect 19740 47058 19796 47068
rect 19516 46564 19572 46574
rect 19516 44210 19572 46508
rect 19628 45668 19684 45678
rect 19628 44322 19684 45612
rect 19628 44270 19630 44322
rect 19682 44270 19684 44322
rect 19628 44258 19684 44270
rect 19740 45444 19796 45454
rect 19516 44158 19518 44210
rect 19570 44158 19572 44210
rect 19516 44146 19572 44158
rect 19404 43820 19684 43876
rect 19180 43710 19182 43762
rect 19234 43710 19236 43762
rect 19180 43698 19236 43710
rect 19404 43652 19460 43662
rect 19404 43558 19460 43596
rect 19292 43540 19348 43550
rect 19292 43446 19348 43484
rect 19292 42980 19348 42990
rect 19068 42978 19348 42980
rect 19068 42926 19294 42978
rect 19346 42926 19348 42978
rect 19068 42924 19348 42926
rect 19292 42914 19348 42924
rect 19516 42756 19572 42766
rect 19292 42754 19572 42756
rect 19292 42702 19518 42754
rect 19570 42702 19572 42754
rect 19292 42700 19572 42702
rect 19180 42532 19236 42542
rect 19180 42194 19236 42476
rect 19180 42142 19182 42194
rect 19234 42142 19236 42194
rect 19180 42130 19236 42142
rect 19292 42082 19348 42700
rect 19516 42690 19572 42700
rect 19628 42196 19684 43820
rect 19516 42140 19684 42196
rect 19740 43538 19796 45388
rect 19740 43486 19742 43538
rect 19794 43486 19796 43538
rect 19292 42030 19294 42082
rect 19346 42030 19348 42082
rect 19292 42018 19348 42030
rect 19404 42084 19460 42094
rect 19404 41990 19460 42028
rect 19068 41972 19124 41982
rect 19068 41878 19124 41916
rect 19516 41636 19572 42140
rect 19292 41580 19572 41636
rect 19628 41970 19684 41982
rect 19628 41918 19630 41970
rect 19682 41918 19684 41970
rect 18900 37660 19012 37716
rect 19068 38722 19124 38734
rect 19068 38670 19070 38722
rect 19122 38670 19124 38722
rect 18844 37490 18900 37660
rect 18844 37438 18846 37490
rect 18898 37438 18900 37490
rect 18844 37426 18900 37438
rect 19068 37490 19124 38670
rect 19068 37438 19070 37490
rect 19122 37438 19124 37490
rect 19068 37426 19124 37438
rect 18956 37266 19012 37278
rect 18956 37214 18958 37266
rect 19010 37214 19012 37266
rect 18844 37156 18900 37166
rect 18844 36484 18900 37100
rect 18956 37044 19012 37214
rect 18956 36978 19012 36988
rect 19180 37266 19236 37278
rect 19180 37214 19182 37266
rect 19234 37214 19236 37266
rect 19180 36820 19236 37214
rect 19180 36754 19236 36764
rect 18956 36484 19012 36494
rect 18844 36482 19012 36484
rect 18844 36430 18958 36482
rect 19010 36430 19012 36482
rect 18844 36428 19012 36430
rect 18732 36418 18788 36428
rect 18732 36260 18788 36270
rect 18732 36258 18900 36260
rect 18732 36206 18734 36258
rect 18786 36206 18900 36258
rect 18732 36204 18900 36206
rect 18732 36194 18788 36204
rect 18172 35588 18228 35598
rect 18060 35586 18228 35588
rect 18060 35534 18174 35586
rect 18226 35534 18228 35586
rect 18060 35532 18228 35534
rect 17836 35476 17892 35486
rect 17836 34692 17892 35420
rect 18060 35026 18116 35532
rect 18172 35522 18228 35532
rect 18222 35308 18486 35318
rect 18278 35252 18326 35308
rect 18382 35252 18430 35308
rect 18222 35242 18486 35252
rect 18732 35308 18788 35318
rect 18060 34974 18062 35026
rect 18114 34974 18116 35026
rect 18060 34962 18116 34974
rect 18620 35138 18676 35150
rect 18620 35086 18622 35138
rect 18674 35086 18676 35138
rect 17948 34916 18004 34926
rect 17948 34822 18004 34860
rect 18172 34914 18228 34926
rect 18172 34862 18174 34914
rect 18226 34862 18228 34914
rect 18172 34804 18228 34862
rect 18508 34916 18564 34926
rect 18620 34916 18676 35086
rect 18508 34914 18676 34916
rect 18508 34862 18510 34914
rect 18562 34862 18676 34914
rect 18508 34860 18676 34862
rect 18508 34850 18564 34860
rect 18172 34738 18228 34748
rect 18620 34692 18676 34702
rect 17836 34636 18004 34692
rect 17724 32722 17780 32732
rect 17388 32676 17444 32686
rect 17388 32582 17444 32620
rect 17724 32562 17780 32574
rect 17724 32510 17726 32562
rect 17778 32510 17780 32562
rect 17276 31726 17278 31778
rect 17330 31726 17332 31778
rect 17276 31220 17332 31726
rect 17500 32450 17556 32462
rect 17500 32398 17502 32450
rect 17554 32398 17556 32450
rect 17500 31444 17556 32398
rect 17724 32452 17780 32510
rect 17724 32386 17780 32396
rect 17836 32562 17892 32574
rect 17836 32510 17838 32562
rect 17890 32510 17892 32562
rect 17500 31378 17556 31388
rect 17836 31220 17892 32510
rect 17276 31154 17332 31164
rect 17724 31164 17892 31220
rect 17948 31218 18004 34636
rect 18620 34354 18676 34636
rect 18620 34302 18622 34354
rect 18674 34302 18676 34354
rect 18620 34290 18676 34302
rect 18060 34020 18116 34030
rect 18060 33926 18116 33964
rect 18222 33740 18486 33750
rect 18278 33684 18326 33740
rect 18382 33684 18430 33740
rect 18222 33674 18486 33684
rect 18060 33572 18116 33582
rect 18060 33458 18116 33516
rect 18060 33406 18062 33458
rect 18114 33406 18116 33458
rect 18060 32564 18116 33406
rect 18508 33122 18564 33134
rect 18508 33070 18510 33122
rect 18562 33070 18564 33122
rect 18508 32788 18564 33070
rect 18508 32722 18564 32732
rect 18732 32786 18788 35252
rect 18732 32734 18734 32786
rect 18786 32734 18788 32786
rect 18732 32722 18788 32734
rect 18844 32788 18900 36204
rect 18956 35364 19012 36428
rect 18956 35298 19012 35308
rect 19068 36258 19124 36270
rect 19068 36206 19070 36258
rect 19122 36206 19124 36258
rect 18956 35140 19012 35150
rect 19068 35140 19124 36206
rect 19180 36258 19236 36270
rect 19180 36206 19182 36258
rect 19234 36206 19236 36258
rect 19180 35588 19236 36206
rect 19180 35522 19236 35532
rect 18956 35138 19124 35140
rect 18956 35086 18958 35138
rect 19010 35086 19124 35138
rect 18956 35084 19124 35086
rect 19180 35140 19236 35150
rect 18956 35074 19012 35084
rect 19180 35046 19236 35084
rect 18844 32722 18900 32732
rect 18956 34916 19012 34926
rect 18956 34690 19012 34860
rect 18956 34638 18958 34690
rect 19010 34638 19012 34690
rect 18060 32498 18116 32508
rect 18396 32562 18452 32574
rect 18396 32510 18398 32562
rect 18450 32510 18452 32562
rect 18396 32452 18452 32510
rect 18396 32340 18452 32396
rect 18060 32284 18452 32340
rect 18620 32562 18676 32574
rect 18620 32510 18622 32562
rect 18674 32510 18676 32562
rect 18060 32004 18116 32284
rect 18222 32172 18486 32182
rect 18278 32116 18326 32172
rect 18382 32116 18430 32172
rect 18222 32106 18486 32116
rect 18060 31948 18228 32004
rect 17948 31166 17950 31218
rect 18002 31166 18004 31218
rect 17388 31108 17444 31118
rect 17388 29988 17444 31052
rect 17388 29922 17444 29932
rect 17612 30994 17668 31006
rect 17612 30942 17614 30994
rect 17666 30942 17668 30994
rect 17612 30324 17668 30942
rect 17724 30436 17780 31164
rect 17948 31154 18004 31166
rect 18172 31108 18228 31948
rect 18172 31014 18228 31052
rect 17836 30996 17892 31006
rect 17836 30902 17892 30940
rect 18060 30994 18116 31006
rect 18060 30942 18062 30994
rect 18114 30942 18116 30994
rect 17724 30380 17892 30436
rect 17612 29652 17668 30268
rect 17724 29652 17780 29662
rect 17612 29650 17780 29652
rect 17612 29598 17726 29650
rect 17778 29598 17780 29650
rect 17612 29596 17780 29598
rect 17724 29586 17780 29596
rect 17836 29650 17892 30380
rect 17836 29598 17838 29650
rect 17890 29598 17892 29650
rect 17836 29586 17892 29598
rect 17388 29426 17444 29438
rect 17948 29428 18004 29438
rect 17388 29374 17390 29426
rect 17442 29374 17444 29426
rect 17388 27636 17444 29374
rect 17836 29426 18004 29428
rect 17836 29374 17950 29426
rect 18002 29374 18004 29426
rect 17836 29372 18004 29374
rect 17836 29316 17892 29372
rect 17948 29362 18004 29372
rect 17612 28532 17668 28542
rect 17612 28530 17780 28532
rect 17612 28478 17614 28530
rect 17666 28478 17780 28530
rect 17612 28476 17780 28478
rect 17612 28466 17668 28476
rect 17724 28082 17780 28476
rect 17836 28420 17892 29260
rect 17836 28354 17892 28364
rect 17724 28030 17726 28082
rect 17778 28030 17780 28082
rect 17724 28018 17780 28030
rect 17836 28084 17892 28094
rect 17836 27970 17892 28028
rect 18060 27972 18116 30942
rect 18620 30996 18676 32510
rect 18844 32564 18900 32574
rect 18844 32470 18900 32508
rect 18620 30930 18676 30940
rect 18732 32004 18788 32014
rect 18732 31106 18788 31948
rect 18732 31054 18734 31106
rect 18786 31054 18788 31106
rect 18222 30604 18486 30614
rect 18278 30548 18326 30604
rect 18382 30548 18430 30604
rect 18222 30538 18486 30548
rect 18396 30324 18452 30334
rect 18396 30230 18452 30268
rect 18732 30212 18788 31054
rect 18844 31106 18900 31118
rect 18844 31054 18846 31106
rect 18898 31054 18900 31106
rect 18844 30434 18900 31054
rect 18956 31108 19012 34638
rect 19068 34356 19124 34366
rect 19068 34262 19124 34300
rect 19068 33236 19124 33246
rect 19068 33142 19124 33180
rect 19068 32562 19124 32574
rect 19068 32510 19070 32562
rect 19122 32510 19124 32562
rect 19068 32228 19124 32510
rect 19068 32162 19124 32172
rect 19180 32002 19236 32014
rect 19180 31950 19182 32002
rect 19234 31950 19236 32002
rect 19068 31780 19124 31790
rect 19068 31218 19124 31724
rect 19180 31332 19236 31950
rect 19292 31948 19348 41580
rect 19404 41412 19460 41422
rect 19404 41186 19460 41356
rect 19516 41300 19572 41310
rect 19516 41206 19572 41244
rect 19404 41134 19406 41186
rect 19458 41134 19460 41186
rect 19404 41122 19460 41134
rect 19628 40962 19684 41918
rect 19628 40910 19630 40962
rect 19682 40910 19684 40962
rect 19404 40852 19460 40862
rect 19404 39842 19460 40796
rect 19628 40292 19684 40910
rect 19740 40964 19796 43486
rect 19740 40898 19796 40908
rect 19852 40740 19908 49644
rect 20076 49028 20132 49038
rect 19964 48130 20020 48142
rect 19964 48078 19966 48130
rect 20018 48078 20020 48130
rect 19964 44436 20020 48078
rect 20076 47570 20132 48972
rect 20188 48916 20244 50316
rect 20188 48850 20244 48860
rect 20076 47518 20078 47570
rect 20130 47518 20132 47570
rect 20076 47506 20132 47518
rect 20300 47346 20356 47358
rect 20300 47294 20302 47346
rect 20354 47294 20356 47346
rect 20188 47236 20244 47246
rect 19964 44380 20132 44436
rect 19964 44210 20020 44222
rect 19964 44158 19966 44210
rect 20018 44158 20020 44210
rect 19964 43314 20020 44158
rect 19964 43262 19966 43314
rect 20018 43262 20020 43314
rect 19964 43250 20020 43262
rect 20076 42980 20132 44380
rect 20188 44324 20244 47180
rect 20300 47124 20356 47294
rect 20300 47058 20356 47068
rect 20412 47068 20468 52780
rect 20748 52386 20804 54012
rect 20860 53956 20916 53966
rect 20860 53060 20916 53900
rect 20860 52994 20916 53004
rect 20748 52334 20750 52386
rect 20802 52334 20804 52386
rect 20748 52322 20804 52334
rect 21084 52946 21140 52958
rect 21084 52894 21086 52946
rect 21138 52894 21140 52946
rect 20524 52164 20580 52174
rect 20524 52070 20580 52108
rect 20748 52052 20804 52062
rect 20748 51492 20804 51996
rect 20860 51492 20916 51502
rect 20748 51490 20916 51492
rect 20748 51438 20862 51490
rect 20914 51438 20916 51490
rect 20748 51436 20916 51438
rect 20860 51426 20916 51436
rect 20748 50818 20804 50830
rect 20748 50766 20750 50818
rect 20802 50766 20804 50818
rect 20524 50370 20580 50382
rect 20524 50318 20526 50370
rect 20578 50318 20580 50370
rect 20524 49924 20580 50318
rect 20524 49858 20580 49868
rect 20636 49140 20692 49150
rect 20636 48914 20692 49084
rect 20636 48862 20638 48914
rect 20690 48862 20692 48914
rect 20524 48356 20580 48366
rect 20636 48356 20692 48862
rect 20524 48354 20692 48356
rect 20524 48302 20526 48354
rect 20578 48302 20692 48354
rect 20524 48300 20692 48302
rect 20524 47796 20580 48300
rect 20524 47730 20580 47740
rect 20524 47572 20580 47582
rect 20580 47516 20692 47572
rect 20524 47506 20580 47516
rect 20524 47236 20580 47246
rect 20636 47236 20692 47516
rect 20748 47460 20804 50766
rect 21084 50484 21140 52894
rect 21196 52052 21252 54236
rect 21308 53170 21364 55020
rect 21308 53118 21310 53170
rect 21362 53118 21364 53170
rect 21308 53106 21364 53118
rect 21308 52836 21364 52846
rect 21420 52836 21476 55132
rect 21644 55094 21700 55132
rect 22204 55076 22260 55086
rect 22204 54982 22260 55020
rect 22428 55074 22484 55916
rect 22428 55022 22430 55074
rect 22482 55022 22484 55074
rect 21624 54908 21888 54918
rect 21680 54852 21728 54908
rect 21784 54852 21832 54908
rect 21624 54842 21888 54852
rect 22428 54740 22484 55022
rect 21756 54684 22484 54740
rect 21644 54628 21700 54638
rect 21532 54572 21644 54628
rect 21532 54290 21588 54572
rect 21644 54562 21700 54572
rect 21532 54238 21534 54290
rect 21586 54238 21588 54290
rect 21532 53730 21588 54238
rect 21532 53678 21534 53730
rect 21586 53678 21588 53730
rect 21532 53666 21588 53678
rect 21644 53842 21700 53854
rect 21644 53790 21646 53842
rect 21698 53790 21700 53842
rect 21644 53620 21700 53790
rect 21756 53730 21812 54684
rect 21980 54402 22036 54414
rect 21980 54350 21982 54402
rect 22034 54350 22036 54402
rect 21980 54180 22036 54350
rect 22428 54404 22484 54414
rect 22428 54310 22484 54348
rect 21980 54114 22036 54124
rect 22540 53956 22596 56028
rect 22652 55076 22708 56140
rect 22764 55970 22820 55982
rect 22764 55918 22766 55970
rect 22818 55918 22820 55970
rect 22764 55412 22820 55918
rect 22764 55346 22820 55356
rect 22876 55298 22932 55310
rect 22876 55246 22878 55298
rect 22930 55246 22932 55298
rect 22876 55188 22932 55246
rect 22876 55122 22932 55132
rect 22652 55020 22820 55076
rect 21756 53678 21758 53730
rect 21810 53678 21812 53730
rect 21756 53666 21812 53678
rect 22316 53900 22596 53956
rect 22652 54852 22708 54862
rect 22204 53620 22260 53630
rect 21644 53554 21700 53564
rect 22092 53564 22204 53620
rect 21980 53508 22036 53518
rect 21980 53414 22036 53452
rect 21624 53340 21888 53350
rect 21680 53284 21728 53340
rect 21784 53284 21832 53340
rect 21624 53274 21888 53284
rect 21644 53060 21700 53070
rect 21364 52780 21476 52836
rect 21532 53004 21644 53060
rect 21308 52770 21364 52780
rect 21532 52162 21588 53004
rect 21644 52994 21700 53004
rect 21756 52836 21812 52846
rect 22092 52836 22148 53564
rect 22204 53526 22260 53564
rect 22316 53396 22372 53900
rect 22652 53508 22708 54796
rect 22764 54740 22820 55020
rect 23100 54852 23156 60396
rect 23212 57876 23268 62188
rect 23324 61572 23380 61582
rect 23324 58828 23380 61516
rect 23436 59444 23492 62860
rect 23548 62244 23604 63870
rect 23772 63924 23828 63934
rect 23660 63810 23716 63822
rect 23660 63758 23662 63810
rect 23714 63758 23716 63810
rect 23660 63028 23716 63758
rect 23660 62962 23716 62972
rect 23548 62178 23604 62188
rect 23772 60228 23828 63868
rect 23772 60162 23828 60172
rect 23436 59378 23492 59388
rect 23660 60116 23716 60126
rect 23660 59442 23716 60060
rect 23772 59892 23828 59902
rect 23772 59798 23828 59836
rect 23660 59390 23662 59442
rect 23714 59390 23716 59442
rect 23660 59378 23716 59390
rect 23436 59218 23492 59230
rect 23436 59166 23438 59218
rect 23490 59166 23492 59218
rect 23436 59108 23492 59166
rect 23548 59220 23604 59230
rect 23548 59126 23604 59164
rect 23436 59042 23492 59052
rect 23324 58772 23492 58828
rect 23324 58658 23380 58670
rect 23324 58606 23326 58658
rect 23378 58606 23380 58658
rect 23324 58546 23380 58606
rect 23324 58494 23326 58546
rect 23378 58494 23380 58546
rect 23324 58482 23380 58494
rect 23436 57988 23492 58772
rect 23772 58548 23828 58558
rect 23772 58454 23828 58492
rect 23884 57988 23940 70030
rect 24332 70812 24500 70868
rect 24220 68740 24276 68750
rect 24220 68516 24276 68684
rect 23996 68514 24276 68516
rect 23996 68462 24222 68514
rect 24274 68462 24276 68514
rect 23996 68460 24276 68462
rect 23996 67058 24052 68460
rect 24220 68450 24276 68460
rect 24220 67956 24276 67966
rect 23996 67006 23998 67058
rect 24050 67006 24052 67058
rect 23996 65828 24052 67006
rect 23996 65762 24052 65772
rect 24108 67954 24276 67956
rect 24108 67902 24222 67954
rect 24274 67902 24276 67954
rect 24108 67900 24276 67902
rect 23996 65492 24052 65502
rect 23996 63698 24052 65436
rect 24108 63812 24164 67900
rect 24220 67890 24276 67900
rect 24332 66948 24388 70812
rect 24780 70756 24836 70766
rect 24780 70662 24836 70700
rect 24444 68516 24500 68526
rect 24444 67732 24500 68460
rect 24444 67170 24500 67676
rect 24444 67118 24446 67170
rect 24498 67118 24500 67170
rect 24444 67106 24500 67118
rect 24556 68404 24612 68414
rect 24556 67170 24612 68348
rect 24556 67118 24558 67170
rect 24610 67118 24612 67170
rect 24556 67106 24612 67118
rect 24668 67172 24724 67182
rect 24668 67078 24724 67116
rect 24332 66892 24612 66948
rect 24444 65492 24500 65530
rect 24444 65426 24500 65436
rect 24444 65268 24500 65278
rect 24220 64820 24276 64830
rect 24220 64726 24276 64764
rect 24220 63924 24276 63934
rect 24220 63830 24276 63868
rect 24108 63746 24164 63756
rect 23996 63646 23998 63698
rect 24050 63646 24052 63698
rect 23996 63250 24052 63646
rect 23996 63198 23998 63250
rect 24050 63198 24052 63250
rect 23996 63186 24052 63198
rect 24332 63028 24388 63038
rect 24220 62244 24276 62282
rect 24220 62178 24276 62188
rect 24108 61684 24164 61694
rect 23996 61570 24052 61582
rect 23996 61518 23998 61570
rect 24050 61518 24052 61570
rect 23996 61460 24052 61518
rect 23996 61394 24052 61404
rect 23436 57922 23492 57932
rect 23548 57932 23940 57988
rect 23996 59218 24052 59230
rect 23996 59166 23998 59218
rect 24050 59166 24052 59218
rect 23212 57820 23380 57876
rect 23212 57650 23268 57662
rect 23212 57598 23214 57650
rect 23266 57598 23268 57650
rect 23212 57540 23268 57598
rect 23212 57204 23268 57484
rect 23212 57138 23268 57148
rect 23324 56308 23380 57820
rect 23436 57652 23492 57662
rect 23436 57558 23492 57596
rect 23436 56308 23492 56318
rect 23324 56306 23492 56308
rect 23324 56254 23438 56306
rect 23490 56254 23492 56306
rect 23324 56252 23492 56254
rect 23436 56242 23492 56252
rect 23324 56082 23380 56094
rect 23324 56030 23326 56082
rect 23378 56030 23380 56082
rect 23324 55748 23380 56030
rect 23436 56084 23492 56094
rect 23436 55970 23492 56028
rect 23436 55918 23438 55970
rect 23490 55918 23492 55970
rect 23436 55906 23492 55918
rect 23324 55692 23492 55748
rect 23212 55412 23268 55422
rect 23212 55318 23268 55356
rect 23100 54786 23156 54796
rect 22876 54740 22932 54750
rect 22764 54738 22932 54740
rect 22764 54686 22878 54738
rect 22930 54686 22932 54738
rect 22764 54684 22932 54686
rect 22876 54674 22932 54684
rect 23436 54740 23492 55692
rect 23436 54674 23492 54684
rect 23324 54404 23380 54414
rect 23212 54402 23380 54404
rect 23212 54350 23326 54402
rect 23378 54350 23380 54402
rect 23212 54348 23380 54350
rect 21756 52834 22148 52836
rect 21756 52782 21758 52834
rect 21810 52782 22148 52834
rect 21756 52780 22148 52782
rect 22204 53340 22372 53396
rect 22428 53452 22708 53508
rect 22764 54290 22820 54302
rect 22764 54238 22766 54290
rect 22818 54238 22820 54290
rect 22764 53618 22820 54238
rect 22764 53566 22766 53618
rect 22818 53566 22820 53618
rect 21756 52770 21812 52780
rect 21868 52388 21924 52398
rect 21868 52386 22036 52388
rect 21868 52334 21870 52386
rect 21922 52334 22036 52386
rect 21868 52332 22036 52334
rect 21868 52322 21924 52332
rect 21532 52110 21534 52162
rect 21586 52110 21588 52162
rect 21532 52098 21588 52110
rect 21868 52162 21924 52174
rect 21868 52110 21870 52162
rect 21922 52110 21924 52162
rect 21308 52052 21364 52062
rect 21196 52050 21364 52052
rect 21196 51998 21310 52050
rect 21362 51998 21364 52050
rect 21196 51996 21364 51998
rect 21308 50932 21364 51996
rect 21644 52052 21700 52062
rect 21644 51938 21700 51996
rect 21868 52052 21924 52110
rect 21868 51986 21924 51996
rect 21644 51886 21646 51938
rect 21698 51886 21700 51938
rect 21644 51874 21700 51886
rect 21624 51772 21888 51782
rect 21680 51716 21728 51772
rect 21784 51716 21832 51772
rect 21624 51706 21888 51716
rect 21980 51716 22036 52332
rect 21980 51650 22036 51660
rect 21308 50866 21364 50876
rect 21420 50594 21476 50606
rect 21420 50542 21422 50594
rect 21474 50542 21476 50594
rect 21084 50428 21364 50484
rect 20972 50036 21028 50046
rect 20860 47908 20916 47918
rect 20972 47908 21028 49980
rect 20916 47852 21028 47908
rect 20860 47842 20916 47852
rect 20860 47684 20916 47694
rect 20972 47684 21028 47852
rect 20972 47628 21140 47684
rect 20860 47590 20916 47628
rect 20748 47404 21028 47460
rect 20748 47236 20804 47246
rect 20636 47234 20804 47236
rect 20636 47182 20750 47234
rect 20802 47182 20804 47234
rect 20636 47180 20804 47182
rect 20524 47142 20580 47180
rect 20748 47124 20804 47180
rect 20412 47012 20692 47068
rect 20748 47012 20916 47068
rect 20300 46676 20356 46686
rect 20300 46582 20356 46620
rect 20524 46674 20580 46686
rect 20524 46622 20526 46674
rect 20578 46622 20580 46674
rect 20412 46562 20468 46574
rect 20412 46510 20414 46562
rect 20466 46510 20468 46562
rect 20412 45892 20468 46510
rect 20300 45836 20468 45892
rect 20300 45332 20356 45836
rect 20412 45668 20468 45678
rect 20412 45574 20468 45612
rect 20300 45276 20468 45332
rect 20188 44322 20356 44324
rect 20188 44270 20190 44322
rect 20242 44270 20356 44322
rect 20188 44268 20356 44270
rect 20188 44258 20244 44268
rect 20188 44100 20244 44110
rect 20188 44006 20244 44044
rect 20188 43764 20244 43774
rect 20188 43670 20244 43708
rect 20300 43316 20356 44268
rect 20412 44322 20468 45276
rect 20524 45220 20580 46622
rect 20524 45154 20580 45164
rect 20412 44270 20414 44322
rect 20466 44270 20468 44322
rect 20412 44258 20468 44270
rect 20524 44994 20580 45006
rect 20524 44942 20526 44994
rect 20578 44942 20580 44994
rect 20524 44100 20580 44942
rect 20524 44034 20580 44044
rect 20300 43250 20356 43260
rect 20636 43426 20692 47012
rect 20860 46900 20916 47012
rect 20860 46834 20916 46844
rect 20860 46674 20916 46686
rect 20860 46622 20862 46674
rect 20914 46622 20916 46674
rect 20860 45444 20916 46622
rect 20972 45892 21028 47404
rect 21084 46676 21140 47628
rect 21308 47682 21364 50428
rect 21420 49140 21476 50542
rect 21624 50204 21888 50214
rect 21680 50148 21728 50204
rect 21784 50148 21832 50204
rect 21624 50138 21888 50148
rect 21868 49812 21924 49822
rect 21868 49810 22036 49812
rect 21868 49758 21870 49810
rect 21922 49758 22036 49810
rect 21868 49756 22036 49758
rect 21868 49746 21924 49756
rect 21420 49046 21476 49084
rect 21868 49026 21924 49038
rect 21868 48974 21870 49026
rect 21922 48974 21924 49026
rect 21868 48916 21924 48974
rect 21868 48850 21924 48860
rect 21624 48636 21888 48646
rect 21680 48580 21728 48636
rect 21784 48580 21832 48636
rect 21624 48570 21888 48580
rect 21644 48244 21700 48254
rect 21644 48150 21700 48188
rect 21308 47630 21310 47682
rect 21362 47630 21364 47682
rect 21308 47618 21364 47630
rect 21532 47684 21588 47694
rect 21588 47628 21700 47684
rect 21532 47618 21588 47628
rect 21644 47570 21700 47628
rect 21644 47518 21646 47570
rect 21698 47518 21700 47570
rect 21644 47506 21700 47518
rect 21420 47460 21476 47470
rect 21420 46900 21476 47404
rect 21868 47458 21924 47470
rect 21868 47406 21870 47458
rect 21922 47406 21924 47458
rect 21868 47236 21924 47406
rect 21980 47460 22036 49756
rect 22204 49252 22260 53340
rect 22428 52388 22484 53452
rect 22316 52332 22484 52388
rect 22540 53284 22596 53294
rect 22316 50820 22372 52332
rect 22428 52164 22484 52174
rect 22428 52070 22484 52108
rect 22316 50818 22484 50820
rect 22316 50766 22318 50818
rect 22370 50766 22484 50818
rect 22316 50764 22484 50766
rect 22316 50754 22372 50764
rect 22204 49186 22260 49196
rect 22316 50596 22372 50606
rect 22316 49140 22372 50540
rect 22428 50484 22484 50764
rect 22428 50418 22484 50428
rect 22540 50428 22596 53228
rect 22652 53172 22708 53182
rect 22764 53172 22820 53566
rect 23100 54180 23156 54190
rect 23100 53730 23156 54124
rect 23100 53678 23102 53730
rect 23154 53678 23156 53730
rect 22988 53508 23044 53518
rect 22988 53414 23044 53452
rect 22708 53116 22820 53172
rect 23100 53172 23156 53678
rect 23212 53732 23268 54348
rect 23324 54338 23380 54348
rect 23212 53666 23268 53676
rect 23324 53844 23380 53854
rect 23324 53730 23380 53788
rect 23324 53678 23326 53730
rect 23378 53678 23380 53730
rect 23324 53666 23380 53678
rect 22652 53106 22708 53116
rect 23100 53106 23156 53116
rect 22652 52612 22708 52622
rect 22652 50820 22708 52556
rect 22652 50754 22708 50764
rect 22764 52162 22820 52174
rect 22764 52110 22766 52162
rect 22818 52110 22820 52162
rect 22540 50372 22708 50428
rect 22540 49700 22596 49710
rect 22540 49606 22596 49644
rect 22316 49084 22596 49140
rect 22204 48804 22260 48814
rect 22092 48468 22148 48478
rect 22092 48354 22148 48412
rect 22092 48302 22094 48354
rect 22146 48302 22148 48354
rect 22092 48290 22148 48302
rect 21980 47394 22036 47404
rect 22204 47236 22260 48748
rect 22428 48692 22484 48702
rect 22316 47348 22372 47358
rect 22316 47254 22372 47292
rect 21868 47180 22260 47236
rect 21624 47068 21888 47078
rect 21680 47012 21728 47068
rect 21784 47012 21832 47068
rect 21624 47002 21888 47012
rect 21644 46900 21700 46910
rect 21420 46844 21588 46900
rect 21196 46676 21252 46686
rect 21084 46674 21252 46676
rect 21084 46622 21198 46674
rect 21250 46622 21252 46674
rect 21084 46620 21252 46622
rect 21196 46116 21252 46620
rect 21420 46676 21476 46686
rect 21420 46582 21476 46620
rect 21532 46562 21588 46844
rect 21644 46806 21700 46844
rect 22092 46788 22148 46798
rect 21532 46510 21534 46562
rect 21586 46510 21588 46562
rect 21532 46498 21588 46510
rect 21980 46732 22092 46788
rect 21196 46060 21476 46116
rect 21308 45892 21364 45902
rect 20972 45890 21364 45892
rect 20972 45838 21310 45890
rect 21362 45838 21364 45890
rect 20972 45836 21364 45838
rect 20860 45378 20916 45388
rect 21196 45108 21252 45118
rect 21196 45014 21252 45052
rect 21196 44210 21252 44222
rect 21196 44158 21198 44210
rect 21250 44158 21252 44210
rect 20636 43374 20638 43426
rect 20690 43374 20692 43426
rect 20076 42924 20244 42980
rect 20076 42756 20132 42766
rect 20076 42662 20132 42700
rect 19964 42642 20020 42654
rect 19964 42590 19966 42642
rect 20018 42590 20020 42642
rect 19964 41972 20020 42590
rect 20188 42532 20244 42924
rect 19964 41906 20020 41916
rect 20076 42476 20244 42532
rect 20300 42754 20356 42766
rect 20300 42702 20302 42754
rect 20354 42702 20356 42754
rect 20076 41970 20132 42476
rect 20300 42196 20356 42702
rect 20636 42196 20692 43374
rect 20860 43540 20916 43550
rect 20860 43314 20916 43484
rect 20860 43262 20862 43314
rect 20914 43262 20916 43314
rect 20748 42756 20804 42766
rect 20748 42662 20804 42700
rect 20636 42140 20804 42196
rect 20300 42130 20356 42140
rect 20076 41918 20078 41970
rect 20130 41918 20132 41970
rect 19964 41186 20020 41198
rect 19964 41134 19966 41186
rect 20018 41134 20020 41186
rect 19964 40964 20020 41134
rect 19964 40898 20020 40908
rect 19628 40226 19684 40236
rect 19740 40684 19908 40740
rect 20076 40852 20132 41918
rect 19740 40068 19796 40684
rect 19404 39790 19406 39842
rect 19458 39790 19460 39842
rect 19404 39730 19460 39790
rect 19404 39678 19406 39730
rect 19458 39678 19460 39730
rect 19404 39666 19460 39678
rect 19516 40012 19796 40068
rect 19964 40516 20020 40526
rect 19404 38834 19460 38846
rect 19404 38782 19406 38834
rect 19458 38782 19460 38834
rect 19404 38724 19460 38782
rect 19404 38658 19460 38668
rect 19516 38388 19572 40012
rect 19628 39842 19684 39854
rect 19628 39790 19630 39842
rect 19682 39790 19684 39842
rect 19628 39058 19684 39790
rect 19852 39396 19908 39406
rect 19852 39302 19908 39340
rect 19628 39006 19630 39058
rect 19682 39006 19684 39058
rect 19628 38668 19684 39006
rect 19964 39058 20020 40460
rect 19964 39006 19966 39058
rect 20018 39006 20020 39058
rect 19852 38948 19908 38958
rect 19852 38854 19908 38892
rect 19740 38836 19796 38846
rect 19740 38742 19796 38780
rect 19628 38612 19908 38668
rect 19516 38332 19796 38388
rect 19404 37268 19460 37278
rect 19404 37266 19572 37268
rect 19404 37214 19406 37266
rect 19458 37214 19572 37266
rect 19404 37212 19572 37214
rect 19404 37202 19460 37212
rect 19516 37156 19572 37212
rect 19404 36932 19460 36942
rect 19404 36370 19460 36876
rect 19404 36318 19406 36370
rect 19458 36318 19460 36370
rect 19404 36306 19460 36318
rect 19516 36148 19572 37100
rect 19404 36092 19572 36148
rect 19404 32116 19460 36092
rect 19516 35588 19572 35598
rect 19516 34132 19572 35532
rect 19740 35028 19796 38332
rect 19852 37940 19908 38612
rect 19852 37874 19908 37884
rect 19740 34962 19796 34972
rect 19852 37492 19908 37502
rect 19964 37492 20020 39006
rect 20076 38836 20132 40796
rect 20076 38770 20132 38780
rect 20188 41970 20244 41982
rect 20188 41918 20190 41970
rect 20242 41918 20244 41970
rect 20188 38500 20244 41918
rect 20300 41972 20356 41982
rect 20300 41878 20356 41916
rect 20412 41972 20468 41982
rect 20412 41970 20580 41972
rect 20412 41918 20414 41970
rect 20466 41918 20580 41970
rect 20412 41916 20580 41918
rect 20412 41906 20468 41916
rect 20412 41748 20468 41758
rect 20412 41298 20468 41692
rect 20412 41246 20414 41298
rect 20466 41246 20468 41298
rect 20188 38434 20244 38444
rect 20300 40628 20356 40638
rect 20076 38220 20244 38276
rect 20076 38164 20132 38220
rect 20076 38098 20132 38108
rect 20188 38162 20244 38220
rect 20188 38110 20190 38162
rect 20242 38110 20244 38162
rect 20188 38098 20244 38110
rect 19852 37490 20020 37492
rect 19852 37438 19854 37490
rect 19906 37438 20020 37490
rect 19852 37436 20020 37438
rect 20300 37604 20356 40572
rect 20412 40516 20468 41246
rect 20412 40450 20468 40460
rect 20412 39732 20468 39742
rect 20524 39732 20580 41916
rect 20636 41970 20692 41982
rect 20636 41918 20638 41970
rect 20690 41918 20692 41970
rect 20636 41860 20692 41918
rect 20636 41794 20692 41804
rect 20748 40404 20804 42140
rect 20860 40740 20916 43262
rect 20972 42084 21028 42094
rect 20972 41636 21028 42028
rect 21084 41972 21140 41982
rect 21084 41878 21140 41916
rect 20972 41570 21028 41580
rect 20860 40684 21140 40740
rect 20748 40338 20804 40348
rect 21084 40626 21140 40684
rect 21084 40574 21086 40626
rect 21138 40574 21140 40626
rect 20636 40292 20692 40302
rect 20636 40198 20692 40236
rect 20468 39676 20580 39732
rect 20412 39638 20468 39676
rect 20748 39394 20804 39406
rect 20748 39342 20750 39394
rect 20802 39342 20804 39394
rect 20748 39172 20804 39342
rect 20748 39106 20804 39116
rect 20636 38834 20692 38846
rect 20636 38782 20638 38834
rect 20690 38782 20692 38834
rect 20636 38724 20692 38782
rect 20636 38658 20692 38668
rect 20748 38500 20804 38510
rect 20748 38162 20804 38444
rect 21084 38276 21140 40574
rect 21196 38500 21252 44158
rect 21308 43876 21364 45836
rect 21420 44996 21476 46060
rect 21624 45500 21888 45510
rect 21680 45444 21728 45500
rect 21784 45444 21832 45500
rect 21624 45434 21888 45444
rect 21980 45332 22036 46732
rect 22092 46694 22148 46732
rect 22092 45780 22148 45790
rect 22092 45778 22260 45780
rect 22092 45726 22094 45778
rect 22146 45726 22260 45778
rect 22092 45724 22260 45726
rect 22092 45714 22148 45724
rect 21868 45276 22036 45332
rect 22092 45444 22148 45454
rect 21756 44996 21812 45006
rect 21420 44940 21756 44996
rect 21756 44902 21812 44940
rect 21420 44324 21476 44334
rect 21420 44230 21476 44268
rect 21756 44212 21812 44222
rect 21868 44212 21924 45276
rect 22092 45218 22148 45388
rect 22204 45330 22260 45724
rect 22204 45278 22206 45330
rect 22258 45278 22260 45330
rect 22204 45266 22260 45278
rect 22092 45166 22094 45218
rect 22146 45166 22148 45218
rect 22092 45154 22148 45166
rect 22428 45218 22484 48636
rect 22428 45166 22430 45218
rect 22482 45166 22484 45218
rect 21756 44210 21868 44212
rect 21756 44158 21758 44210
rect 21810 44158 21868 44210
rect 21756 44156 21868 44158
rect 21756 44146 21812 44156
rect 21868 44118 21924 44156
rect 21980 44996 22036 45006
rect 21624 43932 21888 43942
rect 21680 43876 21728 43932
rect 21784 43876 21832 43932
rect 21308 43820 21476 43876
rect 21624 43866 21888 43876
rect 21308 43652 21364 43662
rect 21308 43558 21364 43596
rect 21308 42866 21364 42878
rect 21308 42814 21310 42866
rect 21362 42814 21364 42866
rect 21308 42532 21364 42814
rect 21308 42466 21364 42476
rect 21308 41970 21364 41982
rect 21308 41918 21310 41970
rect 21362 41918 21364 41970
rect 21308 39396 21364 41918
rect 21420 41972 21476 43820
rect 21980 43764 22036 44940
rect 22316 44884 22372 44894
rect 22316 44210 22372 44828
rect 22316 44158 22318 44210
rect 22370 44158 22372 44210
rect 22316 44146 22372 44158
rect 21644 43708 22036 43764
rect 22092 44100 22148 44110
rect 22092 43762 22148 44044
rect 22092 43710 22094 43762
rect 22146 43710 22148 43762
rect 21644 43426 21700 43708
rect 22092 43652 22148 43710
rect 22092 43586 22148 43596
rect 21644 43374 21646 43426
rect 21698 43374 21700 43426
rect 21644 43204 21700 43374
rect 21644 43138 21700 43148
rect 22316 43314 22372 43326
rect 22316 43262 22318 43314
rect 22370 43262 22372 43314
rect 22204 42532 22260 42542
rect 21624 42364 21888 42374
rect 21680 42308 21728 42364
rect 21784 42308 21832 42364
rect 21624 42298 21888 42308
rect 21868 42196 21924 42206
rect 21868 42102 21924 42140
rect 22092 42084 22148 42094
rect 21420 41906 21476 41916
rect 21868 41970 21924 41982
rect 21868 41918 21870 41970
rect 21922 41918 21924 41970
rect 21644 41748 21700 41758
rect 21644 41654 21700 41692
rect 21420 41412 21476 41422
rect 21420 41298 21476 41356
rect 21420 41246 21422 41298
rect 21474 41246 21476 41298
rect 21420 41234 21476 41246
rect 21868 41188 21924 41918
rect 21868 41122 21924 41132
rect 21868 40964 21924 40974
rect 21868 40962 22036 40964
rect 21868 40910 21870 40962
rect 21922 40910 22036 40962
rect 21868 40908 22036 40910
rect 21868 40898 21924 40908
rect 21420 40852 21476 40862
rect 21980 40852 22036 40908
rect 22092 40852 22148 42028
rect 22204 41970 22260 42476
rect 22204 41918 22206 41970
rect 22258 41918 22260 41970
rect 22204 41906 22260 41918
rect 22204 41748 22260 41758
rect 22204 41654 22260 41692
rect 22316 41636 22372 43262
rect 22316 41188 22372 41580
rect 22428 41410 22484 45166
rect 22540 43652 22596 49084
rect 22652 46228 22708 50372
rect 22764 47572 22820 52110
rect 22988 52162 23044 52174
rect 22988 52110 22990 52162
rect 23042 52110 23044 52162
rect 22988 51604 23044 52110
rect 23548 52164 23604 57932
rect 23996 57876 24052 59166
rect 23996 57810 24052 57820
rect 24108 58212 24164 61628
rect 24220 61572 24276 61582
rect 24332 61572 24388 62972
rect 24220 61570 24388 61572
rect 24220 61518 24222 61570
rect 24274 61518 24388 61570
rect 24220 61516 24388 61518
rect 24220 61506 24276 61516
rect 24332 61348 24388 61358
rect 24332 61254 24388 61292
rect 24444 61346 24500 65212
rect 24444 61294 24446 61346
rect 24498 61294 24500 61346
rect 24108 57876 24164 58156
rect 24332 60676 24388 60686
rect 24444 60676 24500 61294
rect 24332 60674 24500 60676
rect 24332 60622 24334 60674
rect 24386 60622 24500 60674
rect 24332 60620 24500 60622
rect 24220 57876 24276 57886
rect 24108 57874 24276 57876
rect 24108 57822 24222 57874
rect 24274 57822 24276 57874
rect 24108 57820 24276 57822
rect 23884 57764 23940 57774
rect 23884 57670 23940 57708
rect 23772 57650 23828 57662
rect 23772 57598 23774 57650
rect 23826 57598 23828 57650
rect 23772 57428 23828 57598
rect 23772 57362 23828 57372
rect 23996 57650 24052 57662
rect 23996 57598 23998 57650
rect 24050 57598 24052 57650
rect 23996 56980 24052 57598
rect 24108 57316 24164 57820
rect 24220 57810 24276 57820
rect 24108 57250 24164 57260
rect 24332 57092 24388 60620
rect 24556 60228 24612 66892
rect 24668 65828 24724 65838
rect 24668 64818 24724 65772
rect 24668 64766 24670 64818
rect 24722 64766 24724 64818
rect 24668 64148 24724 64766
rect 24668 64054 24724 64092
rect 24780 65492 24836 65502
rect 24668 63698 24724 63710
rect 24668 63646 24670 63698
rect 24722 63646 24724 63698
rect 24668 62578 24724 63646
rect 24780 63588 24836 65436
rect 24780 63522 24836 63532
rect 24668 62526 24670 62578
rect 24722 62526 24724 62578
rect 24668 62514 24724 62526
rect 24668 62244 24724 62254
rect 24668 61570 24724 62188
rect 24668 61518 24670 61570
rect 24722 61518 24724 61570
rect 24668 61506 24724 61518
rect 24780 60228 24836 60238
rect 24556 60172 24724 60228
rect 24556 60004 24612 60014
rect 24556 59910 24612 59948
rect 24556 59444 24612 59454
rect 24444 59108 24500 59118
rect 24556 59108 24612 59388
rect 24500 59052 24612 59108
rect 24444 59014 24500 59052
rect 24444 58324 24500 58334
rect 24444 58210 24500 58268
rect 24444 58158 24446 58210
rect 24498 58158 24500 58210
rect 24444 57876 24500 58158
rect 24444 57810 24500 57820
rect 24444 57428 24500 57438
rect 24556 57428 24612 59052
rect 24500 57372 24612 57428
rect 24444 57362 24500 57372
rect 24668 57204 24724 60172
rect 24780 57204 24836 60172
rect 24892 58548 24948 73836
rect 25340 73892 25396 73902
rect 25340 73332 25396 73836
rect 25452 73556 25508 77308
rect 25564 77028 25620 77420
rect 25564 76962 25620 76972
rect 25676 76020 25732 78542
rect 26124 78594 26180 78606
rect 26124 78542 26126 78594
rect 26178 78542 26180 78594
rect 26012 77924 26068 77934
rect 26012 77830 26068 77868
rect 25900 77140 25956 77150
rect 25900 76466 25956 77084
rect 25900 76414 25902 76466
rect 25954 76414 25956 76466
rect 25900 76402 25956 76414
rect 25564 75964 25732 76020
rect 25564 74228 25620 75964
rect 25676 75796 25732 75806
rect 25676 75702 25732 75740
rect 26124 75236 26180 78542
rect 26236 77140 26292 77150
rect 26236 76690 26292 77084
rect 26460 76804 26516 78878
rect 26908 79548 27412 79604
rect 26908 78930 26964 79548
rect 27580 79490 27636 79502
rect 27580 79438 27582 79490
rect 27634 79438 27636 79490
rect 27356 79378 27412 79390
rect 27356 79326 27358 79378
rect 27410 79326 27412 79378
rect 27356 78932 27412 79326
rect 26908 78878 26910 78930
rect 26962 78878 26964 78930
rect 26684 76916 26740 76926
rect 26516 76748 26628 76804
rect 26460 76738 26516 76748
rect 26236 76638 26238 76690
rect 26290 76638 26292 76690
rect 26236 76626 26292 76638
rect 26348 76468 26404 76478
rect 26348 76374 26404 76412
rect 26460 76466 26516 76478
rect 26460 76414 26462 76466
rect 26514 76414 26516 76466
rect 26460 75794 26516 76414
rect 26460 75742 26462 75794
rect 26514 75742 26516 75794
rect 26460 75730 26516 75742
rect 26572 75684 26628 76748
rect 26572 75618 26628 75628
rect 26348 75458 26404 75470
rect 26572 75460 26628 75470
rect 26348 75406 26350 75458
rect 26402 75406 26404 75458
rect 26124 75180 26292 75236
rect 25788 74786 25844 74798
rect 25788 74734 25790 74786
rect 25842 74734 25844 74786
rect 25676 74228 25732 74238
rect 25564 74172 25676 74228
rect 25676 74162 25732 74172
rect 25676 74004 25732 74042
rect 25676 73938 25732 73948
rect 25452 73490 25508 73500
rect 25564 73890 25620 73902
rect 25564 73838 25566 73890
rect 25618 73838 25620 73890
rect 25340 73330 25508 73332
rect 25340 73278 25342 73330
rect 25394 73278 25508 73330
rect 25340 73276 25508 73278
rect 25340 73266 25396 73276
rect 25026 72940 25290 72950
rect 25082 72884 25130 72940
rect 25186 72884 25234 72940
rect 25026 72874 25290 72884
rect 25004 72322 25060 72334
rect 25004 72270 25006 72322
rect 25058 72270 25060 72322
rect 25004 72212 25060 72270
rect 25004 72146 25060 72156
rect 25340 71650 25396 71662
rect 25340 71598 25342 71650
rect 25394 71598 25396 71650
rect 25340 71540 25396 71598
rect 25340 71474 25396 71484
rect 25026 71372 25290 71382
rect 25082 71316 25130 71372
rect 25186 71316 25234 71372
rect 25026 71306 25290 71316
rect 25340 70980 25396 70990
rect 25452 70980 25508 73276
rect 25564 71876 25620 73838
rect 25788 72884 25844 74734
rect 26124 74788 26180 74798
rect 26124 74694 26180 74732
rect 25788 72818 25844 72828
rect 25900 74674 25956 74686
rect 25900 74622 25902 74674
rect 25954 74622 25956 74674
rect 25900 74114 25956 74622
rect 25900 74062 25902 74114
rect 25954 74062 25956 74114
rect 25564 71810 25620 71820
rect 25676 72546 25732 72558
rect 25676 72494 25678 72546
rect 25730 72494 25732 72546
rect 25676 72100 25732 72494
rect 25340 70978 25508 70980
rect 25340 70926 25342 70978
rect 25394 70926 25508 70978
rect 25340 70924 25508 70926
rect 25340 70914 25396 70924
rect 25676 70420 25732 72044
rect 25452 70418 25732 70420
rect 25452 70366 25678 70418
rect 25730 70366 25732 70418
rect 25452 70364 25732 70366
rect 25026 69804 25290 69814
rect 25082 69748 25130 69804
rect 25186 69748 25234 69804
rect 25026 69738 25290 69748
rect 25340 69524 25396 69534
rect 25452 69524 25508 70364
rect 25676 70354 25732 70364
rect 25900 70194 25956 74062
rect 26236 74114 26292 75180
rect 26348 74900 26404 75406
rect 26348 74834 26404 74844
rect 26460 75458 26628 75460
rect 26460 75406 26574 75458
rect 26626 75406 26628 75458
rect 26460 75404 26628 75406
rect 26236 74062 26238 74114
rect 26290 74062 26292 74114
rect 26124 73890 26180 73902
rect 26124 73838 26126 73890
rect 26178 73838 26180 73890
rect 26012 73444 26068 73454
rect 26124 73444 26180 73838
rect 26012 73442 26180 73444
rect 26012 73390 26014 73442
rect 26066 73390 26180 73442
rect 26012 73388 26180 73390
rect 26012 73378 26068 73388
rect 26012 71650 26068 71662
rect 26012 71598 26014 71650
rect 26066 71598 26068 71650
rect 26012 71092 26068 71598
rect 26012 71026 26068 71036
rect 26012 70866 26068 70878
rect 26012 70814 26014 70866
rect 26066 70814 26068 70866
rect 26012 70420 26068 70814
rect 26124 70420 26180 70430
rect 26012 70418 26180 70420
rect 26012 70366 26126 70418
rect 26178 70366 26180 70418
rect 26012 70364 26180 70366
rect 26124 70354 26180 70364
rect 25900 70142 25902 70194
rect 25954 70142 25956 70194
rect 25340 69522 25508 69524
rect 25340 69470 25342 69522
rect 25394 69470 25508 69522
rect 25340 69468 25508 69470
rect 25788 70084 25844 70094
rect 25788 69522 25844 70028
rect 25788 69470 25790 69522
rect 25842 69470 25844 69522
rect 25340 68740 25396 69468
rect 25788 69458 25844 69470
rect 25340 68674 25396 68684
rect 25788 69300 25844 69310
rect 25900 69300 25956 70142
rect 25844 69244 25956 69300
rect 25228 68516 25284 68526
rect 25228 68422 25284 68460
rect 25026 68236 25290 68246
rect 25082 68180 25130 68236
rect 25186 68180 25234 68236
rect 25026 68170 25290 68180
rect 25340 67172 25396 67182
rect 25396 67116 25508 67172
rect 25340 67106 25396 67116
rect 25228 66946 25284 66958
rect 25228 66894 25230 66946
rect 25282 66894 25284 66946
rect 25228 66836 25284 66894
rect 25228 66770 25284 66780
rect 25026 66668 25290 66678
rect 25082 66612 25130 66668
rect 25186 66612 25234 66668
rect 25026 66602 25290 66612
rect 25452 65828 25508 67116
rect 25340 65772 25732 65828
rect 25340 65490 25396 65772
rect 25340 65438 25342 65490
rect 25394 65438 25396 65490
rect 25340 65426 25396 65438
rect 25452 65604 25508 65614
rect 25026 65100 25290 65110
rect 25082 65044 25130 65100
rect 25186 65044 25234 65100
rect 25026 65034 25290 65044
rect 25340 64708 25396 64718
rect 25452 64708 25508 65548
rect 25340 64706 25508 64708
rect 25340 64654 25342 64706
rect 25394 64654 25508 64706
rect 25340 64652 25508 64654
rect 25564 65380 25620 65390
rect 25340 64642 25396 64652
rect 25564 64484 25620 65324
rect 25676 65268 25732 65772
rect 25788 65492 25844 69244
rect 26012 68740 26068 68750
rect 26012 67844 26068 68684
rect 26012 67750 26068 67788
rect 25788 65398 25844 65436
rect 26124 65490 26180 65502
rect 26124 65438 26126 65490
rect 26178 65438 26180 65490
rect 25900 65380 25956 65390
rect 26124 65380 26180 65438
rect 25900 65378 26068 65380
rect 25900 65326 25902 65378
rect 25954 65326 26068 65378
rect 25900 65324 26068 65326
rect 25900 65314 25956 65324
rect 25676 65212 25844 65268
rect 25564 64418 25620 64428
rect 25228 64204 25620 64260
rect 25116 64148 25172 64158
rect 25116 63922 25172 64092
rect 25116 63870 25118 63922
rect 25170 63870 25172 63922
rect 25116 63858 25172 63870
rect 25228 63700 25284 64204
rect 25564 64146 25620 64204
rect 25564 64094 25566 64146
rect 25618 64094 25620 64146
rect 25564 64082 25620 64094
rect 25676 64148 25732 64158
rect 25676 64054 25732 64092
rect 25788 63924 25844 65212
rect 26012 64818 26068 65324
rect 26124 65314 26180 65324
rect 26012 64766 26014 64818
rect 26066 64766 26068 64818
rect 26012 64754 26068 64766
rect 25788 63830 25844 63868
rect 25900 64484 25956 64494
rect 25676 63812 25732 63822
rect 25228 63644 25508 63700
rect 25026 63532 25290 63542
rect 25082 63476 25130 63532
rect 25186 63476 25234 63532
rect 25026 63466 25290 63476
rect 25228 62244 25284 62254
rect 25452 62244 25508 63644
rect 25284 62188 25508 62244
rect 25228 62150 25284 62188
rect 25026 61964 25290 61974
rect 25082 61908 25130 61964
rect 25186 61908 25234 61964
rect 25026 61898 25290 61908
rect 25340 61796 25396 61806
rect 25116 61346 25172 61358
rect 25116 61294 25118 61346
rect 25170 61294 25172 61346
rect 25116 61236 25172 61294
rect 25116 61170 25172 61180
rect 25340 60564 25396 61740
rect 25676 61572 25732 63756
rect 25900 63700 25956 64428
rect 26012 64148 26068 64158
rect 26068 64092 26180 64148
rect 26012 64082 26068 64092
rect 26124 64034 26180 64092
rect 26124 63982 26126 64034
rect 26178 63982 26180 64034
rect 26124 63970 26180 63982
rect 25452 61570 25732 61572
rect 25452 61518 25678 61570
rect 25730 61518 25732 61570
rect 25452 61516 25732 61518
rect 25452 61010 25508 61516
rect 25676 61506 25732 61516
rect 25788 63644 25956 63700
rect 25452 60958 25454 61010
rect 25506 60958 25508 61010
rect 25452 60946 25508 60958
rect 25676 60900 25732 60910
rect 25340 60508 25620 60564
rect 25026 60396 25290 60406
rect 25082 60340 25130 60396
rect 25186 60340 25234 60396
rect 25026 60330 25290 60340
rect 25340 60004 25396 60014
rect 25340 59108 25396 59948
rect 25340 59106 25508 59108
rect 25340 59054 25342 59106
rect 25394 59054 25508 59106
rect 25340 59052 25508 59054
rect 25340 59042 25396 59052
rect 25452 58884 25508 59052
rect 25026 58828 25290 58838
rect 25082 58772 25130 58828
rect 25186 58772 25234 58828
rect 25026 58762 25290 58772
rect 24892 58482 24948 58492
rect 25340 58436 25396 58446
rect 25452 58436 25508 58828
rect 25340 58434 25508 58436
rect 25340 58382 25342 58434
rect 25394 58382 25508 58434
rect 25340 58380 25508 58382
rect 25340 58370 25396 58380
rect 24892 58212 24948 58222
rect 24892 58118 24948 58156
rect 25340 57538 25396 57550
rect 25340 57486 25342 57538
rect 25394 57486 25396 57538
rect 25340 57428 25396 57486
rect 25340 57362 25396 57372
rect 25026 57260 25290 57270
rect 25082 57204 25130 57260
rect 25186 57204 25234 57260
rect 24780 57148 24948 57204
rect 25026 57194 25290 57204
rect 24668 57138 24724 57148
rect 23884 56196 23940 56206
rect 23996 56196 24052 56924
rect 23884 56194 24052 56196
rect 23884 56142 23886 56194
rect 23938 56142 24052 56194
rect 23884 56140 24052 56142
rect 24108 57036 24388 57092
rect 23884 56130 23940 56140
rect 23660 56084 23716 56094
rect 23660 56082 23828 56084
rect 23660 56030 23662 56082
rect 23714 56030 23828 56082
rect 23660 56028 23828 56030
rect 23660 56018 23716 56028
rect 23660 55074 23716 55086
rect 23660 55022 23662 55074
rect 23714 55022 23716 55074
rect 23660 54516 23716 55022
rect 23772 54628 23828 56028
rect 24108 55074 24164 57036
rect 24556 56980 24612 56990
rect 24780 56980 24836 56990
rect 24612 56978 24836 56980
rect 24612 56926 24782 56978
rect 24834 56926 24836 56978
rect 24612 56924 24836 56926
rect 24556 56914 24612 56924
rect 24780 56914 24836 56924
rect 24332 56644 24388 56654
rect 24332 55970 24388 56588
rect 24332 55918 24334 55970
rect 24386 55918 24388 55970
rect 24108 55022 24110 55074
rect 24162 55022 24164 55074
rect 23772 54562 23828 54572
rect 23884 54852 23940 54862
rect 23660 54450 23716 54460
rect 23772 54402 23828 54414
rect 23772 54350 23774 54402
rect 23826 54350 23828 54402
rect 23772 54068 23828 54350
rect 23772 54002 23828 54012
rect 23884 53732 23940 54796
rect 24108 54740 24164 55022
rect 24108 54674 24164 54684
rect 24220 55748 24276 55758
rect 24332 55748 24388 55918
rect 24276 55692 24388 55748
rect 24220 54738 24276 55692
rect 24220 54686 24222 54738
rect 24274 54686 24276 54738
rect 24220 54674 24276 54686
rect 24556 55188 24612 55198
rect 24556 55074 24612 55132
rect 24556 55022 24558 55074
rect 24610 55022 24612 55074
rect 24556 54290 24612 55022
rect 24668 54964 24724 54974
rect 24668 54738 24724 54908
rect 24668 54686 24670 54738
rect 24722 54686 24724 54738
rect 24668 54674 24724 54686
rect 24556 54238 24558 54290
rect 24610 54238 24612 54290
rect 24556 54226 24612 54238
rect 24108 53844 24164 53854
rect 24108 53750 24164 53788
rect 23772 53676 23940 53732
rect 23772 53618 23828 53676
rect 23772 53566 23774 53618
rect 23826 53566 23828 53618
rect 23772 53554 23828 53566
rect 23996 53620 24052 53630
rect 23996 53526 24052 53564
rect 23884 53508 23940 53518
rect 23884 53058 23940 53452
rect 24220 53508 24276 53518
rect 24220 53414 24276 53452
rect 24668 53506 24724 53518
rect 24668 53454 24670 53506
rect 24722 53454 24724 53506
rect 24556 53396 24612 53406
rect 24668 53396 24724 53454
rect 24612 53340 24724 53396
rect 24556 53330 24612 53340
rect 24892 53172 24948 57148
rect 25340 56084 25396 56094
rect 25452 56084 25508 58380
rect 25564 57764 25620 60508
rect 25564 56980 25620 57708
rect 25564 56886 25620 56924
rect 25676 58660 25732 60844
rect 25676 56196 25732 58604
rect 25676 56130 25732 56140
rect 25340 56082 25508 56084
rect 25340 56030 25342 56082
rect 25394 56030 25508 56082
rect 25340 56028 25508 56030
rect 25788 56084 25844 63644
rect 25900 63252 25956 63262
rect 25900 62188 25956 63196
rect 25900 62132 26180 62188
rect 26012 59890 26068 59902
rect 26012 59838 26014 59890
rect 26066 59838 26068 59890
rect 26012 59442 26068 59838
rect 26012 59390 26014 59442
rect 26066 59390 26068 59442
rect 26012 59378 26068 59390
rect 25900 59330 25956 59342
rect 25900 59278 25902 59330
rect 25954 59278 25956 59330
rect 25900 59108 25956 59278
rect 25900 58548 25956 59052
rect 25900 57762 25956 58492
rect 26012 58322 26068 58334
rect 26012 58270 26014 58322
rect 26066 58270 26068 58322
rect 26012 57874 26068 58270
rect 26012 57822 26014 57874
rect 26066 57822 26068 57874
rect 26012 57810 26068 57822
rect 25900 57710 25902 57762
rect 25954 57710 25956 57762
rect 25900 56756 25956 57710
rect 25900 56690 25956 56700
rect 26012 56644 26068 56654
rect 26012 56550 26068 56588
rect 25340 56018 25396 56028
rect 25788 56018 25844 56028
rect 25676 55972 25732 55982
rect 25452 55916 25676 55972
rect 25026 55692 25290 55702
rect 25082 55636 25130 55692
rect 25186 55636 25234 55692
rect 25026 55626 25290 55636
rect 25116 55298 25172 55310
rect 25116 55246 25118 55298
rect 25170 55246 25172 55298
rect 25116 55188 25172 55246
rect 25116 54290 25172 55132
rect 25340 55300 25396 55310
rect 25340 54740 25396 55244
rect 25452 55074 25508 55916
rect 25676 55906 25732 55916
rect 26012 55972 26068 55982
rect 26012 55878 26068 55916
rect 26124 55748 26180 62132
rect 26236 61796 26292 74062
rect 26460 73556 26516 75404
rect 26572 75394 26628 75404
rect 26684 75122 26740 76860
rect 26908 76690 26964 78878
rect 27020 78930 27412 78932
rect 27020 78878 27358 78930
rect 27410 78878 27412 78930
rect 27020 78876 27412 78878
rect 27020 76916 27076 78876
rect 27356 78866 27412 78876
rect 27356 77140 27412 77150
rect 27356 77046 27412 77084
rect 27020 76850 27076 76860
rect 27132 77028 27188 77038
rect 26908 76638 26910 76690
rect 26962 76638 26964 76690
rect 26684 75070 26686 75122
rect 26738 75070 26740 75122
rect 26684 74674 26740 75070
rect 26684 74622 26686 74674
rect 26738 74622 26740 74674
rect 26684 74610 26740 74622
rect 26796 76468 26852 76478
rect 26796 74452 26852 76412
rect 26796 74386 26852 74396
rect 26908 75460 26964 76638
rect 27020 76692 27076 76702
rect 27020 76598 27076 76636
rect 27132 76466 27188 76972
rect 27132 76414 27134 76466
rect 27186 76414 27188 76466
rect 27020 75684 27076 75694
rect 27020 75590 27076 75628
rect 27132 75572 27188 76414
rect 27132 75506 27188 75516
rect 27356 76578 27412 76590
rect 27356 76526 27358 76578
rect 27410 76526 27412 76578
rect 27356 75794 27412 76526
rect 27580 76468 27636 79438
rect 28028 79378 28084 79774
rect 28028 79326 28030 79378
rect 28082 79326 28084 79378
rect 28028 79314 28084 79326
rect 28140 78932 28196 78942
rect 28028 78876 28140 78932
rect 28028 77250 28084 78876
rect 28140 78838 28196 78876
rect 28428 78428 28692 78438
rect 28484 78372 28532 78428
rect 28588 78372 28636 78428
rect 28428 78362 28692 78372
rect 28028 77198 28030 77250
rect 28082 77198 28084 77250
rect 28028 76692 28084 77198
rect 28140 77922 28196 77934
rect 28140 77870 28142 77922
rect 28194 77870 28196 77922
rect 28140 77028 28196 77870
rect 28140 76962 28196 76972
rect 28428 76860 28692 76870
rect 28484 76804 28532 76860
rect 28588 76804 28636 76860
rect 28428 76794 28692 76804
rect 28140 76692 28196 76702
rect 28028 76690 28196 76692
rect 28028 76638 28142 76690
rect 28194 76638 28196 76690
rect 28028 76636 28196 76638
rect 27580 76402 27636 76412
rect 27356 75742 27358 75794
rect 27410 75742 27412 75794
rect 27356 75684 27412 75742
rect 26572 74116 26628 74126
rect 26572 74022 26628 74060
rect 26908 73892 26964 75404
rect 27132 74786 27188 74798
rect 27132 74734 27134 74786
rect 27186 74734 27188 74786
rect 27132 74674 27188 74734
rect 27132 74622 27134 74674
rect 27186 74622 27188 74674
rect 27132 74610 27188 74622
rect 27020 74116 27076 74126
rect 27020 74022 27076 74060
rect 27132 74004 27188 74042
rect 27356 74004 27412 75628
rect 27804 75460 27860 75470
rect 27804 75366 27860 75404
rect 28140 75124 28196 76636
rect 28428 75292 28692 75302
rect 28484 75236 28532 75292
rect 28588 75236 28636 75292
rect 28428 75226 28692 75236
rect 28140 75122 28308 75124
rect 28140 75070 28142 75122
rect 28194 75070 28308 75122
rect 28140 75068 28308 75070
rect 28140 75058 28196 75068
rect 27580 74786 27636 74798
rect 27580 74734 27582 74786
rect 27634 74734 27636 74786
rect 27580 74674 27636 74734
rect 27580 74622 27582 74674
rect 27634 74622 27636 74674
rect 27580 74610 27636 74622
rect 27132 73938 27188 73948
rect 27244 74002 27412 74004
rect 27244 73950 27358 74002
rect 27410 73950 27412 74002
rect 27244 73948 27412 73950
rect 26460 73490 26516 73500
rect 26572 73890 26964 73892
rect 26572 73838 26910 73890
rect 26962 73838 26964 73890
rect 26572 73836 26964 73838
rect 26460 72884 26516 72894
rect 26460 72212 26516 72828
rect 26348 72156 26516 72212
rect 26348 70308 26404 72156
rect 26460 71988 26516 71998
rect 26572 71988 26628 73836
rect 26908 73826 26964 73836
rect 26460 71986 26628 71988
rect 26460 71934 26462 71986
rect 26514 71934 26628 71986
rect 26460 71932 26628 71934
rect 26684 73668 26740 73678
rect 26684 72100 26740 73612
rect 27244 73668 27300 73948
rect 27356 73938 27412 73948
rect 27580 74340 27636 74350
rect 27580 74116 27636 74284
rect 28028 74228 28084 74238
rect 27916 74116 27972 74126
rect 27580 74114 27972 74116
rect 27580 74062 27918 74114
rect 27970 74062 27972 74114
rect 27580 74060 27972 74062
rect 27244 73602 27300 73612
rect 26684 71988 26740 72044
rect 27468 71988 27524 71998
rect 26684 71932 27188 71988
rect 26460 71922 26516 71932
rect 26684 71764 26740 71774
rect 26684 71762 27076 71764
rect 26684 71710 26686 71762
rect 26738 71710 27076 71762
rect 26684 71708 27076 71710
rect 26684 71698 26740 71708
rect 26572 71650 26628 71662
rect 26572 71598 26574 71650
rect 26626 71598 26628 71650
rect 26348 70306 26516 70308
rect 26348 70254 26350 70306
rect 26402 70254 26516 70306
rect 26348 70252 26516 70254
rect 26348 70242 26404 70252
rect 26348 69300 26404 69310
rect 26348 69206 26404 69244
rect 26460 65828 26516 70252
rect 26572 70306 26628 71598
rect 26572 70254 26574 70306
rect 26626 70254 26628 70306
rect 26572 70242 26628 70254
rect 26684 71092 26740 71102
rect 26684 69410 26740 71036
rect 27020 71092 27076 71708
rect 27020 70306 27076 71036
rect 27132 71762 27188 71932
rect 27468 71894 27524 71932
rect 27132 71710 27134 71762
rect 27186 71710 27188 71762
rect 27132 70420 27188 71710
rect 27132 70354 27188 70364
rect 27020 70254 27022 70306
rect 27074 70254 27076 70306
rect 27020 70242 27076 70254
rect 26684 69358 26686 69410
rect 26738 69358 26740 69410
rect 26572 69186 26628 69198
rect 26572 69134 26574 69186
rect 26626 69134 26628 69186
rect 26572 67396 26628 69134
rect 26572 67330 26628 67340
rect 26460 65772 26628 65828
rect 26348 65492 26404 65502
rect 26348 65490 26516 65492
rect 26348 65438 26350 65490
rect 26402 65438 26516 65490
rect 26348 65436 26516 65438
rect 26348 65426 26404 65436
rect 26348 64708 26404 64718
rect 26348 64034 26404 64652
rect 26348 63982 26350 64034
rect 26402 63982 26404 64034
rect 26348 63252 26404 63982
rect 26460 63700 26516 65436
rect 26572 64148 26628 65772
rect 26572 64082 26628 64092
rect 26460 63634 26516 63644
rect 26572 63810 26628 63822
rect 26572 63758 26574 63810
rect 26626 63758 26628 63810
rect 26348 63186 26404 63196
rect 26572 62916 26628 63758
rect 26572 62850 26628 62860
rect 26236 61730 26292 61740
rect 26684 60900 26740 69358
rect 26796 70084 26852 70094
rect 26796 67228 26852 70028
rect 27468 70084 27524 70094
rect 27468 69990 27524 70028
rect 26908 69972 26964 69982
rect 26908 69878 26964 69916
rect 27580 69410 27636 74060
rect 27916 74050 27972 74060
rect 27580 69358 27582 69410
rect 27634 69358 27636 69410
rect 27580 69346 27636 69358
rect 27692 72660 27748 72670
rect 28028 72660 28084 74172
rect 28140 74004 28196 74014
rect 28140 73218 28196 73948
rect 28140 73166 28142 73218
rect 28194 73166 28196 73218
rect 28140 73154 28196 73166
rect 28252 73892 28308 75068
rect 27692 72658 28084 72660
rect 27692 72606 27694 72658
rect 27746 72606 28084 72658
rect 27692 72604 28084 72606
rect 26908 69300 26964 69310
rect 26908 69298 27076 69300
rect 26908 69246 26910 69298
rect 26962 69246 27076 69298
rect 26908 69244 27076 69246
rect 26908 69234 26964 69244
rect 27020 67954 27076 69244
rect 27244 69298 27300 69310
rect 27244 69246 27246 69298
rect 27298 69246 27300 69298
rect 27244 68404 27300 69246
rect 27580 69186 27636 69198
rect 27580 69134 27582 69186
rect 27634 69134 27636 69186
rect 27580 68852 27636 69134
rect 27356 68796 27636 68852
rect 27356 68738 27412 68796
rect 27356 68686 27358 68738
rect 27410 68686 27412 68738
rect 27356 68674 27412 68686
rect 27244 68338 27300 68348
rect 27020 67902 27022 67954
rect 27074 67902 27076 67954
rect 27020 67890 27076 67902
rect 27356 67844 27412 67854
rect 27356 67730 27412 67788
rect 27356 67678 27358 67730
rect 27410 67678 27412 67730
rect 27356 67666 27412 67678
rect 26908 67618 26964 67630
rect 26908 67566 26910 67618
rect 26962 67566 26964 67618
rect 26908 67228 26964 67566
rect 26796 67172 26964 67228
rect 27132 67618 27188 67630
rect 27132 67566 27134 67618
rect 27186 67566 27188 67618
rect 26796 67096 26852 67116
rect 27132 66836 27188 67566
rect 27356 67396 27412 67406
rect 27356 67170 27412 67340
rect 27356 67118 27358 67170
rect 27410 67118 27412 67170
rect 27356 67106 27412 67118
rect 27132 66770 27188 66780
rect 26908 65492 26964 65502
rect 26796 63924 26852 63934
rect 26908 63924 26964 65436
rect 27356 65380 27412 65390
rect 27356 65286 27412 65324
rect 27020 64932 27076 64942
rect 27020 64148 27076 64876
rect 27020 64146 27412 64148
rect 27020 64094 27022 64146
rect 27074 64094 27412 64146
rect 27020 64092 27412 64094
rect 27020 64082 27076 64092
rect 26796 63922 26964 63924
rect 26796 63870 26798 63922
rect 26850 63870 26964 63922
rect 26796 63868 26964 63870
rect 27244 63922 27300 63934
rect 27244 63870 27246 63922
rect 27298 63870 27300 63922
rect 26796 63858 26852 63868
rect 27132 63812 27188 63822
rect 27132 63718 27188 63756
rect 27244 63700 27300 63870
rect 26796 63588 26852 63598
rect 26796 63140 26852 63532
rect 27020 63252 27076 63262
rect 27020 63158 27076 63196
rect 26796 61012 26852 63084
rect 27244 63028 27300 63644
rect 27356 63252 27412 64092
rect 27468 64036 27524 64046
rect 27468 63942 27524 63980
rect 27468 63252 27524 63262
rect 27356 63250 27524 63252
rect 27356 63198 27470 63250
rect 27522 63198 27524 63250
rect 27356 63196 27524 63198
rect 27468 63186 27524 63196
rect 27244 62962 27300 62972
rect 27356 62916 27412 62926
rect 27356 62466 27412 62860
rect 27356 62414 27358 62466
rect 27410 62414 27412 62466
rect 27356 62402 27412 62414
rect 27692 62188 27748 72604
rect 28140 71988 28196 71998
rect 28252 71988 28308 73836
rect 28428 73724 28692 73734
rect 28484 73668 28532 73724
rect 28588 73668 28636 73724
rect 28428 73658 28692 73668
rect 28428 72156 28692 72166
rect 28484 72100 28532 72156
rect 28588 72100 28636 72156
rect 28428 72090 28692 72100
rect 28140 71986 28308 71988
rect 28140 71934 28142 71986
rect 28194 71934 28308 71986
rect 28140 71932 28308 71934
rect 28140 71922 28196 71932
rect 28140 71092 28196 71102
rect 28140 70998 28196 71036
rect 27916 70420 27972 70430
rect 27916 70326 27972 70364
rect 27804 69300 27860 69310
rect 27804 69206 27860 69244
rect 28140 68628 28196 68638
rect 28252 68628 28308 71932
rect 28428 70588 28692 70598
rect 28484 70532 28532 70588
rect 28588 70532 28636 70588
rect 28428 70522 28692 70532
rect 28428 69020 28692 69030
rect 28484 68964 28532 69020
rect 28588 68964 28636 69020
rect 28428 68954 28692 68964
rect 28140 68626 28308 68628
rect 28140 68574 28142 68626
rect 28194 68574 28308 68626
rect 28140 68572 28308 68574
rect 28140 67954 28196 68572
rect 28140 67902 28142 67954
rect 28194 67902 28196 67954
rect 28140 67060 28196 67902
rect 28428 67452 28692 67462
rect 28484 67396 28532 67452
rect 28588 67396 28636 67452
rect 28428 67386 28692 67396
rect 27916 67058 28196 67060
rect 27916 67006 28142 67058
rect 28194 67006 28196 67058
rect 27916 67004 28196 67006
rect 27916 66386 27972 67004
rect 28140 66994 28196 67004
rect 27916 66334 27918 66386
rect 27970 66334 27972 66386
rect 27916 65604 27972 66334
rect 28428 65884 28692 65894
rect 28484 65828 28532 65884
rect 28588 65828 28636 65884
rect 28428 65818 28692 65828
rect 27804 65492 27860 65502
rect 27804 65398 27860 65436
rect 27916 63252 27972 65548
rect 28140 64818 28196 64830
rect 28140 64766 28142 64818
rect 28194 64766 28196 64818
rect 28028 64036 28084 64046
rect 28028 63942 28084 63980
rect 28140 63700 28196 64766
rect 28428 64316 28692 64326
rect 28484 64260 28532 64316
rect 28588 64260 28636 64316
rect 28428 64250 28692 64260
rect 28140 63634 28196 63644
rect 28140 63252 28196 63262
rect 27916 63250 28196 63252
rect 27916 63198 28142 63250
rect 28194 63198 28196 63250
rect 27916 63196 28196 63198
rect 27580 62132 27748 62188
rect 28028 62354 28084 63196
rect 28140 63186 28196 63196
rect 28428 62748 28692 62758
rect 28484 62692 28532 62748
rect 28588 62692 28636 62748
rect 28428 62682 28692 62692
rect 28028 62302 28030 62354
rect 28082 62302 28084 62354
rect 26908 61796 26964 61806
rect 26908 61682 26964 61740
rect 26908 61630 26910 61682
rect 26962 61630 26964 61682
rect 26908 61618 26964 61630
rect 27580 61012 27636 62132
rect 26796 60956 26964 61012
rect 26684 60834 26740 60844
rect 26572 60786 26628 60798
rect 26572 60734 26574 60786
rect 26626 60734 26628 60786
rect 26236 60676 26292 60686
rect 26572 60676 26628 60734
rect 26796 60786 26852 60798
rect 26796 60734 26798 60786
rect 26850 60734 26852 60786
rect 26236 60674 26628 60676
rect 26236 60622 26238 60674
rect 26290 60622 26628 60674
rect 26236 60620 26628 60622
rect 26684 60674 26740 60686
rect 26684 60622 26686 60674
rect 26738 60622 26740 60674
rect 26236 59444 26292 60620
rect 26684 60452 26740 60622
rect 26460 60396 26740 60452
rect 26236 59378 26292 59388
rect 26348 60116 26404 60126
rect 26236 59220 26292 59230
rect 26236 59126 26292 59164
rect 26236 57764 26292 57774
rect 26236 57670 26292 57708
rect 26348 57428 26404 60060
rect 26460 59330 26516 60396
rect 26460 59278 26462 59330
rect 26514 59278 26516 59330
rect 26460 59266 26516 59278
rect 26684 60228 26740 60238
rect 26572 59220 26628 59230
rect 26460 57652 26516 57662
rect 26460 57558 26516 57596
rect 25900 55692 26180 55748
rect 26236 57372 26404 57428
rect 26460 57428 26516 57438
rect 25564 55300 25620 55310
rect 25564 55206 25620 55244
rect 25788 55188 25844 55198
rect 25788 55094 25844 55132
rect 25452 55022 25454 55074
rect 25506 55022 25508 55074
rect 25452 55010 25508 55022
rect 25340 54674 25396 54684
rect 25788 54852 25844 54862
rect 25788 54738 25844 54796
rect 25788 54686 25790 54738
rect 25842 54686 25844 54738
rect 25788 54674 25844 54686
rect 25676 54628 25732 54638
rect 25340 54404 25396 54414
rect 25340 54310 25396 54348
rect 25116 54238 25118 54290
rect 25170 54238 25172 54290
rect 25116 54226 25172 54238
rect 25452 54290 25508 54302
rect 25452 54238 25454 54290
rect 25506 54238 25508 54290
rect 25026 54124 25290 54134
rect 25082 54068 25130 54124
rect 25186 54068 25234 54124
rect 25026 54058 25290 54068
rect 23884 53006 23886 53058
rect 23938 53006 23940 53058
rect 23884 52994 23940 53006
rect 24668 53116 24948 53172
rect 25116 53506 25172 53518
rect 25116 53454 25118 53506
rect 25170 53454 25172 53506
rect 25116 53172 25172 53454
rect 23660 52948 23716 52958
rect 24556 52948 24612 52958
rect 23716 52892 23828 52948
rect 23660 52882 23716 52892
rect 23772 52276 23828 52892
rect 24556 52854 24612 52892
rect 24332 52388 24388 52398
rect 23884 52276 23940 52286
rect 23772 52274 23940 52276
rect 23772 52222 23886 52274
rect 23938 52222 23940 52274
rect 23772 52220 23940 52222
rect 23884 52210 23940 52220
rect 24332 52274 24388 52332
rect 24332 52222 24334 52274
rect 24386 52222 24388 52274
rect 24332 52210 24388 52222
rect 23996 52164 24052 52174
rect 23548 52108 23828 52164
rect 23436 51940 23492 51950
rect 23436 51846 23492 51884
rect 23212 51604 23268 51614
rect 22988 51602 23268 51604
rect 22988 51550 23214 51602
rect 23266 51550 23268 51602
rect 22988 51548 23268 51550
rect 23212 51538 23268 51548
rect 23324 51490 23380 51502
rect 23324 51438 23326 51490
rect 23378 51438 23380 51490
rect 22988 51380 23044 51390
rect 22988 51266 23044 51324
rect 23212 51268 23268 51278
rect 22988 51214 22990 51266
rect 23042 51214 23044 51266
rect 22988 51202 23044 51214
rect 23100 51212 23212 51268
rect 22764 47506 22820 47516
rect 22876 50820 22932 50830
rect 22652 46162 22708 46172
rect 22764 47348 22820 47358
rect 22876 47348 22932 50764
rect 22764 47346 22932 47348
rect 22764 47294 22766 47346
rect 22818 47294 22932 47346
rect 22764 47292 22932 47294
rect 22988 49252 23044 49262
rect 22764 46116 22820 47292
rect 22876 46900 22932 46910
rect 22988 46900 23044 49196
rect 22876 46898 23044 46900
rect 22876 46846 22878 46898
rect 22930 46846 23044 46898
rect 22876 46844 23044 46846
rect 22876 46834 22932 46844
rect 22988 46788 23044 46844
rect 23100 46900 23156 51212
rect 23212 51202 23268 51212
rect 23324 50932 23380 51438
rect 23548 51380 23604 51390
rect 23548 51286 23604 51324
rect 23212 50876 23380 50932
rect 23436 50932 23492 50942
rect 23212 47124 23268 50876
rect 23436 50428 23492 50876
rect 23324 50372 23492 50428
rect 23324 48914 23380 50372
rect 23436 49700 23492 49710
rect 23436 49138 23492 49644
rect 23436 49086 23438 49138
rect 23490 49086 23492 49138
rect 23436 49074 23492 49086
rect 23660 49028 23716 49038
rect 23660 48934 23716 48972
rect 23324 48862 23326 48914
rect 23378 48862 23380 48914
rect 23324 48356 23380 48862
rect 23324 48300 23716 48356
rect 23212 47058 23268 47068
rect 23324 48130 23380 48142
rect 23324 48078 23326 48130
rect 23378 48078 23380 48130
rect 23324 47348 23380 48078
rect 23436 48130 23492 48142
rect 23436 48078 23438 48130
rect 23490 48078 23492 48130
rect 23436 47572 23492 48078
rect 23436 47506 23492 47516
rect 23548 47460 23604 47470
rect 23548 47366 23604 47404
rect 23324 47012 23380 47292
rect 23324 46956 23604 47012
rect 23100 46834 23156 46844
rect 22988 46722 23044 46732
rect 23100 46676 23156 46686
rect 23100 46582 23156 46620
rect 23324 46674 23380 46686
rect 23324 46622 23326 46674
rect 23378 46622 23380 46674
rect 22764 46050 22820 46060
rect 23212 46562 23268 46574
rect 23212 46510 23214 46562
rect 23266 46510 23268 46562
rect 23212 45892 23268 46510
rect 23324 46564 23380 46622
rect 23324 46498 23380 46508
rect 23548 46340 23604 46956
rect 22652 45836 23268 45892
rect 23324 46284 23604 46340
rect 22652 45218 22708 45836
rect 22652 45166 22654 45218
rect 22706 45166 22708 45218
rect 22652 45154 22708 45166
rect 23100 45668 23156 45678
rect 22988 44324 23044 44334
rect 22764 44212 22820 44222
rect 22540 43596 22708 43652
rect 22540 43426 22596 43438
rect 22540 43374 22542 43426
rect 22594 43374 22596 43426
rect 22540 43316 22596 43374
rect 22540 43250 22596 43260
rect 22540 42756 22596 42766
rect 22540 42082 22596 42700
rect 22540 42030 22542 42082
rect 22594 42030 22596 42082
rect 22540 42018 22596 42030
rect 22652 41748 22708 43596
rect 22428 41358 22430 41410
rect 22482 41358 22484 41410
rect 22428 41346 22484 41358
rect 22540 41692 22708 41748
rect 22316 41132 22484 41188
rect 22316 40964 22372 40974
rect 22316 40870 22372 40908
rect 21420 40628 21476 40796
rect 21624 40796 21888 40806
rect 21980 40796 22148 40852
rect 21680 40740 21728 40796
rect 21784 40740 21832 40796
rect 21624 40730 21888 40740
rect 21532 40628 21588 40638
rect 21420 40626 21588 40628
rect 21420 40574 21534 40626
rect 21586 40574 21588 40626
rect 21420 40572 21588 40574
rect 21532 40562 21588 40572
rect 21980 40516 22036 40526
rect 21980 40422 22036 40460
rect 21308 39330 21364 39340
rect 21420 39394 21476 39406
rect 21420 39342 21422 39394
rect 21474 39342 21476 39394
rect 21420 39284 21476 39342
rect 21868 39396 21924 39434
rect 21868 39330 21924 39340
rect 21420 39218 21476 39228
rect 21624 39228 21888 39238
rect 21680 39172 21728 39228
rect 21784 39172 21832 39228
rect 21624 39162 21888 39172
rect 21756 38836 21812 38846
rect 21308 38722 21364 38734
rect 21308 38670 21310 38722
rect 21362 38670 21364 38722
rect 21308 38668 21364 38670
rect 21308 38612 21588 38668
rect 21196 38434 21252 38444
rect 21084 38220 21252 38276
rect 20748 38110 20750 38162
rect 20802 38110 20804 38162
rect 19852 36260 19908 37436
rect 20076 37380 20132 37390
rect 19964 36932 20020 36942
rect 20076 36932 20132 37324
rect 20020 36876 20132 36932
rect 19964 36594 20020 36876
rect 19964 36542 19966 36594
rect 20018 36542 20020 36594
rect 19964 36530 20020 36542
rect 20300 36260 20356 37548
rect 20524 37604 20580 37614
rect 20412 37380 20468 37390
rect 20412 37286 20468 37324
rect 20412 36260 20468 36270
rect 20300 36258 20468 36260
rect 20300 36206 20414 36258
rect 20466 36206 20468 36258
rect 20300 36204 20468 36206
rect 19628 34914 19684 34926
rect 19628 34862 19630 34914
rect 19682 34862 19684 34914
rect 19628 34356 19684 34862
rect 19740 34802 19796 34814
rect 19740 34750 19742 34802
rect 19794 34750 19796 34802
rect 19740 34580 19796 34750
rect 19852 34692 19908 36204
rect 20300 35588 20356 35598
rect 20300 35494 20356 35532
rect 20188 34916 20244 34954
rect 20188 34850 20244 34860
rect 19852 34626 19908 34636
rect 20076 34802 20132 34814
rect 20076 34750 20078 34802
rect 20130 34750 20132 34802
rect 19740 34514 19796 34524
rect 19964 34356 20020 34366
rect 19628 34354 20020 34356
rect 19628 34302 19966 34354
rect 20018 34302 20020 34354
rect 19628 34300 20020 34302
rect 19964 34290 20020 34300
rect 20076 34356 20132 34750
rect 20076 34290 20132 34300
rect 20188 34692 20244 34702
rect 20188 34354 20244 34636
rect 20188 34302 20190 34354
rect 20242 34302 20244 34354
rect 20188 34290 20244 34302
rect 19628 34132 19684 34142
rect 19516 34130 19684 34132
rect 19516 34078 19630 34130
rect 19682 34078 19684 34130
rect 19516 34076 19684 34078
rect 19628 34066 19684 34076
rect 19852 34132 19908 34142
rect 19852 34038 19908 34076
rect 20076 34130 20132 34142
rect 20076 34078 20078 34130
rect 20130 34078 20132 34130
rect 20076 33796 20132 34078
rect 20076 33740 20244 33796
rect 19964 33684 20020 33694
rect 20020 33628 20132 33684
rect 19964 33618 20020 33628
rect 20076 33346 20132 33628
rect 20188 33572 20244 33740
rect 20188 33506 20244 33516
rect 20076 33294 20078 33346
rect 20130 33294 20132 33346
rect 20076 33282 20132 33294
rect 20188 33348 20244 33386
rect 20188 33282 20244 33292
rect 19516 33122 19572 33134
rect 19516 33070 19518 33122
rect 19570 33070 19572 33122
rect 19516 32564 19572 33070
rect 19964 33122 20020 33134
rect 19964 33070 19966 33122
rect 20018 33070 20020 33122
rect 19964 33012 20020 33070
rect 19964 32946 20020 32956
rect 20188 33124 20244 33134
rect 20188 32786 20244 33068
rect 20188 32734 20190 32786
rect 20242 32734 20244 32786
rect 20188 32722 20244 32734
rect 20300 33122 20356 33134
rect 20300 33070 20302 33122
rect 20354 33070 20356 33122
rect 19516 32470 19572 32508
rect 19964 32562 20020 32574
rect 19964 32510 19966 32562
rect 20018 32510 20020 32562
rect 19964 32452 20020 32510
rect 19964 32386 20020 32396
rect 20076 32562 20132 32574
rect 20076 32510 20078 32562
rect 20130 32510 20132 32562
rect 19404 32060 20020 32116
rect 19292 31892 19684 31948
rect 19404 31780 19460 31790
rect 19404 31686 19460 31724
rect 19516 31668 19572 31678
rect 19516 31574 19572 31612
rect 19180 31266 19236 31276
rect 19068 31166 19070 31218
rect 19122 31166 19124 31218
rect 19068 31154 19124 31166
rect 19516 31220 19572 31230
rect 19516 31126 19572 31164
rect 18956 31042 19012 31052
rect 19068 30996 19124 31006
rect 19628 30996 19684 31892
rect 19852 31332 19908 31342
rect 19852 31106 19908 31276
rect 19852 31054 19854 31106
rect 19906 31054 19908 31106
rect 19852 31042 19908 31054
rect 19124 30940 19236 30996
rect 19068 30930 19124 30940
rect 18844 30382 18846 30434
rect 18898 30382 18900 30434
rect 18844 30370 18900 30382
rect 19068 30434 19124 30446
rect 19068 30382 19070 30434
rect 19122 30382 19124 30434
rect 18844 30212 18900 30222
rect 18732 30210 18900 30212
rect 18732 30158 18846 30210
rect 18898 30158 18900 30210
rect 18732 30156 18900 30158
rect 18844 30146 18900 30156
rect 18844 29428 18900 29438
rect 18844 29426 19012 29428
rect 18844 29374 18846 29426
rect 18898 29374 19012 29426
rect 18844 29372 19012 29374
rect 18844 29362 18900 29372
rect 18508 29204 18564 29242
rect 18508 29138 18564 29148
rect 18844 29202 18900 29214
rect 18844 29150 18846 29202
rect 18898 29150 18900 29202
rect 18222 29036 18486 29046
rect 18278 28980 18326 29036
rect 18382 28980 18430 29036
rect 18222 28970 18486 28980
rect 17836 27918 17838 27970
rect 17890 27918 17892 27970
rect 17836 27906 17892 27918
rect 17948 27916 18116 27972
rect 18396 28756 18452 28766
rect 17388 27570 17444 27580
rect 17612 27858 17668 27870
rect 17612 27806 17614 27858
rect 17666 27806 17668 27858
rect 17612 27412 17668 27806
rect 16380 26852 16436 26862
rect 16380 26514 16436 26796
rect 16380 26462 16382 26514
rect 16434 26462 16436 26514
rect 16380 26450 16436 26462
rect 17052 26852 17220 26908
rect 17388 27356 17668 27412
rect 17724 27524 17780 27534
rect 17388 27076 17444 27356
rect 15820 26014 15822 26066
rect 15874 26014 15876 26066
rect 15820 26002 15876 26014
rect 16716 26180 16772 26190
rect 16716 25618 16772 26124
rect 16716 25566 16718 25618
rect 16770 25566 16772 25618
rect 16716 25554 16772 25566
rect 16828 26180 16884 26190
rect 17052 26180 17108 26852
rect 17388 26404 17444 27020
rect 17388 26310 17444 26348
rect 17612 26290 17668 26302
rect 17612 26238 17614 26290
rect 17666 26238 17668 26290
rect 17500 26180 17556 26190
rect 16828 26178 17332 26180
rect 16828 26126 16830 26178
rect 16882 26126 17332 26178
rect 16828 26124 17332 26126
rect 16044 25506 16100 25518
rect 16044 25454 16046 25506
rect 16098 25454 16100 25506
rect 16044 25284 16100 25454
rect 15708 24948 15764 24958
rect 15596 24892 15708 24948
rect 15708 24854 15764 24892
rect 15932 24612 15988 24622
rect 15820 24610 15988 24612
rect 15820 24558 15934 24610
rect 15986 24558 15988 24610
rect 15820 24556 15988 24558
rect 15820 24162 15876 24556
rect 15932 24546 15988 24556
rect 15820 24110 15822 24162
rect 15874 24110 15876 24162
rect 15820 24098 15876 24110
rect 15484 22866 15540 22876
rect 15708 23828 15764 23838
rect 15260 22754 15316 22764
rect 15596 22820 15652 22830
rect 15596 22484 15652 22764
rect 15708 22708 15764 23772
rect 15708 22642 15764 22652
rect 15820 23714 15876 23726
rect 15820 23662 15822 23714
rect 15874 23662 15876 23714
rect 15820 23156 15876 23662
rect 15708 22484 15764 22494
rect 15596 22482 15764 22484
rect 15596 22430 15710 22482
rect 15762 22430 15764 22482
rect 15596 22428 15764 22430
rect 15708 22418 15764 22428
rect 15820 22370 15876 23100
rect 16044 22932 16100 25228
rect 16268 24948 16324 24958
rect 16268 24834 16324 24892
rect 16268 24782 16270 24834
rect 16322 24782 16324 24834
rect 16268 24770 16324 24782
rect 16156 24722 16212 24734
rect 16156 24670 16158 24722
rect 16210 24670 16212 24722
rect 16156 24164 16212 24670
rect 16604 24722 16660 24734
rect 16604 24670 16606 24722
rect 16658 24670 16660 24722
rect 16156 24098 16212 24108
rect 16268 24612 16324 24622
rect 16268 23826 16324 24556
rect 16604 24162 16660 24670
rect 16604 24110 16606 24162
rect 16658 24110 16660 24162
rect 16604 24098 16660 24110
rect 16716 23940 16772 23950
rect 16716 23846 16772 23884
rect 16268 23774 16270 23826
rect 16322 23774 16324 23826
rect 16268 23762 16324 23774
rect 16604 23828 16660 23838
rect 16492 23714 16548 23726
rect 16492 23662 16494 23714
rect 16546 23662 16548 23714
rect 16380 23156 16436 23166
rect 16380 23042 16436 23100
rect 16380 22990 16382 23042
rect 16434 22990 16436 23042
rect 16380 22978 16436 22990
rect 15820 22318 15822 22370
rect 15874 22318 15876 22370
rect 15820 22306 15876 22318
rect 15932 22876 16100 22932
rect 15148 22082 15204 22092
rect 15596 22148 15652 22158
rect 15596 22054 15652 22092
rect 14820 21980 15084 21990
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 14820 21914 15084 21924
rect 15148 21700 15204 21710
rect 15036 21476 15092 21486
rect 15036 21382 15092 21420
rect 14700 20972 14980 21028
rect 14924 20914 14980 20972
rect 14924 20862 14926 20914
rect 14978 20862 14980 20914
rect 14924 20850 14980 20862
rect 14820 20412 15084 20422
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 14820 20346 15084 20356
rect 13972 20076 14196 20132
rect 13916 20066 13972 20076
rect 12908 19346 13412 19348
rect 12908 19294 12910 19346
rect 12962 19294 13412 19346
rect 12908 19292 13412 19294
rect 12908 19282 12964 19292
rect 13356 19234 13412 19292
rect 13356 19182 13358 19234
rect 13410 19182 13412 19234
rect 13356 19170 13412 19182
rect 13804 19236 13860 19246
rect 13804 19142 13860 19180
rect 13916 19234 13972 19246
rect 13916 19182 13918 19234
rect 13970 19182 13972 19234
rect 12684 17838 12686 17890
rect 12738 17838 12740 17890
rect 12684 17826 12740 17838
rect 12796 19012 12852 19022
rect 12628 17612 12740 17668
rect 12572 17602 12628 17612
rect 12124 16830 12126 16882
rect 12178 16830 12180 16882
rect 12124 16324 12180 16830
rect 12124 16258 12180 16268
rect 12348 17556 12404 17566
rect 12348 16100 12404 17500
rect 12460 17444 12516 17454
rect 12460 17350 12516 17388
rect 12572 16100 12628 16110
rect 11676 12908 11844 12964
rect 11900 15092 12068 15148
rect 12236 16098 12628 16100
rect 12236 16046 12574 16098
rect 12626 16046 12628 16098
rect 12236 16044 12628 16046
rect 12236 15148 12292 16044
rect 12572 16034 12628 16044
rect 12348 15874 12404 15886
rect 12348 15822 12350 15874
rect 12402 15822 12404 15874
rect 12348 15764 12404 15822
rect 12460 15876 12516 15886
rect 12460 15782 12516 15820
rect 12348 15698 12404 15708
rect 12684 15652 12740 17612
rect 12796 16994 12852 18956
rect 13580 19012 13636 19022
rect 13580 18918 13636 18956
rect 13580 18452 13636 18462
rect 13580 18338 13636 18396
rect 13580 18286 13582 18338
rect 13634 18286 13636 18338
rect 12796 16942 12798 16994
rect 12850 16942 12852 16994
rect 12796 16930 12852 16942
rect 12908 17890 12964 17902
rect 12908 17838 12910 17890
rect 12962 17838 12964 17890
rect 12908 17778 12964 17838
rect 12908 17726 12910 17778
rect 12962 17726 12964 17778
rect 12908 17332 12964 17726
rect 12796 16100 12852 16110
rect 12796 15986 12852 16044
rect 12796 15934 12798 15986
rect 12850 15934 12852 15986
rect 12796 15876 12852 15934
rect 12796 15810 12852 15820
rect 12460 15596 12740 15652
rect 12460 15202 12516 15596
rect 12460 15150 12462 15202
rect 12514 15150 12516 15202
rect 12236 15092 12404 15148
rect 12460 15138 12516 15150
rect 12908 15148 12964 17276
rect 13580 16322 13636 18286
rect 13580 16270 13582 16322
rect 13634 16270 13636 16322
rect 13580 16258 13636 16270
rect 13692 18004 13748 18014
rect 13692 16100 13748 17948
rect 13916 17778 13972 19182
rect 13916 17726 13918 17778
rect 13970 17726 13972 17778
rect 13916 17714 13972 17726
rect 14028 19124 14084 19134
rect 14028 17668 14084 19068
rect 14028 17574 14084 17612
rect 13804 17554 13860 17566
rect 13804 17502 13806 17554
rect 13858 17502 13860 17554
rect 13804 16212 13860 17502
rect 14140 16660 14196 20076
rect 14476 20076 14644 20132
rect 14252 17442 14308 17454
rect 14252 17390 14254 17442
rect 14306 17390 14308 17442
rect 14252 17332 14308 17390
rect 14252 16884 14308 17276
rect 14252 16818 14308 16828
rect 14140 16604 14308 16660
rect 13804 16146 13860 16156
rect 14140 16322 14196 16334
rect 14140 16270 14142 16322
rect 14194 16270 14196 16322
rect 14140 16210 14196 16270
rect 14140 16158 14142 16210
rect 14194 16158 14196 16210
rect 13580 16044 13748 16100
rect 13020 15764 13076 15774
rect 13020 15540 13076 15708
rect 13356 15540 13412 15550
rect 13020 15538 13356 15540
rect 13020 15486 13022 15538
rect 13074 15486 13356 15538
rect 13020 15484 13356 15486
rect 13020 15474 13076 15484
rect 13356 15446 13412 15484
rect 13580 15538 13636 16044
rect 13580 15486 13582 15538
rect 13634 15486 13636 15538
rect 11452 12852 11508 12862
rect 11452 12402 11508 12796
rect 11676 12516 11732 12908
rect 11788 12740 11844 12750
rect 11788 12646 11844 12684
rect 11676 12460 11844 12516
rect 11452 12350 11454 12402
rect 11506 12350 11508 12402
rect 11452 12338 11508 12350
rect 11004 12292 11060 12302
rect 11004 12198 11060 12236
rect 11418 11788 11682 11798
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11418 11722 11682 11732
rect 11228 11284 11284 11294
rect 11228 11190 11284 11228
rect 10780 10610 10836 10780
rect 11676 11172 11732 11182
rect 11676 10834 11732 11116
rect 11788 10948 11844 12460
rect 11900 11620 11956 15092
rect 12348 14868 12404 15092
rect 12796 15092 12964 15148
rect 13468 15202 13524 15214
rect 13468 15150 13470 15202
rect 13522 15150 13524 15202
rect 12348 14812 12740 14868
rect 12684 14642 12740 14812
rect 12684 14590 12686 14642
rect 12738 14590 12740 14642
rect 12684 14578 12740 14590
rect 12012 14308 12068 14318
rect 12012 13746 12068 14252
rect 12012 13694 12014 13746
rect 12066 13694 12068 13746
rect 12012 13186 12068 13694
rect 12684 13634 12740 13646
rect 12684 13582 12686 13634
rect 12738 13582 12740 13634
rect 12684 13412 12740 13582
rect 12684 13346 12740 13356
rect 12012 13134 12014 13186
rect 12066 13134 12068 13186
rect 12012 13122 12068 13134
rect 12236 13188 12292 13198
rect 12124 13076 12180 13086
rect 12012 12404 12068 12414
rect 12124 12404 12180 13020
rect 12236 13076 12292 13132
rect 12684 13186 12740 13198
rect 12684 13134 12686 13186
rect 12738 13134 12740 13186
rect 12236 13074 12404 13076
rect 12236 13022 12238 13074
rect 12290 13022 12404 13074
rect 12236 13020 12404 13022
rect 12236 13010 12292 13020
rect 12012 12402 12180 12404
rect 12012 12350 12014 12402
rect 12066 12350 12180 12402
rect 12012 12348 12180 12350
rect 12012 12338 12068 12348
rect 11900 11554 11956 11564
rect 11788 10882 11844 10892
rect 11900 11396 11956 11406
rect 11676 10782 11678 10834
rect 11730 10782 11732 10834
rect 11676 10770 11732 10782
rect 11900 10834 11956 11340
rect 11900 10782 11902 10834
rect 11954 10782 11956 10834
rect 11900 10770 11956 10782
rect 12012 11170 12068 11182
rect 12012 11118 12014 11170
rect 12066 11118 12068 11170
rect 12012 10836 12068 11118
rect 12124 10836 12180 10846
rect 12012 10780 12124 10836
rect 12124 10742 12180 10780
rect 10780 10558 10782 10610
rect 10834 10558 10836 10610
rect 10780 10546 10836 10558
rect 11116 10612 11172 10622
rect 11116 10518 11172 10556
rect 11788 10612 11844 10622
rect 11788 10518 11844 10556
rect 10668 10498 10724 10510
rect 10668 10446 10670 10498
rect 10722 10446 10724 10498
rect 10668 10052 10724 10446
rect 11418 10220 11682 10230
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11418 10154 11682 10164
rect 10444 9996 10724 10052
rect 10444 9938 10500 9996
rect 10444 9886 10446 9938
rect 10498 9886 10500 9938
rect 10444 9874 10500 9886
rect 9772 9828 9828 9838
rect 9772 9734 9828 9772
rect 9212 9550 9214 9602
rect 9266 9550 9268 9602
rect 6524 9044 6580 9054
rect 6412 9042 6580 9044
rect 6412 8990 6526 9042
rect 6578 8990 6580 9042
rect 6412 8988 6580 8990
rect 6524 8978 6580 8988
rect 6636 9042 6692 9054
rect 6636 8990 6638 9042
rect 6690 8990 6692 9042
rect 6300 8484 6356 8494
rect 6636 8484 6692 8990
rect 7756 9042 7812 9054
rect 7756 8990 7758 9042
rect 7810 8990 7812 9042
rect 6860 8484 6916 8494
rect 6356 8428 6804 8484
rect 6300 8418 6356 8428
rect 5516 7494 5572 7532
rect 5852 6914 5908 7532
rect 6188 7474 6244 7644
rect 6188 7422 6190 7474
rect 6242 7422 6244 7474
rect 6188 7410 6244 7422
rect 6300 8146 6356 8158
rect 6300 8094 6302 8146
rect 6354 8094 6356 8146
rect 5852 6862 5854 6914
rect 5906 6862 5908 6914
rect 5852 6802 5908 6862
rect 6300 6914 6356 8094
rect 6300 6862 6302 6914
rect 6354 6862 6356 6914
rect 6300 6850 6356 6862
rect 5852 6750 5854 6802
rect 5906 6750 5908 6802
rect 5852 6738 5908 6750
rect 6188 6692 6244 6702
rect 6412 6692 6468 8428
rect 6636 8258 6692 8270
rect 6636 8206 6638 8258
rect 6690 8206 6692 8258
rect 6636 8148 6692 8206
rect 6748 8260 6804 8428
rect 6860 8482 7028 8484
rect 6860 8430 6862 8482
rect 6914 8430 7028 8482
rect 6860 8428 7028 8430
rect 6860 8418 6916 8428
rect 6972 8372 7028 8428
rect 7532 8372 7588 8382
rect 6972 8370 7588 8372
rect 6972 8318 7534 8370
rect 7586 8318 7588 8370
rect 6972 8316 7588 8318
rect 7532 8306 7588 8316
rect 6860 8260 6916 8270
rect 6748 8258 6916 8260
rect 6748 8206 6862 8258
rect 6914 8206 6916 8258
rect 6748 8204 6916 8206
rect 6860 8194 6916 8204
rect 6636 8082 6692 8092
rect 7420 8146 7476 8158
rect 7420 8094 7422 8146
rect 7474 8094 7476 8146
rect 6748 8036 6804 8046
rect 6748 8034 6916 8036
rect 6748 7982 6750 8034
rect 6802 7982 6916 8034
rect 6748 7980 6916 7982
rect 6748 7970 6804 7980
rect 6860 7586 6916 7980
rect 7420 7924 7476 8094
rect 7420 7858 7476 7868
rect 7644 8036 7700 8046
rect 7756 8036 7812 8990
rect 8092 8148 8148 8158
rect 8092 8054 8148 8092
rect 8204 8146 8260 8158
rect 8204 8094 8206 8146
rect 8258 8094 8260 8146
rect 7644 8034 7812 8036
rect 7644 7982 7646 8034
rect 7698 7982 7812 8034
rect 7644 7980 7812 7982
rect 8204 8036 8260 8094
rect 8652 8036 8708 8046
rect 8204 8034 8708 8036
rect 8204 7982 8654 8034
rect 8706 7982 8708 8034
rect 8204 7980 8708 7982
rect 6860 7534 6862 7586
rect 6914 7534 6916 7586
rect 6860 7522 6916 7534
rect 6636 6914 6692 6926
rect 6636 6862 6638 6914
rect 6690 6862 6692 6914
rect 6636 6802 6692 6862
rect 6636 6750 6638 6802
rect 6690 6750 6692 6802
rect 6636 6738 6692 6750
rect 4844 6638 4846 6690
rect 4898 6638 4900 6690
rect 4844 6626 4900 6638
rect 5180 6636 5404 6692
rect 3836 6466 4004 6468
rect 3836 6414 3838 6466
rect 3890 6414 4004 6466
rect 3836 6412 4004 6414
rect 4060 6580 4116 6590
rect 3836 6132 3892 6412
rect 3836 6066 3892 6076
rect 3388 3332 3556 3388
rect 2940 2770 2996 2782
rect 2940 2718 2942 2770
rect 2994 2718 2996 2770
rect 1932 1988 1988 1998
rect 2716 1988 2772 1998
rect 1932 1986 2772 1988
rect 1932 1934 1934 1986
rect 1986 1934 2718 1986
rect 2770 1934 2772 1986
rect 1932 1932 2772 1934
rect 1932 1922 1988 1932
rect 2380 1764 2436 1774
rect 2380 1670 2436 1708
rect 2716 400 2772 1932
rect 2940 1874 2996 2718
rect 2940 1822 2942 1874
rect 2994 1822 2996 1874
rect 2940 1810 2996 1822
rect 3276 1876 3332 1886
rect 3276 1782 3332 1820
rect 3388 400 3444 3332
rect 4060 2658 4116 6524
rect 4396 6580 4452 6590
rect 4396 6486 4452 6524
rect 5180 6130 5236 6636
rect 5404 6626 5460 6636
rect 5964 6690 6468 6692
rect 5964 6638 6190 6690
rect 6242 6638 6468 6690
rect 5964 6636 6468 6638
rect 5180 6078 5182 6130
rect 5234 6078 5236 6130
rect 5180 6066 5236 6078
rect 5852 6132 5908 6142
rect 5964 6132 6020 6636
rect 6188 6626 6244 6636
rect 7644 6356 7700 7980
rect 8016 7868 8280 7878
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8016 7802 8280 7812
rect 8652 7588 8708 7980
rect 9212 7700 9268 9550
rect 12348 9268 12404 13020
rect 12684 13074 12740 13134
rect 12684 13022 12686 13074
rect 12738 13022 12740 13074
rect 12684 13010 12740 13022
rect 12572 11396 12628 11406
rect 12460 11172 12516 11182
rect 12460 11078 12516 11116
rect 12572 9938 12628 11340
rect 12796 10836 12852 15092
rect 13020 13188 13076 13198
rect 13020 13186 13300 13188
rect 13020 13134 13022 13186
rect 13074 13134 13300 13186
rect 13020 13132 13300 13134
rect 13020 13122 13076 13132
rect 13244 12402 13300 13132
rect 13468 12962 13524 15150
rect 13580 13748 13636 15486
rect 13692 15876 13748 15886
rect 13692 15540 13748 15820
rect 13804 15540 13860 15550
rect 13692 15538 13860 15540
rect 13692 15486 13806 15538
rect 13858 15486 13860 15538
rect 13692 15484 13860 15486
rect 13804 15474 13860 15484
rect 13692 14532 13748 14542
rect 14140 14532 14196 16158
rect 13692 14530 14196 14532
rect 13692 14478 13694 14530
rect 13746 14478 14196 14530
rect 13692 14476 14196 14478
rect 13692 14466 13748 14476
rect 14140 14308 14196 14476
rect 14140 14242 14196 14252
rect 14252 15426 14308 16604
rect 14252 15374 14254 15426
rect 14306 15374 14308 15426
rect 14252 13972 14308 15374
rect 14476 15314 14532 20076
rect 15148 19906 15204 21644
rect 15484 21474 15540 21486
rect 15484 21422 15486 21474
rect 15538 21422 15540 21474
rect 15148 19854 15150 19906
rect 15202 19854 15204 19906
rect 15148 19842 15204 19854
rect 15372 20578 15428 20590
rect 15372 20526 15374 20578
rect 15426 20526 15428 20578
rect 15372 19908 15428 20526
rect 15484 20132 15540 21422
rect 15484 20066 15540 20076
rect 15708 20916 15764 20926
rect 15708 20130 15764 20860
rect 15708 20078 15710 20130
rect 15762 20078 15764 20130
rect 15708 20066 15764 20078
rect 15820 20804 15876 20814
rect 15932 20804 15988 22876
rect 16044 22372 16100 22382
rect 16044 22258 16100 22316
rect 16044 22206 16046 22258
rect 16098 22206 16100 22258
rect 16044 22194 16100 22206
rect 16492 21700 16548 23662
rect 16604 22708 16660 23772
rect 16828 23268 16884 26124
rect 17276 25956 17332 26124
rect 17500 26086 17556 26124
rect 17612 25956 17668 26238
rect 17276 25900 17668 25956
rect 16940 25172 16996 25182
rect 16940 24946 16996 25116
rect 16940 24894 16942 24946
rect 16994 24894 16996 24946
rect 16940 24882 16996 24894
rect 17052 24612 17108 24622
rect 16940 24164 16996 24174
rect 16940 24070 16996 24108
rect 17052 23940 17108 24556
rect 17612 24610 17668 24622
rect 17612 24558 17614 24610
rect 17666 24558 17668 24610
rect 17612 24276 17668 24558
rect 16716 23212 16884 23268
rect 16940 23884 17108 23940
rect 17388 24220 17668 24276
rect 16716 22820 16772 23212
rect 16828 23044 16884 23054
rect 16828 22950 16884 22988
rect 16716 22764 16884 22820
rect 16604 22652 16772 22708
rect 16604 22484 16660 22494
rect 16604 22390 16660 22428
rect 16492 21634 16548 21644
rect 15820 20802 15988 20804
rect 15820 20750 15822 20802
rect 15874 20750 15988 20802
rect 15820 20748 15988 20750
rect 16604 20916 16660 20926
rect 15372 19842 15428 19852
rect 15372 19348 15428 19358
rect 15372 19254 15428 19292
rect 14588 19234 14644 19246
rect 14588 19182 14590 19234
rect 14642 19182 14644 19234
rect 14588 18004 14644 19182
rect 15596 19124 15652 19134
rect 15596 19030 15652 19068
rect 14700 19010 14756 19022
rect 14700 18958 14702 19010
rect 14754 18958 14756 19010
rect 14700 18004 14756 18958
rect 15820 19012 15876 20748
rect 16492 20690 16548 20702
rect 16492 20638 16494 20690
rect 16546 20638 16548 20690
rect 16492 20242 16548 20638
rect 16492 20190 16494 20242
rect 16546 20190 16548 20242
rect 16492 20178 16548 20190
rect 16044 20132 16100 20142
rect 16044 20038 16100 20076
rect 16268 20020 16324 20030
rect 16268 19926 16324 19964
rect 16604 20018 16660 20860
rect 16604 19966 16606 20018
rect 16658 19966 16660 20018
rect 16604 19954 16660 19966
rect 16604 19794 16660 19806
rect 16604 19742 16606 19794
rect 16658 19742 16660 19794
rect 16604 19460 16660 19742
rect 16604 19394 16660 19404
rect 16044 19234 16100 19246
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 16044 19124 16100 19182
rect 16044 19058 16100 19068
rect 16492 19236 16548 19246
rect 16716 19236 16772 22652
rect 16492 19234 16772 19236
rect 16492 19182 16494 19234
rect 16546 19182 16772 19234
rect 16492 19180 16772 19182
rect 16492 19124 16548 19180
rect 16492 19058 16548 19068
rect 15820 18946 15876 18956
rect 14820 18844 15084 18854
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 14820 18778 15084 18788
rect 16268 18340 16324 18350
rect 15820 18228 15876 18238
rect 14700 17948 14980 18004
rect 14588 17938 14644 17948
rect 14588 17668 14644 17678
rect 14588 17108 14644 17612
rect 14924 17668 14980 17948
rect 15260 17780 15316 17790
rect 15260 17686 15316 17724
rect 14924 17574 14980 17612
rect 15372 17666 15428 17678
rect 15372 17614 15374 17666
rect 15426 17614 15428 17666
rect 14700 17556 14756 17566
rect 14700 17462 14756 17500
rect 15148 17444 15204 17454
rect 15148 17442 15316 17444
rect 15148 17390 15150 17442
rect 15202 17390 15316 17442
rect 15148 17388 15316 17390
rect 15148 17378 15204 17388
rect 14820 17276 15084 17286
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 14820 17210 15084 17220
rect 14588 17052 14980 17108
rect 14924 16770 14980 17052
rect 14924 16718 14926 16770
rect 14978 16718 14980 16770
rect 14924 16706 14980 16718
rect 15260 16658 15316 17388
rect 15372 17220 15428 17614
rect 15708 17668 15764 17678
rect 15820 17668 15876 18172
rect 15764 17612 15876 17668
rect 15708 17602 15764 17612
rect 15372 17154 15428 17164
rect 15484 17556 15540 17566
rect 15372 16884 15428 16894
rect 15484 16884 15540 17500
rect 15820 17108 15876 17612
rect 15932 17892 15988 17902
rect 15932 17666 15988 17836
rect 15932 17614 15934 17666
rect 15986 17614 15988 17666
rect 15932 17332 15988 17614
rect 16268 17556 16324 18284
rect 16828 18340 16884 22764
rect 16828 18274 16884 18284
rect 16940 18004 16996 23884
rect 17388 23828 17444 24220
rect 17612 23940 17668 23950
rect 17052 23716 17108 23726
rect 17276 23716 17332 23726
rect 17052 23622 17108 23660
rect 17164 23714 17332 23716
rect 17164 23662 17278 23714
rect 17330 23662 17332 23714
rect 17164 23660 17332 23662
rect 17052 22372 17108 22382
rect 17052 22278 17108 22316
rect 17052 20132 17108 20142
rect 17052 19346 17108 20076
rect 17052 19294 17054 19346
rect 17106 19294 17108 19346
rect 17052 19282 17108 19294
rect 16940 17938 16996 17948
rect 16940 17780 16996 17790
rect 16716 17778 16996 17780
rect 16716 17726 16942 17778
rect 16994 17726 16996 17778
rect 16716 17724 16996 17726
rect 16492 17668 16548 17678
rect 16716 17668 16772 17724
rect 16940 17714 16996 17724
rect 16492 17666 16772 17668
rect 16492 17614 16494 17666
rect 16546 17614 16772 17666
rect 16492 17612 16772 17614
rect 17052 17668 17108 17678
rect 17164 17668 17220 23660
rect 17276 23650 17332 23660
rect 17388 22820 17444 23772
rect 17500 23826 17556 23838
rect 17500 23774 17502 23826
rect 17554 23774 17556 23826
rect 17500 23044 17556 23774
rect 17612 23378 17668 23884
rect 17612 23326 17614 23378
rect 17666 23326 17668 23378
rect 17612 23314 17668 23326
rect 17612 23044 17668 23054
rect 17500 22988 17612 23044
rect 17612 22978 17668 22988
rect 17388 22754 17444 22764
rect 17500 22148 17556 22158
rect 17500 21812 17556 22092
rect 17724 22148 17780 27468
rect 17948 27298 18004 27916
rect 18172 27860 18228 27870
rect 17948 27246 17950 27298
rect 18002 27246 18004 27298
rect 17948 27234 18004 27246
rect 18060 27858 18228 27860
rect 18060 27806 18174 27858
rect 18226 27806 18228 27858
rect 18060 27804 18228 27806
rect 18060 27188 18116 27804
rect 18172 27794 18228 27804
rect 18172 27636 18228 27646
rect 18396 27636 18452 28700
rect 18844 28756 18900 29150
rect 18956 29204 19012 29372
rect 19068 29204 19124 30382
rect 18956 29202 19124 29204
rect 18956 29150 19070 29202
rect 19122 29150 19124 29202
rect 18956 29148 19124 29150
rect 19068 29138 19124 29148
rect 19180 28980 19236 30940
rect 19516 30940 19684 30996
rect 19292 29988 19348 30026
rect 19292 29922 19348 29932
rect 19292 29764 19348 29774
rect 19292 29316 19348 29708
rect 19292 29250 19348 29260
rect 18844 28690 18900 28700
rect 18956 28924 19236 28980
rect 19292 29092 19348 29102
rect 18172 27634 18452 27636
rect 18172 27582 18174 27634
rect 18226 27582 18452 27634
rect 18172 27580 18452 27582
rect 18844 27746 18900 27758
rect 18844 27694 18846 27746
rect 18898 27694 18900 27746
rect 18844 27636 18900 27694
rect 18172 27570 18228 27580
rect 18222 27468 18486 27478
rect 18278 27412 18326 27468
rect 18382 27412 18430 27468
rect 18222 27402 18486 27412
rect 18508 27298 18564 27310
rect 18508 27246 18510 27298
rect 18562 27246 18564 27298
rect 18172 27188 18228 27198
rect 18060 27132 18172 27188
rect 18172 27122 18228 27132
rect 18284 26964 18340 27002
rect 18284 26898 18340 26908
rect 18172 26852 18228 26862
rect 18172 26292 18228 26796
rect 17948 26290 18228 26292
rect 17948 26238 18174 26290
rect 18226 26238 18228 26290
rect 17948 26236 18228 26238
rect 17836 26068 17892 26078
rect 17836 25974 17892 26012
rect 17948 24836 18004 26236
rect 18172 26226 18228 26236
rect 18508 26292 18564 27246
rect 18620 27076 18676 27086
rect 18620 26982 18676 27020
rect 18844 26292 18900 27580
rect 18508 26290 18676 26292
rect 18508 26238 18510 26290
rect 18562 26238 18676 26290
rect 18508 26236 18676 26238
rect 18508 26226 18564 26236
rect 18508 26068 18564 26106
rect 18508 26002 18564 26012
rect 18222 25900 18486 25910
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18222 25834 18486 25844
rect 18620 25732 18676 26236
rect 18732 26236 18900 26292
rect 18732 25956 18788 26236
rect 18732 25890 18788 25900
rect 18844 26066 18900 26078
rect 18844 26014 18846 26066
rect 18898 26014 18900 26066
rect 18844 25844 18900 26014
rect 18844 25778 18900 25788
rect 18620 25676 18788 25732
rect 18732 25620 18788 25676
rect 18844 25620 18900 25630
rect 18732 25618 18900 25620
rect 18732 25566 18846 25618
rect 18898 25566 18900 25618
rect 18732 25564 18900 25566
rect 18844 25554 18900 25564
rect 17836 24780 18004 24836
rect 18620 25396 18676 25406
rect 17836 22484 17892 24780
rect 17948 24610 18004 24622
rect 17948 24558 17950 24610
rect 18002 24558 18004 24610
rect 17948 24500 18004 24558
rect 18396 24612 18452 24622
rect 18396 24518 18452 24556
rect 18004 24444 18116 24500
rect 17948 24434 18004 24444
rect 18060 24164 18116 24444
rect 18222 24332 18486 24342
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18222 24266 18486 24276
rect 18508 24164 18564 24174
rect 18060 24108 18452 24164
rect 17948 23826 18004 23838
rect 17948 23774 17950 23826
rect 18002 23774 18004 23826
rect 17948 23044 18004 23774
rect 18060 23828 18116 23838
rect 18060 23716 18116 23772
rect 18396 23826 18452 24108
rect 18508 24070 18564 24108
rect 18396 23774 18398 23826
rect 18450 23774 18452 23826
rect 18396 23762 18452 23774
rect 18172 23716 18228 23726
rect 18060 23714 18228 23716
rect 18060 23662 18174 23714
rect 18226 23662 18228 23714
rect 18060 23660 18228 23662
rect 18172 23650 18228 23660
rect 17948 22950 18004 22988
rect 18620 23042 18676 25340
rect 18732 24948 18788 24958
rect 18732 24854 18788 24892
rect 18956 24612 19012 28924
rect 19068 28644 19124 28654
rect 19068 27748 19124 28588
rect 19292 27748 19348 29036
rect 19068 27692 19236 27748
rect 19068 27188 19124 27198
rect 19068 27094 19124 27132
rect 19180 26964 19236 27692
rect 19292 27076 19348 27692
rect 19292 27010 19348 27020
rect 19516 27076 19572 30940
rect 19628 30772 19684 30782
rect 19628 29764 19684 30716
rect 19852 30212 19908 30222
rect 19852 30118 19908 30156
rect 19628 29698 19684 29708
rect 19852 29428 19908 29438
rect 19852 29334 19908 29372
rect 19628 29202 19684 29214
rect 19628 29150 19630 29202
rect 19682 29150 19684 29202
rect 19628 28756 19684 29150
rect 19740 28756 19796 28766
rect 19628 28754 19796 28756
rect 19628 28702 19742 28754
rect 19794 28702 19796 28754
rect 19628 28700 19796 28702
rect 19740 28690 19796 28700
rect 19516 27010 19572 27020
rect 19628 27972 19684 27982
rect 19628 27858 19684 27916
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19068 26908 19236 26964
rect 19628 26908 19684 27806
rect 19068 26852 19124 26908
rect 19628 26852 19796 26908
rect 19852 26852 19908 26862
rect 19068 26796 19236 26852
rect 19180 26740 19236 26796
rect 19740 26850 19908 26852
rect 19740 26798 19854 26850
rect 19906 26798 19908 26850
rect 19740 26796 19908 26798
rect 19740 26740 19796 26796
rect 19852 26786 19908 26796
rect 19180 26674 19236 26684
rect 19628 26684 19796 26740
rect 19292 26404 19348 26414
rect 19180 26402 19348 26404
rect 19180 26350 19294 26402
rect 19346 26350 19348 26402
rect 19180 26348 19348 26350
rect 19180 26292 19236 26348
rect 19292 26338 19348 26348
rect 19180 26226 19236 26236
rect 19628 26292 19684 26684
rect 19964 26628 20020 32060
rect 20076 27412 20132 32510
rect 20300 32564 20356 33070
rect 20300 32470 20356 32508
rect 20412 32004 20468 36204
rect 20524 33796 20580 37548
rect 20748 37268 20804 38110
rect 20860 37940 20916 37950
rect 20860 37492 20916 37884
rect 21084 37716 21140 37726
rect 21196 37716 21252 38220
rect 21532 38162 21588 38612
rect 21532 38110 21534 38162
rect 21586 38110 21588 38162
rect 21532 38098 21588 38110
rect 21756 38052 21812 38780
rect 21980 38724 22036 38734
rect 22092 38724 22148 40796
rect 22428 40626 22484 41132
rect 22428 40574 22430 40626
rect 22482 40574 22484 40626
rect 22428 40562 22484 40574
rect 22036 38668 22148 38724
rect 21980 38658 22036 38668
rect 21980 38332 22372 38388
rect 21980 38274 22036 38332
rect 21980 38222 21982 38274
rect 22034 38222 22036 38274
rect 21980 38210 22036 38222
rect 21756 37958 21812 37996
rect 22092 38050 22148 38062
rect 22092 37998 22094 38050
rect 22146 37998 22148 38050
rect 21420 37940 21476 37950
rect 21420 37846 21476 37884
rect 21980 37828 22036 37838
rect 21196 37660 21476 37716
rect 21084 37604 21140 37660
rect 21084 37548 21364 37604
rect 20860 37490 21252 37492
rect 20860 37438 20862 37490
rect 20914 37438 21252 37490
rect 20860 37436 21252 37438
rect 20860 37426 20916 37436
rect 20748 37212 21140 37268
rect 20860 35588 20916 35598
rect 20748 35586 20916 35588
rect 20748 35534 20862 35586
rect 20914 35534 20916 35586
rect 20748 35532 20916 35534
rect 20636 35252 20692 35262
rect 20636 34804 20692 35196
rect 20636 34710 20692 34748
rect 20748 34692 20804 35532
rect 20860 35522 20916 35532
rect 20748 34580 20804 34636
rect 20524 33730 20580 33740
rect 20636 34524 20804 34580
rect 20860 35364 20916 35374
rect 20636 33684 20692 34524
rect 20636 33618 20692 33628
rect 20748 34356 20804 34366
rect 20524 33236 20580 33246
rect 20524 33234 20692 33236
rect 20524 33182 20526 33234
rect 20578 33182 20692 33234
rect 20524 33180 20692 33182
rect 20524 33170 20580 33180
rect 20524 32562 20580 32574
rect 20524 32510 20526 32562
rect 20578 32510 20580 32562
rect 20524 32116 20580 32510
rect 20524 32050 20580 32060
rect 20412 31938 20468 31948
rect 20636 32004 20692 33180
rect 20748 33012 20804 34300
rect 20748 32946 20804 32956
rect 20636 31938 20692 31948
rect 20188 31780 20244 31790
rect 20188 31778 20468 31780
rect 20188 31726 20190 31778
rect 20242 31726 20468 31778
rect 20188 31724 20468 31726
rect 20188 31714 20244 31724
rect 20188 31444 20244 31454
rect 20244 31388 20356 31444
rect 20188 31378 20244 31388
rect 20188 30212 20244 30222
rect 20188 29988 20244 30156
rect 20188 29894 20244 29932
rect 20188 29538 20244 29550
rect 20188 29486 20190 29538
rect 20242 29486 20244 29538
rect 20188 28084 20244 29486
rect 20300 29428 20356 31388
rect 20412 30436 20468 31724
rect 20748 31778 20804 31790
rect 20748 31726 20750 31778
rect 20802 31726 20804 31778
rect 20636 31556 20692 31566
rect 20748 31556 20804 31726
rect 20692 31500 20804 31556
rect 20636 31490 20692 31500
rect 20636 30436 20692 30446
rect 20412 30434 20692 30436
rect 20412 30382 20638 30434
rect 20690 30382 20692 30434
rect 20412 30380 20692 30382
rect 20636 30370 20692 30380
rect 20748 30212 20804 30222
rect 20748 30118 20804 30156
rect 20636 29986 20692 29998
rect 20636 29934 20638 29986
rect 20690 29934 20692 29986
rect 20300 28642 20356 29372
rect 20412 29538 20468 29550
rect 20412 29486 20414 29538
rect 20466 29486 20468 29538
rect 20412 28866 20468 29486
rect 20412 28814 20414 28866
rect 20466 28814 20468 28866
rect 20412 28802 20468 28814
rect 20300 28590 20302 28642
rect 20354 28590 20356 28642
rect 20300 28578 20356 28590
rect 20524 28420 20580 28430
rect 20524 28326 20580 28364
rect 20188 28028 20580 28084
rect 20076 27346 20132 27356
rect 20412 27746 20468 27758
rect 20412 27694 20414 27746
rect 20466 27694 20468 27746
rect 20412 27300 20468 27694
rect 20300 27244 20468 27300
rect 20300 27186 20356 27244
rect 20300 27134 20302 27186
rect 20354 27134 20356 27186
rect 20300 27122 20356 27134
rect 19852 26572 20020 26628
rect 20076 27076 20132 27086
rect 19740 26404 19796 26414
rect 19740 26310 19796 26348
rect 18620 22990 18622 23042
rect 18674 22990 18676 23042
rect 18620 22930 18676 22990
rect 18620 22878 18622 22930
rect 18674 22878 18676 22930
rect 18620 22866 18676 22878
rect 18732 24556 19012 24612
rect 19180 26068 19236 26078
rect 18222 22764 18486 22774
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18222 22698 18486 22708
rect 18620 22484 18676 22494
rect 17892 22428 18004 22484
rect 17836 22418 17892 22428
rect 17724 22082 17780 22092
rect 17948 21812 18004 22428
rect 18620 22390 18676 22428
rect 18172 22148 18228 22158
rect 18172 22054 18228 22092
rect 17500 21756 17780 21812
rect 17612 21588 17668 21598
rect 17612 21494 17668 21532
rect 17612 20018 17668 20030
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 17500 19012 17556 19022
rect 17612 19012 17668 19966
rect 17500 19010 17668 19012
rect 17500 18958 17502 19010
rect 17554 18958 17668 19010
rect 17500 18956 17668 18958
rect 17500 18946 17556 18956
rect 17612 18452 17668 18956
rect 17612 18386 17668 18396
rect 17500 18338 17556 18350
rect 17500 18286 17502 18338
rect 17554 18286 17556 18338
rect 17500 18228 17556 18286
rect 17500 18162 17556 18172
rect 17052 17666 17220 17668
rect 17052 17614 17054 17666
rect 17106 17614 17220 17666
rect 17052 17612 17220 17614
rect 16492 17602 16548 17612
rect 17052 17602 17108 17612
rect 16268 17462 16324 17500
rect 16940 17556 16996 17566
rect 15932 17266 15988 17276
rect 16044 17442 16100 17454
rect 16044 17390 16046 17442
rect 16098 17390 16100 17442
rect 15932 17108 15988 17118
rect 15820 17106 15988 17108
rect 15820 17054 15934 17106
rect 15986 17054 15988 17106
rect 15820 17052 15988 17054
rect 15932 17042 15988 17052
rect 15372 16882 15540 16884
rect 15372 16830 15374 16882
rect 15426 16830 15540 16882
rect 15372 16828 15540 16830
rect 15372 16818 15428 16828
rect 15260 16606 15262 16658
rect 15314 16606 15316 16658
rect 14588 16212 14644 16222
rect 14588 15540 14644 16156
rect 15148 16212 15204 16222
rect 15148 16098 15204 16156
rect 15148 16046 15150 16098
rect 15202 16046 15204 16098
rect 15148 16034 15204 16046
rect 14820 15708 15084 15718
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 14820 15642 15084 15652
rect 15260 15540 15316 16606
rect 15372 15540 15428 15550
rect 14588 15484 15204 15540
rect 15260 15538 15428 15540
rect 15260 15486 15374 15538
rect 15426 15486 15428 15538
rect 15260 15484 15428 15486
rect 15148 15428 15204 15484
rect 15372 15474 15428 15484
rect 14476 15262 14478 15314
rect 14530 15262 14532 15314
rect 14364 15202 14420 15214
rect 14364 15150 14366 15202
rect 14418 15150 14420 15202
rect 14364 14642 14420 15150
rect 14476 15148 14532 15262
rect 14812 15316 14868 15326
rect 14812 15222 14868 15260
rect 15148 15314 15204 15372
rect 15148 15262 15150 15314
rect 15202 15262 15204 15314
rect 14476 15092 14644 15148
rect 14364 14590 14366 14642
rect 14418 14590 14420 14642
rect 14364 14578 14420 14590
rect 14588 14644 14644 15092
rect 14252 13906 14308 13916
rect 13804 13748 13860 13758
rect 13580 13692 13804 13748
rect 13804 13682 13860 13692
rect 13804 13412 13860 13422
rect 13468 12910 13470 12962
rect 13522 12910 13524 12962
rect 13468 12898 13524 12910
rect 13692 13188 13748 13198
rect 13692 12962 13748 13132
rect 13692 12910 13694 12962
rect 13746 12910 13748 12962
rect 13692 12898 13748 12910
rect 13580 12740 13636 12750
rect 13468 12684 13580 12740
rect 13244 12350 13246 12402
rect 13298 12350 13300 12402
rect 12908 11284 12964 11294
rect 12908 11190 12964 11228
rect 12796 10742 12852 10780
rect 12572 9886 12574 9938
rect 12626 9886 12628 9938
rect 12572 9874 12628 9886
rect 12796 9828 12852 9838
rect 13244 9828 13300 12350
rect 13356 12404 13412 12414
rect 13356 10500 13412 12348
rect 13468 11172 13524 12684
rect 13580 12674 13636 12684
rect 13804 12738 13860 13356
rect 14364 13186 14420 13198
rect 14364 13134 14366 13186
rect 14418 13134 14420 13186
rect 14140 13076 14196 13086
rect 14140 12962 14196 13020
rect 14140 12910 14142 12962
rect 14194 12910 14196 12962
rect 14140 12898 14196 12910
rect 13804 12686 13806 12738
rect 13858 12686 13860 12738
rect 13804 12674 13860 12686
rect 14364 12066 14420 13134
rect 14588 13074 14644 14588
rect 14820 14140 15084 14150
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 14820 14074 15084 14084
rect 15036 13972 15092 13982
rect 14924 13860 14980 13870
rect 14812 13748 14868 13758
rect 14812 13634 14868 13692
rect 14812 13582 14814 13634
rect 14866 13582 14868 13634
rect 14812 13570 14868 13582
rect 14588 13022 14590 13074
rect 14642 13022 14644 13074
rect 14588 13010 14644 13022
rect 14924 13076 14980 13804
rect 15036 13186 15092 13916
rect 15036 13134 15038 13186
rect 15090 13134 15092 13186
rect 15036 13122 15092 13134
rect 14924 12982 14980 13020
rect 14820 12572 15084 12582
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 14820 12506 15084 12516
rect 14364 12014 14366 12066
rect 14418 12014 14420 12066
rect 13468 10836 13524 11116
rect 13580 11732 13636 11742
rect 13580 11282 13636 11676
rect 14364 11732 14420 12014
rect 14364 11666 14420 11676
rect 14700 12404 14756 12414
rect 14476 11396 14532 11406
rect 14476 11302 14532 11340
rect 13580 11230 13582 11282
rect 13634 11230 13636 11282
rect 13580 11060 13636 11230
rect 13916 11284 13972 11294
rect 13916 11190 13972 11228
rect 14140 11284 14196 11294
rect 14588 11284 14644 11294
rect 14140 11282 14420 11284
rect 14140 11230 14142 11282
rect 14194 11230 14420 11282
rect 14140 11228 14420 11230
rect 14140 11218 14196 11228
rect 13580 10994 13636 11004
rect 13804 11170 13860 11182
rect 13804 11118 13806 11170
rect 13858 11118 13860 11170
rect 13804 10948 13860 11118
rect 14364 10948 14420 11228
rect 14588 11060 14644 11228
rect 14700 11282 14756 12348
rect 15148 12068 15204 15262
rect 15260 15316 15316 15326
rect 15260 15222 15316 15260
rect 15260 13972 15316 13982
rect 15260 13878 15316 13916
rect 15484 12180 15540 16828
rect 15596 16772 15652 16782
rect 15596 15540 15652 16716
rect 16044 16548 16100 17390
rect 16828 17442 16884 17454
rect 16828 17390 16830 17442
rect 16882 17390 16884 17442
rect 16716 17332 16772 17342
rect 16716 17106 16772 17276
rect 16716 17054 16718 17106
rect 16770 17054 16772 17106
rect 16716 17042 16772 17054
rect 15820 16492 16100 16548
rect 16268 16996 16324 17006
rect 15820 16210 15876 16492
rect 15820 16158 15822 16210
rect 15874 16158 15876 16210
rect 15820 16146 15876 16158
rect 16156 15540 16212 15550
rect 15596 15538 16212 15540
rect 15596 15486 15598 15538
rect 15650 15486 16158 15538
rect 16210 15486 16212 15538
rect 15596 15484 16212 15486
rect 15596 15474 15652 15484
rect 16156 15474 16212 15484
rect 15708 14308 15764 14318
rect 15708 13970 15764 14252
rect 15708 13918 15710 13970
rect 15762 13918 15764 13970
rect 15708 13906 15764 13918
rect 15540 12124 15652 12180
rect 15484 12114 15540 12124
rect 15260 12068 15316 12078
rect 15148 12066 15428 12068
rect 15148 12014 15262 12066
rect 15314 12014 15428 12066
rect 15148 12012 15428 12014
rect 15260 12002 15316 12012
rect 14700 11230 14702 11282
rect 14754 11230 14756 11282
rect 14700 11218 14756 11230
rect 15148 11732 15204 11742
rect 14588 11004 14756 11060
rect 13804 10892 14308 10948
rect 14364 10892 14644 10948
rect 13580 10836 13636 10846
rect 13468 10834 13636 10836
rect 13468 10782 13582 10834
rect 13634 10782 13636 10834
rect 13468 10780 13636 10782
rect 13356 10406 13412 10444
rect 13580 10276 13636 10780
rect 14028 10722 14084 10734
rect 14028 10670 14030 10722
rect 14082 10670 14084 10722
rect 13804 10610 13860 10622
rect 13804 10558 13806 10610
rect 13858 10558 13860 10610
rect 13580 10210 13636 10220
rect 13692 10498 13748 10510
rect 13692 10446 13694 10498
rect 13746 10446 13748 10498
rect 13468 9828 13524 9838
rect 12852 9826 13524 9828
rect 12852 9774 13470 9826
rect 13522 9774 13524 9826
rect 12852 9772 13524 9774
rect 12460 9268 12516 9278
rect 12348 9266 12740 9268
rect 12348 9214 12462 9266
rect 12514 9214 12740 9266
rect 12348 9212 12740 9214
rect 12460 9202 12516 9212
rect 12684 9044 12740 9212
rect 12796 9266 12852 9772
rect 12796 9214 12798 9266
rect 12850 9214 12852 9266
rect 12796 9202 12852 9214
rect 13020 9324 13412 9380
rect 13020 9044 13076 9324
rect 13132 9156 13188 9166
rect 13132 9062 13188 9100
rect 12684 8988 13076 9044
rect 13356 9042 13412 9324
rect 13468 9268 13524 9772
rect 13524 9212 13636 9268
rect 13468 9202 13524 9212
rect 13356 8990 13358 9042
rect 13410 8990 13412 9042
rect 13356 8978 13412 8990
rect 13244 8930 13300 8942
rect 13244 8878 13246 8930
rect 13298 8878 13300 8930
rect 11418 8652 11682 8662
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11418 8586 11682 8596
rect 13244 8372 13300 8878
rect 13244 8306 13300 8316
rect 13580 8258 13636 9212
rect 13692 9154 13748 10446
rect 13804 10388 13860 10558
rect 14028 10612 14084 10670
rect 14028 10546 14084 10556
rect 13804 10322 13860 10332
rect 14252 9938 14308 10892
rect 14588 10834 14644 10892
rect 14588 10782 14590 10834
rect 14642 10782 14644 10834
rect 14588 10770 14644 10782
rect 14700 10834 14756 11004
rect 14820 11004 15084 11014
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 14820 10938 15084 10948
rect 14700 10782 14702 10834
rect 14754 10782 14756 10834
rect 14700 10770 14756 10782
rect 14924 10836 14980 10846
rect 14476 10610 14532 10622
rect 14476 10558 14478 10610
rect 14530 10558 14532 10610
rect 14476 10164 14532 10558
rect 14476 10098 14532 10108
rect 14588 10276 14644 10286
rect 14252 9886 14254 9938
rect 14306 9886 14308 9938
rect 14252 9874 14308 9886
rect 13692 9102 13694 9154
rect 13746 9102 13748 9154
rect 13692 9090 13748 9102
rect 14140 9156 14196 9166
rect 14140 9062 14196 9100
rect 14588 8932 14644 10220
rect 14924 10276 14980 10780
rect 14924 10210 14980 10220
rect 15148 10612 15204 11676
rect 15372 10724 15428 12012
rect 15372 10658 15428 10668
rect 15260 10612 15316 10622
rect 15148 10610 15316 10612
rect 15148 10558 15262 10610
rect 15314 10558 15316 10610
rect 15148 10556 15316 10558
rect 14700 10052 14756 10062
rect 14700 9156 14756 9996
rect 15148 10052 15204 10556
rect 15260 10546 15316 10556
rect 15484 10498 15540 10510
rect 15484 10446 15486 10498
rect 15538 10446 15540 10498
rect 15148 9986 15204 9996
rect 15372 10276 15428 10286
rect 14820 9436 15084 9446
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 14820 9370 15084 9380
rect 14812 9268 14868 9278
rect 15036 9268 15092 9278
rect 14868 9266 15092 9268
rect 14868 9214 15038 9266
rect 15090 9214 15092 9266
rect 14868 9212 15092 9214
rect 14812 9202 14868 9212
rect 14700 9090 14756 9100
rect 14924 9044 14980 9054
rect 14700 8932 14756 8942
rect 14588 8930 14756 8932
rect 14588 8878 14702 8930
rect 14754 8878 14756 8930
rect 14588 8876 14756 8878
rect 14700 8866 14756 8876
rect 14252 8372 14308 8382
rect 14252 8278 14308 8316
rect 13580 8206 13582 8258
rect 13634 8206 13636 8258
rect 9660 7700 9716 7710
rect 9268 7698 9716 7700
rect 9268 7646 9662 7698
rect 9714 7646 9716 7698
rect 9268 7644 9716 7646
rect 9212 7606 9268 7644
rect 9660 7634 9716 7644
rect 13580 7700 13636 8206
rect 14924 8036 14980 8988
rect 15036 8372 15092 9212
rect 15372 9044 15428 10220
rect 15484 9268 15540 10446
rect 15596 9940 15652 12124
rect 16268 12068 16324 16940
rect 16828 16884 16884 17390
rect 16828 16818 16884 16828
rect 16492 16658 16548 16670
rect 16492 16606 16494 16658
rect 16546 16606 16548 16658
rect 16492 14642 16548 16606
rect 16604 15428 16660 15438
rect 16604 15314 16660 15372
rect 16604 15262 16606 15314
rect 16658 15262 16660 15314
rect 16604 15148 16660 15262
rect 16940 15148 16996 17500
rect 17164 16660 17220 17612
rect 17276 17444 17332 17454
rect 17276 17108 17332 17388
rect 17276 17042 17332 17052
rect 17612 16884 17668 16894
rect 17612 16790 17668 16828
rect 17276 16660 17332 16670
rect 17164 16658 17332 16660
rect 17164 16606 17278 16658
rect 17330 16606 17332 16658
rect 17164 16604 17332 16606
rect 17276 16594 17332 16604
rect 16604 15092 16772 15148
rect 16716 15026 16772 15036
rect 16828 15092 16996 15148
rect 17052 16212 17108 16222
rect 16492 14590 16494 14642
rect 16546 14590 16548 14642
rect 16492 14578 16548 14590
rect 16716 13972 16772 13982
rect 16716 12740 16772 13916
rect 16716 12674 16772 12684
rect 16380 12404 16436 12414
rect 16380 12310 16436 12348
rect 16828 12292 16884 15092
rect 16268 11788 16324 12012
rect 16716 12236 16884 12292
rect 16940 14980 16996 14990
rect 16716 11844 16772 12236
rect 16828 12068 16884 12078
rect 16828 11974 16884 12012
rect 16716 11788 16884 11844
rect 15932 11732 16324 11788
rect 15820 11620 15876 11630
rect 15820 11506 15876 11564
rect 15820 11454 15822 11506
rect 15874 11454 15876 11506
rect 15820 11442 15876 11454
rect 15932 11394 15988 11732
rect 15932 11342 15934 11394
rect 15986 11342 15988 11394
rect 15932 11330 15988 11342
rect 16380 11396 16436 11406
rect 16380 11394 16660 11396
rect 16380 11342 16382 11394
rect 16434 11342 16660 11394
rect 16380 11340 16660 11342
rect 16380 11330 16436 11340
rect 15820 11284 15876 11294
rect 15708 11172 15764 11182
rect 15708 10722 15764 11116
rect 15708 10670 15710 10722
rect 15762 10670 15764 10722
rect 15708 10500 15764 10670
rect 15708 10434 15764 10444
rect 15820 9940 15876 11228
rect 16380 10836 16436 10846
rect 15932 10834 16436 10836
rect 15932 10782 16382 10834
rect 16434 10782 16436 10834
rect 15932 10780 16436 10782
rect 15932 10722 15988 10780
rect 16380 10770 16436 10780
rect 15932 10670 15934 10722
rect 15986 10670 15988 10722
rect 15932 10658 15988 10670
rect 16268 10612 16324 10622
rect 16268 10518 16324 10556
rect 16492 10612 16548 10622
rect 16492 10518 16548 10556
rect 16492 10388 16548 10398
rect 16380 9940 16436 9950
rect 15820 9938 16436 9940
rect 15820 9886 16382 9938
rect 16434 9886 16436 9938
rect 15820 9884 16436 9886
rect 15596 9874 15652 9884
rect 16380 9874 16436 9884
rect 15484 9202 15540 9212
rect 15484 9044 15540 9054
rect 15372 9042 15540 9044
rect 15372 8990 15486 9042
rect 15538 8990 15540 9042
rect 15372 8988 15540 8990
rect 15484 8978 15540 8988
rect 16156 8932 16212 8942
rect 16156 8838 16212 8876
rect 15036 8306 15092 8316
rect 16380 8372 16436 8382
rect 16492 8372 16548 10332
rect 16604 10052 16660 11340
rect 16828 10836 16884 11788
rect 16940 11172 16996 14924
rect 17052 14530 17108 16156
rect 17724 14644 17780 21756
rect 17836 21810 18004 21812
rect 17836 21758 17950 21810
rect 18002 21758 18004 21810
rect 17836 21756 18004 21758
rect 17836 20916 17892 21756
rect 17948 21746 18004 21756
rect 17836 20850 17892 20860
rect 17948 21588 18004 21598
rect 17948 20356 18004 21532
rect 17836 20300 18004 20356
rect 18060 21476 18116 21486
rect 18060 20692 18116 21420
rect 18396 21474 18452 21486
rect 18396 21422 18398 21474
rect 18450 21422 18452 21474
rect 18396 21364 18452 21422
rect 18396 21298 18452 21308
rect 18222 21196 18486 21206
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18222 21130 18486 21140
rect 17836 17666 17892 20300
rect 18060 19460 18116 20636
rect 18620 20916 18676 20926
rect 18732 20916 18788 24556
rect 19068 24500 19124 24510
rect 18844 24498 19124 24500
rect 18844 24446 19070 24498
rect 19122 24446 19124 24498
rect 18844 24444 19124 24446
rect 18844 24164 18900 24444
rect 19068 24434 19124 24444
rect 18844 24098 18900 24108
rect 18956 24276 19012 24286
rect 18844 23716 18900 23726
rect 18844 23622 18900 23660
rect 18956 23548 19012 24220
rect 18620 20914 18788 20916
rect 18620 20862 18622 20914
rect 18674 20862 18788 20914
rect 18620 20860 18788 20862
rect 18844 23492 19012 23548
rect 18222 19628 18486 19638
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18222 19562 18486 19572
rect 18172 19460 18228 19470
rect 18060 19458 18228 19460
rect 18060 19406 18174 19458
rect 18226 19406 18228 19458
rect 18060 19404 18228 19406
rect 18172 19394 18228 19404
rect 18284 19460 18340 19470
rect 18284 19346 18340 19404
rect 18284 19294 18286 19346
rect 18338 19294 18340 19346
rect 18284 19282 18340 19294
rect 18508 19236 18564 19246
rect 18620 19236 18676 20860
rect 18508 19234 18676 19236
rect 18508 19182 18510 19234
rect 18562 19182 18676 19234
rect 18508 19180 18676 19182
rect 18508 19170 18564 19180
rect 18620 19012 18676 19022
rect 17836 17614 17838 17666
rect 17890 17614 17892 17666
rect 17836 17602 17892 17614
rect 17948 18452 18004 18462
rect 17948 18338 18004 18396
rect 18508 18452 18564 18462
rect 18620 18452 18676 18956
rect 18508 18450 18676 18452
rect 18508 18398 18510 18450
rect 18562 18398 18676 18450
rect 18508 18396 18676 18398
rect 18508 18386 18564 18396
rect 17948 18286 17950 18338
rect 18002 18286 18004 18338
rect 17948 16884 18004 18286
rect 18222 18060 18486 18070
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18222 17994 18486 18004
rect 18620 17892 18676 18396
rect 18508 17836 18676 17892
rect 18508 17332 18564 17836
rect 18844 17780 18900 23492
rect 19068 23044 19124 23054
rect 19068 22950 19124 22988
rect 18956 22930 19012 22942
rect 18956 22878 18958 22930
rect 19010 22878 19012 22930
rect 18956 21812 19012 22878
rect 19180 22708 19236 26012
rect 19292 25844 19348 25854
rect 19292 25508 19348 25788
rect 19628 25620 19684 26236
rect 19628 25564 19796 25620
rect 19292 25414 19348 25452
rect 19740 25284 19796 25564
rect 19740 25190 19796 25228
rect 19852 25060 19908 26572
rect 20076 26516 20132 27020
rect 20412 27076 20468 27114
rect 20412 27010 20468 27020
rect 20188 26962 20244 26974
rect 20188 26910 20190 26962
rect 20242 26910 20244 26962
rect 20188 26908 20244 26910
rect 20188 26852 20356 26908
rect 20188 26516 20244 26526
rect 20076 26514 20244 26516
rect 20076 26462 20190 26514
rect 20242 26462 20244 26514
rect 20076 26460 20244 26462
rect 19740 25004 19908 25060
rect 19964 26404 20020 26414
rect 19628 24836 19684 24874
rect 19628 24770 19684 24780
rect 19292 24610 19348 24622
rect 19740 24612 19796 25004
rect 19292 24558 19294 24610
rect 19346 24558 19348 24610
rect 19292 24050 19348 24558
rect 19292 23998 19294 24050
rect 19346 23998 19348 24050
rect 19292 23986 19348 23998
rect 19628 24556 19796 24612
rect 19852 24722 19908 24734
rect 19852 24670 19854 24722
rect 19906 24670 19908 24722
rect 19852 24612 19908 24670
rect 19292 23716 19348 23726
rect 19516 23716 19572 23726
rect 19292 23622 19348 23660
rect 19404 23714 19572 23716
rect 19404 23662 19518 23714
rect 19570 23662 19572 23714
rect 19404 23660 19572 23662
rect 19292 22708 19348 22718
rect 19180 22652 19292 22708
rect 19292 22642 19348 22652
rect 19068 22372 19124 22382
rect 19124 22316 19348 22372
rect 19068 22278 19124 22316
rect 19068 21812 19124 21822
rect 18956 21756 19068 21812
rect 18956 21588 19012 21598
rect 18956 21494 19012 21532
rect 18956 20804 19012 20814
rect 19068 20804 19124 21756
rect 18956 20802 19124 20804
rect 18956 20750 18958 20802
rect 19010 20750 19124 20802
rect 18956 20748 19124 20750
rect 19180 21364 19236 21374
rect 19180 20802 19236 21308
rect 19180 20750 19182 20802
rect 19234 20750 19236 20802
rect 18956 20244 19012 20748
rect 19180 20738 19236 20750
rect 18956 20178 19012 20188
rect 19068 20578 19124 20590
rect 19068 20526 19070 20578
rect 19122 20526 19124 20578
rect 18956 19012 19012 19022
rect 18956 18918 19012 18956
rect 19068 18452 19124 20526
rect 19180 18452 19236 18462
rect 19068 18450 19236 18452
rect 19068 18398 19182 18450
rect 19234 18398 19236 18450
rect 19068 18396 19236 18398
rect 19180 18386 19236 18396
rect 18844 17724 19124 17780
rect 18620 17556 18676 17566
rect 18620 17462 18676 17500
rect 18956 17556 19012 17566
rect 18844 17332 18900 17342
rect 18508 17276 18788 17332
rect 18060 17108 18116 17118
rect 18060 17014 18116 17052
rect 18508 17106 18564 17118
rect 18508 17054 18510 17106
rect 18562 17054 18564 17106
rect 18508 16996 18564 17054
rect 18620 16996 18676 17006
rect 18508 16940 18620 16996
rect 18620 16930 18676 16940
rect 17948 16828 18116 16884
rect 17836 16658 17892 16670
rect 17836 16606 17838 16658
rect 17890 16606 17892 16658
rect 17836 16212 17892 16606
rect 17948 16212 18004 16222
rect 17836 16210 18004 16212
rect 17836 16158 17950 16210
rect 18002 16158 18004 16210
rect 17836 16156 18004 16158
rect 17948 16146 18004 16156
rect 18060 16100 18116 16828
rect 18222 16492 18486 16502
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18222 16426 18486 16436
rect 18396 16212 18452 16222
rect 18396 16118 18452 16156
rect 18732 16212 18788 17276
rect 18844 16994 18900 17276
rect 18956 17106 19012 17500
rect 19068 17332 19124 17724
rect 19068 17266 19124 17276
rect 18956 17054 18958 17106
rect 19010 17054 19012 17106
rect 18956 17042 19012 17054
rect 18844 16942 18846 16994
rect 18898 16942 18900 16994
rect 18844 16930 18900 16942
rect 19180 16996 19236 17006
rect 19292 16996 19348 22316
rect 19404 20132 19460 23660
rect 19516 23650 19572 23660
rect 19516 23044 19572 23054
rect 19516 22950 19572 22988
rect 19628 22484 19684 24556
rect 19852 24546 19908 24556
rect 19852 24388 19908 24398
rect 19852 23938 19908 24332
rect 19852 23886 19854 23938
rect 19906 23886 19908 23938
rect 19852 23548 19908 23886
rect 19740 23492 19908 23548
rect 19740 23044 19796 23492
rect 19740 22978 19796 22988
rect 19852 23380 19908 23390
rect 19516 22428 19684 22484
rect 19516 21252 19572 22428
rect 19852 22372 19908 23324
rect 19852 22278 19908 22316
rect 19628 22258 19684 22270
rect 19628 22206 19630 22258
rect 19682 22206 19684 22258
rect 19628 21812 19684 22206
rect 19628 21746 19684 21756
rect 19740 22146 19796 22158
rect 19740 22094 19742 22146
rect 19794 22094 19796 22146
rect 19740 21698 19796 22094
rect 19740 21646 19742 21698
rect 19794 21646 19796 21698
rect 19740 21634 19796 21646
rect 19516 21196 19684 21252
rect 19516 21028 19572 21038
rect 19516 20934 19572 20972
rect 19516 20804 19572 20814
rect 19516 20710 19572 20748
rect 19628 20244 19684 21196
rect 19964 20804 20020 26348
rect 20076 25396 20132 26460
rect 20188 26450 20244 26460
rect 20300 25844 20356 26852
rect 20300 25778 20356 25788
rect 20412 26852 20468 26862
rect 20188 25620 20244 25630
rect 20412 25620 20468 26796
rect 20188 25618 20468 25620
rect 20188 25566 20190 25618
rect 20242 25566 20468 25618
rect 20188 25564 20468 25566
rect 20188 25554 20244 25564
rect 20076 25340 20356 25396
rect 20188 24948 20244 24958
rect 20188 24854 20244 24892
rect 20076 24834 20132 24846
rect 20076 24782 20078 24834
rect 20130 24782 20132 24834
rect 20076 24500 20132 24782
rect 20076 24052 20132 24444
rect 20188 24052 20244 24062
rect 20076 23996 20188 24052
rect 20188 23958 20244 23996
rect 20076 23716 20132 23726
rect 20076 23378 20132 23660
rect 20076 23326 20078 23378
rect 20130 23326 20132 23378
rect 20076 23314 20132 23326
rect 20300 23380 20356 25340
rect 20412 24834 20468 25564
rect 20524 25396 20580 28028
rect 20636 26292 20692 29934
rect 20748 29876 20804 29886
rect 20748 28530 20804 29820
rect 20748 28478 20750 28530
rect 20802 28478 20804 28530
rect 20748 27524 20804 28478
rect 20748 27458 20804 27468
rect 20748 27076 20804 27086
rect 20748 26962 20804 27020
rect 20748 26910 20750 26962
rect 20802 26910 20804 26962
rect 20748 26898 20804 26910
rect 20636 26226 20692 26236
rect 20748 25956 20804 25966
rect 20748 25618 20804 25900
rect 20748 25566 20750 25618
rect 20802 25566 20804 25618
rect 20748 25554 20804 25566
rect 20748 25396 20804 25406
rect 20524 25340 20748 25396
rect 20748 25330 20804 25340
rect 20860 25060 20916 35308
rect 20972 32452 21028 32462
rect 20972 32358 21028 32396
rect 21084 32228 21140 37212
rect 21196 34356 21252 37436
rect 21308 37154 21364 37548
rect 21308 37102 21310 37154
rect 21362 37102 21364 37154
rect 21308 37042 21364 37102
rect 21308 36990 21310 37042
rect 21362 36990 21364 37042
rect 21308 36978 21364 36990
rect 21420 36820 21476 37660
rect 21624 37660 21888 37670
rect 21680 37604 21728 37660
rect 21784 37604 21832 37660
rect 21624 37594 21888 37604
rect 21980 37380 22036 37772
rect 22092 37492 22148 37998
rect 22092 37426 22148 37436
rect 22204 38052 22260 38062
rect 21868 37324 22036 37380
rect 21756 37156 21812 37166
rect 21756 37062 21812 37100
rect 21308 36764 21476 36820
rect 21308 36482 21364 36764
rect 21868 36596 21924 37324
rect 22204 37268 22260 37996
rect 22316 37490 22372 38332
rect 22540 38164 22596 41692
rect 22764 41636 22820 44156
rect 22988 42196 23044 44268
rect 23100 43650 23156 45612
rect 23212 45332 23268 45342
rect 23324 45332 23380 46284
rect 23212 45330 23380 45332
rect 23212 45278 23214 45330
rect 23266 45278 23380 45330
rect 23212 45276 23380 45278
rect 23548 45444 23604 45454
rect 23212 45266 23268 45276
rect 23548 44996 23604 45388
rect 23660 45330 23716 48300
rect 23660 45278 23662 45330
rect 23714 45278 23716 45330
rect 23660 45266 23716 45278
rect 23100 43598 23102 43650
rect 23154 43598 23156 43650
rect 23100 43586 23156 43598
rect 23324 44940 23604 44996
rect 23100 42196 23156 42206
rect 22988 42194 23156 42196
rect 22988 42142 23102 42194
rect 23154 42142 23156 42194
rect 22988 42140 23156 42142
rect 23100 42130 23156 42140
rect 23324 41972 23380 44940
rect 23772 44548 23828 52108
rect 23884 51492 23940 51502
rect 23884 51378 23940 51436
rect 23884 51326 23886 51378
rect 23938 51326 23940 51378
rect 23884 51314 23940 51326
rect 23996 50428 24052 52108
rect 24220 51716 24276 51726
rect 24276 51660 24388 51716
rect 24220 51650 24276 51660
rect 24332 51602 24388 51660
rect 24332 51550 24334 51602
rect 24386 51550 24388 51602
rect 24332 51538 24388 51550
rect 24220 51492 24276 51502
rect 24108 51380 24164 51418
rect 24108 51314 24164 51324
rect 23996 50372 24164 50428
rect 24108 49588 24164 50372
rect 24220 50036 24276 51436
rect 24444 51156 24500 51166
rect 24332 50708 24388 50718
rect 24332 50614 24388 50652
rect 24444 50596 24500 51100
rect 24444 50530 24500 50540
rect 24332 50484 24388 50494
rect 24332 50372 24500 50428
rect 24276 49980 24388 50036
rect 24220 49970 24276 49980
rect 23884 49252 23940 49290
rect 23884 49186 23940 49196
rect 23996 49028 24052 49038
rect 23996 46900 24052 48972
rect 23996 46834 24052 46844
rect 24108 49026 24164 49532
rect 24108 48974 24110 49026
rect 24162 48974 24164 49026
rect 23884 46674 23940 46686
rect 23884 46622 23886 46674
rect 23938 46622 23940 46674
rect 23884 45444 23940 46622
rect 23884 45378 23940 45388
rect 23996 45332 24052 45342
rect 23996 45238 24052 45276
rect 23660 44492 23828 44548
rect 23436 43876 23492 43886
rect 23436 43762 23492 43820
rect 23436 43710 23438 43762
rect 23490 43710 23492 43762
rect 23436 43314 23492 43710
rect 23436 43262 23438 43314
rect 23490 43262 23492 43314
rect 23436 43250 23492 43262
rect 23436 42642 23492 42654
rect 23436 42590 23438 42642
rect 23490 42590 23492 42642
rect 23436 42196 23492 42590
rect 23660 42532 23716 44492
rect 23772 44324 23828 44334
rect 23772 44230 23828 44268
rect 24108 43708 24164 48974
rect 24332 49028 24388 49980
rect 24332 48962 24388 48972
rect 24220 48916 24276 48926
rect 24220 48132 24276 48860
rect 24444 48914 24500 50372
rect 24668 49924 24724 53116
rect 25116 53106 25172 53116
rect 24892 52948 24948 52958
rect 24780 52612 24836 52622
rect 24780 52274 24836 52556
rect 24780 52222 24782 52274
rect 24834 52222 24836 52274
rect 24780 52210 24836 52222
rect 24892 50594 24948 52892
rect 25228 52948 25284 52958
rect 25228 52854 25284 52892
rect 25026 52556 25290 52566
rect 25082 52500 25130 52556
rect 25186 52500 25234 52556
rect 25026 52490 25290 52500
rect 25228 52164 25284 52174
rect 25228 52070 25284 52108
rect 25340 51266 25396 51278
rect 25340 51214 25342 51266
rect 25394 51214 25396 51266
rect 25340 51156 25396 51214
rect 25340 51090 25396 51100
rect 25026 50988 25290 50998
rect 25082 50932 25130 50988
rect 25186 50932 25234 50988
rect 25026 50922 25290 50932
rect 25452 50820 25508 54238
rect 25676 52164 25732 54572
rect 25788 54290 25844 54302
rect 25788 54238 25790 54290
rect 25842 54238 25844 54290
rect 25788 53730 25844 54238
rect 25788 53678 25790 53730
rect 25842 53678 25844 53730
rect 25788 53666 25844 53678
rect 25676 52098 25732 52108
rect 25788 53172 25844 53182
rect 25676 51940 25732 51950
rect 25788 51940 25844 53116
rect 25676 51938 25844 51940
rect 25676 51886 25678 51938
rect 25730 51886 25844 51938
rect 25676 51884 25844 51886
rect 25676 51874 25732 51884
rect 25788 51492 25844 51502
rect 25788 51398 25844 51436
rect 25452 50764 25620 50820
rect 24892 50542 24894 50594
rect 24946 50542 24948 50594
rect 24668 49868 24836 49924
rect 24668 49698 24724 49710
rect 24668 49646 24670 49698
rect 24722 49646 24724 49698
rect 24668 49028 24724 49646
rect 24668 48934 24724 48972
rect 24444 48862 24446 48914
rect 24498 48862 24500 48914
rect 24444 48850 24500 48862
rect 24332 48804 24388 48814
rect 24332 48710 24388 48748
rect 24556 48132 24612 48142
rect 24220 48130 24612 48132
rect 24220 48078 24558 48130
rect 24610 48078 24612 48130
rect 24220 48076 24612 48078
rect 24556 48066 24612 48076
rect 24220 47346 24276 47358
rect 24220 47294 24222 47346
rect 24274 47294 24276 47346
rect 24220 46898 24276 47294
rect 24220 46846 24222 46898
rect 24274 46846 24276 46898
rect 24220 46834 24276 46846
rect 24332 46900 24388 46910
rect 24220 46676 24276 46686
rect 24220 46002 24276 46620
rect 24220 45950 24222 46002
rect 24274 45950 24276 46002
rect 24220 45938 24276 45950
rect 24332 46674 24388 46844
rect 24332 46622 24334 46674
rect 24386 46622 24388 46674
rect 24332 45668 24388 46622
rect 24332 45602 24388 45612
rect 24444 46788 24500 46798
rect 24444 45220 24500 46732
rect 24556 46676 24612 46686
rect 24556 46582 24612 46620
rect 24668 45668 24724 45678
rect 24668 45574 24724 45612
rect 24444 45164 24612 45220
rect 24444 44996 24500 45006
rect 24444 44902 24500 44940
rect 23660 42466 23716 42476
rect 23772 43652 24164 43708
rect 23436 42130 23492 42140
rect 23548 41972 23604 41982
rect 23324 41970 23604 41972
rect 23324 41918 23550 41970
rect 23602 41918 23604 41970
rect 23324 41916 23604 41918
rect 22652 41580 22820 41636
rect 22876 41746 22932 41758
rect 22876 41694 22878 41746
rect 22930 41694 22932 41746
rect 22652 39730 22708 41580
rect 22652 39678 22654 39730
rect 22706 39678 22708 39730
rect 22652 38612 22708 39678
rect 22764 41410 22820 41422
rect 22764 41358 22766 41410
rect 22818 41358 22820 41410
rect 22764 41298 22820 41358
rect 22764 41246 22766 41298
rect 22818 41246 22820 41298
rect 22764 38836 22820 41246
rect 22876 41300 22932 41694
rect 23324 41746 23380 41916
rect 23492 41804 23604 41916
rect 23324 41694 23326 41746
rect 23378 41694 23380 41746
rect 23324 41682 23380 41694
rect 22876 40626 22932 41244
rect 22876 40574 22878 40626
rect 22930 40574 22932 40626
rect 22876 40516 22932 40574
rect 22876 40450 22932 40460
rect 23212 41188 23268 41198
rect 23548 41188 23604 41198
rect 23212 40180 23268 41132
rect 23324 41132 23548 41188
rect 23324 40628 23380 41132
rect 23548 41122 23604 41132
rect 23548 40964 23604 40974
rect 23548 40870 23604 40908
rect 23324 40534 23380 40572
rect 23660 40516 23716 40526
rect 22764 38770 22820 38780
rect 22988 39844 23044 39854
rect 22988 39730 23044 39788
rect 22988 39678 22990 39730
rect 23042 39678 23044 39730
rect 22652 38546 22708 38556
rect 22316 37438 22318 37490
rect 22370 37438 22372 37490
rect 22316 37426 22372 37438
rect 22428 38108 22596 38164
rect 22204 37212 22372 37268
rect 21980 37156 22036 37166
rect 21980 37062 22036 37100
rect 22204 37042 22260 37054
rect 22204 36990 22206 37042
rect 22258 36990 22260 37042
rect 22204 36596 22260 36990
rect 21756 36540 21924 36596
rect 22092 36540 22260 36596
rect 22316 36596 22372 37212
rect 22428 36820 22484 38108
rect 22764 38052 22820 38062
rect 22540 37996 22764 38052
rect 22988 38052 23044 39678
rect 23212 39060 23268 40124
rect 23100 38052 23156 38062
rect 22988 38050 23156 38052
rect 22988 37998 23102 38050
rect 23154 37998 23156 38050
rect 22988 37996 23156 37998
rect 22540 37266 22596 37996
rect 22764 37958 22820 37996
rect 23100 37986 23156 37996
rect 22540 37214 22542 37266
rect 22594 37214 22596 37266
rect 22540 37202 22596 37214
rect 22652 37826 22708 37838
rect 22652 37774 22654 37826
rect 22706 37774 22708 37826
rect 22652 37156 22708 37774
rect 22876 37826 22932 37838
rect 22876 37774 22878 37826
rect 22930 37774 22932 37826
rect 22652 37090 22708 37100
rect 22764 37380 22820 37390
rect 22428 36764 22596 36820
rect 22428 36596 22484 36606
rect 22316 36594 22484 36596
rect 22316 36542 22430 36594
rect 22482 36542 22484 36594
rect 22316 36540 22484 36542
rect 21308 36430 21310 36482
rect 21362 36430 21364 36482
rect 21308 35924 21364 36430
rect 21532 36484 21588 36494
rect 21420 36372 21476 36382
rect 21532 36372 21588 36428
rect 21420 36370 21588 36372
rect 21420 36318 21422 36370
rect 21474 36318 21588 36370
rect 21420 36316 21588 36318
rect 21644 36372 21700 36382
rect 21756 36372 21812 36540
rect 21644 36370 21812 36372
rect 21644 36318 21646 36370
rect 21698 36318 21812 36370
rect 21644 36316 21812 36318
rect 21868 36372 21924 36382
rect 21868 36370 22036 36372
rect 21868 36318 21870 36370
rect 21922 36318 22036 36370
rect 21868 36316 22036 36318
rect 21420 36306 21476 36316
rect 21644 36260 21700 36316
rect 21868 36306 21924 36316
rect 21644 36194 21700 36204
rect 21308 35858 21364 35868
rect 21420 36148 21476 36158
rect 21420 35028 21476 36092
rect 21624 36092 21888 36102
rect 21680 36036 21728 36092
rect 21784 36036 21832 36092
rect 21624 36026 21888 36036
rect 21532 35028 21588 35038
rect 21420 35026 21588 35028
rect 21420 34974 21534 35026
rect 21586 34974 21588 35026
rect 21420 34972 21588 34974
rect 21532 34962 21588 34972
rect 21980 35026 22036 36316
rect 22092 35252 22148 36540
rect 22428 36530 22484 36540
rect 22540 36372 22596 36764
rect 22764 36596 22820 37324
rect 22876 37268 22932 37774
rect 22988 37828 23044 37838
rect 22988 37826 23156 37828
rect 22988 37774 22990 37826
rect 23042 37774 23156 37826
rect 22988 37772 23156 37774
rect 22988 37762 23044 37772
rect 22988 37492 23044 37502
rect 22988 37398 23044 37436
rect 22876 37202 22932 37212
rect 23100 36708 23156 37772
rect 23212 37492 23268 39004
rect 23548 40292 23604 40302
rect 23436 38722 23492 38734
rect 23436 38670 23438 38722
rect 23490 38670 23492 38722
rect 23436 38052 23492 38670
rect 23548 38274 23604 40236
rect 23660 38836 23716 40460
rect 23660 38742 23716 38780
rect 23772 38724 23828 43652
rect 23996 43538 24052 43550
rect 23996 43486 23998 43538
rect 24050 43486 24052 43538
rect 23884 42644 23940 42654
rect 23884 42194 23940 42588
rect 23884 42142 23886 42194
rect 23938 42142 23940 42194
rect 23884 42130 23940 42142
rect 23996 42196 24052 43486
rect 24220 43538 24276 43550
rect 24220 43486 24222 43538
rect 24274 43486 24276 43538
rect 24108 43426 24164 43438
rect 24108 43374 24110 43426
rect 24162 43374 24164 43426
rect 24108 42980 24164 43374
rect 24220 43204 24276 43486
rect 24556 43540 24612 45164
rect 24556 43538 24724 43540
rect 24556 43486 24558 43538
rect 24610 43486 24724 43538
rect 24556 43484 24724 43486
rect 24556 43474 24612 43484
rect 24220 43148 24500 43204
rect 24108 42924 24276 42980
rect 23996 42130 24052 42140
rect 24108 42754 24164 42766
rect 24108 42702 24110 42754
rect 24162 42702 24164 42754
rect 24108 42084 24164 42702
rect 24108 42018 24164 42028
rect 24220 42082 24276 42924
rect 24444 42868 24500 43148
rect 24556 42868 24612 42878
rect 24444 42866 24612 42868
rect 24444 42814 24558 42866
rect 24610 42814 24612 42866
rect 24444 42812 24612 42814
rect 24220 42030 24222 42082
rect 24274 42030 24276 42082
rect 24220 42018 24276 42030
rect 24444 42532 24500 42542
rect 23884 41972 23940 41982
rect 23884 40626 23940 41916
rect 23996 41970 24052 41982
rect 23996 41918 23998 41970
rect 24050 41918 24052 41970
rect 23996 41860 24052 41918
rect 23996 41804 24164 41860
rect 23996 41636 24052 41646
rect 23996 41298 24052 41580
rect 23996 41246 23998 41298
rect 24050 41246 24052 41298
rect 23996 41234 24052 41246
rect 24108 40964 24164 41804
rect 24444 41636 24500 42476
rect 24556 41860 24612 42812
rect 24668 42196 24724 43484
rect 24668 42130 24724 42140
rect 24668 41972 24724 41982
rect 24668 41878 24724 41916
rect 24556 41794 24612 41804
rect 24668 41636 24724 41646
rect 24444 41580 24612 41636
rect 24220 40964 24276 40974
rect 24108 40908 24220 40964
rect 24220 40898 24276 40908
rect 23884 40574 23886 40626
rect 23938 40574 23940 40626
rect 23884 40562 23940 40574
rect 24108 40516 24164 40526
rect 24108 40422 24164 40460
rect 24332 40404 24388 40414
rect 24332 40402 24500 40404
rect 24332 40350 24334 40402
rect 24386 40350 24500 40402
rect 24332 40348 24500 40350
rect 24332 40338 24388 40348
rect 24220 40290 24276 40302
rect 24220 40238 24222 40290
rect 24274 40238 24276 40290
rect 24220 40180 24276 40238
rect 24220 40124 24388 40180
rect 24108 39508 24164 39518
rect 23996 39452 24108 39508
rect 23996 39058 24052 39452
rect 24108 39442 24164 39452
rect 23996 39006 23998 39058
rect 24050 39006 24052 39058
rect 23996 38994 24052 39006
rect 24108 39060 24164 39070
rect 24108 38946 24164 39004
rect 24108 38894 24110 38946
rect 24162 38894 24164 38946
rect 24108 38882 24164 38894
rect 24332 38946 24388 40124
rect 24444 39844 24500 40348
rect 24444 39778 24500 39788
rect 24556 39620 24612 41580
rect 24332 38894 24334 38946
rect 24386 38894 24388 38946
rect 24332 38882 24388 38894
rect 24444 39564 24612 39620
rect 24668 41298 24724 41580
rect 24668 41246 24670 41298
rect 24722 41246 24724 41298
rect 24668 40402 24724 41246
rect 24668 40350 24670 40402
rect 24722 40350 24724 40402
rect 23996 38836 24052 38846
rect 23772 38668 23940 38724
rect 23548 38222 23550 38274
rect 23602 38222 23604 38274
rect 23548 38210 23604 38222
rect 23436 37986 23492 37996
rect 23660 38052 23716 38062
rect 23660 37958 23716 37996
rect 23212 37426 23268 37436
rect 23436 37716 23492 37726
rect 23436 37490 23492 37660
rect 23436 37438 23438 37490
rect 23490 37438 23492 37490
rect 23436 37426 23492 37438
rect 22092 35186 22148 35196
rect 22204 36316 22596 36372
rect 22652 36594 22820 36596
rect 22652 36542 22766 36594
rect 22818 36542 22820 36594
rect 22652 36540 22820 36542
rect 21980 34974 21982 35026
rect 22034 34974 22036 35026
rect 21980 34962 22036 34974
rect 21868 34804 21924 34814
rect 21868 34692 21924 34748
rect 22092 34692 22148 34702
rect 21868 34690 22036 34692
rect 21868 34638 21870 34690
rect 21922 34638 22036 34690
rect 21868 34636 22036 34638
rect 21868 34626 21924 34636
rect 21624 34524 21888 34534
rect 21680 34468 21728 34524
rect 21784 34468 21832 34524
rect 21624 34458 21888 34468
rect 21980 34468 22036 34636
rect 22092 34598 22148 34636
rect 22204 34580 22260 36316
rect 22204 34514 22260 34524
rect 22316 35924 22372 35934
rect 21980 34402 22036 34412
rect 21196 34262 21252 34300
rect 21756 34356 21812 34366
rect 21756 34262 21812 34300
rect 21980 34244 22036 34254
rect 21420 33572 21476 33582
rect 20972 32172 21140 32228
rect 21196 33570 21476 33572
rect 21196 33518 21422 33570
rect 21474 33518 21476 33570
rect 21196 33516 21476 33518
rect 20972 27300 21028 32172
rect 21196 32004 21252 33516
rect 21420 33506 21476 33516
rect 21308 33348 21364 33358
rect 21308 33254 21364 33292
rect 21420 33124 21476 33134
rect 21420 33030 21476 33068
rect 21624 32956 21888 32966
rect 21680 32900 21728 32956
rect 21784 32900 21832 32956
rect 21624 32890 21888 32900
rect 21868 32564 21924 32574
rect 21980 32564 22036 34188
rect 21868 32562 22036 32564
rect 21868 32510 21870 32562
rect 21922 32510 22036 32562
rect 21868 32508 22036 32510
rect 22092 34020 22148 34030
rect 22316 34020 22372 35868
rect 22540 34916 22596 34926
rect 22652 34916 22708 36540
rect 22764 36530 22820 36540
rect 22876 36652 23156 36708
rect 23212 36820 23268 36830
rect 22540 34914 22708 34916
rect 22540 34862 22542 34914
rect 22594 34862 22708 34914
rect 22540 34860 22708 34862
rect 22764 35252 22820 35262
rect 22764 34916 22820 35196
rect 22540 34356 22596 34860
rect 22540 34290 22596 34300
rect 22764 34354 22820 34860
rect 22764 34302 22766 34354
rect 22818 34302 22820 34354
rect 22764 34290 22820 34302
rect 22876 34690 22932 36652
rect 23212 36596 23268 36764
rect 23100 36540 23268 36596
rect 22988 36484 23044 36494
rect 22988 35810 23044 36428
rect 22988 35758 22990 35810
rect 23042 35758 23044 35810
rect 22988 35746 23044 35758
rect 22876 34638 22878 34690
rect 22930 34638 22932 34690
rect 22092 34018 22372 34020
rect 22092 33966 22094 34018
rect 22146 33966 22372 34018
rect 22092 33964 22372 33966
rect 21868 32498 21924 32508
rect 21420 32452 21476 32462
rect 21420 32358 21476 32396
rect 21196 31948 21476 32004
rect 21084 31892 21140 31902
rect 21140 31836 21252 31892
rect 21084 31826 21140 31836
rect 21196 31108 21252 31836
rect 21308 31780 21364 31790
rect 21308 31686 21364 31724
rect 21084 30996 21140 31006
rect 21084 29538 21140 30940
rect 21196 30548 21252 31052
rect 21420 30996 21476 31948
rect 21532 31666 21588 31678
rect 21532 31614 21534 31666
rect 21586 31614 21588 31666
rect 21532 31556 21588 31614
rect 21532 31490 21588 31500
rect 21624 31388 21888 31398
rect 21680 31332 21728 31388
rect 21784 31332 21832 31388
rect 21624 31322 21888 31332
rect 21644 31220 21700 31230
rect 21644 31126 21700 31164
rect 21532 30996 21588 31006
rect 21420 30994 21588 30996
rect 21420 30942 21534 30994
rect 21586 30942 21588 30994
rect 21420 30940 21588 30942
rect 21532 30930 21588 30940
rect 21980 30996 22036 31006
rect 21980 30902 22036 30940
rect 21196 30492 21364 30548
rect 21308 29652 21364 30492
rect 21420 30436 21476 30446
rect 21420 30322 21476 30380
rect 21420 30270 21422 30322
rect 21474 30270 21476 30322
rect 21420 29876 21476 30270
rect 21868 29988 21924 30026
rect 21868 29922 21924 29932
rect 21420 29810 21476 29820
rect 21624 29820 21888 29830
rect 21680 29764 21728 29820
rect 21784 29764 21832 29820
rect 21624 29754 21888 29764
rect 21868 29652 21924 29662
rect 21308 29596 21812 29652
rect 21084 29486 21086 29538
rect 21138 29486 21140 29538
rect 21084 29474 21140 29486
rect 21308 29428 21364 29438
rect 21364 29372 21476 29428
rect 21308 27412 21364 29372
rect 21420 29314 21476 29372
rect 21420 29262 21422 29314
rect 21474 29262 21476 29314
rect 21420 29250 21476 29262
rect 21756 29314 21812 29596
rect 21756 29262 21758 29314
rect 21810 29262 21812 29314
rect 21756 29250 21812 29262
rect 21868 28754 21924 29596
rect 21868 28702 21870 28754
rect 21922 28702 21924 28754
rect 21868 28690 21924 28702
rect 21980 28420 22036 28430
rect 21624 28252 21888 28262
rect 21680 28196 21728 28252
rect 21784 28196 21832 28252
rect 21624 28186 21888 28196
rect 21308 27346 21364 27356
rect 20972 27234 21028 27244
rect 21308 27076 21364 27086
rect 21308 26908 21364 27020
rect 21308 26852 21476 26908
rect 21308 26516 21364 26526
rect 21308 26422 21364 26460
rect 21420 26514 21476 26852
rect 21624 26684 21888 26694
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21624 26618 21888 26628
rect 21420 26462 21422 26514
rect 21474 26462 21476 26514
rect 21420 26450 21476 26462
rect 21532 26516 21588 26526
rect 21980 26516 22036 28364
rect 21532 26514 22036 26516
rect 21532 26462 21534 26514
rect 21586 26462 22036 26514
rect 21532 26460 22036 26462
rect 21532 26450 21588 26460
rect 21644 26292 21700 26302
rect 20972 26178 21028 26190
rect 20972 26126 20974 26178
rect 21026 26126 21028 26178
rect 20972 25956 21028 26126
rect 20972 25890 21028 25900
rect 20412 24782 20414 24834
rect 20466 24782 20468 24834
rect 20412 23940 20468 24782
rect 20412 23874 20468 23884
rect 20524 25004 20916 25060
rect 20972 25620 21028 25630
rect 20524 23492 20580 25004
rect 20972 24946 21028 25564
rect 21644 25618 21700 26236
rect 21980 26290 22036 26302
rect 21980 26238 21982 26290
rect 22034 26238 22036 26290
rect 21980 26068 22036 26238
rect 21980 26002 22036 26012
rect 21644 25566 21646 25618
rect 21698 25566 21700 25618
rect 21644 25554 21700 25566
rect 21420 25396 21476 25406
rect 20972 24894 20974 24946
rect 21026 24894 21028 24946
rect 20972 24882 21028 24894
rect 21084 25172 21140 25182
rect 20860 24834 20916 24846
rect 20860 24782 20862 24834
rect 20914 24782 20916 24834
rect 20636 24724 20692 24734
rect 20636 24722 20804 24724
rect 20636 24670 20638 24722
rect 20690 24670 20804 24722
rect 20636 24668 20804 24670
rect 20636 24658 20692 24668
rect 20636 24052 20692 24062
rect 20636 23958 20692 23996
rect 20524 23436 20692 23492
rect 20300 23314 20356 23324
rect 20524 23156 20580 23166
rect 20188 23154 20580 23156
rect 20188 23102 20526 23154
rect 20578 23102 20580 23154
rect 20188 23100 20580 23102
rect 20188 22594 20244 23100
rect 20524 23090 20580 23100
rect 20636 23156 20692 23436
rect 20636 23090 20692 23100
rect 20748 23154 20804 24668
rect 20860 24052 20916 24782
rect 20860 23986 20916 23996
rect 20972 24724 21028 24734
rect 20748 23102 20750 23154
rect 20802 23102 20804 23154
rect 20188 22542 20190 22594
rect 20242 22542 20244 22594
rect 20188 22530 20244 22542
rect 20412 22932 20468 22942
rect 20300 22484 20356 22494
rect 20300 22370 20356 22428
rect 20300 22318 20302 22370
rect 20354 22318 20356 22370
rect 20300 22306 20356 22318
rect 20076 21028 20132 21038
rect 20076 20934 20132 20972
rect 20076 20804 20132 20814
rect 19964 20802 20132 20804
rect 19964 20750 20078 20802
rect 20130 20750 20132 20802
rect 19964 20748 20132 20750
rect 19628 20188 19908 20244
rect 19404 20076 19796 20132
rect 19404 19906 19460 19918
rect 19404 19854 19406 19906
rect 19458 19854 19460 19906
rect 19404 19012 19460 19854
rect 19516 19460 19572 19470
rect 19516 19234 19572 19404
rect 19516 19182 19518 19234
rect 19570 19182 19572 19234
rect 19516 19170 19572 19182
rect 19740 19234 19796 20076
rect 19740 19182 19742 19234
rect 19794 19182 19796 19234
rect 19404 18946 19460 18956
rect 19628 19010 19684 19022
rect 19628 18958 19630 19010
rect 19682 18958 19684 19010
rect 19236 16940 19348 16996
rect 19404 16996 19460 17006
rect 19628 16996 19684 18958
rect 19740 18452 19796 19182
rect 19740 18386 19796 18396
rect 19404 16994 19684 16996
rect 19404 16942 19406 16994
rect 19458 16942 19684 16994
rect 19404 16940 19684 16942
rect 19740 17332 19796 17342
rect 18732 16146 18788 16156
rect 18060 16034 18116 16044
rect 18956 15540 19012 15550
rect 18956 15446 19012 15484
rect 18732 15316 18788 15326
rect 18732 15222 18788 15260
rect 18844 15202 18900 15214
rect 18844 15150 18846 15202
rect 18898 15150 18900 15202
rect 18844 15148 18900 15150
rect 18620 15092 18900 15148
rect 18222 14924 18486 14934
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18222 14858 18486 14868
rect 17724 14588 18340 14644
rect 17052 14478 17054 14530
rect 17106 14478 17108 14530
rect 17052 14466 17108 14478
rect 17724 14420 17780 14430
rect 17724 14418 18228 14420
rect 17724 14366 17726 14418
rect 17778 14366 18228 14418
rect 17724 14364 18228 14366
rect 17724 14354 17780 14364
rect 18172 13970 18228 14364
rect 18172 13918 18174 13970
rect 18226 13918 18228 13970
rect 18172 13906 18228 13918
rect 17948 13860 18004 13870
rect 17948 13746 18004 13804
rect 18284 13748 18340 14588
rect 18620 13858 18676 15092
rect 19180 14756 19236 16940
rect 19404 16930 19460 16940
rect 19740 16772 19796 17276
rect 19852 16996 19908 20188
rect 20076 19908 20132 20748
rect 20412 20692 20468 22876
rect 20748 21476 20804 23102
rect 20972 21700 21028 24668
rect 20972 21634 21028 21644
rect 20748 21410 20804 21420
rect 20468 20636 20580 20692
rect 20412 20598 20468 20636
rect 20076 19842 20132 19852
rect 20300 19460 20356 19470
rect 20076 19234 20132 19246
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 20076 19012 20132 19182
rect 20076 18946 20132 18956
rect 20300 17106 20356 19404
rect 20524 19348 20580 20636
rect 20524 19254 20580 19292
rect 20636 19012 20692 19022
rect 20300 17054 20302 17106
rect 20354 17054 20356 17106
rect 20300 16996 20356 17054
rect 19852 16940 20020 16996
rect 19852 16772 19908 16782
rect 19740 16770 19908 16772
rect 19740 16718 19854 16770
rect 19906 16718 19908 16770
rect 19740 16716 19908 16718
rect 19852 16706 19908 16716
rect 19292 15876 19348 15886
rect 19292 15428 19348 15820
rect 19964 15540 20020 16940
rect 20300 16930 20356 16940
rect 20524 17108 20580 17118
rect 20636 17108 20692 18956
rect 20748 18452 20804 18462
rect 20748 17778 20804 18396
rect 20748 17726 20750 17778
rect 20802 17726 20804 17778
rect 20748 17714 20804 17726
rect 20748 17108 20804 17118
rect 20972 17108 21028 17118
rect 20580 17106 20804 17108
rect 20580 17054 20750 17106
rect 20802 17054 20804 17106
rect 20580 17052 20804 17054
rect 20188 16884 20244 16894
rect 19292 15314 19348 15372
rect 19740 15428 19796 15438
rect 19740 15334 19796 15372
rect 19292 15262 19294 15314
rect 19346 15262 19348 15314
rect 19292 15250 19348 15262
rect 19964 15148 20020 15484
rect 19180 14690 19236 14700
rect 19852 15092 20020 15148
rect 20076 16212 20132 16222
rect 20188 16212 20244 16828
rect 20132 16156 20244 16212
rect 20076 15148 20132 16156
rect 20300 16100 20356 16110
rect 20300 16006 20356 16044
rect 20188 15316 20244 15354
rect 20188 15250 20244 15260
rect 20524 15148 20580 17052
rect 20748 17042 20804 17052
rect 20860 17052 20972 17108
rect 20748 16212 20804 16222
rect 20860 16212 20916 17052
rect 20972 17042 21028 17052
rect 20748 16210 20916 16212
rect 20748 16158 20750 16210
rect 20802 16158 20916 16210
rect 20748 16156 20916 16158
rect 20748 16146 20804 16156
rect 20636 15540 20692 15550
rect 20636 15446 20692 15484
rect 20076 15092 20356 15148
rect 19852 14642 19908 15092
rect 19852 14590 19854 14642
rect 19906 14590 19908 14642
rect 19852 14578 19908 14590
rect 18620 13806 18622 13858
rect 18674 13806 18676 13858
rect 18620 13794 18676 13806
rect 19068 14420 19124 14430
rect 19068 13860 19124 14364
rect 19068 13766 19124 13804
rect 20300 14306 20356 15092
rect 20300 14254 20302 14306
rect 20354 14254 20356 14306
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 13682 18004 13694
rect 18060 13692 18340 13748
rect 18396 13746 18452 13758
rect 18396 13694 18398 13746
rect 18450 13694 18452 13746
rect 17052 13636 17108 13646
rect 17052 13076 17108 13580
rect 17724 13636 17780 13646
rect 17724 13076 17780 13580
rect 18060 13188 18116 13692
rect 18396 13636 18452 13694
rect 18396 13570 18452 13580
rect 20188 13746 20244 13758
rect 20188 13694 20190 13746
rect 20242 13694 20244 13746
rect 18222 13356 18486 13366
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18222 13290 18486 13300
rect 18060 13132 18340 13188
rect 17052 13074 17780 13076
rect 17052 13022 17054 13074
rect 17106 13022 17780 13074
rect 17052 13020 17780 13022
rect 17052 13010 17108 13020
rect 17612 12962 17668 13020
rect 17612 12910 17614 12962
rect 17666 12910 17668 12962
rect 17612 12898 17668 12910
rect 17388 12850 17444 12862
rect 17388 12798 17390 12850
rect 17442 12798 17444 12850
rect 17388 12740 17444 12798
rect 17948 12852 18004 12862
rect 17948 12758 18004 12796
rect 17388 12674 17444 12684
rect 17500 12738 17556 12750
rect 17500 12686 17502 12738
rect 17554 12686 17556 12738
rect 17500 12068 17556 12686
rect 18172 12740 18228 12750
rect 17724 12404 17780 12414
rect 17724 12310 17780 12348
rect 18172 12402 18228 12684
rect 18284 12738 18340 13132
rect 18956 12964 19012 12974
rect 19740 12964 19796 12974
rect 18956 12962 19796 12964
rect 18956 12910 18958 12962
rect 19010 12910 19742 12962
rect 19794 12910 19796 12962
rect 18956 12908 19796 12910
rect 18956 12898 19012 12908
rect 18396 12852 18452 12862
rect 18396 12758 18452 12796
rect 18284 12686 18286 12738
rect 18338 12686 18340 12738
rect 18284 12628 18340 12686
rect 18284 12562 18340 12572
rect 18508 12738 18564 12750
rect 18508 12686 18510 12738
rect 18562 12686 18564 12738
rect 18172 12350 18174 12402
rect 18226 12350 18228 12402
rect 18172 12338 18228 12350
rect 17052 12012 17556 12068
rect 17724 12180 17780 12190
rect 17052 11506 17108 12012
rect 17052 11454 17054 11506
rect 17106 11454 17108 11506
rect 17052 11442 17108 11454
rect 17388 11844 17444 11854
rect 16940 11106 16996 11116
rect 16828 10780 17332 10836
rect 16716 10724 16772 10734
rect 16716 10612 16772 10668
rect 16828 10612 16884 10622
rect 16716 10610 16884 10612
rect 16716 10558 16830 10610
rect 16882 10558 16884 10610
rect 16716 10556 16884 10558
rect 16716 10276 16772 10556
rect 16716 10210 16772 10220
rect 16604 9986 16660 9996
rect 16716 9826 16772 9838
rect 16716 9774 16718 9826
rect 16770 9774 16772 9826
rect 16716 8932 16772 9774
rect 16828 9492 16884 10556
rect 16828 9426 16884 9436
rect 16940 10612 16996 10622
rect 16828 9156 16884 9166
rect 16828 9062 16884 9100
rect 16716 8866 16772 8876
rect 16940 8708 16996 10556
rect 17052 9940 17108 9950
rect 17052 9828 17108 9884
rect 17052 9826 17220 9828
rect 17052 9774 17054 9826
rect 17106 9774 17220 9826
rect 17052 9772 17220 9774
rect 17052 9762 17108 9772
rect 16380 8370 16548 8372
rect 16380 8318 16382 8370
rect 16434 8318 16548 8370
rect 16380 8316 16548 8318
rect 16828 8652 16996 8708
rect 17052 9602 17108 9614
rect 17052 9550 17054 9602
rect 17106 9550 17108 9602
rect 16380 8306 16436 8316
rect 14700 7980 14980 8036
rect 13580 7698 13972 7700
rect 13580 7646 13582 7698
rect 13634 7646 13972 7698
rect 13580 7644 13972 7646
rect 13580 7634 13636 7644
rect 8988 7588 9044 7598
rect 8652 7532 8988 7588
rect 8988 7362 9044 7532
rect 13916 7474 13972 7644
rect 14700 7586 14756 7980
rect 14820 7868 15084 7878
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 14820 7802 15084 7812
rect 14700 7534 14702 7586
rect 14754 7534 14756 7586
rect 14700 7522 14756 7534
rect 13916 7422 13918 7474
rect 13970 7422 13972 7474
rect 13916 7410 13972 7422
rect 8988 7310 8990 7362
rect 9042 7310 9044 7362
rect 8988 7298 9044 7310
rect 16156 7364 16212 7374
rect 11418 7084 11682 7094
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11418 7018 11682 7028
rect 16156 6690 16212 7308
rect 16828 7362 16884 8652
rect 16940 8482 16996 8494
rect 16940 8430 16942 8482
rect 16994 8430 16996 8482
rect 16940 8370 16996 8430
rect 16940 8318 16942 8370
rect 16994 8318 16996 8370
rect 16940 8306 16996 8318
rect 16828 7310 16830 7362
rect 16882 7310 16884 7362
rect 16828 7298 16884 7310
rect 17052 7140 17108 9550
rect 17164 8482 17220 9772
rect 17164 8430 17166 8482
rect 17218 8430 17220 8482
rect 17164 8418 17220 8430
rect 17276 8036 17332 10780
rect 17388 10610 17444 11788
rect 17388 10558 17390 10610
rect 17442 10558 17444 10610
rect 17388 10500 17444 10558
rect 17612 10722 17668 10734
rect 17612 10670 17614 10722
rect 17666 10670 17668 10722
rect 17612 10612 17668 10670
rect 17612 10546 17668 10556
rect 17388 10434 17444 10444
rect 17388 9716 17444 9754
rect 17388 9650 17444 9660
rect 17388 9492 17444 9502
rect 17388 8370 17444 9436
rect 17612 9492 17668 9502
rect 17612 9266 17668 9436
rect 17612 9214 17614 9266
rect 17666 9214 17668 9266
rect 17612 9202 17668 9214
rect 17388 8318 17390 8370
rect 17442 8318 17444 8370
rect 17388 8260 17444 8318
rect 17388 8194 17444 8204
rect 17276 7970 17332 7980
rect 17724 7588 17780 12124
rect 18508 12068 18564 12686
rect 18956 12404 19012 12414
rect 18956 12310 19012 12348
rect 18508 12002 18564 12012
rect 18620 12292 18676 12302
rect 18620 12178 18676 12236
rect 18620 12126 18622 12178
rect 18674 12126 18676 12178
rect 18620 11956 18676 12126
rect 18620 11890 18676 11900
rect 18732 12290 18788 12302
rect 18732 12238 18734 12290
rect 18786 12238 18788 12290
rect 18222 11788 18486 11798
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18222 11722 18486 11732
rect 18620 11732 18676 11742
rect 17948 10836 18004 10846
rect 17948 10742 18004 10780
rect 18620 10834 18676 11676
rect 18620 10782 18622 10834
rect 18674 10782 18676 10834
rect 18620 10770 18676 10782
rect 18508 10610 18564 10622
rect 18508 10558 18510 10610
rect 18562 10558 18564 10610
rect 18508 10388 18564 10558
rect 18508 10322 18564 10332
rect 18222 10220 18486 10230
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18222 10154 18486 10164
rect 17836 10052 17892 10062
rect 17836 9826 17892 9996
rect 18620 9940 18676 9950
rect 18620 9846 18676 9884
rect 17836 9774 17838 9826
rect 17890 9774 17892 9826
rect 17836 9762 17892 9774
rect 18060 9716 18116 9726
rect 18060 9266 18116 9660
rect 18732 9380 18788 12238
rect 19068 10724 19124 12908
rect 19740 12898 19796 12908
rect 20188 12964 20244 13694
rect 20188 12898 20244 12908
rect 19292 12738 19348 12750
rect 19292 12686 19294 12738
rect 19346 12686 19348 12738
rect 19292 12292 19348 12686
rect 19292 12226 19348 12236
rect 19628 12740 19684 12750
rect 19516 12178 19572 12190
rect 19516 12126 19518 12178
rect 19570 12126 19572 12178
rect 19292 12068 19348 12078
rect 19516 12068 19572 12126
rect 19180 12012 19292 12068
rect 19348 12012 19572 12068
rect 19180 11506 19236 12012
rect 19292 12002 19348 12012
rect 19180 11454 19182 11506
rect 19234 11454 19236 11506
rect 19180 11442 19236 11454
rect 19628 11394 19684 12684
rect 20188 12738 20244 12750
rect 20188 12686 20190 12738
rect 20242 12686 20244 12738
rect 20188 12628 20244 12686
rect 19852 12290 19908 12302
rect 19852 12238 19854 12290
rect 19906 12238 19908 12290
rect 19628 11342 19630 11394
rect 19682 11342 19684 11394
rect 19628 11330 19684 11342
rect 19740 11844 19796 11854
rect 19852 11844 19908 12238
rect 19796 11788 19908 11844
rect 20188 11844 20244 12572
rect 19068 10658 19124 10668
rect 19628 10836 19684 10846
rect 19740 10836 19796 11788
rect 20188 11778 20244 11788
rect 19964 11508 20020 11518
rect 20300 11508 20356 14254
rect 20412 15092 20580 15148
rect 20412 11954 20468 15092
rect 20748 14644 20804 14654
rect 20748 14550 20804 14588
rect 20860 14308 20916 16156
rect 20748 14252 20916 14308
rect 20524 12964 20580 12974
rect 20524 12068 20580 12908
rect 20524 12066 20692 12068
rect 20524 12014 20526 12066
rect 20578 12014 20692 12066
rect 20524 12012 20692 12014
rect 20524 12002 20580 12012
rect 20412 11902 20414 11954
rect 20466 11902 20468 11954
rect 20412 11890 20468 11902
rect 20300 11452 20580 11508
rect 19628 10834 19796 10836
rect 19628 10782 19630 10834
rect 19682 10782 19796 10834
rect 19628 10780 19796 10782
rect 19852 11170 19908 11182
rect 19852 11118 19854 11170
rect 19906 11118 19908 11170
rect 19516 10164 19572 10174
rect 19068 9492 19124 9502
rect 18060 9214 18062 9266
rect 18114 9214 18116 9266
rect 18060 9202 18116 9214
rect 18172 9324 19012 9380
rect 18172 9266 18228 9324
rect 18172 9214 18174 9266
rect 18226 9214 18228 9266
rect 18172 9202 18228 9214
rect 17948 9156 18004 9166
rect 17948 9062 18004 9100
rect 18844 9156 18900 9166
rect 18620 9042 18676 9054
rect 18620 8990 18622 9042
rect 18674 8990 18676 9042
rect 17836 8932 17892 8942
rect 17836 8370 17892 8876
rect 18222 8652 18486 8662
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18222 8586 18486 8596
rect 17836 8318 17838 8370
rect 17890 8318 17892 8370
rect 17836 8306 17892 8318
rect 18172 8372 18228 8382
rect 18172 8278 18228 8316
rect 18620 8260 18676 8990
rect 18844 8370 18900 9100
rect 18844 8318 18846 8370
rect 18898 8318 18900 8370
rect 18844 8306 18900 8318
rect 18620 8194 18676 8204
rect 17724 7522 17780 7532
rect 16156 6638 16158 6690
rect 16210 6638 16212 6690
rect 16156 6626 16212 6638
rect 16828 7084 17108 7140
rect 18222 7084 18486 7094
rect 16828 6690 16884 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18222 7018 18486 7028
rect 18956 6802 19012 9324
rect 19068 9266 19124 9436
rect 19068 9214 19070 9266
rect 19122 9214 19124 9266
rect 19068 9202 19124 9214
rect 19516 9268 19572 10108
rect 19628 9492 19684 10780
rect 19852 9940 19908 11118
rect 19964 10610 20020 11452
rect 20076 11396 20132 11406
rect 20076 11302 20132 11340
rect 20188 11394 20244 11406
rect 20188 11342 20190 11394
rect 20242 11342 20244 11394
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19964 10546 20020 10558
rect 20188 10612 20244 11342
rect 20300 10836 20356 10846
rect 20300 10742 20356 10780
rect 20188 10546 20244 10556
rect 20300 10610 20356 10622
rect 20300 10558 20302 10610
rect 20354 10558 20356 10610
rect 20300 10500 20356 10558
rect 20524 10500 20580 11452
rect 20300 10434 20356 10444
rect 20412 10444 20580 10500
rect 19852 9874 19908 9884
rect 19628 9426 19684 9436
rect 19964 9268 20020 9278
rect 19516 9266 20020 9268
rect 19516 9214 19518 9266
rect 19570 9214 19966 9266
rect 20018 9214 20020 9266
rect 19516 9212 20020 9214
rect 19516 9202 19572 9212
rect 19964 9202 20020 9212
rect 19292 8260 19348 8270
rect 19292 8166 19348 8204
rect 20076 8258 20132 8270
rect 20076 8206 20078 8258
rect 20130 8206 20132 8258
rect 19740 8148 19796 8158
rect 19740 8054 19796 8092
rect 19852 7588 19908 7598
rect 20076 7588 20132 8206
rect 20300 8146 20356 8158
rect 20300 8094 20302 8146
rect 20354 8094 20356 8146
rect 20300 7700 20356 8094
rect 20300 7634 20356 7644
rect 19852 7586 20132 7588
rect 19852 7534 19854 7586
rect 19906 7534 20132 7586
rect 19852 7532 20132 7534
rect 19852 7522 19908 7532
rect 19068 7364 19124 7374
rect 19068 7270 19124 7308
rect 18956 6750 18958 6802
rect 19010 6750 19012 6802
rect 18956 6738 19012 6750
rect 19516 6802 19572 6814
rect 19516 6750 19518 6802
rect 19570 6750 19572 6802
rect 16828 6638 16830 6690
rect 16882 6638 16884 6690
rect 16828 6626 16884 6638
rect 19516 6692 19572 6750
rect 19516 6626 19572 6636
rect 7644 6290 7700 6300
rect 8016 6300 8280 6310
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8016 6234 8280 6244
rect 14820 6300 15084 6310
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 14820 6234 15084 6244
rect 5852 6130 6020 6132
rect 5852 6078 5854 6130
rect 5906 6078 6020 6130
rect 5852 6076 6020 6078
rect 18732 6132 18788 6142
rect 5852 6066 5908 6076
rect 18732 6038 18788 6076
rect 19852 5906 19908 5918
rect 19852 5854 19854 5906
rect 19906 5854 19908 5906
rect 19852 5796 19908 5854
rect 19852 5730 19908 5740
rect 4614 5516 4878 5526
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4614 5450 4878 5460
rect 11418 5516 11682 5526
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11418 5450 11682 5460
rect 18222 5516 18486 5526
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18222 5450 18486 5460
rect 18732 5124 18788 5134
rect 18732 5030 18788 5068
rect 19740 5012 19796 5022
rect 19180 5010 19796 5012
rect 19180 4958 19742 5010
rect 19794 4958 19796 5010
rect 19180 4956 19796 4958
rect 19068 4900 19124 4910
rect 18844 4898 19124 4900
rect 18844 4846 19070 4898
rect 19122 4846 19124 4898
rect 18844 4844 19124 4846
rect 8016 4732 8280 4742
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8016 4666 8280 4676
rect 14820 4732 15084 4742
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 14820 4666 15084 4676
rect 11788 4452 11844 4462
rect 18508 4452 18564 4462
rect 18844 4452 18900 4844
rect 19068 4834 19124 4844
rect 11788 4450 12404 4452
rect 11788 4398 11790 4450
rect 11842 4398 12404 4450
rect 11788 4396 12404 4398
rect 11788 4386 11844 4396
rect 11228 4338 11284 4350
rect 11228 4286 11230 4338
rect 11282 4286 11284 4338
rect 10780 4226 10836 4238
rect 10780 4174 10782 4226
rect 10834 4174 10836 4226
rect 4614 3948 4878 3958
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4614 3882 4878 3892
rect 7644 3556 7700 3566
rect 6972 3554 7700 3556
rect 6972 3502 7646 3554
rect 7698 3502 7700 3554
rect 6972 3500 7700 3502
rect 4956 3444 5012 3454
rect 4620 3330 4676 3342
rect 4620 3278 4622 3330
rect 4674 3278 4676 3330
rect 4060 2606 4062 2658
rect 4114 2606 4116 2658
rect 4060 2594 4116 2606
rect 4284 2772 4340 2782
rect 3612 2212 3668 2222
rect 3612 1874 3668 2156
rect 4060 1986 4116 1998
rect 4060 1934 4062 1986
rect 4114 1934 4116 1986
rect 3612 1822 3614 1874
rect 3666 1822 3668 1874
rect 3612 1810 3668 1822
rect 3948 1876 4004 1886
rect 3948 1204 4004 1820
rect 4060 1652 4116 1934
rect 4284 1874 4340 2716
rect 4620 2548 4676 3278
rect 4284 1822 4286 1874
rect 4338 1822 4340 1874
rect 4284 1810 4340 1822
rect 4396 2492 4676 2548
rect 4396 1652 4452 2492
rect 4614 2380 4878 2390
rect 4670 2324 4718 2380
rect 4774 2324 4822 2380
rect 4614 2314 4878 2324
rect 4732 1986 4788 1998
rect 4732 1934 4734 1986
rect 4786 1934 4788 1986
rect 4732 1876 4788 1934
rect 4732 1810 4788 1820
rect 4956 1874 5012 3388
rect 4956 1822 4958 1874
rect 5010 1822 5012 1874
rect 4956 1810 5012 1822
rect 5180 3442 5236 3454
rect 5180 3390 5182 3442
rect 5234 3390 5236 3442
rect 5180 1876 5236 3390
rect 5628 3442 5684 3454
rect 5628 3390 5630 3442
rect 5682 3390 5684 3442
rect 5404 1876 5460 1886
rect 5180 1820 5404 1876
rect 5628 1876 5684 3390
rect 5740 3444 5796 3482
rect 5740 3378 5796 3388
rect 6412 3444 6468 3454
rect 5964 3330 6020 3342
rect 6300 3332 6356 3342
rect 5964 3278 5966 3330
rect 6018 3278 6020 3330
rect 5964 2658 6020 3278
rect 5964 2606 5966 2658
rect 6018 2606 6020 2658
rect 5964 2594 6020 2606
rect 6076 3330 6356 3332
rect 6076 3278 6302 3330
rect 6354 3278 6356 3330
rect 6076 3276 6356 3278
rect 6076 1986 6132 3276
rect 6300 3266 6356 3276
rect 6188 2996 6244 3006
rect 6412 2996 6468 3388
rect 6860 3332 6916 3342
rect 6188 2994 6468 2996
rect 6188 2942 6190 2994
rect 6242 2942 6468 2994
rect 6188 2940 6468 2942
rect 6524 3330 6916 3332
rect 6524 3278 6862 3330
rect 6914 3278 6916 3330
rect 6524 3276 6916 3278
rect 6188 2930 6244 2940
rect 6188 2772 6244 2782
rect 6188 2678 6244 2716
rect 6300 2770 6356 2782
rect 6300 2718 6302 2770
rect 6354 2718 6356 2770
rect 6300 2212 6356 2718
rect 6300 2146 6356 2156
rect 6076 1934 6078 1986
rect 6130 1934 6132 1986
rect 5740 1876 5796 1886
rect 5628 1874 5796 1876
rect 5628 1822 5742 1874
rect 5794 1822 5796 1874
rect 5628 1820 5796 1822
rect 4060 1596 4788 1652
rect 3948 1148 4116 1204
rect 4060 400 4116 1148
rect 4732 400 4788 1596
rect 5404 400 5460 1820
rect 5740 1810 5796 1820
rect 6076 400 6132 1934
rect 6524 1988 6580 3276
rect 6860 3266 6916 3276
rect 6524 1986 6692 1988
rect 6524 1934 6526 1986
rect 6578 1934 6692 1986
rect 6524 1932 6692 1934
rect 6524 1922 6580 1932
rect 6636 1540 6692 1932
rect 6748 1876 6804 1886
rect 6972 1876 7028 3500
rect 7644 3490 7700 3500
rect 8764 3556 8820 3566
rect 7756 3442 7812 3454
rect 7756 3390 7758 3442
rect 7810 3390 7812 3442
rect 7420 3332 7476 3342
rect 7196 3330 7476 3332
rect 7196 3278 7422 3330
rect 7474 3278 7476 3330
rect 7196 3276 7476 3278
rect 7196 1988 7252 3276
rect 7420 3266 7476 3276
rect 7756 2884 7812 3390
rect 8016 3164 8280 3174
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8016 3098 8280 3108
rect 7420 2828 7812 2884
rect 8092 2996 8148 3006
rect 7196 1986 7364 1988
rect 7196 1934 7198 1986
rect 7250 1934 7364 1986
rect 7196 1932 7364 1934
rect 7196 1922 7252 1932
rect 6748 1874 7028 1876
rect 6748 1822 6750 1874
rect 6802 1822 7028 1874
rect 6748 1820 7028 1822
rect 6748 1810 6804 1820
rect 7308 1540 7364 1932
rect 7420 1874 7476 2828
rect 7756 2658 7812 2670
rect 7756 2606 7758 2658
rect 7810 2606 7812 2658
rect 7756 1988 7812 2606
rect 7868 1988 7924 1998
rect 7756 1986 7924 1988
rect 7756 1934 7870 1986
rect 7922 1934 7924 1986
rect 7756 1932 7924 1934
rect 7420 1822 7422 1874
rect 7474 1822 7476 1874
rect 7420 1810 7476 1822
rect 6636 1484 6804 1540
rect 7308 1484 7476 1540
rect 6748 400 6804 1484
rect 7420 400 7476 1484
rect 7868 1428 7924 1932
rect 8092 1874 8148 2940
rect 8204 2658 8260 2670
rect 8204 2606 8206 2658
rect 8258 2606 8260 2658
rect 8204 1988 8260 2606
rect 8652 2658 8708 2670
rect 8652 2606 8654 2658
rect 8706 2606 8708 2658
rect 8540 1988 8596 1998
rect 8204 1986 8596 1988
rect 8204 1934 8542 1986
rect 8594 1934 8596 1986
rect 8204 1932 8596 1934
rect 8092 1822 8094 1874
rect 8146 1822 8148 1874
rect 8092 1810 8148 1822
rect 8016 1596 8280 1606
rect 8072 1540 8120 1596
rect 8176 1540 8224 1596
rect 8016 1530 8280 1540
rect 7868 1372 8148 1428
rect 8092 400 8148 1372
rect 8540 1316 8596 1932
rect 8652 1652 8708 2606
rect 8764 1874 8820 3500
rect 9660 3556 9716 3566
rect 9660 3462 9716 3500
rect 10220 3442 10276 3454
rect 10220 3390 10222 3442
rect 10274 3390 10276 3442
rect 10220 3220 10276 3390
rect 10780 3388 10836 4174
rect 11004 3668 11060 3678
rect 11228 3668 11284 4286
rect 11564 4338 11620 4350
rect 11564 4286 11566 4338
rect 11618 4286 11620 4338
rect 11564 4116 11620 4286
rect 11676 4228 11732 4238
rect 12236 4228 12292 4238
rect 11676 4134 11732 4172
rect 12012 4226 12292 4228
rect 12012 4174 12238 4226
rect 12290 4174 12292 4226
rect 12012 4172 12292 4174
rect 11564 4050 11620 4060
rect 11418 3948 11682 3958
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11418 3882 11682 3892
rect 11004 3666 11284 3668
rect 11004 3614 11006 3666
rect 11058 3614 11284 3666
rect 11004 3612 11284 3614
rect 11004 3556 11060 3612
rect 11004 3490 11060 3500
rect 11788 3556 11844 3566
rect 11788 3462 11844 3500
rect 12012 3388 12068 4172
rect 12236 4162 12292 4172
rect 10220 3154 10276 3164
rect 10668 3332 10836 3388
rect 11900 3332 12068 3388
rect 12124 4004 12180 4014
rect 12124 3444 12180 3948
rect 12348 3442 12404 4396
rect 18060 4450 18564 4452
rect 18060 4398 18510 4450
rect 18562 4398 18564 4450
rect 18060 4396 18564 4398
rect 17836 4228 17892 4238
rect 17836 4226 18004 4228
rect 17836 4174 17838 4226
rect 17890 4174 18004 4226
rect 17836 4172 18004 4174
rect 17836 4162 17892 4172
rect 13020 3780 13076 3790
rect 13020 3666 13076 3724
rect 13020 3614 13022 3666
rect 13074 3614 13076 3666
rect 13020 3602 13076 3614
rect 17612 3612 17892 3668
rect 12348 3390 12350 3442
rect 12402 3390 12404 3442
rect 12348 3388 12404 3390
rect 12124 3378 12180 3388
rect 12236 3332 12404 3388
rect 15148 3554 15204 3566
rect 15148 3502 15150 3554
rect 15202 3502 15204 3554
rect 9100 2996 9156 3006
rect 9100 2994 9828 2996
rect 9100 2942 9102 2994
rect 9154 2942 9828 2994
rect 9100 2940 9828 2942
rect 9100 2930 9156 2940
rect 9660 2770 9716 2782
rect 9660 2718 9662 2770
rect 9714 2718 9716 2770
rect 9660 2212 9716 2718
rect 8764 1822 8766 1874
rect 8818 1822 8820 1874
rect 8764 1810 8820 1822
rect 9436 2156 9716 2212
rect 9436 1652 9492 2156
rect 9660 1988 9716 1998
rect 9772 1988 9828 2940
rect 9996 2882 10052 2894
rect 9996 2830 9998 2882
rect 10050 2830 10052 2882
rect 9996 2772 10052 2830
rect 9996 2706 10052 2716
rect 10556 2772 10612 2782
rect 10556 2678 10612 2716
rect 10444 2548 10500 2558
rect 10668 2548 10724 3332
rect 11676 2996 11732 3006
rect 11676 2770 11732 2940
rect 11900 2884 11956 3332
rect 12012 2996 12068 3006
rect 12236 2996 12292 3332
rect 13580 3330 13636 3342
rect 13580 3278 13582 3330
rect 13634 3278 13636 3330
rect 12012 2994 12292 2996
rect 12012 2942 12014 2994
rect 12066 2942 12292 2994
rect 12012 2940 12292 2942
rect 12572 2996 12628 3006
rect 12012 2930 12068 2940
rect 12572 2902 12628 2940
rect 11676 2718 11678 2770
rect 11730 2718 11732 2770
rect 11676 2706 11732 2718
rect 11788 2828 11956 2884
rect 11116 2660 11172 2670
rect 11452 2660 11508 2670
rect 11116 2658 11508 2660
rect 11116 2606 11118 2658
rect 11170 2606 11454 2658
rect 11506 2606 11508 2658
rect 11116 2604 11508 2606
rect 11116 2594 11172 2604
rect 11452 2594 11508 2604
rect 9660 1986 9828 1988
rect 9660 1934 9662 1986
rect 9714 1934 9828 1986
rect 9660 1932 9828 1934
rect 9660 1922 9716 1932
rect 8652 1596 9492 1652
rect 9772 1652 9828 1932
rect 9884 2546 10500 2548
rect 9884 2494 10446 2546
rect 10498 2494 10500 2546
rect 9884 2492 10500 2494
rect 9884 1874 9940 2492
rect 10444 2482 10500 2492
rect 10556 2492 10724 2548
rect 10780 2546 10836 2558
rect 10780 2494 10782 2546
rect 10834 2494 10836 2546
rect 10556 2100 10612 2492
rect 10780 2212 10836 2494
rect 10780 2146 10836 2156
rect 11004 2546 11060 2558
rect 11004 2494 11006 2546
rect 11058 2494 11060 2546
rect 10332 2044 10612 2100
rect 10332 1986 10388 2044
rect 10332 1934 10334 1986
rect 10386 1934 10388 1986
rect 10332 1922 10388 1934
rect 9884 1822 9886 1874
rect 9938 1822 9940 1874
rect 9884 1810 9940 1822
rect 10444 1652 10500 2044
rect 11004 1988 11060 2494
rect 10556 1932 11060 1988
rect 11228 2436 11284 2446
rect 11228 1988 11284 2380
rect 11418 2380 11682 2390
rect 11474 2324 11522 2380
rect 11578 2324 11626 2380
rect 11418 2314 11682 2324
rect 11676 1988 11732 1998
rect 11788 1988 11844 2828
rect 12684 2772 12740 2782
rect 11228 1986 11508 1988
rect 11228 1934 11230 1986
rect 11282 1934 11508 1986
rect 11228 1932 11508 1934
rect 10556 1874 10612 1932
rect 11228 1922 11284 1932
rect 10556 1822 10558 1874
rect 10610 1822 10612 1874
rect 10556 1810 10612 1822
rect 10892 1764 10948 1802
rect 10892 1698 10948 1708
rect 9772 1596 10164 1652
rect 10444 1596 10836 1652
rect 8540 1260 8820 1316
rect 8764 400 8820 1260
rect 9436 400 9492 1596
rect 10108 400 10164 1596
rect 10780 400 10836 1596
rect 11452 400 11508 1932
rect 11676 1986 11844 1988
rect 11676 1934 11678 1986
rect 11730 1934 11844 1986
rect 11676 1932 11844 1934
rect 11676 1922 11732 1932
rect 11788 1652 11844 1932
rect 11900 2770 12740 2772
rect 11900 2718 12686 2770
rect 12738 2718 12740 2770
rect 11900 2716 12740 2718
rect 11900 1874 11956 2716
rect 12684 2706 12740 2716
rect 13580 2660 13636 3278
rect 14820 3164 15084 3174
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 14820 3098 15084 3108
rect 13580 2594 13636 2604
rect 13692 2660 13748 2670
rect 13692 2658 13860 2660
rect 13692 2606 13694 2658
rect 13746 2606 13860 2658
rect 13692 2604 13860 2606
rect 13692 2594 13748 2604
rect 12572 2546 12628 2558
rect 12572 2494 12574 2546
rect 12626 2494 12628 2546
rect 12348 2212 12404 2222
rect 12348 1986 12404 2156
rect 12348 1934 12350 1986
rect 12402 1934 12404 1986
rect 12348 1922 12404 1934
rect 11900 1822 11902 1874
rect 11954 1822 11956 1874
rect 11900 1810 11956 1822
rect 12572 1874 12628 2494
rect 12908 2548 12964 2558
rect 12908 2454 12964 2492
rect 13132 2546 13188 2558
rect 13132 2494 13134 2546
rect 13186 2494 13188 2546
rect 12572 1822 12574 1874
rect 12626 1822 12628 1874
rect 12572 1810 12628 1822
rect 12796 2212 12852 2222
rect 13132 2212 13188 2494
rect 13132 2156 13748 2212
rect 11788 1596 12180 1652
rect 12124 400 12180 1596
rect 12796 400 12852 2156
rect 13468 1988 13524 1998
rect 13468 1894 13524 1932
rect 13692 1874 13748 2156
rect 13804 1988 13860 2604
rect 14140 2658 14196 2670
rect 14140 2606 14142 2658
rect 14194 2606 14196 2658
rect 14140 2212 14196 2606
rect 14812 2658 14868 2670
rect 14812 2606 14814 2658
rect 14866 2606 14868 2658
rect 14140 2146 14196 2156
rect 14364 2548 14420 2558
rect 13916 1988 13972 1998
rect 13804 1986 13972 1988
rect 13804 1934 13918 1986
rect 13970 1934 13972 1986
rect 13804 1932 13972 1934
rect 13692 1822 13694 1874
rect 13746 1822 13748 1874
rect 13692 1810 13748 1822
rect 13916 1540 13972 1932
rect 13468 1484 13972 1540
rect 14140 1988 14196 1998
rect 13468 400 13524 1484
rect 14140 400 14196 1932
rect 14364 1874 14420 2492
rect 14700 1988 14756 1998
rect 14700 1894 14756 1932
rect 14364 1822 14366 1874
rect 14418 1822 14420 1874
rect 14364 1810 14420 1822
rect 14812 1764 14868 2606
rect 15036 1874 15092 1886
rect 15036 1822 15038 1874
rect 15090 1822 15092 1874
rect 15036 1764 15092 1822
rect 15148 1876 15204 3502
rect 17276 3556 17332 3566
rect 17612 3556 17668 3612
rect 17276 3554 17668 3556
rect 17276 3502 17278 3554
rect 17330 3502 17668 3554
rect 17276 3500 17668 3502
rect 17276 3490 17332 3500
rect 16268 3442 16324 3454
rect 16268 3390 16270 3442
rect 16322 3390 16324 3442
rect 16268 2884 16324 3390
rect 17724 3442 17780 3454
rect 17724 3390 17726 3442
rect 17778 3390 17780 3442
rect 17724 3388 17780 3390
rect 16044 2828 16324 2884
rect 17276 3332 17780 3388
rect 15484 2658 15540 2670
rect 15484 2606 15486 2658
rect 15538 2606 15540 2658
rect 15372 1876 15428 1886
rect 15148 1874 15428 1876
rect 15148 1822 15374 1874
rect 15426 1822 15428 1874
rect 15148 1820 15428 1822
rect 15372 1810 15428 1820
rect 15484 1876 15540 2606
rect 15708 1876 15764 1886
rect 15484 1874 15764 1876
rect 15484 1822 15710 1874
rect 15762 1822 15764 1874
rect 15484 1820 15764 1822
rect 14700 1708 15092 1764
rect 14700 1428 14756 1708
rect 14820 1596 15084 1606
rect 14876 1540 14924 1596
rect 14980 1540 15028 1596
rect 14820 1530 15084 1540
rect 14700 1372 14868 1428
rect 14812 400 14868 1372
rect 15484 400 15540 1820
rect 15708 1810 15764 1820
rect 16044 1874 16100 2828
rect 16268 2660 16324 2670
rect 16268 2566 16324 2604
rect 16716 2658 16772 2670
rect 16716 2606 16718 2658
rect 16770 2606 16772 2658
rect 16044 1822 16046 1874
rect 16098 1822 16100 1874
rect 16044 1810 16100 1822
rect 16156 1876 16212 1886
rect 16716 1876 16772 2606
rect 17052 2660 17108 2670
rect 16940 1876 16996 1886
rect 16716 1820 16940 1876
rect 16156 400 16212 1820
rect 16940 1782 16996 1820
rect 17052 1540 17108 2604
rect 17276 1874 17332 3332
rect 17500 3220 17556 3230
rect 17500 2994 17556 3164
rect 17500 2942 17502 2994
rect 17554 2942 17556 2994
rect 17500 2930 17556 2942
rect 17724 3108 17780 3118
rect 17388 2772 17444 2782
rect 17388 2678 17444 2716
rect 17612 2660 17668 2670
rect 17612 1986 17668 2604
rect 17612 1934 17614 1986
rect 17666 1934 17668 1986
rect 17612 1922 17668 1934
rect 17276 1822 17278 1874
rect 17330 1822 17332 1874
rect 17276 1810 17332 1822
rect 17724 1764 17780 3052
rect 17836 1876 17892 3612
rect 17948 3108 18004 4172
rect 17948 3042 18004 3052
rect 17948 2884 18004 2894
rect 18060 2884 18116 4396
rect 18508 4386 18564 4396
rect 18732 4450 18900 4452
rect 18732 4398 18846 4450
rect 18898 4398 18900 4450
rect 18732 4396 18900 4398
rect 18284 4226 18340 4238
rect 18284 4174 18286 4226
rect 18338 4174 18340 4226
rect 18284 4116 18340 4174
rect 18284 4050 18340 4060
rect 18222 3948 18486 3958
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18222 3882 18486 3892
rect 17948 2882 18116 2884
rect 17948 2830 17950 2882
rect 18002 2830 18116 2882
rect 17948 2828 18116 2830
rect 18396 2884 18452 2894
rect 17948 2818 18004 2828
rect 18396 2770 18452 2828
rect 18396 2718 18398 2770
rect 18450 2718 18452 2770
rect 18396 2706 18452 2718
rect 18620 2658 18676 2670
rect 18620 2606 18622 2658
rect 18674 2606 18676 2658
rect 18222 2380 18486 2390
rect 18278 2324 18326 2380
rect 18382 2324 18430 2380
rect 18222 2314 18486 2324
rect 18172 2212 18228 2222
rect 17948 1876 18004 1886
rect 17836 1874 18004 1876
rect 17836 1822 17950 1874
rect 18002 1822 18004 1874
rect 17836 1820 18004 1822
rect 17948 1810 18004 1820
rect 16828 1484 17108 1540
rect 17500 1708 17780 1764
rect 16828 400 16884 1484
rect 17500 400 17556 1708
rect 18172 400 18228 2156
rect 18620 1986 18676 2606
rect 18620 1934 18622 1986
rect 18674 1934 18676 1986
rect 18620 1922 18676 1934
rect 18508 1876 18564 1886
rect 18508 1782 18564 1820
rect 18732 1540 18788 4396
rect 18844 4386 18900 4396
rect 19180 4450 19236 4956
rect 19740 4946 19796 4956
rect 19852 4900 19908 4910
rect 19628 4788 19684 4798
rect 19628 4562 19684 4732
rect 19628 4510 19630 4562
rect 19682 4510 19684 4562
rect 19628 4498 19684 4510
rect 19180 4398 19182 4450
rect 19234 4398 19236 4450
rect 18844 3330 18900 3342
rect 18844 3278 18846 3330
rect 18898 3278 18900 3330
rect 18844 1876 18900 3278
rect 19180 3220 19236 4398
rect 19404 4338 19460 4350
rect 19404 4286 19406 4338
rect 19458 4286 19460 4338
rect 19292 4116 19348 4126
rect 19292 3554 19348 4060
rect 19292 3502 19294 3554
rect 19346 3502 19348 3554
rect 19292 3490 19348 3502
rect 19404 3444 19460 4286
rect 19740 4114 19796 4126
rect 19740 4062 19742 4114
rect 19794 4062 19796 4114
rect 19740 3668 19796 4062
rect 19740 3602 19796 3612
rect 19852 3556 19908 4844
rect 19964 3780 20020 7532
rect 20300 7364 20356 7374
rect 20412 7364 20468 10444
rect 20636 10388 20692 12012
rect 20748 11396 20804 14252
rect 21084 14196 21140 25116
rect 21196 24948 21252 24958
rect 21420 24948 21476 25340
rect 21624 25116 21888 25126
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21624 25050 21888 25060
rect 22092 25060 22148 33964
rect 22428 33908 22484 33918
rect 22876 33908 22932 34638
rect 22484 33852 22932 33908
rect 22988 35588 23044 35598
rect 22428 33842 22484 33852
rect 22316 33460 22372 33470
rect 22316 33236 22372 33404
rect 22428 33348 22484 33358
rect 22428 33254 22484 33292
rect 22652 33346 22708 33852
rect 22652 33294 22654 33346
rect 22706 33294 22708 33346
rect 22316 33122 22372 33180
rect 22652 33236 22708 33294
rect 22652 33170 22708 33180
rect 22876 33234 22932 33246
rect 22876 33182 22878 33234
rect 22930 33182 22932 33234
rect 22316 33070 22318 33122
rect 22370 33070 22372 33122
rect 22316 32004 22372 33070
rect 22540 33124 22596 33134
rect 22540 33030 22596 33068
rect 22876 33124 22932 33182
rect 22876 33058 22932 33068
rect 22988 32900 23044 35532
rect 22428 32844 23044 32900
rect 23100 32900 23156 36540
rect 23436 36482 23492 36494
rect 23436 36430 23438 36482
rect 23490 36430 23492 36482
rect 23436 35700 23492 36430
rect 23772 35700 23828 35710
rect 23436 35698 23828 35700
rect 23436 35646 23774 35698
rect 23826 35646 23828 35698
rect 23436 35644 23828 35646
rect 23660 35476 23716 35486
rect 22428 32228 22484 32844
rect 23100 32834 23156 32844
rect 23212 35364 23268 35374
rect 22540 32452 22596 32462
rect 22540 32450 23156 32452
rect 22540 32398 22542 32450
rect 22594 32398 23156 32450
rect 22540 32396 23156 32398
rect 22540 32386 22596 32396
rect 22428 32172 22708 32228
rect 22316 31938 22372 31948
rect 22204 31666 22260 31678
rect 22204 31614 22206 31666
rect 22258 31614 22260 31666
rect 22204 25620 22260 31614
rect 22540 31666 22596 31678
rect 22540 31614 22542 31666
rect 22594 31614 22596 31666
rect 22540 31106 22596 31614
rect 22540 31054 22542 31106
rect 22594 31054 22596 31106
rect 22540 31042 22596 31054
rect 22540 29986 22596 29998
rect 22540 29934 22542 29986
rect 22594 29934 22596 29986
rect 22540 29876 22596 29934
rect 22540 29810 22596 29820
rect 22540 29652 22596 29662
rect 22428 29596 22540 29652
rect 22316 29540 22372 29550
rect 22316 27186 22372 29484
rect 22316 27134 22318 27186
rect 22370 27134 22372 27186
rect 22316 27122 22372 27134
rect 22428 26908 22484 29596
rect 22540 29586 22596 29596
rect 22540 28420 22596 28430
rect 22540 27746 22596 28364
rect 22540 27694 22542 27746
rect 22594 27694 22596 27746
rect 22540 27682 22596 27694
rect 22428 26852 22596 26908
rect 22204 25554 22260 25564
rect 22316 26180 22372 26190
rect 22316 25284 22372 26124
rect 22316 25218 22372 25228
rect 22092 25004 22484 25060
rect 21420 24892 21588 24948
rect 21196 23716 21252 24892
rect 21420 24724 21476 24734
rect 21196 23650 21252 23660
rect 21308 24722 21476 24724
rect 21308 24670 21422 24722
rect 21474 24670 21476 24722
rect 21308 24668 21476 24670
rect 21196 23042 21252 23054
rect 21196 22990 21198 23042
rect 21250 22990 21252 23042
rect 21196 22932 21252 22990
rect 21196 22866 21252 22876
rect 21308 20132 21364 24668
rect 21420 24658 21476 24668
rect 21532 24610 21588 24892
rect 21532 24558 21534 24610
rect 21586 24558 21588 24610
rect 21532 24546 21588 24558
rect 21644 24722 21700 24734
rect 21644 24670 21646 24722
rect 21698 24670 21700 24722
rect 21420 24388 21476 24398
rect 21644 24388 21700 24670
rect 21476 24332 21700 24388
rect 22204 24722 22260 24734
rect 22204 24670 22206 24722
rect 22258 24670 22260 24722
rect 21420 24050 21476 24332
rect 21420 23998 21422 24050
rect 21474 23998 21476 24050
rect 21420 23986 21476 23998
rect 22092 24162 22148 24174
rect 22092 24110 22094 24162
rect 22146 24110 22148 24162
rect 21868 23716 21924 23726
rect 22092 23716 22148 24110
rect 21868 23714 22148 23716
rect 21868 23662 21870 23714
rect 21922 23662 22148 23714
rect 21868 23660 22148 23662
rect 21868 23650 21924 23660
rect 21624 23548 21888 23558
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21624 23482 21888 23492
rect 21420 23380 21476 23390
rect 21420 22146 21476 23324
rect 21980 23268 22036 23278
rect 21868 23042 21924 23054
rect 21868 22990 21870 23042
rect 21922 22990 21924 23042
rect 21868 22930 21924 22990
rect 21868 22878 21870 22930
rect 21922 22878 21924 22930
rect 21868 22866 21924 22878
rect 21868 22484 21924 22494
rect 21980 22484 22036 23212
rect 21868 22482 22036 22484
rect 21868 22430 21870 22482
rect 21922 22430 22036 22482
rect 21868 22428 22036 22430
rect 21868 22418 21924 22428
rect 21420 22094 21422 22146
rect 21474 22094 21476 22146
rect 21420 21812 21476 22094
rect 21624 21980 21888 21990
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21624 21914 21888 21924
rect 21420 20580 21476 21756
rect 21868 21476 21924 21486
rect 21868 21382 21924 21420
rect 21420 20486 21476 20524
rect 21624 20412 21888 20422
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21624 20346 21888 20356
rect 21196 20076 21924 20132
rect 21196 17780 21252 20076
rect 21308 19908 21364 19918
rect 21308 18338 21364 19852
rect 21644 19460 21700 19470
rect 21644 19234 21700 19404
rect 21644 19182 21646 19234
rect 21698 19182 21700 19234
rect 21644 19170 21700 19182
rect 21868 19234 21924 20076
rect 21868 19182 21870 19234
rect 21922 19182 21924 19234
rect 21868 19170 21924 19182
rect 21532 19124 21588 19134
rect 21308 18286 21310 18338
rect 21362 18286 21364 18338
rect 21308 18274 21364 18286
rect 21420 19068 21532 19124
rect 21308 17780 21364 17790
rect 21196 17778 21364 17780
rect 21196 17726 21310 17778
rect 21362 17726 21364 17778
rect 21196 17724 21364 17726
rect 21308 17714 21364 17724
rect 21308 17556 21364 17566
rect 21196 17332 21252 17342
rect 21196 16994 21252 17276
rect 21308 17106 21364 17500
rect 21308 17054 21310 17106
rect 21362 17054 21364 17106
rect 21308 17042 21364 17054
rect 21420 17108 21476 19068
rect 21532 19058 21588 19068
rect 21756 19124 21812 19134
rect 21756 19030 21812 19068
rect 21624 18844 21888 18854
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21624 18778 21888 18788
rect 21624 17276 21888 17286
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21624 17210 21888 17220
rect 21756 17108 21812 17118
rect 21980 17108 22036 22428
rect 22092 22484 22148 23660
rect 22204 23380 22260 24670
rect 22204 23314 22260 23324
rect 22316 23714 22372 23726
rect 22316 23662 22318 23714
rect 22370 23662 22372 23714
rect 22316 23604 22372 23662
rect 22316 23044 22372 23548
rect 22428 23548 22484 25004
rect 22540 24722 22596 26852
rect 22652 26852 22708 32172
rect 22988 32116 23044 32126
rect 22652 26786 22708 26796
rect 22876 32004 22932 32014
rect 22876 27858 22932 31948
rect 22988 31778 23044 32060
rect 23100 31890 23156 32396
rect 23100 31838 23102 31890
rect 23154 31838 23156 31890
rect 23100 31826 23156 31838
rect 22988 31726 22990 31778
rect 23042 31726 23044 31778
rect 22988 29876 23044 31726
rect 22988 28644 23044 29820
rect 23212 29652 23268 35308
rect 23548 35364 23604 35374
rect 23324 34692 23380 34702
rect 23324 34690 23492 34692
rect 23324 34638 23326 34690
rect 23378 34638 23492 34690
rect 23324 34636 23492 34638
rect 23324 34626 23380 34636
rect 23324 34468 23380 34478
rect 23324 34354 23380 34412
rect 23324 34302 23326 34354
rect 23378 34302 23380 34354
rect 23324 34290 23380 34302
rect 23436 34132 23492 34636
rect 23324 33684 23380 33694
rect 23436 33684 23492 34076
rect 23380 33628 23492 33684
rect 23324 33618 23380 33628
rect 23548 33572 23604 35308
rect 23660 34020 23716 35420
rect 23772 35140 23828 35644
rect 23772 35074 23828 35084
rect 23884 34916 23940 38668
rect 23996 38164 24052 38780
rect 23996 37378 24052 38108
rect 24108 38274 24164 38286
rect 24108 38222 24110 38274
rect 24162 38222 24164 38274
rect 24108 38162 24164 38222
rect 24108 38110 24110 38162
rect 24162 38110 24164 38162
rect 24108 38098 24164 38110
rect 24332 37604 24388 37614
rect 24332 37380 24388 37548
rect 23996 37326 23998 37378
rect 24050 37326 24052 37378
rect 23996 35252 24052 37326
rect 24220 37378 24388 37380
rect 24220 37326 24334 37378
rect 24386 37326 24388 37378
rect 24220 37324 24388 37326
rect 24108 37154 24164 37166
rect 24108 37102 24110 37154
rect 24162 37102 24164 37154
rect 24108 36594 24164 37102
rect 24108 36542 24110 36594
rect 24162 36542 24164 36594
rect 24108 36530 24164 36542
rect 24220 36484 24276 37324
rect 24332 37314 24388 37324
rect 24220 35812 24276 36428
rect 24108 35756 24276 35812
rect 24332 37156 24388 37166
rect 24108 35476 24164 35756
rect 24332 35700 24388 37100
rect 24108 35410 24164 35420
rect 24220 35644 24388 35700
rect 24220 35586 24276 35644
rect 24220 35534 24222 35586
rect 24274 35534 24276 35586
rect 24220 35364 24276 35534
rect 24220 35298 24276 35308
rect 24332 35476 24388 35486
rect 23996 35186 24052 35196
rect 23660 33926 23716 33964
rect 23772 34860 23940 34916
rect 23996 35028 24052 35038
rect 23436 33516 23604 33572
rect 23660 33684 23716 33694
rect 23324 33460 23380 33470
rect 23436 33460 23492 33516
rect 23380 33404 23492 33460
rect 23324 33394 23380 33404
rect 23660 33348 23716 33628
rect 23436 33292 23716 33348
rect 23436 33124 23492 33292
rect 23324 33122 23492 33124
rect 23324 33070 23438 33122
rect 23490 33070 23492 33122
rect 23324 33068 23492 33070
rect 23324 31892 23380 33068
rect 23436 33058 23492 33068
rect 23548 33122 23604 33134
rect 23548 33070 23550 33122
rect 23602 33070 23604 33122
rect 23324 31826 23380 31836
rect 23436 32900 23492 32910
rect 23324 31668 23380 31678
rect 23324 31574 23380 31612
rect 23436 31444 23492 32844
rect 23548 31778 23604 33070
rect 23660 33124 23716 33134
rect 23660 32452 23716 33068
rect 23660 32386 23716 32396
rect 23548 31726 23550 31778
rect 23602 31726 23604 31778
rect 23548 31714 23604 31726
rect 23212 29586 23268 29596
rect 23324 31388 23492 31444
rect 22988 28578 23044 28588
rect 22876 27806 22878 27858
rect 22930 27806 22932 27858
rect 22876 26516 22932 27806
rect 22988 28084 23044 28094
rect 22988 27746 23044 28028
rect 22988 27694 22990 27746
rect 23042 27694 23044 27746
rect 22988 27682 23044 27694
rect 23100 27858 23156 27870
rect 23100 27806 23102 27858
rect 23154 27806 23156 27858
rect 23100 27300 23156 27806
rect 23100 27234 23156 27244
rect 23324 27858 23380 31388
rect 23660 30212 23716 30222
rect 23660 29988 23716 30156
rect 23660 28642 23716 29932
rect 23660 28590 23662 28642
rect 23714 28590 23716 28642
rect 23548 28532 23604 28542
rect 23548 28084 23604 28476
rect 23324 27806 23326 27858
rect 23378 27806 23380 27858
rect 23212 27076 23268 27086
rect 22876 26450 22932 26460
rect 23100 26740 23156 26750
rect 22652 26292 22708 26302
rect 22652 26198 22708 26236
rect 22540 24670 22542 24722
rect 22594 24670 22596 24722
rect 22540 24612 22596 24670
rect 22764 26178 22820 26190
rect 22764 26126 22766 26178
rect 22818 26126 22820 26178
rect 22540 24556 22708 24612
rect 22428 23492 22596 23548
rect 22428 23380 22484 23390
rect 22428 23266 22484 23324
rect 22428 23214 22430 23266
rect 22482 23214 22484 23266
rect 22428 23202 22484 23214
rect 22316 22988 22484 23044
rect 22092 22418 22148 22428
rect 22204 22932 22260 22942
rect 22204 22260 22260 22876
rect 22316 22484 22372 22494
rect 22316 22390 22372 22428
rect 22204 22204 22372 22260
rect 22092 20578 22148 20590
rect 22092 20526 22094 20578
rect 22146 20526 22148 20578
rect 22092 20244 22148 20526
rect 22092 18228 22148 20188
rect 22204 20580 22260 20590
rect 22204 18338 22260 20524
rect 22316 20356 22372 22204
rect 22428 20580 22484 22988
rect 22428 20514 22484 20524
rect 22316 20300 22484 20356
rect 22316 20132 22372 20142
rect 22316 19234 22372 20076
rect 22316 19182 22318 19234
rect 22370 19182 22372 19234
rect 22316 19012 22372 19182
rect 22428 19236 22484 20300
rect 22540 19460 22596 23492
rect 22652 23492 22708 24556
rect 22764 24498 22820 26126
rect 22988 26068 23044 26078
rect 23100 26068 23156 26684
rect 23212 26180 23268 27020
rect 23324 26908 23380 27806
rect 23436 28028 23604 28084
rect 23436 27636 23492 28028
rect 23548 27860 23604 27870
rect 23548 27766 23604 27804
rect 23436 27580 23604 27636
rect 23324 26852 23492 26908
rect 23212 26114 23268 26124
rect 23436 26178 23492 26852
rect 23548 26292 23604 27580
rect 23660 27076 23716 28590
rect 23772 28196 23828 34860
rect 23884 34692 23940 34702
rect 23996 34692 24052 34972
rect 23884 34690 24052 34692
rect 23884 34638 23886 34690
rect 23938 34638 24052 34690
rect 23884 34636 24052 34638
rect 24108 34804 24164 34814
rect 23884 34626 23940 34636
rect 24108 34132 24164 34748
rect 24220 34690 24276 34702
rect 24220 34638 24222 34690
rect 24274 34638 24276 34690
rect 24220 34244 24276 34638
rect 24220 34178 24276 34188
rect 23884 34076 24164 34132
rect 23884 32676 23940 34076
rect 24220 34020 24276 34030
rect 24332 34020 24388 35420
rect 24220 34018 24388 34020
rect 24220 33966 24222 34018
rect 24274 33966 24388 34018
rect 24220 33964 24388 33966
rect 23884 32116 23940 32620
rect 23884 32050 23940 32060
rect 23996 33906 24052 33918
rect 23996 33854 23998 33906
rect 24050 33854 24052 33906
rect 23996 33346 24052 33854
rect 23996 33294 23998 33346
rect 24050 33294 24052 33346
rect 23996 30884 24052 33294
rect 24220 32564 24276 33964
rect 24444 33460 24500 39564
rect 24668 39172 24724 40350
rect 24668 38276 24724 39116
rect 24668 38210 24724 38220
rect 24780 38052 24836 49868
rect 24892 49140 24948 50542
rect 25452 50596 25508 50606
rect 25026 49420 25290 49430
rect 25082 49364 25130 49420
rect 25186 49364 25234 49420
rect 25026 49354 25290 49364
rect 25452 49364 25508 50540
rect 25564 49810 25620 50764
rect 25788 50596 25844 50606
rect 25676 50482 25732 50494
rect 25676 50430 25678 50482
rect 25730 50430 25732 50482
rect 25676 50034 25732 50430
rect 25676 49982 25678 50034
rect 25730 49982 25732 50034
rect 25676 49970 25732 49982
rect 25564 49758 25566 49810
rect 25618 49758 25620 49810
rect 25564 49700 25620 49758
rect 25564 49476 25620 49644
rect 25564 49410 25620 49420
rect 25228 49252 25284 49290
rect 25228 49186 25284 49196
rect 24892 49084 25060 49140
rect 24892 48916 24948 48926
rect 24892 48822 24948 48860
rect 24668 37996 24836 38052
rect 24892 48692 24948 48702
rect 24556 37268 24612 37278
rect 24556 37174 24612 37212
rect 24668 37044 24724 37996
rect 24780 37828 24836 37838
rect 24780 37734 24836 37772
rect 24444 33394 24500 33404
rect 24556 36988 24724 37044
rect 24780 37604 24836 37614
rect 24444 33124 24500 33134
rect 24444 33030 24500 33068
rect 24108 32508 24276 32564
rect 24108 31220 24164 32508
rect 24220 31892 24276 31902
rect 24220 31798 24276 31836
rect 24108 31126 24164 31164
rect 24332 31108 24388 31118
rect 24332 31014 24388 31052
rect 23996 30818 24052 30828
rect 24220 30882 24276 30894
rect 24220 30830 24222 30882
rect 24274 30830 24276 30882
rect 23996 30210 24052 30222
rect 23996 30158 23998 30210
rect 24050 30158 24052 30210
rect 23996 30100 24052 30158
rect 23884 29316 23940 29326
rect 23884 29222 23940 29260
rect 23772 28130 23828 28140
rect 23996 28082 24052 30044
rect 24220 28642 24276 30830
rect 24556 29540 24612 36988
rect 24668 35588 24724 35598
rect 24668 35494 24724 35532
rect 24668 35252 24724 35262
rect 24668 35026 24724 35196
rect 24780 35138 24836 37548
rect 24780 35086 24782 35138
rect 24834 35086 24836 35138
rect 24780 35074 24836 35086
rect 24668 34974 24670 35026
rect 24722 34974 24724 35026
rect 24668 34962 24724 34974
rect 24892 34916 24948 48636
rect 25004 48244 25060 49084
rect 25228 49028 25284 49038
rect 25228 48934 25284 48972
rect 25452 48916 25508 49308
rect 25564 48916 25620 48926
rect 25452 48914 25732 48916
rect 25452 48862 25566 48914
rect 25618 48862 25732 48914
rect 25452 48860 25732 48862
rect 25564 48850 25620 48860
rect 25340 48244 25396 48254
rect 25004 48242 25396 48244
rect 25004 48190 25342 48242
rect 25394 48190 25396 48242
rect 25004 48188 25396 48190
rect 25340 48020 25396 48188
rect 25340 47964 25620 48020
rect 25026 47852 25290 47862
rect 25082 47796 25130 47852
rect 25186 47796 25234 47852
rect 25026 47786 25290 47796
rect 25564 47460 25620 47964
rect 25452 47236 25508 47246
rect 25452 46898 25508 47180
rect 25452 46846 25454 46898
rect 25506 46846 25508 46898
rect 25452 46834 25508 46846
rect 25228 46674 25284 46686
rect 25228 46622 25230 46674
rect 25282 46622 25284 46674
rect 25228 46564 25284 46622
rect 25340 46676 25396 46686
rect 25340 46582 25396 46620
rect 25228 46498 25284 46508
rect 25026 46284 25290 46294
rect 25082 46228 25130 46284
rect 25186 46228 25234 46284
rect 25026 46218 25290 46228
rect 25116 46004 25172 46014
rect 25116 45910 25172 45948
rect 25564 45108 25620 47404
rect 25676 47124 25732 48860
rect 25676 47058 25732 47068
rect 25788 46900 25844 50540
rect 25900 49810 25956 55692
rect 26236 55636 26292 57372
rect 26124 55580 26292 55636
rect 26348 57092 26404 57102
rect 26012 55412 26068 55422
rect 26012 55076 26068 55356
rect 26012 54404 26068 55020
rect 26012 54338 26068 54348
rect 26124 54180 26180 55580
rect 26348 55298 26404 57036
rect 26460 56642 26516 57372
rect 26572 56756 26628 59164
rect 26684 58884 26740 60172
rect 26796 60116 26852 60734
rect 26796 60050 26852 60060
rect 26908 59444 26964 60956
rect 26908 59330 26964 59388
rect 26908 59278 26910 59330
rect 26962 59278 26964 59330
rect 26908 59266 26964 59278
rect 27244 61010 27636 61012
rect 27244 60958 27582 61010
rect 27634 60958 27636 61010
rect 27244 60956 27636 60958
rect 27244 60786 27300 60956
rect 27580 60946 27636 60956
rect 27244 60734 27246 60786
rect 27298 60734 27300 60786
rect 26684 56980 26740 58828
rect 27244 58324 27300 60734
rect 28028 60228 28084 62302
rect 28428 61180 28692 61190
rect 28484 61124 28532 61180
rect 28588 61124 28636 61180
rect 28428 61114 28692 61124
rect 28028 59444 28084 60172
rect 28140 60116 28196 60126
rect 28140 60022 28196 60060
rect 28428 59612 28692 59622
rect 28484 59556 28532 59612
rect 28588 59556 28636 59612
rect 28428 59546 28692 59556
rect 28140 59444 28196 59454
rect 28028 59442 28196 59444
rect 28028 59390 28142 59442
rect 28194 59390 28196 59442
rect 28028 59388 28196 59390
rect 28140 59378 28196 59388
rect 27356 59332 27412 59342
rect 27356 59238 27412 59276
rect 28140 58548 28196 58558
rect 27244 57876 27300 58268
rect 28028 58546 28196 58548
rect 28028 58494 28142 58546
rect 28194 58494 28196 58546
rect 28028 58492 28196 58494
rect 27804 57876 27860 57886
rect 27244 57874 27860 57876
rect 27244 57822 27246 57874
rect 27298 57822 27806 57874
rect 27858 57822 27860 57874
rect 27244 57820 27860 57822
rect 27244 57810 27300 57820
rect 26796 57650 26852 57662
rect 26796 57598 26798 57650
rect 26850 57598 26852 57650
rect 26796 57428 26852 57598
rect 26908 57652 26964 57662
rect 26908 57558 26964 57596
rect 27020 57650 27076 57662
rect 27020 57598 27022 57650
rect 27074 57598 27076 57650
rect 26796 57362 26852 57372
rect 26796 57092 26852 57102
rect 27020 57092 27076 57598
rect 26852 57036 27020 57092
rect 26796 57026 26852 57036
rect 27020 56998 27076 57036
rect 26684 56914 26740 56924
rect 27692 56980 27748 56990
rect 27692 56886 27748 56924
rect 26908 56756 26964 56766
rect 26572 56700 26740 56756
rect 26460 56590 26462 56642
rect 26514 56590 26516 56642
rect 26460 55412 26516 56590
rect 26460 55346 26516 55356
rect 26348 55246 26350 55298
rect 26402 55246 26404 55298
rect 26348 55234 26404 55246
rect 26236 55074 26292 55086
rect 26236 55022 26238 55074
rect 26290 55022 26292 55074
rect 26236 54628 26292 55022
rect 26460 55074 26516 55086
rect 26460 55022 26462 55074
rect 26514 55022 26516 55074
rect 26236 54562 26292 54572
rect 26348 54740 26404 54750
rect 26236 54404 26292 54414
rect 26348 54404 26404 54684
rect 26236 54402 26404 54404
rect 26236 54350 26238 54402
rect 26290 54350 26404 54402
rect 26236 54348 26404 54350
rect 26236 54338 26292 54348
rect 26124 54124 26292 54180
rect 26124 53620 26180 53630
rect 26124 53526 26180 53564
rect 26012 53506 26068 53518
rect 26012 53454 26014 53506
rect 26066 53454 26068 53506
rect 26012 53058 26068 53454
rect 26236 53508 26292 54124
rect 26460 53956 26516 55022
rect 26572 55076 26628 55086
rect 26572 54982 26628 55020
rect 26684 54852 26740 56700
rect 26964 56700 27076 56756
rect 26908 56662 26964 56700
rect 27020 55412 27076 56700
rect 27020 55346 27076 55356
rect 27468 56644 27524 56654
rect 26796 55300 26852 55310
rect 26796 55206 26852 55244
rect 27356 55300 27412 55310
rect 27356 55206 27412 55244
rect 27244 55188 27300 55198
rect 27244 55094 27300 55132
rect 27132 55076 27188 55086
rect 26460 53890 26516 53900
rect 26572 54796 26740 54852
rect 27020 55074 27188 55076
rect 27020 55022 27134 55074
rect 27186 55022 27188 55074
rect 27020 55020 27188 55022
rect 26348 53732 26404 53742
rect 26348 53638 26404 53676
rect 26572 53620 26628 54796
rect 26684 54402 26740 54414
rect 26684 54350 26686 54402
rect 26738 54350 26740 54402
rect 26684 54290 26740 54350
rect 26684 54238 26686 54290
rect 26738 54238 26740 54290
rect 26684 54226 26740 54238
rect 26796 53732 26852 53742
rect 26460 53564 26628 53620
rect 26684 53620 26740 53658
rect 26796 53638 26852 53676
rect 26236 53452 26404 53508
rect 26012 53006 26014 53058
rect 26066 53006 26068 53058
rect 26012 52994 26068 53006
rect 26236 52276 26292 52286
rect 26236 52182 26292 52220
rect 26348 52162 26404 53452
rect 26348 52110 26350 52162
rect 26402 52110 26404 52162
rect 26348 52098 26404 52110
rect 26236 52052 26292 52062
rect 26236 51958 26292 51996
rect 25900 49758 25902 49810
rect 25954 49758 25956 49810
rect 25900 49140 25956 49758
rect 26012 51940 26068 51950
rect 26012 49700 26068 51884
rect 26348 51940 26404 51950
rect 26460 51940 26516 53564
rect 26684 53554 26740 53564
rect 26908 53508 26964 53518
rect 26796 53506 26964 53508
rect 26796 53454 26910 53506
rect 26962 53454 26964 53506
rect 26796 53452 26964 53454
rect 26684 53396 26740 53406
rect 26572 53284 26628 53294
rect 26572 52052 26628 53228
rect 26572 51958 26628 51996
rect 26404 51884 26516 51940
rect 26348 51874 26404 51884
rect 26236 51492 26292 51502
rect 26236 51044 26292 51436
rect 26460 51380 26516 51390
rect 26460 51286 26516 51324
rect 26236 50978 26292 50988
rect 26348 51266 26404 51278
rect 26348 51214 26350 51266
rect 26402 51214 26404 51266
rect 26348 50428 26404 51214
rect 26124 50372 26404 50428
rect 26684 50428 26740 53340
rect 26796 52836 26852 53452
rect 26908 53442 26964 53452
rect 27020 53508 27076 55020
rect 27132 55010 27188 55020
rect 26796 52162 26852 52780
rect 26796 52110 26798 52162
rect 26850 52110 26852 52162
rect 26796 52098 26852 52110
rect 26908 51492 26964 51502
rect 27020 51492 27076 53452
rect 27132 54852 27188 54862
rect 27132 54402 27188 54796
rect 27132 54350 27134 54402
rect 27186 54350 27188 54402
rect 27132 53284 27188 54350
rect 27132 53218 27188 53228
rect 27244 53730 27300 53742
rect 27244 53678 27246 53730
rect 27298 53678 27300 53730
rect 27244 53620 27300 53678
rect 27132 52164 27188 52174
rect 27132 52070 27188 52108
rect 27244 51716 27300 53564
rect 27468 53284 27524 56588
rect 27804 55468 27860 57820
rect 27916 57092 27972 57102
rect 28028 57092 28084 58492
rect 28140 58482 28196 58492
rect 28428 58044 28692 58054
rect 28484 57988 28532 58044
rect 28588 57988 28636 58044
rect 28428 57978 28692 57988
rect 27972 57036 28084 57092
rect 27916 57026 27972 57036
rect 28140 56980 28196 56990
rect 28140 56886 28196 56924
rect 28428 56476 28692 56486
rect 28484 56420 28532 56476
rect 28588 56420 28636 56476
rect 28428 56410 28692 56420
rect 28140 55970 28196 55982
rect 28140 55918 28142 55970
rect 28194 55918 28196 55970
rect 27804 55412 27972 55468
rect 27692 55298 27748 55310
rect 27692 55246 27694 55298
rect 27746 55246 27748 55298
rect 27692 54516 27748 55246
rect 27580 54402 27636 54414
rect 27580 54350 27582 54402
rect 27634 54350 27636 54402
rect 27580 53508 27636 54350
rect 27692 53620 27748 54460
rect 27692 53526 27748 53564
rect 27580 53442 27636 53452
rect 27468 53228 27748 53284
rect 27468 52724 27524 52734
rect 27468 52274 27524 52668
rect 27468 52222 27470 52274
rect 27522 52222 27524 52274
rect 27468 52210 27524 52222
rect 27580 52052 27636 52062
rect 26964 51436 27076 51492
rect 27132 51660 27300 51716
rect 27356 51938 27412 51950
rect 27356 51886 27358 51938
rect 27410 51886 27412 51938
rect 26908 51426 26964 51436
rect 26796 51378 26852 51390
rect 26796 51326 26798 51378
rect 26850 51326 26852 51378
rect 26796 51268 26852 51326
rect 27132 51268 27188 51660
rect 26796 51212 27188 51268
rect 27244 51266 27300 51278
rect 27244 51214 27246 51266
rect 27298 51214 27300 51266
rect 26684 50372 26852 50428
rect 26124 49922 26180 50372
rect 26124 49870 26126 49922
rect 26178 49870 26180 49922
rect 26124 49858 26180 49870
rect 26012 49644 26180 49700
rect 25900 49074 25956 49084
rect 26012 49476 26068 49486
rect 26012 49026 26068 49420
rect 26012 48974 26014 49026
rect 26066 48974 26068 49026
rect 26012 48962 26068 48974
rect 26124 48692 26180 49644
rect 26572 49698 26628 49710
rect 26572 49646 26574 49698
rect 26626 49646 26628 49698
rect 26572 49364 26628 49646
rect 26572 49298 26628 49308
rect 26348 49028 26404 49038
rect 26348 48934 26404 48972
rect 26572 49028 26628 49038
rect 25564 45042 25620 45052
rect 25676 46844 25844 46900
rect 25900 48636 26180 48692
rect 26236 48802 26292 48814
rect 26236 48750 26238 48802
rect 26290 48750 26292 48802
rect 25228 44994 25284 45006
rect 25228 44942 25230 44994
rect 25282 44942 25284 44994
rect 25228 44884 25284 44942
rect 25228 44818 25284 44828
rect 25026 44716 25290 44726
rect 25082 44660 25130 44716
rect 25186 44660 25234 44716
rect 25026 44650 25290 44660
rect 25676 44548 25732 46844
rect 25788 46676 25844 46686
rect 25788 46582 25844 46620
rect 25452 44492 25732 44548
rect 25788 45444 25844 45454
rect 25026 43148 25290 43158
rect 25082 43092 25130 43148
rect 25186 43092 25234 43148
rect 25026 43082 25290 43092
rect 25228 41860 25284 41870
rect 25228 41766 25284 41804
rect 25026 41580 25290 41590
rect 25082 41524 25130 41580
rect 25186 41524 25234 41580
rect 25026 41514 25290 41524
rect 25116 41300 25172 41310
rect 25116 41206 25172 41244
rect 25340 40852 25396 40862
rect 25340 40626 25396 40796
rect 25340 40574 25342 40626
rect 25394 40574 25396 40626
rect 25340 40562 25396 40574
rect 25026 40012 25290 40022
rect 25082 39956 25130 40012
rect 25186 39956 25234 40012
rect 25026 39946 25290 39956
rect 25116 39508 25172 39518
rect 25116 39414 25172 39452
rect 25228 38948 25284 38958
rect 25228 38722 25284 38892
rect 25228 38670 25230 38722
rect 25282 38670 25284 38722
rect 25228 38658 25284 38670
rect 25026 38444 25290 38454
rect 25082 38388 25130 38444
rect 25186 38388 25234 38444
rect 25026 38378 25290 38388
rect 25228 38276 25284 38286
rect 25228 38164 25284 38220
rect 25116 38162 25284 38164
rect 25116 38110 25230 38162
rect 25282 38110 25284 38162
rect 25116 38108 25284 38110
rect 25116 37604 25172 38108
rect 25228 38098 25284 38108
rect 25116 37538 25172 37548
rect 25228 37492 25284 37502
rect 25452 37492 25508 44492
rect 25788 44436 25844 45388
rect 25676 44380 25844 44436
rect 25564 43876 25620 43886
rect 25564 43652 25620 43820
rect 25564 43586 25620 43596
rect 25564 43314 25620 43326
rect 25564 43262 25566 43314
rect 25618 43262 25620 43314
rect 25564 42756 25620 43262
rect 25564 42690 25620 42700
rect 25564 41972 25620 41982
rect 25564 41636 25620 41916
rect 25564 41570 25620 41580
rect 25676 40404 25732 44380
rect 25788 43764 25844 43774
rect 25788 43670 25844 43708
rect 25900 43540 25956 48636
rect 26012 48356 26068 48366
rect 26236 48356 26292 48750
rect 26572 48692 26628 48972
rect 26684 48916 26740 48926
rect 26684 48822 26740 48860
rect 26012 48354 26292 48356
rect 26012 48302 26014 48354
rect 26066 48302 26292 48354
rect 26012 48300 26292 48302
rect 26460 48636 26628 48692
rect 26012 48290 26068 48300
rect 26124 48132 26180 48142
rect 26012 47124 26068 47134
rect 26012 43764 26068 47068
rect 26012 43698 26068 43708
rect 25788 43484 25956 43540
rect 25788 41188 25844 43484
rect 25900 43316 25956 43326
rect 25900 43222 25956 43260
rect 26124 42084 26180 48076
rect 26348 47570 26404 47582
rect 26348 47518 26350 47570
rect 26402 47518 26404 47570
rect 26348 47236 26404 47518
rect 26348 47170 26404 47180
rect 26236 46562 26292 46574
rect 26236 46510 26238 46562
rect 26290 46510 26292 46562
rect 26236 45892 26292 46510
rect 26236 45444 26292 45836
rect 26236 45378 26292 45388
rect 26460 45220 26516 48636
rect 26796 47796 26852 50372
rect 26908 49586 26964 51212
rect 26908 49534 26910 49586
rect 26962 49534 26964 49586
rect 26908 49522 26964 49534
rect 27020 51044 27076 51054
rect 27020 49698 27076 50988
rect 27244 50708 27300 51214
rect 27356 51154 27412 51886
rect 27356 51102 27358 51154
rect 27410 51102 27412 51154
rect 27356 51090 27412 51102
rect 27244 50642 27300 50652
rect 27020 49646 27022 49698
rect 27074 49646 27076 49698
rect 26684 47740 26852 47796
rect 26908 48916 26964 48926
rect 26684 47460 26740 47740
rect 26796 47572 26852 47582
rect 26908 47572 26964 48860
rect 27020 48020 27076 49646
rect 27468 49700 27524 49710
rect 27132 49588 27188 49598
rect 27132 49138 27188 49532
rect 27132 49086 27134 49138
rect 27186 49086 27188 49138
rect 27132 49074 27188 49086
rect 27020 47964 27412 48020
rect 27244 47572 27300 47582
rect 26796 47570 26964 47572
rect 26796 47518 26798 47570
rect 26850 47518 26964 47570
rect 26796 47516 26964 47518
rect 27020 47570 27300 47572
rect 27020 47518 27246 47570
rect 27298 47518 27300 47570
rect 27020 47516 27300 47518
rect 26796 47506 26852 47516
rect 26572 47458 26740 47460
rect 26572 47406 26686 47458
rect 26738 47406 26740 47458
rect 26572 47404 26740 47406
rect 26572 46452 26628 47404
rect 26684 47394 26740 47404
rect 26908 47348 26964 47358
rect 27020 47348 27076 47516
rect 27244 47506 27300 47516
rect 26908 47346 27076 47348
rect 26908 47294 26910 47346
rect 26962 47294 27076 47346
rect 26908 47292 27076 47294
rect 26908 47282 26964 47292
rect 27132 47236 27188 47246
rect 27132 47234 27300 47236
rect 27132 47182 27134 47234
rect 27186 47182 27300 47234
rect 27132 47180 27300 47182
rect 27132 47170 27188 47180
rect 26684 47012 26740 47022
rect 26684 46898 26740 46956
rect 27244 47012 27300 47180
rect 26684 46846 26686 46898
rect 26738 46846 26740 46898
rect 26684 46834 26740 46846
rect 27132 46900 27188 46910
rect 27132 46806 27188 46844
rect 26572 46004 26628 46396
rect 27244 46004 27300 46956
rect 26572 46002 26740 46004
rect 26572 45950 26574 46002
rect 26626 45950 26740 46002
rect 26572 45948 26740 45950
rect 26572 45938 26628 45948
rect 26460 45164 26628 45220
rect 26460 44996 26516 45006
rect 26460 43762 26516 44940
rect 26460 43710 26462 43762
rect 26514 43710 26516 43762
rect 26460 43698 26516 43710
rect 26572 43708 26628 45164
rect 26684 43876 26740 45948
rect 27244 45332 27300 45948
rect 27356 45892 27412 47964
rect 27468 46228 27524 49644
rect 27580 49140 27636 51996
rect 27692 51602 27748 53228
rect 27692 51550 27694 51602
rect 27746 51550 27748 51602
rect 27692 51538 27748 51550
rect 27804 52050 27860 52062
rect 27804 51998 27806 52050
rect 27858 51998 27860 52050
rect 27804 51380 27860 51998
rect 27804 50706 27860 51324
rect 27804 50654 27806 50706
rect 27858 50654 27860 50706
rect 27804 50642 27860 50654
rect 27916 50428 27972 55412
rect 28028 55412 28084 55422
rect 28028 55076 28084 55356
rect 28140 55300 28196 55918
rect 28140 55234 28196 55244
rect 28140 55076 28196 55086
rect 28028 55074 28196 55076
rect 28028 55022 28142 55074
rect 28194 55022 28196 55074
rect 28028 55020 28196 55022
rect 28028 54402 28084 54414
rect 28028 54350 28030 54402
rect 28082 54350 28084 54402
rect 28028 53844 28084 54350
rect 28140 54290 28196 55020
rect 28428 54908 28692 54918
rect 28484 54852 28532 54908
rect 28588 54852 28636 54908
rect 28428 54842 28692 54852
rect 28140 54238 28142 54290
rect 28194 54238 28196 54290
rect 28140 54226 28196 54238
rect 28028 53778 28084 53788
rect 28140 53508 28196 53518
rect 28140 53414 28196 53452
rect 28428 53340 28692 53350
rect 28484 53284 28532 53340
rect 28588 53284 28636 53340
rect 28428 53274 28692 53284
rect 28140 52836 28196 52846
rect 28140 52742 28196 52780
rect 28428 51772 28692 51782
rect 28484 51716 28532 51772
rect 28588 51716 28636 51772
rect 28428 51706 28692 51716
rect 28140 51268 28196 51278
rect 28140 51266 28308 51268
rect 28140 51214 28142 51266
rect 28194 51214 28308 51266
rect 28140 51212 28308 51214
rect 28140 51202 28196 51212
rect 27804 50372 27972 50428
rect 28028 51154 28084 51166
rect 28028 51102 28030 51154
rect 28082 51102 28084 51154
rect 28028 50428 28084 51102
rect 28028 50372 28196 50428
rect 27580 49138 27748 49140
rect 27580 49086 27582 49138
rect 27634 49086 27748 49138
rect 27580 49084 27748 49086
rect 27580 49074 27636 49084
rect 27692 47570 27748 49084
rect 27692 47518 27694 47570
rect 27746 47518 27748 47570
rect 27692 47506 27748 47518
rect 27804 47012 27860 50372
rect 27804 46946 27860 46956
rect 27916 49698 27972 49710
rect 27916 49646 27918 49698
rect 27970 49646 27972 49698
rect 27916 49586 27972 49646
rect 27916 49534 27918 49586
rect 27970 49534 27972 49586
rect 27916 48804 27972 49534
rect 28028 48804 28084 48814
rect 27916 48802 28084 48804
rect 27916 48750 28030 48802
rect 28082 48750 28084 48802
rect 27916 48748 28084 48750
rect 27580 46562 27636 46574
rect 27580 46510 27582 46562
rect 27634 46510 27636 46562
rect 27580 46340 27636 46510
rect 27916 46340 27972 48748
rect 28028 48738 28084 48748
rect 28140 48132 28196 50372
rect 28028 48130 28196 48132
rect 28028 48078 28142 48130
rect 28194 48078 28196 48130
rect 28028 48076 28196 48078
rect 28028 47682 28084 48076
rect 28140 48066 28196 48076
rect 28028 47630 28030 47682
rect 28082 47630 28084 47682
rect 28028 47618 28084 47630
rect 28140 47572 28196 47582
rect 28252 47572 28308 51212
rect 28428 50204 28692 50214
rect 28484 50148 28532 50204
rect 28588 50148 28636 50204
rect 28428 50138 28692 50148
rect 28428 48636 28692 48646
rect 28484 48580 28532 48636
rect 28588 48580 28636 48636
rect 28428 48570 28692 48580
rect 28140 47570 28308 47572
rect 28140 47518 28142 47570
rect 28194 47518 28308 47570
rect 28140 47516 28308 47518
rect 28140 46898 28196 47516
rect 28428 47068 28692 47078
rect 28484 47012 28532 47068
rect 28588 47012 28636 47068
rect 28428 47002 28692 47012
rect 28140 46846 28142 46898
rect 28194 46846 28196 46898
rect 27580 46284 28084 46340
rect 27468 46172 27636 46228
rect 27580 46004 27636 46172
rect 27580 45948 27748 46004
rect 27356 45826 27412 45836
rect 27244 45276 27636 45332
rect 26796 45108 26852 45118
rect 26796 44434 26852 45052
rect 27468 45108 27524 45118
rect 27356 44996 27412 45006
rect 27356 44902 27412 44940
rect 27132 44884 27188 44894
rect 27188 44828 27300 44884
rect 27132 44818 27188 44828
rect 26796 44382 26798 44434
rect 26850 44382 26852 44434
rect 26796 44370 26852 44382
rect 26740 43820 26852 43876
rect 26684 43810 26740 43820
rect 26796 43708 26852 43820
rect 27244 43708 27300 44828
rect 26572 43652 26740 43708
rect 26796 43652 27076 43708
rect 27244 43652 27412 43708
rect 26236 43538 26292 43550
rect 26236 43486 26238 43538
rect 26290 43486 26292 43538
rect 26236 43428 26292 43486
rect 26236 43362 26292 43372
rect 26460 43540 26516 43550
rect 26124 42018 26180 42028
rect 26348 43316 26404 43326
rect 26012 41636 26068 41646
rect 25788 41132 25956 41188
rect 25788 40964 25844 40974
rect 25788 40870 25844 40908
rect 25788 40404 25844 40414
rect 25676 40402 25844 40404
rect 25676 40350 25790 40402
rect 25842 40350 25844 40402
rect 25676 40348 25844 40350
rect 25676 38612 25732 38622
rect 25676 38162 25732 38556
rect 25676 38110 25678 38162
rect 25730 38110 25732 38162
rect 25676 37828 25732 38110
rect 25676 37762 25732 37772
rect 25676 37604 25732 37614
rect 25452 37436 25620 37492
rect 25228 37398 25284 37436
rect 25340 37268 25396 37278
rect 25340 37174 25396 37212
rect 25452 37266 25508 37278
rect 25452 37214 25454 37266
rect 25506 37214 25508 37266
rect 25026 36876 25290 36886
rect 25082 36820 25130 36876
rect 25186 36820 25234 36876
rect 25026 36810 25290 36820
rect 25452 36708 25508 37214
rect 25452 36642 25508 36652
rect 25228 36596 25284 36606
rect 25228 35586 25284 36540
rect 25228 35534 25230 35586
rect 25282 35534 25284 35586
rect 25228 35522 25284 35534
rect 25026 35308 25290 35318
rect 25082 35252 25130 35308
rect 25186 35252 25234 35308
rect 25026 35242 25290 35252
rect 24780 34860 24948 34916
rect 25004 35140 25060 35150
rect 24668 34692 24724 34702
rect 24668 34018 24724 34636
rect 24668 33966 24670 34018
rect 24722 33966 24724 34018
rect 24668 33906 24724 33966
rect 24668 33854 24670 33906
rect 24722 33854 24724 33906
rect 24668 33842 24724 33854
rect 24668 32452 24724 32462
rect 24668 32358 24724 32396
rect 24668 31668 24724 31706
rect 24668 31602 24724 31612
rect 24668 30994 24724 31006
rect 24668 30942 24670 30994
rect 24722 30942 24724 30994
rect 24668 30884 24724 30942
rect 24668 30818 24724 30828
rect 24220 28590 24222 28642
rect 24274 28590 24276 28642
rect 24220 28578 24276 28590
rect 24332 29484 24612 29540
rect 24668 30100 24724 30110
rect 23996 28030 23998 28082
rect 24050 28030 24052 28082
rect 23996 28018 24052 28030
rect 24332 27748 24388 29484
rect 24668 29426 24724 30044
rect 24780 29876 24836 34860
rect 25004 34804 25060 35084
rect 24892 34748 25060 34804
rect 25116 35138 25172 35150
rect 25116 35086 25118 35138
rect 25170 35086 25172 35138
rect 24892 33458 24948 34748
rect 25116 34692 25172 35086
rect 25116 34598 25172 34636
rect 25340 34804 25396 34814
rect 25340 34354 25396 34748
rect 25340 34302 25342 34354
rect 25394 34302 25396 34354
rect 25340 34290 25396 34302
rect 25026 33740 25290 33750
rect 25082 33684 25130 33740
rect 25186 33684 25234 33740
rect 25026 33674 25290 33684
rect 25340 33572 25396 33582
rect 25396 33516 25508 33572
rect 25340 33506 25396 33516
rect 24892 33406 24894 33458
rect 24946 33406 24948 33458
rect 24892 33394 24948 33406
rect 25228 33458 25284 33470
rect 25228 33406 25230 33458
rect 25282 33406 25284 33458
rect 25228 33348 25284 33406
rect 25228 33282 25284 33292
rect 25452 32788 25508 33516
rect 25026 32172 25290 32182
rect 25082 32116 25130 32172
rect 25186 32116 25234 32172
rect 25026 32106 25290 32116
rect 25452 32004 25508 32732
rect 25564 32676 25620 37436
rect 25676 37490 25732 37548
rect 25676 37438 25678 37490
rect 25730 37438 25732 37490
rect 25676 37426 25732 37438
rect 25788 37492 25844 40348
rect 25900 40292 25956 41132
rect 25900 40226 25956 40236
rect 25788 37426 25844 37436
rect 25900 39618 25956 39630
rect 25900 39566 25902 39618
rect 25954 39566 25956 39618
rect 25676 35588 25732 35598
rect 25676 34690 25732 35532
rect 25900 35140 25956 39566
rect 25900 35046 25956 35084
rect 25676 34638 25678 34690
rect 25730 34638 25732 34690
rect 25676 34356 25732 34638
rect 25676 34290 25732 34300
rect 25900 34692 25956 34702
rect 25900 34132 25956 34636
rect 26012 34132 26068 41580
rect 26348 41410 26404 43260
rect 26348 41358 26350 41410
rect 26402 41358 26404 41410
rect 26348 41346 26404 41358
rect 26236 41188 26292 41198
rect 26124 41132 26236 41188
rect 26124 37826 26180 41132
rect 26236 41122 26292 41132
rect 26348 41186 26404 41198
rect 26348 41134 26350 41186
rect 26402 41134 26404 41186
rect 26348 40740 26404 41134
rect 26460 40964 26516 43484
rect 26572 43538 26628 43550
rect 26572 43486 26574 43538
rect 26626 43486 26628 43538
rect 26572 43316 26628 43486
rect 26572 41188 26628 43260
rect 26684 42868 26740 43652
rect 26796 43540 26852 43550
rect 27020 43540 27076 43652
rect 27356 43650 27412 43652
rect 27356 43598 27358 43650
rect 27410 43598 27412 43650
rect 27356 43586 27412 43598
rect 27132 43540 27188 43550
rect 27020 43538 27188 43540
rect 27020 43486 27134 43538
rect 27186 43486 27188 43538
rect 27020 43484 27188 43486
rect 26796 43446 26852 43484
rect 26684 42812 26852 42868
rect 26684 42644 26740 42654
rect 26684 42550 26740 42588
rect 26572 41122 26628 41132
rect 26684 41188 26740 41198
rect 26796 41188 26852 42812
rect 26684 41186 26796 41188
rect 26684 41134 26686 41186
rect 26738 41134 26796 41186
rect 26684 41132 26796 41134
rect 26684 41122 26740 41132
rect 26796 41122 26852 41132
rect 27020 41860 27076 41870
rect 26908 41074 26964 41086
rect 26908 41022 26910 41074
rect 26962 41022 26964 41074
rect 26796 40964 26852 40974
rect 26460 40908 26740 40964
rect 26348 40684 26628 40740
rect 26236 40628 26292 40638
rect 26236 39620 26292 40572
rect 26348 40516 26404 40526
rect 26348 40422 26404 40460
rect 26460 40292 26516 40302
rect 26460 39620 26516 40236
rect 26572 40180 26628 40684
rect 26572 40114 26628 40124
rect 26236 39618 26404 39620
rect 26236 39566 26238 39618
rect 26290 39566 26404 39618
rect 26236 39564 26404 39566
rect 26236 39554 26292 39564
rect 26124 37774 26126 37826
rect 26178 37774 26180 37826
rect 26124 34468 26180 37774
rect 26236 38724 26292 38734
rect 26236 37154 26292 38668
rect 26348 38388 26404 39564
rect 26460 39618 26628 39620
rect 26460 39566 26462 39618
rect 26514 39566 26628 39618
rect 26460 39564 26628 39566
rect 26460 39554 26516 39564
rect 26572 39060 26628 39564
rect 26348 38332 26516 38388
rect 26460 38274 26516 38332
rect 26460 38222 26462 38274
rect 26514 38222 26516 38274
rect 26348 38164 26404 38174
rect 26348 37828 26404 38108
rect 26460 38052 26516 38222
rect 26572 38052 26628 39004
rect 26684 38668 26740 40908
rect 26796 40870 26852 40908
rect 26908 40628 26964 41022
rect 27020 40964 27076 41804
rect 27020 40898 27076 40908
rect 26908 40562 26964 40572
rect 27132 40516 27188 43484
rect 27244 43540 27300 43550
rect 27244 43446 27300 43484
rect 27356 43428 27412 43438
rect 27356 42084 27412 43372
rect 26796 40404 26852 40414
rect 26796 40310 26852 40348
rect 26908 40180 26964 40190
rect 26796 39844 26852 39854
rect 26796 39750 26852 39788
rect 26908 39618 26964 40124
rect 26908 39566 26910 39618
rect 26962 39566 26964 39618
rect 26908 38836 26964 39566
rect 27020 39396 27076 39406
rect 27020 39302 27076 39340
rect 26908 38770 26964 38780
rect 27132 38668 27188 40460
rect 26684 38612 26852 38668
rect 26572 37996 26740 38052
rect 26460 37986 26516 37996
rect 26572 37828 26628 37838
rect 26348 37826 26628 37828
rect 26348 37774 26574 37826
rect 26626 37774 26628 37826
rect 26348 37772 26628 37774
rect 26572 37762 26628 37772
rect 26236 37102 26238 37154
rect 26290 37102 26292 37154
rect 26236 36932 26292 37102
rect 26236 36866 26292 36876
rect 26348 37492 26404 37502
rect 26236 36708 26292 36718
rect 26236 36594 26292 36652
rect 26236 36542 26238 36594
rect 26290 36542 26292 36594
rect 26236 36530 26292 36542
rect 26236 35028 26292 35038
rect 26236 34934 26292 34972
rect 26348 34580 26404 37436
rect 26572 37044 26628 37054
rect 26460 37042 26628 37044
rect 26460 36990 26574 37042
rect 26626 36990 26628 37042
rect 26460 36988 26628 36990
rect 26460 34916 26516 36988
rect 26572 36978 26628 36988
rect 26572 36820 26628 36830
rect 26572 36482 26628 36764
rect 26572 36430 26574 36482
rect 26626 36430 26628 36482
rect 26572 35588 26628 36430
rect 26572 35522 26628 35532
rect 26460 34850 26516 34860
rect 26572 35138 26628 35150
rect 26572 35086 26574 35138
rect 26626 35086 26628 35138
rect 26572 35026 26628 35086
rect 26572 34974 26574 35026
rect 26626 34974 26628 35026
rect 26572 34804 26628 34974
rect 26684 35028 26740 37996
rect 26796 37380 26852 38612
rect 26908 38612 27188 38668
rect 27244 42028 27412 42084
rect 27468 42754 27524 45052
rect 27468 42702 27470 42754
rect 27522 42702 27524 42754
rect 27244 41300 27300 42028
rect 27468 41972 27524 42702
rect 27468 41906 27524 41916
rect 27356 41860 27412 41870
rect 27356 41766 27412 41804
rect 27356 41300 27412 41310
rect 27580 41300 27636 45276
rect 27692 43708 27748 45948
rect 27804 45892 27860 45902
rect 27804 45798 27860 45836
rect 27692 43652 27972 43708
rect 27692 43428 27748 43652
rect 27692 43362 27748 43372
rect 27804 43538 27860 43550
rect 27804 43486 27806 43538
rect 27858 43486 27860 43538
rect 27244 41298 27412 41300
rect 27244 41246 27358 41298
rect 27410 41246 27412 41298
rect 27244 41244 27412 41246
rect 27244 38668 27300 41244
rect 27356 41234 27412 41244
rect 27468 41244 27580 41300
rect 27468 40626 27524 41244
rect 27580 41234 27636 41244
rect 27692 42756 27748 42766
rect 27468 40574 27470 40626
rect 27522 40574 27524 40626
rect 27468 40562 27524 40574
rect 27580 41076 27636 41086
rect 27356 39844 27412 39854
rect 27356 39750 27412 39788
rect 27356 39396 27412 39406
rect 27356 38946 27412 39340
rect 27356 38894 27358 38946
rect 27410 38894 27412 38946
rect 27356 38882 27412 38894
rect 27468 39394 27524 39406
rect 27468 39342 27470 39394
rect 27522 39342 27524 39394
rect 27468 38948 27524 39342
rect 27468 38882 27524 38892
rect 27244 38612 27524 38668
rect 26908 38164 26964 38612
rect 27244 38274 27300 38286
rect 27244 38222 27246 38274
rect 27298 38222 27300 38274
rect 27020 38164 27076 38174
rect 26908 38162 27076 38164
rect 26908 38110 27022 38162
rect 27074 38110 27076 38162
rect 26908 38108 27076 38110
rect 27020 38098 27076 38108
rect 26796 37314 26852 37324
rect 26908 37266 26964 37278
rect 26908 37214 26910 37266
rect 26962 37214 26964 37266
rect 26796 37154 26852 37166
rect 26796 37102 26798 37154
rect 26850 37102 26852 37154
rect 26796 36706 26852 37102
rect 26796 36654 26798 36706
rect 26850 36654 26852 36706
rect 26796 36642 26852 36654
rect 26908 36596 26964 37214
rect 26908 36530 26964 36540
rect 27020 36484 27076 36494
rect 27244 36484 27300 38222
rect 27468 38162 27524 38612
rect 27468 38110 27470 38162
rect 27522 38110 27524 38162
rect 27468 38098 27524 38110
rect 27356 37940 27412 37950
rect 27356 37490 27412 37884
rect 27580 37716 27636 41020
rect 27692 39844 27748 42700
rect 27804 42644 27860 43486
rect 27916 42866 27972 43652
rect 27916 42814 27918 42866
rect 27970 42814 27972 42866
rect 27916 42802 27972 42814
rect 28028 42644 28084 46284
rect 28140 45108 28196 46846
rect 28428 45500 28692 45510
rect 28484 45444 28532 45500
rect 28588 45444 28636 45500
rect 28428 45434 28692 45444
rect 28140 45014 28196 45052
rect 28428 43932 28692 43942
rect 28484 43876 28532 43932
rect 28588 43876 28636 43932
rect 28428 43866 28692 43876
rect 28140 43652 28196 43662
rect 28140 43558 28196 43596
rect 27804 42588 28084 42644
rect 27692 39750 27748 39788
rect 27692 37716 27748 37726
rect 27580 37660 27692 37716
rect 27356 37438 27358 37490
rect 27410 37438 27412 37490
rect 27356 37426 27412 37438
rect 27692 36596 27748 37660
rect 27916 37154 27972 42588
rect 28428 42364 28692 42374
rect 28484 42308 28532 42364
rect 28588 42308 28636 42364
rect 28428 42298 28692 42308
rect 28028 41972 28084 41982
rect 28028 41300 28084 41916
rect 28028 41298 28196 41300
rect 28028 41246 28030 41298
rect 28082 41246 28196 41298
rect 28028 41244 28196 41246
rect 28028 41234 28084 41244
rect 28140 40628 28196 41244
rect 28428 40796 28692 40806
rect 28484 40740 28532 40796
rect 28588 40740 28636 40796
rect 28428 40730 28692 40740
rect 28028 40572 28140 40628
rect 28028 38834 28084 40572
rect 28140 40534 28196 40572
rect 28140 39844 28196 39854
rect 28140 39730 28196 39788
rect 28140 39678 28142 39730
rect 28194 39678 28196 39730
rect 28140 39666 28196 39678
rect 28428 39228 28692 39238
rect 28484 39172 28532 39228
rect 28588 39172 28636 39228
rect 28428 39162 28692 39172
rect 28028 38782 28030 38834
rect 28082 38782 28084 38834
rect 28028 38668 28084 38782
rect 28028 38612 28196 38668
rect 27916 37102 27918 37154
rect 27970 37102 27972 37154
rect 27804 36596 27860 36606
rect 27692 36594 27860 36596
rect 27692 36542 27806 36594
rect 27858 36542 27860 36594
rect 27692 36540 27860 36542
rect 27804 36530 27860 36540
rect 27356 36484 27412 36494
rect 27020 36390 27076 36428
rect 27132 36482 27412 36484
rect 27132 36430 27358 36482
rect 27410 36430 27412 36482
rect 27132 36428 27412 36430
rect 26684 34962 26740 34972
rect 26796 36372 26852 36382
rect 26572 34738 26628 34748
rect 26348 34524 26628 34580
rect 26124 34402 26180 34412
rect 26348 34356 26404 34366
rect 26124 34132 26180 34142
rect 26012 34130 26180 34132
rect 26012 34078 26126 34130
rect 26178 34078 26180 34130
rect 26012 34076 26180 34078
rect 25900 34038 25956 34076
rect 25676 34020 25732 34030
rect 25676 32786 25732 33964
rect 26124 32788 26180 34076
rect 26348 34132 26404 34300
rect 26460 34132 26516 34142
rect 26348 34130 26516 34132
rect 26348 34078 26462 34130
rect 26514 34078 26516 34130
rect 26348 34076 26516 34078
rect 26348 33684 26404 34076
rect 26460 34066 26516 34076
rect 26460 33908 26516 33918
rect 26460 33814 26516 33852
rect 26348 33628 26516 33684
rect 25676 32734 25678 32786
rect 25730 32734 25732 32786
rect 25676 32722 25732 32734
rect 25900 32732 26180 32788
rect 26348 32788 26404 32798
rect 25564 32610 25620 32620
rect 25900 32228 25956 32732
rect 26012 32562 26068 32574
rect 26012 32510 26014 32562
rect 26066 32510 26068 32562
rect 26012 32452 26068 32510
rect 26348 32562 26404 32732
rect 26348 32510 26350 32562
rect 26402 32510 26404 32562
rect 26348 32498 26404 32510
rect 26124 32452 26180 32462
rect 26012 32396 26124 32452
rect 26124 32386 26180 32396
rect 26460 32452 26516 33628
rect 25228 31948 25508 32004
rect 25564 32172 25956 32228
rect 26348 32338 26404 32350
rect 26348 32286 26350 32338
rect 26402 32286 26404 32338
rect 25228 31890 25284 31948
rect 25228 31838 25230 31890
rect 25282 31838 25284 31890
rect 25228 31826 25284 31838
rect 24780 29810 24836 29820
rect 24892 31220 24948 31230
rect 24668 29374 24670 29426
rect 24722 29374 24724 29426
rect 24668 29362 24724 29374
rect 24556 29316 24612 29326
rect 24108 27692 24388 27748
rect 24444 28868 24500 28878
rect 24444 28642 24500 28812
rect 24556 28756 24612 29260
rect 24668 28756 24724 28766
rect 24556 28754 24724 28756
rect 24556 28702 24670 28754
rect 24722 28702 24724 28754
rect 24556 28700 24724 28702
rect 24668 28690 24724 28700
rect 24444 28590 24446 28642
rect 24498 28590 24500 28642
rect 23660 26982 23716 27020
rect 23996 27186 24052 27198
rect 23996 27134 23998 27186
rect 24050 27134 24052 27186
rect 23548 26226 23604 26236
rect 23660 26516 23716 26526
rect 23436 26126 23438 26178
rect 23490 26126 23492 26178
rect 22988 26066 23156 26068
rect 22988 26014 22990 26066
rect 23042 26014 23156 26066
rect 22988 26012 23156 26014
rect 22988 26002 23044 26012
rect 23100 25508 23156 26012
rect 22988 25396 23044 25406
rect 22988 24946 23044 25340
rect 22988 24894 22990 24946
rect 23042 24894 23044 24946
rect 22988 24882 23044 24894
rect 22764 24446 22766 24498
rect 22818 24446 22820 24498
rect 22764 24434 22820 24446
rect 22876 24722 22932 24734
rect 22876 24670 22878 24722
rect 22930 24670 22932 24722
rect 22876 24164 22932 24670
rect 23100 24498 23156 25452
rect 23436 24836 23492 26126
rect 23100 24446 23102 24498
rect 23154 24446 23156 24498
rect 23100 24434 23156 24446
rect 23212 24780 23492 24836
rect 23548 25956 23604 25966
rect 23212 24500 23268 24780
rect 23436 24610 23492 24622
rect 23436 24558 23438 24610
rect 23490 24558 23492 24610
rect 23212 24444 23380 24500
rect 22876 24162 23044 24164
rect 22876 24110 22878 24162
rect 22930 24110 23044 24162
rect 22876 24108 23044 24110
rect 22876 24098 22932 24108
rect 22764 23716 22820 23726
rect 22764 23622 22820 23660
rect 22652 23436 22820 23492
rect 22652 23268 22708 23278
rect 22652 23174 22708 23212
rect 22652 22932 22708 22942
rect 22764 22932 22820 23436
rect 22988 23154 23044 24108
rect 23212 23714 23268 23726
rect 23212 23662 23214 23714
rect 23266 23662 23268 23714
rect 23212 23548 23268 23662
rect 23100 23492 23268 23548
rect 23324 23492 23380 24444
rect 23436 24498 23492 24558
rect 23436 24446 23438 24498
rect 23490 24446 23492 24498
rect 23436 23716 23492 24446
rect 23436 23650 23492 23660
rect 23100 23380 23156 23492
rect 23324 23436 23492 23492
rect 23100 23314 23156 23324
rect 23212 23380 23268 23390
rect 23212 23378 23380 23380
rect 23212 23326 23214 23378
rect 23266 23326 23380 23378
rect 23212 23324 23380 23326
rect 23212 23314 23268 23324
rect 22988 23102 22990 23154
rect 23042 23102 23044 23154
rect 22988 23090 23044 23102
rect 22708 22876 22820 22932
rect 22988 22932 23044 22942
rect 22988 22930 23156 22932
rect 22988 22878 22990 22930
rect 23042 22878 23156 22930
rect 22988 22876 23156 22878
rect 22652 22866 22708 22876
rect 22988 22866 23044 22876
rect 22988 22708 23044 22718
rect 22876 22484 22932 22494
rect 22876 22146 22932 22428
rect 22876 22094 22878 22146
rect 22930 22094 22932 22146
rect 22764 21924 22820 21934
rect 22652 21588 22708 21598
rect 22652 20804 22708 21532
rect 22652 20710 22708 20748
rect 22764 21586 22820 21868
rect 22764 21534 22766 21586
rect 22818 21534 22820 21586
rect 22540 19394 22596 19404
rect 22652 19348 22708 19358
rect 22652 19254 22708 19292
rect 22428 19170 22484 19180
rect 22316 18946 22372 18956
rect 22764 18788 22820 21534
rect 22876 21252 22932 22094
rect 22988 22146 23044 22652
rect 22988 22094 22990 22146
rect 23042 22094 23044 22146
rect 22988 22082 23044 22094
rect 23100 21812 23156 22876
rect 23100 21746 23156 21756
rect 23212 22370 23268 22382
rect 23212 22318 23214 22370
rect 23266 22318 23268 22370
rect 22876 21196 23156 21252
rect 22876 20804 22932 20814
rect 22932 20748 23044 20804
rect 22876 20738 22932 20748
rect 22204 18286 22206 18338
rect 22258 18286 22260 18338
rect 22204 18274 22260 18286
rect 22316 18732 22820 18788
rect 22876 20580 22932 20590
rect 22092 18162 22148 18172
rect 21420 17052 21700 17108
rect 21196 16942 21198 16994
rect 21250 16942 21252 16994
rect 21196 15764 21252 16942
rect 21532 16882 21588 16894
rect 21532 16830 21534 16882
rect 21586 16830 21588 16882
rect 21532 16660 21588 16830
rect 21644 16882 21700 17052
rect 21644 16830 21646 16882
rect 21698 16830 21700 16882
rect 21644 16818 21700 16830
rect 21812 17052 22036 17108
rect 21756 16660 21812 17052
rect 22204 16884 22260 16922
rect 22204 16818 22260 16828
rect 21532 16604 21812 16660
rect 22204 16658 22260 16670
rect 22204 16606 22206 16658
rect 22258 16606 22260 16658
rect 21308 16100 21364 16110
rect 21308 16006 21364 16044
rect 21196 15708 21476 15764
rect 21420 15540 21476 15708
rect 21624 15708 21888 15718
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21624 15642 21888 15652
rect 21756 15540 21812 15550
rect 21420 15538 21812 15540
rect 21420 15486 21758 15538
rect 21810 15486 21812 15538
rect 21420 15484 21812 15486
rect 21756 15474 21812 15484
rect 22204 15538 22260 16606
rect 22204 15486 22206 15538
rect 22258 15486 22260 15538
rect 22204 15474 22260 15486
rect 21980 15314 22036 15326
rect 21980 15262 21982 15314
rect 22034 15262 22036 15314
rect 21196 15204 21252 15242
rect 21196 15138 21252 15148
rect 21980 14756 22036 15262
rect 21756 14700 22036 14756
rect 22092 15202 22148 15214
rect 22092 15150 22094 15202
rect 22146 15150 22148 15202
rect 21532 14644 21588 14654
rect 21196 14530 21252 14542
rect 21196 14478 21198 14530
rect 21250 14478 21252 14530
rect 21196 14420 21252 14478
rect 21532 14530 21588 14588
rect 21532 14478 21534 14530
rect 21586 14478 21588 14530
rect 21532 14466 21588 14478
rect 21196 14354 21252 14364
rect 20860 14140 21140 14196
rect 21420 14306 21476 14318
rect 21420 14254 21422 14306
rect 21474 14254 21476 14306
rect 20860 13636 20916 14140
rect 21420 14084 21476 14254
rect 21756 14308 21812 14700
rect 22092 14644 22148 15150
rect 21868 14588 22148 14644
rect 22204 15204 22260 15214
rect 21868 14530 21924 14588
rect 21868 14478 21870 14530
rect 21922 14478 21924 14530
rect 21868 14466 21924 14478
rect 22092 14308 22148 14318
rect 21756 14252 22036 14308
rect 20972 14028 21476 14084
rect 21624 14140 21888 14150
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21624 14074 21888 14084
rect 20972 13858 21028 14028
rect 20972 13806 20974 13858
rect 21026 13806 21028 13858
rect 20972 13794 21028 13806
rect 21980 13748 22036 14252
rect 20860 13580 21140 13636
rect 20972 12740 21028 12750
rect 20972 12402 21028 12684
rect 20972 12350 20974 12402
rect 21026 12350 21028 12402
rect 20972 12338 21028 12350
rect 20748 11302 20804 11340
rect 20860 11954 20916 11966
rect 20860 11902 20862 11954
rect 20914 11902 20916 11954
rect 20860 10948 20916 11902
rect 20524 10332 20692 10388
rect 20748 10892 20916 10948
rect 21084 10948 21140 13580
rect 21624 12572 21888 12582
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21624 12506 21888 12516
rect 21756 12404 21812 12414
rect 21756 12310 21812 12348
rect 21980 12180 22036 13692
rect 22092 13074 22148 14252
rect 22092 13022 22094 13074
rect 22146 13022 22148 13074
rect 22092 13010 22148 13022
rect 22204 12404 22260 15148
rect 22204 12290 22260 12348
rect 22204 12238 22206 12290
rect 22258 12238 22260 12290
rect 22204 12226 22260 12238
rect 21980 12114 22036 12124
rect 22092 12178 22148 12190
rect 22092 12126 22094 12178
rect 22146 12126 22148 12178
rect 21308 11508 21364 11518
rect 21308 11414 21364 11452
rect 22092 11172 22148 12126
rect 22316 11620 22372 18732
rect 22764 17220 22820 17230
rect 22652 16996 22708 17006
rect 22652 16902 22708 16940
rect 22652 15764 22708 15774
rect 22652 15314 22708 15708
rect 22652 15262 22654 15314
rect 22706 15262 22708 15314
rect 22652 15148 22708 15262
rect 22428 15092 22708 15148
rect 22428 14642 22484 15092
rect 22764 14756 22820 17164
rect 22876 15092 22932 20524
rect 22988 17668 23044 20748
rect 23100 20244 23156 21196
rect 23100 20150 23156 20188
rect 23100 19346 23156 19358
rect 23100 19294 23102 19346
rect 23154 19294 23156 19346
rect 23100 18676 23156 19294
rect 23100 18610 23156 18620
rect 22988 17108 23044 17612
rect 23100 17108 23156 17118
rect 22988 17106 23156 17108
rect 22988 17054 23102 17106
rect 23154 17054 23156 17106
rect 22988 17052 23156 17054
rect 23100 17042 23156 17052
rect 23212 16658 23268 22318
rect 23324 20914 23380 23324
rect 23436 22484 23492 23436
rect 23436 22418 23492 22428
rect 23548 21924 23604 25900
rect 23548 21858 23604 21868
rect 23660 23378 23716 26460
rect 23884 26516 23940 26526
rect 23884 26422 23940 26460
rect 23772 25396 23828 25406
rect 23772 25302 23828 25340
rect 23772 25172 23828 25182
rect 23772 23492 23828 25116
rect 23996 23940 24052 27134
rect 24108 25060 24164 27692
rect 24444 27636 24500 28590
rect 24780 28644 24836 28654
rect 24780 28550 24836 28588
rect 24332 27580 24500 27636
rect 24668 28084 24724 28094
rect 24892 28084 24948 31164
rect 25340 30884 25396 30894
rect 25340 30790 25396 30828
rect 25026 30604 25290 30614
rect 25082 30548 25130 30604
rect 25186 30548 25234 30604
rect 25026 30538 25290 30548
rect 25340 29876 25396 29886
rect 25396 29820 25508 29876
rect 25340 29810 25396 29820
rect 25228 29316 25284 29326
rect 25228 29222 25284 29260
rect 25026 29036 25290 29046
rect 25082 28980 25130 29036
rect 25186 28980 25234 29036
rect 25026 28970 25290 28980
rect 25340 28756 25396 28766
rect 24668 28082 24948 28084
rect 24668 28030 24670 28082
rect 24722 28030 24948 28082
rect 24668 28028 24948 28030
rect 25004 28644 25060 28654
rect 24108 24994 24164 25004
rect 24220 27524 24276 27534
rect 24220 24836 24276 27468
rect 23884 23884 24052 23940
rect 24108 24780 24276 24836
rect 24332 26514 24388 27580
rect 24668 27298 24724 28028
rect 25004 27972 25060 28588
rect 25228 28644 25284 28654
rect 25340 28644 25396 28700
rect 25228 28642 25396 28644
rect 25228 28590 25230 28642
rect 25282 28590 25396 28642
rect 25228 28588 25396 28590
rect 25452 28642 25508 29820
rect 25452 28590 25454 28642
rect 25506 28590 25508 28642
rect 25228 28578 25284 28588
rect 24668 27246 24670 27298
rect 24722 27246 24724 27298
rect 24668 27234 24724 27246
rect 24780 27916 25060 27972
rect 24444 27188 24500 27198
rect 24444 27094 24500 27132
rect 24332 26462 24334 26514
rect 24386 26462 24388 26514
rect 23884 23492 23940 23884
rect 23996 23716 24052 23754
rect 23996 23650 24052 23660
rect 23996 23492 24052 23502
rect 23884 23436 23996 23492
rect 23772 23426 23828 23436
rect 23996 23426 24052 23436
rect 23660 23326 23662 23378
rect 23714 23326 23716 23378
rect 23660 22370 23716 23326
rect 23772 23268 23828 23306
rect 23772 23202 23828 23212
rect 23996 23154 24052 23166
rect 23996 23102 23998 23154
rect 24050 23102 24052 23154
rect 23884 23042 23940 23054
rect 23884 22990 23886 23042
rect 23938 22990 23940 23042
rect 23884 22708 23940 22990
rect 23884 22642 23940 22652
rect 23996 22484 24052 23102
rect 23996 22418 24052 22428
rect 23660 22318 23662 22370
rect 23714 22318 23716 22370
rect 23436 21700 23492 21710
rect 23436 21474 23492 21644
rect 23436 21422 23438 21474
rect 23490 21422 23492 21474
rect 23436 21410 23492 21422
rect 23324 20862 23326 20914
rect 23378 20862 23380 20914
rect 23324 20850 23380 20862
rect 23548 20244 23604 20254
rect 23436 18452 23492 18462
rect 23212 16606 23214 16658
rect 23266 16606 23268 16658
rect 23212 15652 23268 16606
rect 22876 15026 22932 15036
rect 23100 15596 23268 15652
rect 23324 18396 23436 18452
rect 22764 14700 22932 14756
rect 22428 14590 22430 14642
rect 22482 14590 22484 14642
rect 22428 14578 22484 14590
rect 22764 14530 22820 14542
rect 22764 14478 22766 14530
rect 22818 14478 22820 14530
rect 22764 12964 22820 14478
rect 22764 12870 22820 12908
rect 22540 12740 22596 12750
rect 22540 12290 22596 12684
rect 22540 12238 22542 12290
rect 22594 12238 22596 12290
rect 22540 12226 22596 12238
rect 22428 12066 22484 12078
rect 22428 12014 22430 12066
rect 22482 12014 22484 12066
rect 22428 11956 22484 12014
rect 22764 11956 22820 11966
rect 22428 11954 22820 11956
rect 22428 11902 22766 11954
rect 22818 11902 22820 11954
rect 22428 11900 22820 11902
rect 22764 11890 22820 11900
rect 22316 11554 22372 11564
rect 22540 11732 22596 11742
rect 22428 11508 22484 11518
rect 22092 11106 22148 11116
rect 22316 11172 22372 11182
rect 21624 11004 21888 11014
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21084 10892 21252 10948
rect 21624 10938 21888 10948
rect 20524 10052 20580 10332
rect 20748 10276 20804 10892
rect 21196 10836 21252 10892
rect 21196 10780 21588 10836
rect 20524 9986 20580 9996
rect 20636 10220 20804 10276
rect 20860 10722 20916 10734
rect 20860 10670 20862 10722
rect 20914 10670 20916 10722
rect 20860 10276 20916 10670
rect 21196 10610 21252 10622
rect 21196 10558 21198 10610
rect 21250 10558 21252 10610
rect 21196 10500 21252 10558
rect 21308 10612 21364 10622
rect 21308 10518 21364 10556
rect 21420 10610 21476 10622
rect 21420 10558 21422 10610
rect 21474 10558 21476 10610
rect 21196 10434 21252 10444
rect 21420 10388 21476 10558
rect 21308 10332 21476 10388
rect 21308 10276 21364 10332
rect 21532 10276 21588 10780
rect 22316 10834 22372 11116
rect 22316 10782 22318 10834
rect 22370 10782 22372 10834
rect 22316 10770 22372 10782
rect 22428 10834 22484 11452
rect 22428 10782 22430 10834
rect 22482 10782 22484 10834
rect 22428 10770 22484 10782
rect 22540 10836 22596 11676
rect 21644 10724 21700 10734
rect 21644 10630 21700 10668
rect 22204 10612 22260 10622
rect 22540 10612 22596 10780
rect 22652 10724 22708 10734
rect 22652 10630 22708 10668
rect 22204 10610 22596 10612
rect 22204 10558 22206 10610
rect 22258 10558 22596 10610
rect 22204 10556 22596 10558
rect 22204 10546 22260 10556
rect 20860 10220 21364 10276
rect 21420 10220 21588 10276
rect 21980 10500 22036 10510
rect 20636 8372 20692 10220
rect 20748 9964 20804 9976
rect 20748 9912 20750 9964
rect 20802 9940 20804 9964
rect 20860 9940 20916 10220
rect 20802 9912 20916 9940
rect 20748 9884 20916 9912
rect 21420 9268 21476 10220
rect 21532 10052 21588 10062
rect 21532 9938 21588 9996
rect 21532 9886 21534 9938
rect 21586 9886 21588 9938
rect 21532 9874 21588 9886
rect 21980 9938 22036 10444
rect 21980 9886 21982 9938
rect 22034 9886 22036 9938
rect 21624 9436 21888 9446
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21624 9370 21888 9380
rect 21420 9212 21588 9268
rect 20636 8258 20692 8316
rect 20636 8206 20638 8258
rect 20690 8206 20692 8258
rect 20636 8194 20692 8206
rect 20972 8932 21028 8942
rect 20748 8146 20804 8158
rect 20748 8094 20750 8146
rect 20802 8094 20804 8146
rect 20636 8036 20692 8046
rect 20524 7700 20580 7710
rect 20524 7474 20580 7644
rect 20636 7698 20692 7980
rect 20636 7646 20638 7698
rect 20690 7646 20692 7698
rect 20636 7634 20692 7646
rect 20524 7422 20526 7474
rect 20578 7422 20580 7474
rect 20524 7410 20580 7422
rect 20356 7308 20468 7364
rect 20300 7298 20356 7308
rect 20748 6804 20804 8094
rect 20412 6748 20804 6804
rect 20076 6690 20132 6702
rect 20076 6638 20078 6690
rect 20130 6638 20132 6690
rect 20076 6020 20132 6638
rect 20076 5926 20132 5964
rect 20412 5348 20468 6748
rect 20972 6692 21028 8876
rect 21196 8372 21252 8382
rect 21420 8372 21476 8382
rect 21252 8370 21476 8372
rect 21252 8318 21422 8370
rect 21474 8318 21476 8370
rect 21252 8316 21476 8318
rect 21196 8306 21252 8316
rect 21420 8306 21476 8316
rect 21532 8148 21588 9212
rect 21980 9156 22036 9886
rect 21980 9090 22036 9100
rect 22652 9044 22708 9054
rect 22652 8370 22708 8988
rect 22652 8318 22654 8370
rect 22706 8318 22708 8370
rect 22652 8306 22708 8318
rect 21420 8092 21588 8148
rect 22092 8258 22148 8270
rect 22092 8206 22094 8258
rect 22146 8206 22148 8258
rect 20972 6626 21028 6636
rect 21196 7474 21252 7486
rect 21196 7422 21198 7474
rect 21250 7422 21252 7474
rect 20524 6580 20580 6590
rect 20524 6486 20580 6524
rect 20412 5282 20468 5292
rect 20860 5908 20916 5918
rect 21196 5908 21252 7422
rect 21308 6580 21364 6590
rect 21308 6486 21364 6524
rect 21420 6130 21476 8092
rect 21624 7868 21888 7878
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21624 7802 21888 7812
rect 22092 7700 22148 8206
rect 22092 7634 22148 7644
rect 22316 8258 22372 8270
rect 22316 8206 22318 8258
rect 22370 8206 22372 8258
rect 21644 6692 21700 6702
rect 21644 6598 21700 6636
rect 22092 6690 22148 6702
rect 22092 6638 22094 6690
rect 22146 6638 22148 6690
rect 21624 6300 21888 6310
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21624 6234 21888 6244
rect 21420 6078 21422 6130
rect 21474 6078 21476 6130
rect 21420 6066 21476 6078
rect 21868 6020 21924 6030
rect 22092 6020 22148 6638
rect 21868 6018 22148 6020
rect 21868 5966 21870 6018
rect 21922 5966 22148 6018
rect 21868 5964 22148 5966
rect 21756 5908 21812 5918
rect 21196 5906 21812 5908
rect 21196 5854 21758 5906
rect 21810 5854 21812 5906
rect 21196 5852 21812 5854
rect 20636 5122 20692 5134
rect 20636 5070 20638 5122
rect 20690 5070 20692 5122
rect 20412 5012 20468 5022
rect 20412 4918 20468 4956
rect 20076 4898 20132 4910
rect 20076 4846 20078 4898
rect 20130 4846 20132 4898
rect 20076 4676 20132 4846
rect 20524 4898 20580 4910
rect 20524 4846 20526 4898
rect 20578 4846 20580 4898
rect 20524 4676 20580 4846
rect 20636 4900 20692 5070
rect 20636 4834 20692 4844
rect 20748 5124 20804 5134
rect 20076 4610 20132 4620
rect 20188 4620 20580 4676
rect 20636 4676 20692 4686
rect 20076 3780 20132 3790
rect 19964 3778 20132 3780
rect 19964 3726 20078 3778
rect 20130 3726 20132 3778
rect 19964 3724 20132 3726
rect 20076 3714 20132 3724
rect 19852 3500 20020 3556
rect 19404 3378 19460 3388
rect 19628 3442 19684 3454
rect 19628 3390 19630 3442
rect 19682 3390 19684 3442
rect 19180 3154 19236 3164
rect 19292 3108 19348 3118
rect 19348 3052 19460 3108
rect 19292 3042 19348 3052
rect 18956 2772 19012 2782
rect 18956 2770 19348 2772
rect 18956 2718 18958 2770
rect 19010 2718 19348 2770
rect 18956 2716 19348 2718
rect 18956 2706 19012 2716
rect 18956 2100 19012 2110
rect 18956 2006 19012 2044
rect 18844 1810 18900 1820
rect 19292 1874 19348 2716
rect 19292 1822 19294 1874
rect 19346 1822 19348 1874
rect 19292 1810 19348 1822
rect 19404 1876 19460 3052
rect 19516 2884 19572 2894
rect 19628 2884 19684 3390
rect 19964 3444 20020 3500
rect 19964 3378 20020 3388
rect 20076 3554 20132 3566
rect 20076 3502 20078 3554
rect 20130 3502 20132 3554
rect 19516 2882 19684 2884
rect 19516 2830 19518 2882
rect 19570 2830 19684 2882
rect 19516 2828 19684 2830
rect 19516 2818 19572 2828
rect 20076 2660 20132 3502
rect 20188 3388 20244 4620
rect 20636 4450 20692 4620
rect 20636 4398 20638 4450
rect 20690 4398 20692 4450
rect 20636 4386 20692 4398
rect 20748 4228 20804 5068
rect 20412 4172 20804 4228
rect 20300 3780 20356 3790
rect 20300 3554 20356 3724
rect 20300 3502 20302 3554
rect 20354 3502 20356 3554
rect 20300 3490 20356 3502
rect 20188 3332 20356 3388
rect 19852 2604 20132 2660
rect 19404 1810 19460 1820
rect 19516 1988 19572 1998
rect 18732 1484 18900 1540
rect 18844 400 18900 1484
rect 19516 400 19572 1932
rect 19852 1986 19908 2604
rect 19852 1934 19854 1986
rect 19906 1934 19908 1986
rect 19852 1922 19908 1934
rect 20076 2212 20132 2222
rect 19628 1876 19684 1886
rect 19628 1782 19684 1820
rect 20076 1874 20132 2156
rect 20188 1988 20244 1998
rect 20300 1988 20356 3332
rect 20188 1986 20356 1988
rect 20188 1934 20190 1986
rect 20242 1934 20356 1986
rect 20188 1932 20356 1934
rect 20188 1922 20244 1932
rect 20076 1822 20078 1874
rect 20130 1822 20132 1874
rect 20076 1810 20132 1822
rect 20412 1764 20468 4172
rect 20524 4004 20580 4014
rect 20524 1988 20580 3948
rect 20524 1922 20580 1932
rect 20636 3892 20692 3902
rect 20636 1876 20692 3836
rect 20748 3220 20804 3230
rect 20748 2882 20804 3164
rect 20748 2830 20750 2882
rect 20802 2830 20804 2882
rect 20748 2212 20804 2830
rect 20860 2658 20916 5852
rect 21756 5236 21812 5852
rect 21868 5908 21924 5964
rect 21868 5842 21924 5852
rect 21756 5170 21812 5180
rect 22204 5684 22260 5694
rect 22316 5684 22372 8206
rect 22764 7700 22820 7710
rect 22876 7700 22932 14700
rect 23100 13634 23156 15596
rect 23324 15540 23380 18396
rect 23436 18386 23492 18396
rect 23436 17556 23492 17566
rect 23436 17462 23492 17500
rect 23548 17106 23604 20188
rect 23660 20130 23716 22318
rect 23772 22372 23828 22382
rect 23772 20244 23828 22316
rect 23996 22258 24052 22270
rect 23996 22206 23998 22258
rect 24050 22206 24052 22258
rect 23996 20804 24052 22206
rect 23996 20738 24052 20748
rect 23772 20178 23828 20188
rect 23660 20078 23662 20130
rect 23714 20078 23716 20130
rect 23660 20020 23716 20078
rect 24108 20132 24164 24780
rect 24220 24612 24276 24622
rect 24220 24518 24276 24556
rect 24220 24388 24276 24398
rect 24220 23380 24276 24332
rect 24332 23716 24388 26462
rect 24556 26964 24612 26974
rect 24556 25506 24612 26908
rect 24556 25454 24558 25506
rect 24610 25454 24612 25506
rect 24332 23650 24388 23660
rect 24444 25060 24500 25070
rect 24220 23324 24388 23380
rect 24220 23154 24276 23166
rect 24220 23102 24222 23154
rect 24274 23102 24276 23154
rect 24220 22036 24276 23102
rect 24332 22596 24388 23324
rect 24444 22820 24500 25004
rect 24556 24388 24612 25454
rect 24780 24724 24836 27916
rect 25026 27468 25290 27478
rect 25082 27412 25130 27468
rect 25186 27412 25234 27468
rect 25026 27402 25290 27412
rect 25228 27300 25284 27310
rect 25228 27186 25284 27244
rect 25228 27134 25230 27186
rect 25282 27134 25284 27186
rect 25228 27122 25284 27134
rect 25340 27076 25396 27086
rect 24892 26852 24948 26862
rect 24892 26758 24948 26796
rect 25228 26516 25284 26526
rect 25340 26516 25396 27020
rect 25452 26908 25508 28590
rect 25564 28084 25620 32172
rect 26236 32004 26292 32014
rect 26124 31668 26180 31678
rect 26124 31108 26180 31612
rect 26124 31014 26180 31052
rect 25900 30996 25956 31006
rect 25900 30902 25956 30940
rect 26236 30212 26292 31948
rect 26348 30994 26404 32286
rect 26348 30942 26350 30994
rect 26402 30942 26404 30994
rect 26348 30930 26404 30942
rect 26460 30994 26516 32396
rect 26460 30942 26462 30994
rect 26514 30942 26516 30994
rect 26460 30772 26516 30942
rect 26572 30996 26628 34524
rect 26684 34354 26740 34366
rect 26684 34302 26686 34354
rect 26738 34302 26740 34354
rect 26684 33460 26740 34302
rect 26684 33394 26740 33404
rect 26684 32340 26740 32350
rect 26684 31948 26740 32284
rect 26796 32116 26852 36316
rect 27132 35026 27188 36428
rect 27356 36418 27412 36428
rect 27244 36258 27300 36270
rect 27244 36206 27246 36258
rect 27298 36206 27300 36258
rect 27244 35812 27300 36206
rect 27356 35812 27412 35822
rect 27244 35810 27412 35812
rect 27244 35758 27358 35810
rect 27410 35758 27412 35810
rect 27244 35756 27412 35758
rect 27356 35746 27412 35756
rect 27132 34974 27134 35026
rect 27186 34974 27188 35026
rect 27132 34692 27188 34974
rect 27132 34626 27188 34636
rect 27356 34916 27412 34926
rect 27132 34242 27188 34254
rect 27356 34244 27412 34860
rect 27692 34690 27748 34702
rect 27692 34638 27694 34690
rect 27746 34638 27748 34690
rect 27692 34468 27748 34638
rect 27692 34402 27748 34412
rect 27804 34692 27860 34702
rect 27804 34354 27860 34636
rect 27804 34302 27806 34354
rect 27858 34302 27860 34354
rect 27804 34244 27860 34302
rect 27132 34190 27134 34242
rect 27186 34190 27188 34242
rect 27020 33908 27076 33918
rect 27020 33814 27076 33852
rect 27020 33348 27076 33358
rect 27132 33348 27188 34190
rect 27076 33292 27188 33348
rect 27244 34242 27412 34244
rect 27244 34190 27358 34242
rect 27410 34190 27412 34242
rect 27244 34188 27412 34190
rect 27020 33282 27076 33292
rect 27132 32788 27188 32798
rect 27244 32788 27300 34188
rect 27356 34178 27412 34188
rect 27580 34188 27860 34244
rect 27356 33460 27412 33470
rect 27356 33366 27412 33404
rect 27132 32786 27300 32788
rect 27132 32734 27134 32786
rect 27186 32734 27300 32786
rect 27132 32732 27300 32734
rect 27132 32722 27188 32732
rect 26796 32050 26852 32060
rect 27244 31948 27300 32732
rect 26684 31892 26964 31948
rect 27244 31892 27524 31948
rect 26684 31668 26740 31678
rect 26684 31218 26740 31612
rect 26684 31166 26686 31218
rect 26738 31166 26740 31218
rect 26684 31154 26740 31166
rect 26572 30940 26852 30996
rect 26460 30716 26740 30772
rect 26236 30146 26292 30156
rect 25676 28644 25732 28654
rect 25676 28550 25732 28588
rect 26460 28644 26516 28654
rect 26460 28550 26516 28588
rect 26124 28532 26180 28542
rect 26348 28532 26404 28542
rect 26124 28530 26292 28532
rect 26124 28478 26126 28530
rect 26178 28478 26292 28530
rect 26124 28476 26292 28478
rect 26124 28466 26180 28476
rect 25788 28420 25844 28430
rect 25676 28084 25732 28094
rect 25564 28082 25732 28084
rect 25564 28030 25678 28082
rect 25730 28030 25732 28082
rect 25564 28028 25732 28030
rect 25676 28018 25732 28028
rect 25452 26852 25620 26908
rect 25228 26514 25396 26516
rect 25228 26462 25230 26514
rect 25282 26462 25396 26514
rect 25228 26460 25396 26462
rect 25228 26450 25284 26460
rect 24892 26292 24948 26302
rect 24892 25618 24948 26236
rect 25452 26292 25508 26302
rect 25452 26198 25508 26236
rect 25340 26178 25396 26190
rect 25340 26126 25342 26178
rect 25394 26126 25396 26178
rect 25340 26068 25396 26126
rect 25340 26012 25508 26068
rect 25026 25900 25290 25910
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25026 25834 25290 25844
rect 24892 25566 24894 25618
rect 24946 25566 24948 25618
rect 24892 25554 24948 25566
rect 25452 25396 25508 26012
rect 24780 24658 24836 24668
rect 25340 25340 25508 25396
rect 25340 24722 25396 25340
rect 25340 24670 25342 24722
rect 25394 24670 25396 24722
rect 25340 24658 25396 24670
rect 25452 24948 25508 24958
rect 25452 24834 25508 24892
rect 25452 24782 25454 24834
rect 25506 24782 25508 24834
rect 24668 24612 24724 24622
rect 24668 24518 24724 24556
rect 24556 24332 24724 24388
rect 24556 24164 24612 24174
rect 24556 24050 24612 24108
rect 24556 23998 24558 24050
rect 24610 23998 24612 24050
rect 24556 23986 24612 23998
rect 24668 23044 24724 24332
rect 25026 24332 25290 24342
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25026 24266 25290 24276
rect 25340 24052 25396 24062
rect 25340 23958 25396 23996
rect 25004 23940 25060 23950
rect 24668 22950 24724 22988
rect 24892 23884 25004 23940
rect 24444 22764 24836 22820
rect 24332 22540 24612 22596
rect 24556 22482 24612 22540
rect 24556 22430 24558 22482
rect 24610 22430 24612 22482
rect 24220 21980 24500 22036
rect 24332 21812 24388 21822
rect 24332 21718 24388 21756
rect 24220 21698 24276 21710
rect 24220 21646 24222 21698
rect 24274 21646 24276 21698
rect 24220 21588 24276 21646
rect 24444 21588 24500 21980
rect 24220 21522 24276 21532
rect 24332 21532 24500 21588
rect 24108 20076 24276 20132
rect 23660 19964 24164 20020
rect 24108 19906 24164 19964
rect 24108 19854 24110 19906
rect 24162 19854 24164 19906
rect 24108 19842 24164 19854
rect 23996 18450 24052 18462
rect 23996 18398 23998 18450
rect 24050 18398 24052 18450
rect 23996 17220 24052 18398
rect 23996 17154 24052 17164
rect 24108 17668 24164 17678
rect 23548 17054 23550 17106
rect 23602 17054 23604 17106
rect 23548 17042 23604 17054
rect 24108 16212 24164 17612
rect 24220 16548 24276 20076
rect 24332 18676 24388 21532
rect 24444 21362 24500 21374
rect 24444 21310 24446 21362
rect 24498 21310 24500 21362
rect 24444 20692 24500 21310
rect 24444 19348 24500 20636
rect 24444 19282 24500 19292
rect 24332 18610 24388 18620
rect 24444 19012 24500 19022
rect 24332 17108 24388 17118
rect 24444 17108 24500 18956
rect 24332 17106 24500 17108
rect 24332 17054 24334 17106
rect 24386 17054 24500 17106
rect 24332 17052 24500 17054
rect 24332 17042 24388 17052
rect 24220 16492 24388 16548
rect 23212 15484 23380 15540
rect 23660 16210 24164 16212
rect 23660 16158 24110 16210
rect 24162 16158 24164 16210
rect 23660 16156 24164 16158
rect 23212 15314 23268 15484
rect 23212 15262 23214 15314
rect 23266 15262 23268 15314
rect 23212 14420 23268 15262
rect 23324 15316 23380 15326
rect 23324 15314 23492 15316
rect 23324 15262 23326 15314
rect 23378 15262 23492 15314
rect 23324 15260 23492 15262
rect 23324 15250 23380 15260
rect 23436 14644 23492 15260
rect 23548 15314 23604 15326
rect 23548 15262 23550 15314
rect 23602 15262 23604 15314
rect 23548 15204 23604 15262
rect 23548 15138 23604 15148
rect 23548 14644 23604 14654
rect 23436 14642 23604 14644
rect 23436 14590 23550 14642
rect 23602 14590 23604 14642
rect 23436 14588 23604 14590
rect 23548 14578 23604 14588
rect 23212 14354 23268 14364
rect 23548 13748 23604 13758
rect 23548 13654 23604 13692
rect 23100 13582 23102 13634
rect 23154 13582 23156 13634
rect 23100 13570 23156 13582
rect 23436 12962 23492 12974
rect 23436 12910 23438 12962
rect 23490 12910 23492 12962
rect 22988 12740 23044 12750
rect 22988 12402 23044 12684
rect 22988 12350 22990 12402
rect 23042 12350 23044 12402
rect 22988 9938 23044 12350
rect 23436 12180 23492 12910
rect 23548 12964 23604 12974
rect 23660 12964 23716 16156
rect 24108 16146 24164 16156
rect 24220 15540 24276 15550
rect 23772 15538 24276 15540
rect 23772 15486 24222 15538
rect 24274 15486 24276 15538
rect 23772 15484 24276 15486
rect 23772 15426 23828 15484
rect 24220 15474 24276 15484
rect 24332 15538 24388 16492
rect 24332 15486 24334 15538
rect 24386 15486 24388 15538
rect 23772 15374 23774 15426
rect 23826 15374 23828 15426
rect 23772 15362 23828 15374
rect 24108 15316 24164 15326
rect 24108 15222 24164 15260
rect 24332 14756 24388 15486
rect 24556 15316 24612 22430
rect 24668 20132 24724 20142
rect 24668 20038 24724 20076
rect 24668 19348 24724 19358
rect 24668 18564 24724 19292
rect 24668 18450 24724 18508
rect 24668 18398 24670 18450
rect 24722 18398 24724 18450
rect 24668 18386 24724 18398
rect 24668 17220 24724 17230
rect 24668 17106 24724 17164
rect 24668 17054 24670 17106
rect 24722 17054 24724 17106
rect 24668 17042 24724 17054
rect 24556 15250 24612 15260
rect 24668 15540 24724 15550
rect 24668 15314 24724 15484
rect 24668 15262 24670 15314
rect 24722 15262 24724 15314
rect 24668 15250 24724 15262
rect 24332 14690 24388 14700
rect 24444 14420 24500 14430
rect 24220 13636 24276 13646
rect 23604 12908 23716 12964
rect 24108 13076 24164 13086
rect 23548 12404 23604 12908
rect 23548 12402 24052 12404
rect 23548 12350 23550 12402
rect 23602 12350 24052 12402
rect 23548 12348 24052 12350
rect 23548 12338 23604 12348
rect 23436 12114 23492 12124
rect 23436 11954 23492 11966
rect 23436 11902 23438 11954
rect 23490 11902 23492 11954
rect 23436 11506 23492 11902
rect 23436 11454 23438 11506
rect 23490 11454 23492 11506
rect 23436 11442 23492 11454
rect 23996 11396 24052 12348
rect 24108 12402 24164 13020
rect 24108 12350 24110 12402
rect 24162 12350 24164 12402
rect 24108 12338 24164 12350
rect 24108 11396 24164 11406
rect 23996 11394 24164 11396
rect 23996 11342 24110 11394
rect 24162 11342 24164 11394
rect 23996 11340 24164 11342
rect 24108 11330 24164 11340
rect 24108 10836 24164 10846
rect 24108 10742 24164 10780
rect 23212 10724 23268 10734
rect 23212 10630 23268 10668
rect 23660 10724 23716 10734
rect 23660 10630 23716 10668
rect 22988 9886 22990 9938
rect 23042 9886 23044 9938
rect 22988 9874 23044 9886
rect 24220 9266 24276 13580
rect 24444 13636 24500 14364
rect 24668 13636 24724 13646
rect 24444 13634 24724 13636
rect 24444 13582 24670 13634
rect 24722 13582 24724 13634
rect 24444 13580 24724 13582
rect 24444 13076 24500 13580
rect 24668 13570 24724 13580
rect 24444 12982 24500 13020
rect 24668 12180 24724 12190
rect 24668 12068 24724 12124
rect 24220 9214 24222 9266
rect 24274 9214 24276 9266
rect 24220 9202 24276 9214
rect 24444 12066 24724 12068
rect 24444 12014 24670 12066
rect 24722 12014 24724 12066
rect 24444 12012 24724 12014
rect 23436 9044 23492 9054
rect 23436 8950 23492 8988
rect 23996 8146 24052 8158
rect 23996 8094 23998 8146
rect 24050 8094 24052 8146
rect 22764 7698 22932 7700
rect 22764 7646 22766 7698
rect 22818 7646 22932 7698
rect 22764 7644 22932 7646
rect 23212 7700 23268 7710
rect 22764 7634 22820 7644
rect 23212 7606 23268 7644
rect 22428 7474 22484 7486
rect 22428 7422 22430 7474
rect 22482 7422 22484 7474
rect 22428 6914 22484 7422
rect 22428 6862 22430 6914
rect 22482 6862 22484 6914
rect 22428 6850 22484 6862
rect 23660 7474 23716 7486
rect 23660 7422 23662 7474
rect 23714 7422 23716 7474
rect 22540 6580 22596 6590
rect 22260 5628 22372 5684
rect 22428 6578 22596 6580
rect 22428 6526 22542 6578
rect 22594 6526 22596 6578
rect 22428 6524 22596 6526
rect 22428 5796 22484 6524
rect 22540 6514 22596 6524
rect 23660 6132 23716 7422
rect 23772 7474 23828 7486
rect 23772 7422 23774 7474
rect 23826 7422 23828 7474
rect 23772 6692 23828 7422
rect 23884 7476 23940 7486
rect 23884 7382 23940 7420
rect 23772 6626 23828 6636
rect 23884 6580 23940 6590
rect 23996 6580 24052 8094
rect 24444 8034 24500 12012
rect 24668 12002 24724 12012
rect 24668 11396 24724 11406
rect 24780 11396 24836 22764
rect 24892 22484 24948 23884
rect 25004 23874 25060 23884
rect 25452 23828 25508 24782
rect 25564 24612 25620 26852
rect 25788 26852 25844 28364
rect 26236 28420 26292 28476
rect 26348 28438 26404 28476
rect 26572 28420 26628 28430
rect 26236 28354 26292 28364
rect 26460 28418 26628 28420
rect 26460 28366 26574 28418
rect 26626 28366 26628 28418
rect 26460 28364 26628 28366
rect 26124 28308 26180 28318
rect 25900 27972 25956 27982
rect 25900 27878 25956 27916
rect 26124 27970 26180 28252
rect 26460 28084 26516 28364
rect 26572 28354 26628 28364
rect 26684 28308 26740 30716
rect 26684 28242 26740 28252
rect 26124 27918 26126 27970
rect 26178 27918 26180 27970
rect 26124 27906 26180 27918
rect 26236 28028 26516 28084
rect 26572 28196 26628 28206
rect 26124 27412 26180 27422
rect 26124 26908 26180 27356
rect 26236 27076 26292 28028
rect 26460 27860 26516 27870
rect 26348 27636 26404 27646
rect 26348 27542 26404 27580
rect 26236 27010 26292 27020
rect 26460 27188 26516 27804
rect 25900 26852 25956 26862
rect 26124 26852 26292 26908
rect 25788 26796 25900 26852
rect 25900 26290 25956 26796
rect 26236 26514 26292 26852
rect 26236 26462 26238 26514
rect 26290 26462 26292 26514
rect 26236 26450 26292 26462
rect 25900 26238 25902 26290
rect 25954 26238 25956 26290
rect 25900 26180 25956 26238
rect 25956 26124 26292 26180
rect 25900 26086 25956 26124
rect 25676 25396 25732 25406
rect 25676 24946 25732 25340
rect 25676 24894 25678 24946
rect 25730 24894 25732 24946
rect 25676 24882 25732 24894
rect 25900 24724 25956 24734
rect 25900 24630 25956 24668
rect 25564 24546 25620 24556
rect 26124 24612 26180 24622
rect 25452 23762 25508 23772
rect 25004 23716 25060 23726
rect 25004 23622 25060 23660
rect 26012 23716 26068 23726
rect 25676 23492 25732 23502
rect 25228 23268 25284 23278
rect 25228 23044 25284 23212
rect 25228 23042 25508 23044
rect 25228 22990 25230 23042
rect 25282 22990 25508 23042
rect 25228 22988 25508 22990
rect 25228 22978 25284 22988
rect 25026 22764 25290 22774
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25026 22698 25290 22708
rect 25116 22596 25172 22606
rect 25004 22484 25060 22494
rect 24892 22482 25060 22484
rect 24892 22430 25006 22482
rect 25058 22430 25060 22482
rect 24892 22428 25060 22430
rect 25004 22418 25060 22428
rect 24892 22260 24948 22270
rect 25116 22260 25172 22540
rect 25228 22372 25284 22382
rect 25452 22372 25508 22988
rect 25228 22370 25508 22372
rect 25228 22318 25230 22370
rect 25282 22318 25508 22370
rect 25228 22316 25508 22318
rect 25228 22306 25284 22316
rect 24892 22258 25116 22260
rect 24892 22206 24894 22258
rect 24946 22206 25116 22258
rect 24892 22204 25116 22206
rect 24892 22194 24948 22204
rect 25116 22166 25172 22204
rect 25452 21588 25508 21598
rect 25026 21196 25290 21206
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25026 21130 25290 21140
rect 25452 20914 25508 21532
rect 25452 20862 25454 20914
rect 25506 20862 25508 20914
rect 25452 20356 25508 20862
rect 25452 20290 25508 20300
rect 25340 20020 25396 20030
rect 25340 19926 25396 19964
rect 25026 19628 25290 19638
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25026 19562 25290 19572
rect 25452 19236 25508 19246
rect 25228 19124 25284 19134
rect 25228 19122 25396 19124
rect 25228 19070 25230 19122
rect 25282 19070 25396 19122
rect 25228 19068 25396 19070
rect 25228 19058 25284 19068
rect 25340 18674 25396 19068
rect 25340 18622 25342 18674
rect 25394 18622 25396 18674
rect 25340 18610 25396 18622
rect 25228 18452 25284 18462
rect 25228 18358 25284 18396
rect 25452 18452 25508 19180
rect 25676 19012 25732 23436
rect 26012 22370 26068 23660
rect 26012 22318 26014 22370
rect 26066 22318 26068 22370
rect 26012 21586 26068 22318
rect 26012 21534 26014 21586
rect 26066 21534 26068 21586
rect 25788 21364 25844 21374
rect 25788 20692 25844 21308
rect 25788 20598 25844 20636
rect 25900 20578 25956 20590
rect 25900 20526 25902 20578
rect 25954 20526 25956 20578
rect 25900 20132 25956 20526
rect 26012 20356 26068 21534
rect 26124 20802 26180 24556
rect 26236 24610 26292 26124
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 24388 26292 24558
rect 26236 24322 26292 24332
rect 26460 24164 26516 27132
rect 26572 24276 26628 28140
rect 26684 28082 26740 28094
rect 26684 28030 26686 28082
rect 26738 28030 26740 28082
rect 26684 27188 26740 28030
rect 26684 27122 26740 27132
rect 26796 26908 26852 30940
rect 26572 24210 26628 24220
rect 26684 26852 26852 26908
rect 26124 20750 26126 20802
rect 26178 20750 26180 20802
rect 26124 20692 26180 20750
rect 26236 24108 26516 24164
rect 26236 24052 26292 24108
rect 26684 24052 26740 26852
rect 26908 26514 26964 31892
rect 27356 31668 27412 31678
rect 27356 31574 27412 31612
rect 27132 30882 27188 30894
rect 27132 30830 27134 30882
rect 27186 30830 27188 30882
rect 27132 30100 27188 30830
rect 27132 30034 27188 30044
rect 27244 30770 27300 30782
rect 27244 30718 27246 30770
rect 27298 30718 27300 30770
rect 27132 28756 27188 28766
rect 27244 28756 27300 30718
rect 27132 28754 27300 28756
rect 27132 28702 27134 28754
rect 27186 28702 27300 28754
rect 27132 28700 27300 28702
rect 27356 29314 27412 29326
rect 27356 29262 27358 29314
rect 27410 29262 27412 29314
rect 27356 28756 27412 29262
rect 27132 28690 27188 28700
rect 27356 28690 27412 28700
rect 27468 28754 27524 31892
rect 27468 28702 27470 28754
rect 27522 28702 27524 28754
rect 27132 27970 27188 27982
rect 27132 27918 27134 27970
rect 27186 27918 27188 27970
rect 27020 27636 27076 27646
rect 27020 27542 27076 27580
rect 27020 27300 27076 27310
rect 27132 27300 27188 27918
rect 27356 27972 27412 27982
rect 27468 27972 27524 28702
rect 27356 27970 27524 27972
rect 27356 27918 27358 27970
rect 27410 27918 27524 27970
rect 27356 27916 27524 27918
rect 27580 30884 27636 34188
rect 27916 34132 27972 37102
rect 28140 37828 28196 38612
rect 27580 27972 27636 30828
rect 27804 34076 27972 34132
rect 28028 35698 28084 35710
rect 28028 35646 28030 35698
rect 28082 35646 28084 35698
rect 28028 34804 28084 35646
rect 27804 28196 27860 34076
rect 28028 33346 28084 34748
rect 28028 33294 28030 33346
rect 28082 33294 28084 33346
rect 27916 32452 27972 32462
rect 27916 32358 27972 32396
rect 28028 31778 28084 33294
rect 28028 31726 28030 31778
rect 28082 31726 28084 31778
rect 27916 30100 27972 30110
rect 28028 30100 28084 31726
rect 28140 34690 28196 37772
rect 28428 37660 28692 37670
rect 28484 37604 28532 37660
rect 28588 37604 28636 37660
rect 28428 37594 28692 37604
rect 28428 36092 28692 36102
rect 28484 36036 28532 36092
rect 28588 36036 28636 36092
rect 28428 36026 28692 36036
rect 28140 34638 28142 34690
rect 28194 34638 28196 34690
rect 28140 34468 28196 34638
rect 28428 34524 28692 34534
rect 28484 34468 28532 34524
rect 28588 34468 28636 34524
rect 28428 34458 28692 34468
rect 28140 30882 28196 34412
rect 28428 32956 28692 32966
rect 28484 32900 28532 32956
rect 28588 32900 28636 32956
rect 28428 32890 28692 32900
rect 28428 31388 28692 31398
rect 28484 31332 28532 31388
rect 28588 31332 28636 31388
rect 28428 31322 28692 31332
rect 28140 30830 28142 30882
rect 28194 30830 28196 30882
rect 28140 30770 28196 30830
rect 28140 30718 28142 30770
rect 28194 30718 28196 30770
rect 28140 30706 28196 30718
rect 27972 30044 28084 30100
rect 27916 29428 27972 30044
rect 28428 29820 28692 29830
rect 28484 29764 28532 29820
rect 28588 29764 28636 29820
rect 28428 29754 28692 29764
rect 28140 29428 28196 29438
rect 27916 29426 28196 29428
rect 27916 29374 28142 29426
rect 28194 29374 28196 29426
rect 27916 29372 28196 29374
rect 27804 28130 27860 28140
rect 28140 28418 28196 29372
rect 28140 28366 28142 28418
rect 28194 28366 28196 28418
rect 27804 27972 27860 27982
rect 27580 27916 27804 27972
rect 27356 27906 27412 27916
rect 27076 27244 27188 27300
rect 27020 27234 27076 27244
rect 27356 27188 27412 27198
rect 27356 27094 27412 27132
rect 26908 26462 26910 26514
rect 26962 26462 26964 26514
rect 26908 24836 26964 26462
rect 27244 27076 27300 27086
rect 27020 25396 27076 25406
rect 27020 25302 27076 25340
rect 26908 24780 27076 24836
rect 26236 23938 26292 23996
rect 26460 23996 26740 24052
rect 26908 24610 26964 24622
rect 26908 24558 26910 24610
rect 26962 24558 26964 24610
rect 26236 23886 26238 23938
rect 26290 23886 26292 23938
rect 26236 21700 26292 23886
rect 26348 23940 26404 23950
rect 26348 23846 26404 23884
rect 26236 20804 26292 21644
rect 26348 21028 26404 21038
rect 26348 20934 26404 20972
rect 26348 20804 26404 20814
rect 26236 20802 26404 20804
rect 26236 20750 26350 20802
rect 26402 20750 26404 20802
rect 26236 20748 26404 20750
rect 26124 20626 26180 20636
rect 26012 20300 26180 20356
rect 26012 20132 26068 20142
rect 25900 20130 26068 20132
rect 25900 20078 26014 20130
rect 26066 20078 26068 20130
rect 25900 20076 26068 20078
rect 26012 20066 26068 20076
rect 25900 19234 25956 19246
rect 25900 19182 25902 19234
rect 25954 19182 25956 19234
rect 25676 18956 25844 19012
rect 25676 18452 25732 18462
rect 25452 18450 25620 18452
rect 25452 18398 25454 18450
rect 25506 18398 25620 18450
rect 25452 18396 25620 18398
rect 25452 18386 25508 18396
rect 25026 18060 25290 18070
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25026 17994 25290 18004
rect 25228 17778 25284 17790
rect 25228 17726 25230 17778
rect 25282 17726 25284 17778
rect 25228 17444 25284 17726
rect 25228 17378 25284 17388
rect 25026 16492 25290 16502
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25026 16426 25290 16436
rect 25026 14924 25290 14934
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25026 14858 25290 14868
rect 25452 13972 25508 13982
rect 25564 13972 25620 18396
rect 25676 18358 25732 18396
rect 25788 15314 25844 18956
rect 25900 17668 25956 19182
rect 26124 19124 26180 20300
rect 25900 17602 25956 17612
rect 26012 19068 26180 19124
rect 26012 17220 26068 19068
rect 26348 19012 26404 20748
rect 26460 19236 26516 23996
rect 26572 23828 26628 23838
rect 26572 20132 26628 23772
rect 26796 23828 26852 23838
rect 26908 23828 26964 24558
rect 26796 23826 26964 23828
rect 26796 23774 26798 23826
rect 26850 23774 26964 23826
rect 26796 23772 26964 23774
rect 26684 23714 26740 23726
rect 26684 23662 26686 23714
rect 26738 23662 26740 23714
rect 26684 23156 26740 23662
rect 26796 23604 26852 23772
rect 26796 23538 26852 23548
rect 26684 23090 26740 23100
rect 26796 23380 26852 23390
rect 26572 20066 26628 20076
rect 26460 19180 26628 19236
rect 26460 19012 26516 19022
rect 26404 19010 26516 19012
rect 26404 18958 26462 19010
rect 26514 18958 26516 19010
rect 26404 18956 26516 18958
rect 26348 18918 26404 18956
rect 26460 18946 26516 18956
rect 26124 18788 26180 18798
rect 26124 18674 26180 18732
rect 26124 18622 26126 18674
rect 26178 18622 26180 18674
rect 26124 18610 26180 18622
rect 26348 18676 26404 18686
rect 26348 18582 26404 18620
rect 26236 18452 26292 18462
rect 26236 18358 26292 18396
rect 26012 17154 26068 17164
rect 26572 17666 26628 19180
rect 26572 17614 26574 17666
rect 26626 17614 26628 17666
rect 26348 16996 26404 17006
rect 26348 16902 26404 16940
rect 26572 16884 26628 17614
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 25788 15148 25844 15262
rect 26348 15316 26404 15326
rect 26348 15202 26404 15260
rect 26348 15150 26350 15202
rect 26402 15150 26404 15202
rect 25788 15092 26292 15148
rect 25676 14756 25732 14766
rect 25676 14642 25732 14700
rect 25676 14590 25678 14642
rect 25730 14590 25732 14642
rect 25676 14578 25732 14590
rect 25452 13970 25620 13972
rect 25452 13918 25454 13970
rect 25506 13918 25620 13970
rect 25452 13916 25620 13918
rect 26124 14306 26180 14318
rect 26124 14254 26126 14306
rect 26178 14254 26180 14306
rect 25452 13906 25508 13916
rect 25788 13636 25844 13646
rect 25788 13542 25844 13580
rect 25026 13356 25290 13366
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25026 13290 25290 13300
rect 26124 12964 26180 14254
rect 26236 13634 26292 15092
rect 26236 13582 26238 13634
rect 26290 13582 26292 13634
rect 26236 13300 26292 13582
rect 26236 13234 26292 13244
rect 26236 13076 26292 13086
rect 26348 13076 26404 15150
rect 26572 15148 26628 16828
rect 26460 15092 26628 15148
rect 26796 18450 26852 23324
rect 26908 22482 26964 23772
rect 26908 22430 26910 22482
rect 26962 22430 26964 22482
rect 26908 21364 26964 22430
rect 27020 22260 27076 24780
rect 27244 24500 27300 27020
rect 27356 26516 27412 26526
rect 27356 26422 27412 26460
rect 27468 25172 27524 27916
rect 27804 27878 27860 27916
rect 28140 27074 28196 28366
rect 28428 28252 28692 28262
rect 28484 28196 28532 28252
rect 28588 28196 28636 28252
rect 28428 28186 28692 28196
rect 28140 27022 28142 27074
rect 28194 27022 28196 27074
rect 28140 26516 28196 27022
rect 28428 26684 28692 26694
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28428 26618 28692 26628
rect 28140 26178 28196 26460
rect 28140 26126 28142 26178
rect 28194 26126 28196 26178
rect 27804 25506 27860 25518
rect 27804 25454 27806 25506
rect 27858 25454 27860 25506
rect 27468 25116 27748 25172
rect 27356 24724 27412 24734
rect 27356 24610 27412 24668
rect 27356 24558 27358 24610
rect 27410 24558 27412 24610
rect 27356 24500 27412 24558
rect 27356 24444 27636 24500
rect 27244 24050 27300 24444
rect 27244 23998 27246 24050
rect 27298 23998 27300 24050
rect 27244 23986 27300 23998
rect 27356 23156 27412 23166
rect 27356 23062 27412 23100
rect 27020 21476 27076 22204
rect 27020 21474 27524 21476
rect 27020 21422 27022 21474
rect 27074 21422 27524 21474
rect 27020 21420 27524 21422
rect 27020 21410 27076 21420
rect 26908 21298 26964 21308
rect 27132 21028 27188 21038
rect 27132 20934 27188 20972
rect 27132 20804 27188 20814
rect 27132 20710 27188 20748
rect 27244 20188 27300 21420
rect 27468 21026 27524 21420
rect 27468 20974 27470 21026
rect 27522 20974 27524 21026
rect 27468 20962 27524 20974
rect 27020 20132 27076 20142
rect 27020 19346 27076 20076
rect 27020 19294 27022 19346
rect 27074 19294 27076 19346
rect 27020 19282 27076 19294
rect 27132 20132 27300 20188
rect 27468 20692 27524 20702
rect 27020 18788 27076 18798
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 15540 26852 18398
rect 26460 13636 26516 15092
rect 26796 14980 26852 15484
rect 26908 18732 27020 18788
rect 26908 15092 26964 18732
rect 27020 18722 27076 18732
rect 27132 18338 27188 20132
rect 27132 18286 27134 18338
rect 27186 18286 27188 18338
rect 27132 18226 27188 18286
rect 27132 18174 27134 18226
rect 27186 18174 27188 18226
rect 27132 18162 27188 18174
rect 27356 19010 27412 19022
rect 27356 18958 27358 19010
rect 27410 18958 27412 19010
rect 27020 17220 27076 17230
rect 27356 17220 27412 18958
rect 27468 17780 27524 20636
rect 27580 20580 27636 24444
rect 27692 24050 27748 25116
rect 27804 24612 27860 25454
rect 28140 24612 28196 26126
rect 28428 25116 28692 25126
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28428 25050 28692 25060
rect 27804 24610 28196 24612
rect 27804 24558 28142 24610
rect 28194 24558 28196 24610
rect 27804 24556 28196 24558
rect 27692 23998 27694 24050
rect 27746 23998 27748 24050
rect 27692 23716 27748 23998
rect 27692 23650 27748 23660
rect 28140 23714 28196 24556
rect 28140 23662 28142 23714
rect 28194 23662 28196 23714
rect 28028 23156 28084 23166
rect 28140 23156 28196 23662
rect 28428 23548 28692 23558
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28428 23482 28692 23492
rect 28028 23154 28196 23156
rect 28028 23102 28030 23154
rect 28082 23102 28196 23154
rect 28028 23100 28196 23102
rect 28028 23044 28084 23100
rect 27916 20580 27972 20590
rect 27580 20578 27972 20580
rect 27580 20526 27918 20578
rect 27970 20526 27972 20578
rect 27580 20524 27972 20526
rect 27804 18788 27860 20524
rect 27916 20514 27972 20524
rect 27804 18722 27860 18732
rect 27916 20356 27972 20366
rect 27580 18564 27636 18574
rect 27580 18340 27636 18508
rect 27916 18452 27972 20300
rect 28028 20020 28084 22988
rect 28428 21980 28692 21990
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28428 21914 28692 21924
rect 28028 19348 28084 19964
rect 28140 20804 28196 20814
rect 28140 19906 28196 20748
rect 28428 20412 28692 20422
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28428 20346 28692 20356
rect 28140 19854 28142 19906
rect 28194 19854 28196 19906
rect 28140 19842 28196 19854
rect 28028 19346 28196 19348
rect 28028 19294 28030 19346
rect 28082 19294 28196 19346
rect 28028 19292 28196 19294
rect 28028 19282 28084 19292
rect 28028 18452 28084 18462
rect 27916 18450 28084 18452
rect 27916 18398 28030 18450
rect 28082 18398 28084 18450
rect 27916 18396 28084 18398
rect 28028 18386 28084 18396
rect 27580 18338 27748 18340
rect 27580 18286 27582 18338
rect 27634 18286 27748 18338
rect 27580 18284 27748 18286
rect 27580 18274 27636 18284
rect 27580 17780 27636 17790
rect 27468 17778 27636 17780
rect 27468 17726 27582 17778
rect 27634 17726 27636 17778
rect 27468 17724 27636 17726
rect 27580 17714 27636 17724
rect 27076 17164 27412 17220
rect 27020 16210 27076 17164
rect 27580 16884 27636 16894
rect 27580 16790 27636 16828
rect 27020 16158 27022 16210
rect 27074 16158 27076 16210
rect 27020 16146 27076 16158
rect 27580 16212 27636 16222
rect 27692 16212 27748 18284
rect 27580 16210 27748 16212
rect 27580 16158 27582 16210
rect 27634 16158 27748 16210
rect 27580 16156 27748 16158
rect 27804 18226 27860 18238
rect 27804 18174 27806 18226
rect 27858 18174 27860 18226
rect 27580 16146 27636 16156
rect 26908 15036 27188 15092
rect 26684 14924 27076 14980
rect 26460 13570 26516 13580
rect 26572 14306 26628 14318
rect 26572 14254 26574 14306
rect 26626 14254 26628 14306
rect 26236 13074 26404 13076
rect 26236 13022 26238 13074
rect 26290 13022 26404 13074
rect 26236 13020 26404 13022
rect 26460 13188 26516 13198
rect 26236 13010 26292 13020
rect 26124 12898 26180 12908
rect 25228 12180 25284 12190
rect 25228 12086 25284 12124
rect 26460 12180 26516 13132
rect 26572 12964 26628 14254
rect 26684 13970 26740 14924
rect 27020 14642 27076 14924
rect 27020 14590 27022 14642
rect 27074 14590 27076 14642
rect 27020 14578 27076 14590
rect 26684 13918 26686 13970
rect 26738 13918 26740 13970
rect 26684 13906 26740 13918
rect 27132 13970 27188 15036
rect 27804 14642 27860 18174
rect 28028 17444 28084 17454
rect 28028 17350 28084 17388
rect 27804 14590 27806 14642
rect 27858 14590 27860 14642
rect 27804 14578 27860 14590
rect 28140 16210 28196 19292
rect 28428 18844 28692 18854
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28428 18778 28692 18788
rect 28428 17276 28692 17286
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28428 17210 28692 17220
rect 28140 16158 28142 16210
rect 28194 16158 28196 16210
rect 28140 14642 28196 16158
rect 28428 15708 28692 15718
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28428 15642 28692 15652
rect 28140 14590 28142 14642
rect 28194 14590 28196 14642
rect 28140 14578 28196 14590
rect 28428 14140 28692 14150
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28428 14074 28692 14084
rect 27132 13918 27134 13970
rect 27186 13918 27188 13970
rect 27132 13860 27188 13918
rect 27020 13186 27076 13198
rect 27020 13134 27022 13186
rect 27074 13134 27076 13186
rect 27020 13074 27076 13134
rect 27020 13022 27022 13074
rect 27074 13022 27076 13074
rect 27020 13010 27076 13022
rect 26572 12870 26628 12908
rect 26460 12114 26516 12124
rect 27132 12066 27188 13804
rect 28428 12572 28692 12582
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28428 12506 28692 12516
rect 27132 12014 27134 12066
rect 27186 12014 27188 12066
rect 27132 12002 27188 12014
rect 25026 11788 25290 11798
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25026 11722 25290 11732
rect 24668 11394 24836 11396
rect 24668 11342 24670 11394
rect 24722 11342 24836 11394
rect 24668 11340 24836 11342
rect 25788 11506 25844 11518
rect 25788 11454 25790 11506
rect 25842 11454 25844 11506
rect 24556 10500 24612 10510
rect 24668 10500 24724 11340
rect 25788 10836 25844 11454
rect 28428 11004 28692 11014
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28428 10938 28692 10948
rect 25788 10770 25844 10780
rect 24556 10498 24724 10500
rect 24556 10446 24558 10498
rect 24610 10446 24724 10498
rect 24556 10444 24724 10446
rect 25564 10610 25620 10622
rect 25564 10558 25566 10610
rect 25618 10558 25620 10610
rect 24556 9828 24612 10444
rect 25026 10220 25290 10230
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25026 10154 25290 10164
rect 24892 9828 24948 9838
rect 24556 9772 24892 9828
rect 24444 7982 24446 8034
rect 24498 7982 24500 8034
rect 24444 7970 24500 7982
rect 24556 8258 24612 8270
rect 24556 8206 24558 8258
rect 24610 8206 24612 8258
rect 24444 6692 24500 6702
rect 23884 6578 24164 6580
rect 23884 6526 23886 6578
rect 23938 6526 24164 6578
rect 23884 6524 24164 6526
rect 23884 6514 23940 6524
rect 22988 6076 23268 6132
rect 23660 6076 24052 6132
rect 22540 6020 22596 6030
rect 22540 5926 22596 5964
rect 22988 5906 23044 6076
rect 22988 5854 22990 5906
rect 23042 5854 23044 5906
rect 22988 5842 23044 5854
rect 23100 5906 23156 5918
rect 23100 5854 23102 5906
rect 23154 5854 23156 5906
rect 21532 5124 21588 5134
rect 21532 5030 21588 5068
rect 21980 5012 22036 5022
rect 21308 4900 21364 4910
rect 21084 4898 21364 4900
rect 21084 4846 21310 4898
rect 21362 4846 21364 4898
rect 21084 4844 21364 4846
rect 20860 2606 20862 2658
rect 20914 2606 20916 2658
rect 20860 2594 20916 2606
rect 20972 3444 21028 3454
rect 20748 2098 20804 2156
rect 20748 2046 20750 2098
rect 20802 2046 20804 2098
rect 20748 2034 20804 2046
rect 20972 2098 21028 3388
rect 20972 2046 20974 2098
rect 21026 2046 21028 2098
rect 20972 2034 21028 2046
rect 21084 1986 21140 4844
rect 21308 4834 21364 4844
rect 21624 4732 21888 4742
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21624 4666 21888 4676
rect 21980 4564 22036 4956
rect 21868 4508 22036 4564
rect 21532 4340 21588 4350
rect 21420 4338 21588 4340
rect 21420 4286 21534 4338
rect 21586 4286 21588 4338
rect 21420 4284 21588 4286
rect 21420 3666 21476 4284
rect 21532 4274 21588 4284
rect 21420 3614 21422 3666
rect 21474 3614 21476 3666
rect 21308 3332 21364 3342
rect 21196 3330 21364 3332
rect 21196 3278 21310 3330
rect 21362 3278 21364 3330
rect 21196 3276 21364 3278
rect 21196 2770 21252 3276
rect 21308 3266 21364 3276
rect 21420 3332 21476 3614
rect 21868 4226 21924 4508
rect 21868 4174 21870 4226
rect 21922 4174 21924 4226
rect 21868 3332 21924 4174
rect 22204 3778 22260 5628
rect 22428 4562 22484 5740
rect 22540 5236 22596 5246
rect 22540 5142 22596 5180
rect 22428 4510 22430 4562
rect 22482 4510 22484 4562
rect 22428 4498 22484 4510
rect 22988 5124 23044 5134
rect 23100 5124 23156 5854
rect 22988 5122 23156 5124
rect 22988 5070 22990 5122
rect 23042 5070 23156 5122
rect 22988 5068 23156 5070
rect 22988 4450 23044 5068
rect 22988 4398 22990 4450
rect 23042 4398 23044 4450
rect 22988 4386 23044 4398
rect 23212 5010 23268 6076
rect 23436 6020 23492 6030
rect 23436 5906 23492 5964
rect 23436 5854 23438 5906
rect 23490 5854 23492 5906
rect 23436 5842 23492 5854
rect 23660 5908 23716 5918
rect 23716 5852 23828 5908
rect 23660 5814 23716 5852
rect 23212 4958 23214 5010
rect 23266 4958 23268 5010
rect 23212 4452 23268 4958
rect 23772 5012 23828 5852
rect 23884 5906 23940 5918
rect 23884 5854 23886 5906
rect 23938 5854 23940 5906
rect 23884 5684 23940 5854
rect 23884 5618 23940 5628
rect 23996 5572 24052 6076
rect 24108 5794 24164 6524
rect 24444 6132 24500 6636
rect 24444 6066 24500 6076
rect 24220 6020 24276 6030
rect 24556 6020 24612 8206
rect 24780 8258 24836 8270
rect 24780 8206 24782 8258
rect 24834 8206 24836 8258
rect 24780 7476 24836 8206
rect 24668 6804 24724 6814
rect 24780 6804 24836 7420
rect 24668 6802 24836 6804
rect 24668 6750 24670 6802
rect 24722 6750 24836 6802
rect 24668 6748 24836 6750
rect 24668 6738 24724 6748
rect 24220 6018 24388 6020
rect 24220 5966 24222 6018
rect 24274 5966 24388 6018
rect 24220 5964 24388 5966
rect 24220 5954 24276 5964
rect 24108 5742 24110 5794
rect 24162 5742 24164 5794
rect 24108 5730 24164 5742
rect 24332 5572 24388 5964
rect 24556 5796 24612 5964
rect 24556 5730 24612 5740
rect 24780 6020 24836 6748
rect 24892 6466 24948 9772
rect 25564 9828 25620 10558
rect 26348 10500 26404 10510
rect 26348 10406 26404 10444
rect 25564 9734 25620 9772
rect 26012 9828 26068 9838
rect 26012 9734 26068 9772
rect 28428 9436 28692 9446
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28428 9370 28692 9380
rect 25026 8652 25290 8662
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25026 8586 25290 8596
rect 28428 7868 28692 7878
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28428 7802 28692 7812
rect 25026 7084 25290 7094
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25026 7018 25290 7028
rect 24892 6414 24894 6466
rect 24946 6414 24948 6466
rect 24892 6402 24948 6414
rect 28428 6300 28692 6310
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28428 6234 28692 6244
rect 23996 5516 24388 5572
rect 23884 5012 23940 5022
rect 23772 5010 23940 5012
rect 23772 4958 23886 5010
rect 23938 4958 23940 5010
rect 23772 4956 23940 4958
rect 23884 4946 23940 4956
rect 23212 4386 23268 4396
rect 23996 4900 24052 4910
rect 23436 4338 23492 4350
rect 23436 4286 23438 4338
rect 23490 4286 23492 4338
rect 23212 4228 23268 4238
rect 23212 4134 23268 4172
rect 22204 3726 22206 3778
rect 22258 3726 22260 3778
rect 22204 3714 22260 3726
rect 22316 3780 22372 3790
rect 21980 3668 22036 3678
rect 21980 3574 22036 3612
rect 22316 3554 22372 3724
rect 22764 3780 22820 3790
rect 22316 3502 22318 3554
rect 22370 3502 22372 3554
rect 22316 3490 22372 3502
rect 22652 3554 22708 3566
rect 22652 3502 22654 3554
rect 22706 3502 22708 3554
rect 21868 3276 22036 3332
rect 21196 2718 21198 2770
rect 21250 2718 21252 2770
rect 21196 2706 21252 2718
rect 21420 2212 21476 3276
rect 21624 3164 21888 3174
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21624 3098 21888 3108
rect 21644 2884 21700 2894
rect 21980 2884 22036 3276
rect 22652 2996 22708 3502
rect 22652 2930 22708 2940
rect 21644 2882 22036 2884
rect 21644 2830 21646 2882
rect 21698 2830 22036 2882
rect 21644 2828 22036 2830
rect 21644 2818 21700 2828
rect 21420 2146 21476 2156
rect 21868 2098 21924 2828
rect 21868 2046 21870 2098
rect 21922 2046 21924 2098
rect 21868 2034 21924 2046
rect 22428 2660 22484 2670
rect 21532 1988 21588 1998
rect 21084 1934 21086 1986
rect 21138 1934 21140 1986
rect 21084 1922 21140 1934
rect 21420 1932 21532 1988
rect 20636 1820 20916 1876
rect 20188 1708 20468 1764
rect 20188 400 20244 1708
rect 20860 400 20916 1820
rect 21420 1428 21476 1932
rect 21532 1922 21588 1932
rect 22428 1988 22484 2604
rect 22428 1894 22484 1932
rect 21624 1596 21888 1606
rect 21680 1540 21728 1596
rect 21784 1540 21832 1596
rect 21624 1530 21888 1540
rect 21420 1372 21588 1428
rect 21532 400 21588 1372
rect 22764 644 22820 3724
rect 23212 3668 23268 3678
rect 22876 2772 22932 2782
rect 22988 2772 23044 2782
rect 22932 2770 23044 2772
rect 22932 2718 22990 2770
rect 23042 2718 23044 2770
rect 22932 2716 23044 2718
rect 22876 2098 22932 2716
rect 22988 2706 23044 2716
rect 22876 2046 22878 2098
rect 22930 2046 22932 2098
rect 22876 2034 22932 2046
rect 23212 1986 23268 3612
rect 23324 3444 23380 3482
rect 23324 3378 23380 3388
rect 23436 2996 23492 4286
rect 23660 4116 23716 4126
rect 23660 3892 23716 4060
rect 23660 3554 23716 3836
rect 23660 3502 23662 3554
rect 23714 3502 23716 3554
rect 23660 3490 23716 3502
rect 23996 4004 24052 4844
rect 24220 4340 24276 4350
rect 24220 4246 24276 4284
rect 23436 2930 23492 2940
rect 23772 3332 23828 3342
rect 23660 2884 23716 2894
rect 23212 1934 23214 1986
rect 23266 1934 23268 1986
rect 22764 588 22932 644
rect 22428 532 22484 542
rect 22204 476 22428 532
rect 22204 400 22260 476
rect 22428 466 22484 476
rect 22876 400 22932 588
rect 23212 532 23268 1934
rect 23212 466 23268 476
rect 23548 1988 23604 1998
rect 23548 400 23604 1932
rect 23660 1874 23716 2828
rect 23772 2658 23828 3276
rect 23772 2606 23774 2658
rect 23826 2606 23828 2658
rect 23772 2594 23828 2606
rect 23996 1986 24052 3948
rect 24108 4226 24164 4238
rect 24108 4174 24110 4226
rect 24162 4174 24164 4226
rect 24108 3780 24164 4174
rect 24108 3724 24276 3780
rect 24108 3556 24164 3566
rect 24108 3462 24164 3500
rect 24108 2772 24164 2782
rect 24220 2772 24276 3724
rect 24332 2994 24388 5516
rect 24668 4226 24724 4238
rect 24668 4174 24670 4226
rect 24722 4174 24724 4226
rect 24556 4114 24612 4126
rect 24556 4062 24558 4114
rect 24610 4062 24612 4114
rect 24556 3554 24612 4062
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24332 2942 24334 2994
rect 24386 2942 24388 2994
rect 24332 2930 24388 2942
rect 24668 2884 24724 4174
rect 24668 2818 24724 2828
rect 24332 2772 24388 2782
rect 24220 2770 24388 2772
rect 24220 2718 24334 2770
rect 24386 2718 24388 2770
rect 24220 2716 24388 2718
rect 24108 2678 24164 2716
rect 23996 1934 23998 1986
rect 24050 1934 24052 1986
rect 23996 1922 24052 1934
rect 24220 2100 24276 2110
rect 23660 1822 23662 1874
rect 23714 1822 23716 1874
rect 23660 1810 23716 1822
rect 24220 400 24276 2044
rect 24332 1876 24388 2716
rect 24668 2100 24724 2110
rect 24780 2100 24836 5964
rect 25452 6132 25508 6142
rect 25026 5516 25290 5526
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25026 5450 25290 5460
rect 25452 5122 25508 6076
rect 26012 6020 26068 6030
rect 26012 5926 26068 5964
rect 25900 5908 25956 5918
rect 25900 5814 25956 5852
rect 25452 5070 25454 5122
rect 25506 5070 25508 5122
rect 25452 5058 25508 5070
rect 25564 5796 25620 5806
rect 25228 4452 25284 4462
rect 25228 4358 25284 4396
rect 25340 4340 25396 4350
rect 25340 4246 25396 4284
rect 24668 2098 24836 2100
rect 24668 2046 24670 2098
rect 24722 2046 24836 2098
rect 24668 2044 24836 2046
rect 24892 4228 24948 4238
rect 24892 3780 24948 4172
rect 25026 3948 25290 3958
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25026 3882 25290 3892
rect 24668 2034 24724 2044
rect 24892 1988 24948 3724
rect 25564 3388 25620 5740
rect 25228 3332 25620 3388
rect 25676 5348 25732 5358
rect 25676 3442 25732 5292
rect 26908 5122 26964 5134
rect 26908 5070 26910 5122
rect 26962 5070 26964 5122
rect 26012 4900 26068 4910
rect 26460 4900 26516 4910
rect 26012 4806 26068 4844
rect 26124 4898 26516 4900
rect 26124 4846 26462 4898
rect 26514 4846 26516 4898
rect 26124 4844 26516 4846
rect 25788 4340 25844 4350
rect 25788 4338 25956 4340
rect 25788 4286 25790 4338
rect 25842 4286 25956 4338
rect 25788 4284 25956 4286
rect 25788 4274 25844 4284
rect 25676 3390 25678 3442
rect 25730 3390 25732 3442
rect 25228 2548 25284 3332
rect 25340 2996 25396 3034
rect 25340 2930 25396 2940
rect 25676 2996 25732 3390
rect 25452 2884 25508 2894
rect 25452 2790 25508 2828
rect 25340 2770 25396 2782
rect 25340 2718 25342 2770
rect 25394 2718 25396 2770
rect 25340 2660 25396 2718
rect 25676 2660 25732 2940
rect 25340 2604 25732 2660
rect 25788 3556 25844 3566
rect 25788 2548 25844 3500
rect 25900 2772 25956 4284
rect 26124 4004 26180 4844
rect 26460 4834 26516 4844
rect 26908 4452 26964 5070
rect 27356 5124 27412 5134
rect 27804 5124 27860 5134
rect 27356 5122 27636 5124
rect 27356 5070 27358 5122
rect 27410 5070 27636 5122
rect 27356 5068 27636 5070
rect 27356 5058 27412 5068
rect 26908 4396 27300 4452
rect 26460 4226 26516 4238
rect 26460 4174 26462 4226
rect 26514 4174 26516 4226
rect 26460 4116 26516 4174
rect 26908 4228 26964 4238
rect 26908 4134 26964 4172
rect 26460 4050 26516 4060
rect 27020 4114 27076 4126
rect 27020 4062 27022 4114
rect 27074 4062 27076 4114
rect 25900 2706 25956 2716
rect 26012 3948 26180 4004
rect 25228 2492 25508 2548
rect 25026 2380 25290 2390
rect 25082 2324 25130 2380
rect 25186 2324 25234 2380
rect 25026 2314 25290 2324
rect 25452 2098 25508 2492
rect 25452 2046 25454 2098
rect 25506 2046 25508 2098
rect 25452 2034 25508 2046
rect 25564 2492 25844 2548
rect 25004 1988 25060 1998
rect 24892 1986 25060 1988
rect 24892 1934 25006 1986
rect 25058 1934 25060 1986
rect 24892 1932 25060 1934
rect 25004 1922 25060 1932
rect 24332 1810 24388 1820
rect 24892 1764 24948 1774
rect 24892 400 24948 1708
rect 25564 400 25620 2492
rect 25676 1988 25732 1998
rect 25900 1988 25956 1998
rect 26012 1988 26068 3948
rect 26124 3554 26180 3566
rect 26124 3502 26126 3554
rect 26178 3502 26180 3554
rect 26124 3444 26180 3502
rect 26124 2882 26180 3388
rect 26236 2996 26292 3006
rect 27020 2996 27076 4062
rect 27132 3444 27188 3454
rect 27132 3350 27188 3388
rect 26292 2940 26516 2996
rect 26236 2930 26292 2940
rect 26124 2830 26126 2882
rect 26178 2830 26180 2882
rect 26124 2818 26180 2830
rect 26460 2098 26516 2940
rect 26908 2940 27076 2996
rect 26684 2882 26740 2894
rect 26684 2830 26686 2882
rect 26738 2830 26740 2882
rect 26684 2772 26740 2830
rect 26684 2706 26740 2716
rect 26460 2046 26462 2098
rect 26514 2046 26516 2098
rect 26460 2034 26516 2046
rect 26908 1988 26964 2940
rect 25732 1986 26068 1988
rect 25732 1934 25902 1986
rect 25954 1934 26068 1986
rect 25732 1932 26068 1934
rect 26572 1986 26964 1988
rect 26572 1934 26910 1986
rect 26962 1934 26964 1986
rect 26572 1932 26964 1934
rect 25676 1922 25732 1932
rect 25900 1922 25956 1932
rect 26572 1876 26628 1932
rect 26908 1922 26964 1932
rect 27020 2772 27076 2782
rect 27244 2772 27300 4396
rect 27356 4226 27412 4238
rect 27356 4174 27358 4226
rect 27410 4174 27412 4226
rect 27356 3444 27412 4174
rect 27580 3556 27636 5068
rect 27468 3444 27524 3454
rect 27356 3442 27524 3444
rect 27356 3390 27470 3442
rect 27522 3390 27524 3442
rect 27356 3388 27524 3390
rect 27356 2884 27412 2894
rect 27356 2790 27412 2828
rect 27020 2770 27300 2772
rect 27020 2718 27022 2770
rect 27074 2718 27300 2770
rect 27020 2716 27300 2718
rect 26236 1820 26628 1876
rect 26236 400 26292 1820
rect 26908 1764 26964 1774
rect 27020 1764 27076 2716
rect 27356 1876 27412 1886
rect 27356 1782 27412 1820
rect 26964 1708 27076 1764
rect 26908 1698 26964 1708
rect 27468 1540 27524 3388
rect 27580 2770 27636 3500
rect 27580 2718 27582 2770
rect 27634 2718 27636 2770
rect 27580 2706 27636 2718
rect 27692 5122 27860 5124
rect 27692 5070 27806 5122
rect 27858 5070 27860 5122
rect 27692 5068 27860 5070
rect 27580 2100 27636 2110
rect 27692 2100 27748 5068
rect 27804 5058 27860 5068
rect 28428 4732 28692 4742
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28428 4666 28692 4676
rect 27804 4226 27860 4238
rect 27804 4174 27806 4226
rect 27858 4174 27860 4226
rect 27804 4114 27860 4174
rect 27804 4062 27806 4114
rect 27858 4062 27860 4114
rect 27804 4050 27860 4062
rect 27916 3668 27972 3678
rect 27916 3574 27972 3612
rect 28428 3164 28692 3174
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28428 3098 28692 3108
rect 28140 2660 28196 2670
rect 28140 2566 28196 2604
rect 27636 2044 27748 2100
rect 27580 1986 27636 2044
rect 27580 1934 27582 1986
rect 27634 1934 27636 1986
rect 27580 1922 27636 1934
rect 26908 1484 27524 1540
rect 28428 1596 28692 1606
rect 28484 1540 28532 1596
rect 28588 1540 28636 1596
rect 28428 1530 28692 1540
rect 26908 400 26964 1484
rect 2688 0 2800 400
rect 3360 0 3472 400
rect 4032 0 4144 400
rect 4704 0 4816 400
rect 5376 0 5488 400
rect 6048 0 6160 400
rect 6720 0 6832 400
rect 7392 0 7504 400
rect 8064 0 8176 400
rect 8736 0 8848 400
rect 9408 0 9520 400
rect 10080 0 10192 400
rect 10752 0 10864 400
rect 11424 0 11536 400
rect 12096 0 12208 400
rect 12768 0 12880 400
rect 13440 0 13552 400
rect 14112 0 14224 400
rect 14784 0 14896 400
rect 15456 0 15568 400
rect 16128 0 16240 400
rect 16800 0 16912 400
rect 17472 0 17584 400
rect 18144 0 18256 400
rect 18816 0 18928 400
rect 19488 0 19600 400
rect 20160 0 20272 400
rect 20832 0 20944 400
rect 21504 0 21616 400
rect 22176 0 22288 400
rect 22848 0 22960 400
rect 23520 0 23632 400
rect 24192 0 24304 400
rect 24864 0 24976 400
rect 25536 0 25648 400
rect 26208 0 26320 400
rect 26880 0 26992 400
<< via2 >>
rect 4614 118410 4670 118412
rect 4614 118358 4616 118410
rect 4616 118358 4668 118410
rect 4668 118358 4670 118410
rect 4614 118356 4670 118358
rect 4718 118410 4774 118412
rect 4718 118358 4720 118410
rect 4720 118358 4772 118410
rect 4772 118358 4774 118410
rect 4718 118356 4774 118358
rect 4822 118410 4878 118412
rect 4822 118358 4824 118410
rect 4824 118358 4876 118410
rect 4876 118358 4878 118410
rect 4822 118356 4878 118358
rect 11418 118410 11474 118412
rect 11418 118358 11420 118410
rect 11420 118358 11472 118410
rect 11472 118358 11474 118410
rect 11418 118356 11474 118358
rect 11522 118410 11578 118412
rect 11522 118358 11524 118410
rect 11524 118358 11576 118410
rect 11576 118358 11578 118410
rect 11522 118356 11578 118358
rect 11626 118410 11682 118412
rect 11626 118358 11628 118410
rect 11628 118358 11680 118410
rect 11680 118358 11682 118410
rect 11626 118356 11682 118358
rect 8016 117626 8072 117628
rect 8016 117574 8018 117626
rect 8018 117574 8070 117626
rect 8070 117574 8072 117626
rect 8016 117572 8072 117574
rect 8120 117626 8176 117628
rect 8120 117574 8122 117626
rect 8122 117574 8174 117626
rect 8174 117574 8176 117626
rect 8120 117572 8176 117574
rect 8224 117626 8280 117628
rect 8224 117574 8226 117626
rect 8226 117574 8278 117626
rect 8278 117574 8280 117626
rect 8224 117572 8280 117574
rect 4614 116842 4670 116844
rect 4614 116790 4616 116842
rect 4616 116790 4668 116842
rect 4668 116790 4670 116842
rect 4614 116788 4670 116790
rect 4718 116842 4774 116844
rect 4718 116790 4720 116842
rect 4720 116790 4772 116842
rect 4772 116790 4774 116842
rect 4718 116788 4774 116790
rect 4822 116842 4878 116844
rect 4822 116790 4824 116842
rect 4824 116790 4876 116842
rect 4876 116790 4878 116842
rect 4822 116788 4878 116790
rect 11418 116842 11474 116844
rect 11418 116790 11420 116842
rect 11420 116790 11472 116842
rect 11472 116790 11474 116842
rect 11418 116788 11474 116790
rect 11522 116842 11578 116844
rect 11522 116790 11524 116842
rect 11524 116790 11576 116842
rect 11576 116790 11578 116842
rect 11522 116788 11578 116790
rect 11626 116842 11682 116844
rect 11626 116790 11628 116842
rect 11628 116790 11680 116842
rect 11680 116790 11682 116842
rect 11626 116788 11682 116790
rect 8016 116058 8072 116060
rect 8016 116006 8018 116058
rect 8018 116006 8070 116058
rect 8070 116006 8072 116058
rect 8016 116004 8072 116006
rect 8120 116058 8176 116060
rect 8120 116006 8122 116058
rect 8122 116006 8174 116058
rect 8174 116006 8176 116058
rect 8120 116004 8176 116006
rect 8224 116058 8280 116060
rect 8224 116006 8226 116058
rect 8226 116006 8278 116058
rect 8278 116006 8280 116058
rect 8224 116004 8280 116006
rect 10780 115612 10836 115668
rect 12236 115666 12292 115668
rect 12236 115614 12238 115666
rect 12238 115614 12290 115666
rect 12290 115614 12292 115666
rect 12236 115612 12292 115614
rect 4614 115274 4670 115276
rect 4614 115222 4616 115274
rect 4616 115222 4668 115274
rect 4668 115222 4670 115274
rect 4614 115220 4670 115222
rect 4718 115274 4774 115276
rect 4718 115222 4720 115274
rect 4720 115222 4772 115274
rect 4772 115222 4774 115274
rect 4718 115220 4774 115222
rect 4822 115274 4878 115276
rect 4822 115222 4824 115274
rect 4824 115222 4876 115274
rect 4876 115222 4878 115274
rect 4822 115220 4878 115222
rect 1708 114940 1764 114996
rect 8016 114490 8072 114492
rect 8016 114438 8018 114490
rect 8018 114438 8070 114490
rect 8070 114438 8072 114490
rect 8016 114436 8072 114438
rect 8120 114490 8176 114492
rect 8120 114438 8122 114490
rect 8122 114438 8174 114490
rect 8174 114438 8176 114490
rect 8120 114436 8176 114438
rect 8224 114490 8280 114492
rect 8224 114438 8226 114490
rect 8226 114438 8278 114490
rect 8278 114438 8280 114490
rect 8224 114436 8280 114438
rect 13356 115612 13412 115668
rect 11418 115274 11474 115276
rect 11418 115222 11420 115274
rect 11420 115222 11472 115274
rect 11472 115222 11474 115274
rect 11418 115220 11474 115222
rect 11522 115274 11578 115276
rect 11522 115222 11524 115274
rect 11524 115222 11576 115274
rect 11576 115222 11578 115274
rect 11522 115220 11578 115222
rect 11626 115274 11682 115276
rect 11626 115222 11628 115274
rect 11628 115222 11680 115274
rect 11680 115222 11682 115274
rect 11626 115220 11682 115222
rect 10108 114156 10164 114212
rect 11116 114156 11172 114212
rect 4614 113706 4670 113708
rect 4614 113654 4616 113706
rect 4616 113654 4668 113706
rect 4668 113654 4670 113706
rect 4614 113652 4670 113654
rect 4718 113706 4774 113708
rect 4718 113654 4720 113706
rect 4720 113654 4772 113706
rect 4772 113654 4774 113706
rect 4718 113652 4774 113654
rect 4822 113706 4878 113708
rect 4822 113654 4824 113706
rect 4824 113654 4876 113706
rect 4876 113654 4878 113706
rect 4822 113652 4878 113654
rect 7980 113148 8036 113204
rect 8016 112922 8072 112924
rect 8016 112870 8018 112922
rect 8018 112870 8070 112922
rect 8070 112870 8072 112922
rect 8016 112868 8072 112870
rect 8120 112922 8176 112924
rect 8120 112870 8122 112922
rect 8122 112870 8174 112922
rect 8174 112870 8176 112922
rect 8120 112868 8176 112870
rect 8224 112922 8280 112924
rect 8224 112870 8226 112922
rect 8226 112870 8278 112922
rect 8278 112870 8280 112922
rect 8224 112868 8280 112870
rect 8428 112588 8484 112644
rect 8876 112588 8932 112644
rect 9212 113148 9268 113204
rect 3948 112252 4004 112308
rect 1708 109564 1764 109620
rect 4614 112138 4670 112140
rect 4614 112086 4616 112138
rect 4616 112086 4668 112138
rect 4668 112086 4670 112138
rect 4614 112084 4670 112086
rect 4718 112138 4774 112140
rect 4718 112086 4720 112138
rect 4720 112086 4772 112138
rect 4772 112086 4774 112138
rect 4718 112084 4774 112086
rect 4822 112138 4878 112140
rect 4822 112086 4824 112138
rect 4824 112086 4876 112138
rect 4876 112086 4878 112138
rect 4822 112084 4878 112086
rect 10556 114044 10612 114100
rect 10556 113148 10612 113204
rect 12124 114098 12180 114100
rect 12124 114046 12126 114098
rect 12126 114046 12178 114098
rect 12178 114046 12180 114098
rect 12124 114044 12180 114046
rect 12684 114044 12740 114100
rect 11418 113706 11474 113708
rect 11418 113654 11420 113706
rect 11420 113654 11472 113706
rect 11472 113654 11474 113706
rect 11418 113652 11474 113654
rect 11522 113706 11578 113708
rect 11522 113654 11524 113706
rect 11524 113654 11576 113706
rect 11576 113654 11578 113706
rect 11522 113652 11578 113654
rect 11626 113706 11682 113708
rect 11626 113654 11628 113706
rect 11628 113654 11680 113706
rect 11680 113654 11682 113706
rect 11626 113652 11682 113654
rect 8016 111354 8072 111356
rect 8016 111302 8018 111354
rect 8018 111302 8070 111354
rect 8070 111302 8072 111354
rect 8016 111300 8072 111302
rect 8120 111354 8176 111356
rect 8120 111302 8122 111354
rect 8122 111302 8174 111354
rect 8174 111302 8176 111354
rect 8120 111300 8176 111302
rect 8224 111354 8280 111356
rect 8224 111302 8226 111354
rect 8226 111302 8278 111354
rect 8278 111302 8280 111354
rect 8224 111300 8280 111302
rect 6860 110908 6916 110964
rect 4614 110570 4670 110572
rect 4614 110518 4616 110570
rect 4616 110518 4668 110570
rect 4668 110518 4670 110570
rect 4614 110516 4670 110518
rect 4718 110570 4774 110572
rect 4718 110518 4720 110570
rect 4720 110518 4772 110570
rect 4772 110518 4774 110570
rect 4718 110516 4774 110518
rect 4822 110570 4878 110572
rect 4822 110518 4824 110570
rect 4824 110518 4876 110570
rect 4876 110518 4878 110570
rect 4822 110516 4878 110518
rect 9548 110684 9604 110740
rect 8988 110124 9044 110180
rect 8016 109786 8072 109788
rect 8016 109734 8018 109786
rect 8018 109734 8070 109786
rect 8070 109734 8072 109786
rect 8016 109732 8072 109734
rect 8120 109786 8176 109788
rect 8120 109734 8122 109786
rect 8122 109734 8174 109786
rect 8174 109734 8176 109786
rect 8120 109732 8176 109734
rect 8224 109786 8280 109788
rect 8224 109734 8226 109786
rect 8226 109734 8278 109786
rect 8278 109734 8280 109786
rect 8224 109732 8280 109734
rect 4614 109002 4670 109004
rect 4614 108950 4616 109002
rect 4616 108950 4668 109002
rect 4668 108950 4670 109002
rect 4614 108948 4670 108950
rect 4718 109002 4774 109004
rect 4718 108950 4720 109002
rect 4720 108950 4772 109002
rect 4772 108950 4774 109002
rect 4718 108948 4774 108950
rect 4822 109002 4878 109004
rect 4822 108950 4824 109002
rect 4824 108950 4876 109002
rect 4876 108950 4878 109002
rect 4822 108948 4878 108950
rect 10220 110684 10276 110740
rect 10332 112588 10388 112644
rect 11228 112588 11284 112644
rect 12124 113036 12180 113092
rect 11452 112530 11508 112532
rect 11452 112478 11454 112530
rect 11454 112478 11506 112530
rect 11506 112478 11508 112530
rect 11452 112476 11508 112478
rect 11418 112138 11474 112140
rect 11418 112086 11420 112138
rect 11420 112086 11472 112138
rect 11472 112086 11474 112138
rect 11418 112084 11474 112086
rect 11522 112138 11578 112140
rect 11522 112086 11524 112138
rect 11524 112086 11576 112138
rect 11576 112086 11578 112138
rect 11522 112084 11578 112086
rect 11626 112138 11682 112140
rect 11626 112086 11628 112138
rect 11628 112086 11680 112138
rect 11680 112086 11682 112138
rect 11626 112084 11682 112086
rect 9660 110178 9716 110180
rect 9660 110126 9662 110178
rect 9662 110126 9714 110178
rect 9714 110126 9716 110178
rect 9660 110124 9716 110126
rect 11004 110684 11060 110740
rect 11676 110738 11732 110740
rect 11676 110686 11678 110738
rect 11678 110686 11730 110738
rect 11730 110686 11732 110738
rect 11676 110684 11732 110686
rect 11788 110796 11844 110852
rect 11418 110570 11474 110572
rect 11418 110518 11420 110570
rect 11420 110518 11472 110570
rect 11472 110518 11474 110570
rect 11418 110516 11474 110518
rect 11522 110570 11578 110572
rect 11522 110518 11524 110570
rect 11524 110518 11576 110570
rect 11576 110518 11578 110570
rect 11522 110516 11578 110518
rect 11626 110570 11682 110572
rect 11626 110518 11628 110570
rect 11628 110518 11680 110570
rect 11680 110518 11682 110570
rect 11626 110516 11682 110518
rect 11452 110290 11508 110292
rect 11452 110238 11454 110290
rect 11454 110238 11506 110290
rect 11506 110238 11508 110290
rect 11452 110236 11508 110238
rect 10332 110124 10388 110180
rect 10780 110124 10836 110180
rect 11676 110178 11732 110180
rect 11676 110126 11678 110178
rect 11678 110126 11730 110178
rect 11730 110126 11732 110178
rect 11676 110124 11732 110126
rect 12796 113090 12852 113092
rect 12796 113038 12798 113090
rect 12798 113038 12850 113090
rect 12850 113038 12852 113090
rect 12796 113036 12852 113038
rect 12684 110796 12740 110852
rect 14820 117626 14876 117628
rect 14820 117574 14822 117626
rect 14822 117574 14874 117626
rect 14874 117574 14876 117626
rect 14820 117572 14876 117574
rect 14924 117626 14980 117628
rect 14924 117574 14926 117626
rect 14926 117574 14978 117626
rect 14978 117574 14980 117626
rect 14924 117572 14980 117574
rect 15028 117626 15084 117628
rect 15028 117574 15030 117626
rect 15030 117574 15082 117626
rect 15082 117574 15084 117626
rect 15028 117572 15084 117574
rect 15148 116396 15204 116452
rect 13916 115612 13972 115668
rect 14820 116058 14876 116060
rect 14820 116006 14822 116058
rect 14822 116006 14874 116058
rect 14874 116006 14876 116058
rect 14820 116004 14876 116006
rect 14924 116058 14980 116060
rect 14924 116006 14926 116058
rect 14926 116006 14978 116058
rect 14978 116006 14980 116058
rect 14924 116004 14980 116006
rect 15028 116058 15084 116060
rect 15028 116006 15030 116058
rect 15030 116006 15082 116058
rect 15082 116006 15084 116058
rect 15028 116004 15084 116006
rect 14820 114490 14876 114492
rect 14820 114438 14822 114490
rect 14822 114438 14874 114490
rect 14874 114438 14876 114490
rect 14820 114436 14876 114438
rect 14924 114490 14980 114492
rect 14924 114438 14926 114490
rect 14926 114438 14978 114490
rect 14978 114438 14980 114490
rect 14924 114436 14980 114438
rect 15028 114490 15084 114492
rect 15028 114438 15030 114490
rect 15030 114438 15082 114490
rect 15082 114438 15084 114490
rect 15028 114436 15084 114438
rect 16828 116508 16884 116564
rect 16268 116396 16324 116452
rect 16716 116450 16772 116452
rect 16716 116398 16718 116450
rect 16718 116398 16770 116450
rect 16770 116398 16772 116450
rect 16716 116396 16772 116398
rect 18222 118410 18278 118412
rect 18222 118358 18224 118410
rect 18224 118358 18276 118410
rect 18276 118358 18278 118410
rect 18222 118356 18278 118358
rect 18326 118410 18382 118412
rect 18326 118358 18328 118410
rect 18328 118358 18380 118410
rect 18380 118358 18382 118410
rect 18326 118356 18382 118358
rect 18430 118410 18486 118412
rect 18430 118358 18432 118410
rect 18432 118358 18484 118410
rect 18484 118358 18486 118410
rect 18430 118356 18486 118358
rect 17388 116396 17444 116452
rect 13356 113036 13412 113092
rect 13020 112476 13076 112532
rect 12460 110236 12516 110292
rect 11418 109002 11474 109004
rect 11418 108950 11420 109002
rect 11420 108950 11472 109002
rect 11472 108950 11474 109002
rect 11418 108948 11474 108950
rect 11522 109002 11578 109004
rect 11522 108950 11524 109002
rect 11524 108950 11576 109002
rect 11576 108950 11578 109002
rect 11522 108948 11578 108950
rect 11626 109002 11682 109004
rect 11626 108950 11628 109002
rect 11628 108950 11680 109002
rect 11680 108950 11682 109002
rect 11626 108948 11682 108950
rect 9212 108498 9268 108500
rect 9212 108446 9214 108498
rect 9214 108446 9266 108498
rect 9266 108446 9268 108498
rect 9212 108444 9268 108446
rect 8016 108218 8072 108220
rect 8016 108166 8018 108218
rect 8018 108166 8070 108218
rect 8070 108166 8072 108218
rect 8016 108164 8072 108166
rect 8120 108218 8176 108220
rect 8120 108166 8122 108218
rect 8122 108166 8174 108218
rect 8174 108166 8176 108218
rect 8120 108164 8176 108166
rect 8224 108218 8280 108220
rect 8224 108166 8226 108218
rect 8226 108166 8278 108218
rect 8278 108166 8280 108218
rect 8224 108164 8280 108166
rect 7532 107660 7588 107716
rect 4614 107434 4670 107436
rect 4614 107382 4616 107434
rect 4616 107382 4668 107434
rect 4668 107382 4670 107434
rect 4614 107380 4670 107382
rect 4718 107434 4774 107436
rect 4718 107382 4720 107434
rect 4720 107382 4772 107434
rect 4772 107382 4774 107434
rect 4718 107380 4774 107382
rect 4822 107434 4878 107436
rect 4822 107382 4824 107434
rect 4824 107382 4876 107434
rect 4876 107382 4878 107434
rect 4822 107380 4878 107382
rect 3948 106428 4004 106484
rect 4284 106876 4340 106932
rect 3164 106092 3220 106148
rect 3836 106146 3892 106148
rect 3836 106094 3838 106146
rect 3838 106094 3890 106146
rect 3890 106094 3892 106146
rect 3836 106092 3892 106094
rect 1708 104860 1764 104916
rect 3836 104914 3892 104916
rect 3836 104862 3838 104914
rect 3838 104862 3890 104914
rect 3890 104862 3892 104914
rect 3836 104860 3892 104862
rect 4060 105644 4116 105700
rect 5628 106428 5684 106484
rect 4956 106092 5012 106148
rect 4844 105980 4900 106036
rect 4614 105866 4670 105868
rect 4614 105814 4616 105866
rect 4616 105814 4668 105866
rect 4668 105814 4670 105866
rect 4614 105812 4670 105814
rect 4718 105866 4774 105868
rect 4718 105814 4720 105866
rect 4720 105814 4772 105866
rect 4772 105814 4774 105866
rect 4718 105812 4774 105814
rect 4822 105866 4878 105868
rect 4822 105814 4824 105866
rect 4824 105814 4876 105866
rect 4876 105814 4878 105866
rect 4822 105812 4878 105814
rect 4284 105196 4340 105252
rect 4508 105474 4564 105476
rect 4508 105422 4510 105474
rect 4510 105422 4562 105474
rect 4562 105422 4564 105474
rect 4508 105420 4564 105422
rect 4284 104802 4340 104804
rect 4284 104750 4286 104802
rect 4286 104750 4338 104802
rect 4338 104750 4340 104802
rect 4284 104748 4340 104750
rect 3724 104690 3780 104692
rect 3724 104638 3726 104690
rect 3726 104638 3778 104690
rect 3778 104638 3780 104690
rect 3724 104636 3780 104638
rect 3276 104578 3332 104580
rect 3276 104526 3278 104578
rect 3278 104526 3330 104578
rect 3330 104526 3332 104578
rect 3276 104524 3332 104526
rect 1708 104018 1764 104020
rect 1708 103966 1710 104018
rect 1710 103966 1762 104018
rect 1762 103966 1764 104018
rect 1708 103964 1764 103966
rect 1708 103292 1764 103348
rect 2604 103122 2660 103124
rect 2604 103070 2606 103122
rect 2606 103070 2658 103122
rect 2658 103070 2660 103122
rect 2604 103068 2660 103070
rect 1708 101612 1764 101668
rect 4396 104524 4452 104580
rect 5740 106146 5796 106148
rect 5740 106094 5742 106146
rect 5742 106094 5794 106146
rect 5794 106094 5796 106146
rect 5740 106092 5796 106094
rect 5292 105420 5348 105476
rect 5180 104690 5236 104692
rect 5180 104638 5182 104690
rect 5182 104638 5234 104690
rect 5234 104638 5236 104690
rect 5180 104636 5236 104638
rect 5852 105196 5908 105252
rect 4614 104298 4670 104300
rect 4614 104246 4616 104298
rect 4616 104246 4668 104298
rect 4668 104246 4670 104298
rect 4614 104244 4670 104246
rect 4718 104298 4774 104300
rect 4718 104246 4720 104298
rect 4720 104246 4772 104298
rect 4772 104246 4774 104298
rect 4718 104244 4774 104246
rect 4822 104298 4878 104300
rect 4822 104246 4824 104298
rect 4824 104246 4876 104298
rect 4876 104246 4878 104298
rect 4822 104244 4878 104246
rect 4844 103964 4900 104020
rect 3276 103628 3332 103684
rect 3500 103234 3556 103236
rect 3500 103182 3502 103234
rect 3502 103182 3554 103234
rect 3554 103182 3556 103234
rect 3500 103180 3556 103182
rect 4284 103346 4340 103348
rect 4284 103294 4286 103346
rect 4286 103294 4338 103346
rect 4338 103294 4340 103346
rect 4284 103292 4340 103294
rect 4060 103234 4116 103236
rect 4060 103182 4062 103234
rect 4062 103182 4114 103234
rect 4114 103182 4116 103234
rect 4060 103180 4116 103182
rect 2716 102172 2772 102228
rect 2604 100658 2660 100660
rect 2604 100606 2606 100658
rect 2606 100606 2658 100658
rect 2658 100606 2660 100658
rect 2604 100604 2660 100606
rect 1708 98812 1764 98868
rect 2380 98364 2436 98420
rect 3052 101500 3108 101556
rect 3948 103122 4004 103124
rect 3948 103070 3950 103122
rect 3950 103070 4002 103122
rect 4002 103070 4004 103122
rect 3948 103068 4004 103070
rect 3612 102956 3668 103012
rect 3388 102338 3444 102340
rect 3388 102286 3390 102338
rect 3390 102286 3442 102338
rect 3442 102286 3444 102338
rect 3388 102284 3444 102286
rect 3500 101612 3556 101668
rect 2828 98700 2884 98756
rect 2716 98364 2772 98420
rect 2604 97692 2660 97748
rect 3948 100492 4004 100548
rect 4956 103628 5012 103684
rect 4956 103292 5012 103348
rect 5068 104076 5124 104132
rect 4844 103068 4900 103124
rect 5292 103852 5348 103908
rect 5852 104412 5908 104468
rect 6300 105532 6356 105588
rect 6860 104860 6916 104916
rect 6524 104690 6580 104692
rect 6524 104638 6526 104690
rect 6526 104638 6578 104690
rect 6578 104638 6580 104690
rect 6524 104636 6580 104638
rect 7084 104524 7140 104580
rect 6412 103180 6468 103236
rect 4614 102730 4670 102732
rect 4614 102678 4616 102730
rect 4616 102678 4668 102730
rect 4668 102678 4670 102730
rect 4614 102676 4670 102678
rect 4718 102730 4774 102732
rect 4718 102678 4720 102730
rect 4720 102678 4772 102730
rect 4772 102678 4774 102730
rect 4718 102676 4774 102678
rect 4822 102730 4878 102732
rect 4822 102678 4824 102730
rect 4824 102678 4876 102730
rect 4876 102678 4878 102730
rect 4822 102676 4878 102678
rect 4284 102284 4340 102340
rect 4284 102114 4340 102116
rect 4284 102062 4286 102114
rect 4286 102062 4338 102114
rect 4338 102062 4340 102114
rect 4284 102060 4340 102062
rect 4396 101500 4452 101556
rect 4732 102114 4788 102116
rect 4732 102062 4734 102114
rect 4734 102062 4786 102114
rect 4786 102062 4788 102114
rect 4732 102060 4788 102062
rect 5068 101500 5124 101556
rect 7084 103740 7140 103796
rect 6972 103346 7028 103348
rect 6972 103294 6974 103346
rect 6974 103294 7026 103346
rect 7026 103294 7028 103346
rect 6972 103292 7028 103294
rect 6524 102508 6580 102564
rect 6860 102844 6916 102900
rect 8016 106650 8072 106652
rect 8016 106598 8018 106650
rect 8018 106598 8070 106650
rect 8070 106598 8072 106650
rect 8016 106596 8072 106598
rect 8120 106650 8176 106652
rect 8120 106598 8122 106650
rect 8122 106598 8174 106650
rect 8174 106598 8176 106650
rect 8120 106596 8176 106598
rect 8224 106650 8280 106652
rect 8224 106598 8226 106650
rect 8226 106598 8278 106650
rect 8278 106598 8280 106650
rect 8224 106596 8280 106598
rect 8092 106258 8148 106260
rect 8092 106206 8094 106258
rect 8094 106206 8146 106258
rect 8146 106206 8148 106258
rect 8092 106204 8148 106206
rect 7644 106146 7700 106148
rect 7644 106094 7646 106146
rect 7646 106094 7698 106146
rect 7698 106094 7700 106146
rect 7644 106092 7700 106094
rect 8540 106146 8596 106148
rect 8540 106094 8542 106146
rect 8542 106094 8594 106146
rect 8594 106094 8596 106146
rect 8540 106092 8596 106094
rect 7532 105756 7588 105812
rect 7756 105586 7812 105588
rect 7756 105534 7758 105586
rect 7758 105534 7810 105586
rect 7810 105534 7812 105586
rect 7756 105532 7812 105534
rect 7532 105084 7588 105140
rect 8016 105082 8072 105084
rect 8016 105030 8018 105082
rect 8018 105030 8070 105082
rect 8070 105030 8072 105082
rect 8016 105028 8072 105030
rect 8120 105082 8176 105084
rect 8120 105030 8122 105082
rect 8122 105030 8174 105082
rect 8174 105030 8176 105082
rect 8120 105028 8176 105030
rect 8224 105082 8280 105084
rect 8224 105030 8226 105082
rect 8226 105030 8278 105082
rect 8278 105030 8280 105082
rect 8224 105028 8280 105030
rect 8092 104914 8148 104916
rect 8092 104862 8094 104914
rect 8094 104862 8146 104914
rect 8146 104862 8148 104914
rect 8092 104860 8148 104862
rect 8316 104860 8372 104916
rect 7644 104690 7700 104692
rect 7644 104638 7646 104690
rect 7646 104638 7698 104690
rect 7698 104638 7700 104690
rect 7644 104636 7700 104638
rect 7532 104412 7588 104468
rect 7868 104412 7924 104468
rect 7644 103628 7700 103684
rect 8540 104300 8596 104356
rect 8316 104188 8372 104244
rect 7980 103794 8036 103796
rect 7980 103742 7982 103794
rect 7982 103742 8034 103794
rect 8034 103742 8036 103794
rect 7980 103740 8036 103742
rect 8652 104188 8708 104244
rect 9100 106370 9156 106372
rect 9100 106318 9102 106370
rect 9102 106318 9154 106370
rect 9154 106318 9156 106370
rect 9100 106316 9156 106318
rect 8876 105362 8932 105364
rect 8876 105310 8878 105362
rect 8878 105310 8930 105362
rect 8930 105310 8932 105362
rect 8876 105308 8932 105310
rect 8988 104636 9044 104692
rect 8988 104076 9044 104132
rect 8876 103852 8932 103908
rect 8540 103740 8596 103796
rect 8016 103514 8072 103516
rect 8016 103462 8018 103514
rect 8018 103462 8070 103514
rect 8070 103462 8072 103514
rect 8016 103460 8072 103462
rect 8120 103514 8176 103516
rect 8120 103462 8122 103514
rect 8122 103462 8174 103514
rect 8174 103462 8176 103514
rect 8120 103460 8176 103462
rect 8224 103514 8280 103516
rect 8224 103462 8226 103514
rect 8226 103462 8278 103514
rect 8278 103462 8280 103514
rect 8224 103460 8280 103462
rect 8204 103292 8260 103348
rect 7756 103234 7812 103236
rect 7756 103182 7758 103234
rect 7758 103182 7810 103234
rect 7810 103182 7812 103234
rect 7756 103180 7812 103182
rect 5852 101554 5908 101556
rect 5852 101502 5854 101554
rect 5854 101502 5906 101554
rect 5906 101502 5908 101554
rect 5852 101500 5908 101502
rect 5180 101442 5236 101444
rect 5180 101390 5182 101442
rect 5182 101390 5234 101442
rect 5234 101390 5236 101442
rect 5180 101388 5236 101390
rect 4614 101162 4670 101164
rect 4614 101110 4616 101162
rect 4616 101110 4668 101162
rect 4668 101110 4670 101162
rect 4614 101108 4670 101110
rect 4718 101162 4774 101164
rect 4718 101110 4720 101162
rect 4720 101110 4772 101162
rect 4772 101110 4774 101162
rect 4718 101108 4774 101110
rect 4822 101162 4878 101164
rect 4822 101110 4824 101162
rect 4824 101110 4876 101162
rect 4876 101110 4878 101162
rect 4822 101108 4878 101110
rect 4844 100658 4900 100660
rect 4844 100606 4846 100658
rect 4846 100606 4898 100658
rect 4898 100606 4900 100658
rect 4844 100604 4900 100606
rect 4284 100210 4340 100212
rect 4284 100158 4286 100210
rect 4286 100158 4338 100210
rect 4338 100158 4340 100210
rect 4284 100156 4340 100158
rect 4956 100380 5012 100436
rect 4614 99594 4670 99596
rect 4614 99542 4616 99594
rect 4616 99542 4668 99594
rect 4668 99542 4670 99594
rect 4614 99540 4670 99542
rect 4718 99594 4774 99596
rect 4718 99542 4720 99594
rect 4720 99542 4772 99594
rect 4772 99542 4774 99594
rect 4718 99540 4774 99542
rect 4822 99594 4878 99596
rect 4822 99542 4824 99594
rect 4824 99542 4876 99594
rect 4876 99542 4878 99594
rect 4822 99540 4878 99542
rect 3164 98700 3220 98756
rect 3276 98812 3332 98868
rect 4396 98642 4452 98644
rect 4396 98590 4398 98642
rect 4398 98590 4450 98642
rect 4450 98590 4452 98642
rect 4396 98588 4452 98590
rect 4060 98530 4116 98532
rect 4060 98478 4062 98530
rect 4062 98478 4114 98530
rect 4114 98478 4116 98530
rect 4060 98476 4116 98478
rect 3388 98418 3444 98420
rect 3388 98366 3390 98418
rect 3390 98366 3442 98418
rect 3442 98366 3444 98418
rect 3388 98364 3444 98366
rect 5628 100716 5684 100772
rect 5740 100604 5796 100660
rect 5180 99372 5236 99428
rect 4956 98252 5012 98308
rect 4614 98026 4670 98028
rect 4614 97974 4616 98026
rect 4616 97974 4668 98026
rect 4668 97974 4670 98026
rect 4614 97972 4670 97974
rect 4718 98026 4774 98028
rect 4718 97974 4720 98026
rect 4720 97974 4772 98026
rect 4772 97974 4774 98026
rect 4718 97972 4774 97974
rect 4822 98026 4878 98028
rect 4822 97974 4824 98026
rect 4824 97974 4876 98026
rect 4876 97974 4878 98026
rect 4822 97972 4878 97974
rect 4620 97804 4676 97860
rect 3276 97746 3332 97748
rect 3276 97694 3278 97746
rect 3278 97694 3330 97746
rect 3330 97694 3332 97746
rect 3276 97692 3332 97694
rect 3836 97634 3892 97636
rect 3836 97582 3838 97634
rect 3838 97582 3890 97634
rect 3890 97582 3892 97634
rect 3836 97580 3892 97582
rect 1708 96178 1764 96180
rect 1708 96126 1710 96178
rect 1710 96126 1762 96178
rect 1762 96126 1764 96178
rect 1708 96124 1764 96126
rect 3164 96738 3220 96740
rect 3164 96686 3166 96738
rect 3166 96686 3218 96738
rect 3218 96686 3220 96738
rect 3164 96684 3220 96686
rect 2268 96124 2324 96180
rect 2380 95506 2436 95508
rect 2380 95454 2382 95506
rect 2382 95454 2434 95506
rect 2434 95454 2436 95506
rect 2380 95452 2436 95454
rect 2828 95394 2884 95396
rect 2828 95342 2830 95394
rect 2830 95342 2882 95394
rect 2882 95342 2884 95394
rect 2828 95340 2884 95342
rect 2492 93996 2548 94052
rect 3836 96684 3892 96740
rect 3276 95676 3332 95732
rect 3388 96572 3444 96628
rect 4172 96738 4228 96740
rect 4172 96686 4174 96738
rect 4174 96686 4226 96738
rect 4226 96686 4228 96738
rect 4172 96684 4228 96686
rect 4956 97692 5012 97748
rect 3724 95170 3780 95172
rect 3724 95118 3726 95170
rect 3726 95118 3778 95170
rect 3778 95118 3780 95170
rect 3724 95116 3780 95118
rect 3948 95004 4004 95060
rect 3052 94610 3108 94612
rect 3052 94558 3054 94610
rect 3054 94558 3106 94610
rect 3106 94558 3108 94610
rect 3052 94556 3108 94558
rect 1708 93436 1764 93492
rect 3724 94556 3780 94612
rect 3276 93996 3332 94052
rect 3052 93602 3108 93604
rect 3052 93550 3054 93602
rect 3054 93550 3106 93602
rect 3106 93550 3108 93602
rect 3052 93548 3108 93550
rect 4614 96458 4670 96460
rect 4614 96406 4616 96458
rect 4616 96406 4668 96458
rect 4668 96406 4670 96458
rect 4614 96404 4670 96406
rect 4718 96458 4774 96460
rect 4718 96406 4720 96458
rect 4720 96406 4772 96458
rect 4772 96406 4774 96458
rect 4718 96404 4774 96406
rect 4822 96458 4878 96460
rect 4822 96406 4824 96458
rect 4824 96406 4876 96458
rect 4876 96406 4878 96458
rect 4822 96404 4878 96406
rect 5180 98418 5236 98420
rect 5180 98366 5182 98418
rect 5182 98366 5234 98418
rect 5234 98366 5236 98418
rect 5180 98364 5236 98366
rect 5068 97522 5124 97524
rect 5068 97470 5070 97522
rect 5070 97470 5122 97522
rect 5122 97470 5124 97522
rect 5068 97468 5124 97470
rect 4508 95170 4564 95172
rect 4508 95118 4510 95170
rect 4510 95118 4562 95170
rect 4562 95118 4564 95170
rect 4508 95116 4564 95118
rect 4614 94890 4670 94892
rect 4614 94838 4616 94890
rect 4616 94838 4668 94890
rect 4668 94838 4670 94890
rect 4614 94836 4670 94838
rect 4718 94890 4774 94892
rect 4718 94838 4720 94890
rect 4720 94838 4772 94890
rect 4772 94838 4774 94890
rect 4718 94836 4774 94838
rect 4822 94890 4878 94892
rect 4822 94838 4824 94890
rect 4824 94838 4876 94890
rect 4876 94838 4878 94890
rect 4822 94836 4878 94838
rect 4844 94668 4900 94724
rect 4060 94220 4116 94276
rect 5180 95116 5236 95172
rect 5180 94780 5236 94836
rect 3500 93436 3556 93492
rect 3836 93548 3892 93604
rect 4508 93602 4564 93604
rect 4508 93550 4510 93602
rect 4510 93550 4562 93602
rect 4562 93550 4564 93602
rect 4508 93548 4564 93550
rect 4614 93322 4670 93324
rect 4614 93270 4616 93322
rect 4616 93270 4668 93322
rect 4668 93270 4670 93322
rect 4614 93268 4670 93270
rect 4718 93322 4774 93324
rect 4718 93270 4720 93322
rect 4720 93270 4772 93322
rect 4772 93270 4774 93322
rect 4718 93268 4774 93270
rect 4822 93322 4878 93324
rect 4822 93270 4824 93322
rect 4824 93270 4876 93322
rect 4876 93270 4878 93322
rect 4822 93268 4878 93270
rect 6524 100716 6580 100772
rect 5964 100604 6020 100660
rect 6412 100658 6468 100660
rect 6412 100606 6414 100658
rect 6414 100606 6466 100658
rect 6466 100606 6468 100658
rect 6412 100604 6468 100606
rect 6188 100268 6244 100324
rect 5740 99148 5796 99204
rect 5852 98476 5908 98532
rect 5964 98252 6020 98308
rect 6188 98588 6244 98644
rect 5516 96124 5572 96180
rect 5628 97580 5684 97636
rect 5404 95788 5460 95844
rect 5852 97634 5908 97636
rect 5852 97582 5854 97634
rect 5854 97582 5906 97634
rect 5906 97582 5908 97634
rect 5852 97580 5908 97582
rect 6076 97634 6132 97636
rect 6076 97582 6078 97634
rect 6078 97582 6130 97634
rect 6130 97582 6132 97634
rect 6076 97580 6132 97582
rect 5740 96684 5796 96740
rect 5964 96348 6020 96404
rect 5628 95340 5684 95396
rect 5292 93548 5348 93604
rect 5180 93042 5236 93044
rect 5180 92990 5182 93042
rect 5182 92990 5234 93042
rect 5234 92990 5236 93042
rect 5180 92988 5236 92990
rect 2940 92316 2996 92372
rect 4284 92316 4340 92372
rect 2492 92258 2548 92260
rect 2492 92206 2494 92258
rect 2494 92206 2546 92258
rect 2546 92206 2548 92258
rect 2492 92204 2548 92206
rect 3276 92258 3332 92260
rect 3276 92206 3278 92258
rect 3278 92206 3330 92258
rect 3330 92206 3332 92258
rect 3276 92204 3332 92206
rect 1820 91980 1876 92036
rect 2828 92034 2884 92036
rect 2828 91982 2830 92034
rect 2830 91982 2882 92034
rect 2882 91982 2884 92034
rect 2828 91980 2884 91982
rect 3388 91532 3444 91588
rect 1708 90524 1764 90580
rect 2492 88844 2548 88900
rect 1708 88114 1764 88116
rect 1708 88062 1710 88114
rect 1710 88062 1762 88114
rect 1762 88062 1764 88114
rect 1708 88060 1764 88062
rect 3836 88898 3892 88900
rect 3836 88846 3838 88898
rect 3838 88846 3890 88898
rect 3890 88846 3892 88898
rect 3836 88844 3892 88846
rect 2828 87948 2884 88004
rect 3388 88002 3444 88004
rect 3388 87950 3390 88002
rect 3390 87950 3442 88002
rect 3442 87950 3444 88002
rect 3388 87948 3444 87950
rect 2044 87500 2100 87556
rect 3052 87388 3108 87444
rect 2044 85986 2100 85988
rect 2044 85934 2046 85986
rect 2046 85934 2098 85986
rect 2098 85934 2100 85986
rect 2044 85932 2100 85934
rect 1708 85372 1764 85428
rect 4620 91980 4676 92036
rect 4614 91754 4670 91756
rect 4614 91702 4616 91754
rect 4616 91702 4668 91754
rect 4668 91702 4670 91754
rect 4614 91700 4670 91702
rect 4718 91754 4774 91756
rect 4718 91702 4720 91754
rect 4720 91702 4772 91754
rect 4772 91702 4774 91754
rect 4718 91700 4774 91702
rect 4822 91754 4878 91756
rect 4822 91702 4824 91754
rect 4824 91702 4876 91754
rect 4876 91702 4878 91754
rect 4822 91700 4878 91702
rect 4508 90690 4564 90692
rect 4508 90638 4510 90690
rect 4510 90638 4562 90690
rect 4562 90638 4564 90690
rect 4508 90636 4564 90638
rect 4614 90186 4670 90188
rect 4614 90134 4616 90186
rect 4616 90134 4668 90186
rect 4668 90134 4670 90186
rect 4614 90132 4670 90134
rect 4718 90186 4774 90188
rect 4718 90134 4720 90186
rect 4720 90134 4772 90186
rect 4772 90134 4774 90186
rect 4718 90132 4774 90134
rect 4822 90186 4878 90188
rect 4822 90134 4824 90186
rect 4824 90134 4876 90186
rect 4876 90134 4878 90186
rect 4822 90132 4878 90134
rect 5068 91138 5124 91140
rect 5068 91086 5070 91138
rect 5070 91086 5122 91138
rect 5122 91086 5124 91138
rect 5068 91084 5124 91086
rect 5404 95228 5460 95284
rect 6076 95954 6132 95956
rect 6076 95902 6078 95954
rect 6078 95902 6130 95954
rect 6130 95902 6132 95954
rect 6076 95900 6132 95902
rect 6076 95452 6132 95508
rect 6300 97692 6356 97748
rect 8316 103180 8372 103236
rect 8316 102732 8372 102788
rect 6860 102114 6916 102116
rect 6860 102062 6862 102114
rect 6862 102062 6914 102114
rect 6914 102062 6916 102114
rect 6860 102060 6916 102062
rect 6860 101500 6916 101556
rect 7084 99820 7140 99876
rect 6636 99202 6692 99204
rect 6636 99150 6638 99202
rect 6638 99150 6690 99202
rect 6690 99150 6692 99202
rect 6636 99148 6692 99150
rect 6860 99036 6916 99092
rect 8876 103516 8932 103572
rect 8988 103068 9044 103124
rect 8988 102732 9044 102788
rect 8764 102284 8820 102340
rect 8652 102060 8708 102116
rect 8016 101946 8072 101948
rect 8016 101894 8018 101946
rect 8018 101894 8070 101946
rect 8070 101894 8072 101946
rect 8016 101892 8072 101894
rect 8120 101946 8176 101948
rect 8120 101894 8122 101946
rect 8122 101894 8174 101946
rect 8174 101894 8176 101946
rect 8120 101892 8176 101894
rect 8224 101946 8280 101948
rect 8224 101894 8226 101946
rect 8226 101894 8278 101946
rect 8278 101894 8280 101946
rect 8224 101892 8280 101894
rect 7756 101276 7812 101332
rect 8540 101836 8596 101892
rect 7420 100882 7476 100884
rect 7420 100830 7422 100882
rect 7422 100830 7474 100882
rect 7474 100830 7476 100882
rect 7420 100828 7476 100830
rect 7420 100604 7476 100660
rect 7308 100380 7364 100436
rect 7756 100268 7812 100324
rect 8016 100378 8072 100380
rect 8016 100326 8018 100378
rect 8018 100326 8070 100378
rect 8070 100326 8072 100378
rect 8016 100324 8072 100326
rect 8120 100378 8176 100380
rect 8120 100326 8122 100378
rect 8122 100326 8174 100378
rect 8174 100326 8176 100378
rect 8120 100324 8176 100326
rect 8224 100378 8280 100380
rect 8224 100326 8226 100378
rect 8226 100326 8278 100378
rect 8278 100326 8280 100378
rect 8224 100324 8280 100326
rect 7532 99932 7588 99988
rect 8876 100940 8932 100996
rect 8988 102172 9044 102228
rect 8764 100828 8820 100884
rect 9212 104076 9268 104132
rect 9660 106764 9716 106820
rect 9772 107772 9828 107828
rect 9884 107548 9940 107604
rect 9996 106988 10052 107044
rect 12460 109228 12516 109284
rect 11418 107434 11474 107436
rect 11418 107382 11420 107434
rect 11420 107382 11472 107434
rect 11472 107382 11474 107434
rect 11418 107380 11474 107382
rect 11522 107434 11578 107436
rect 11522 107382 11524 107434
rect 11524 107382 11576 107434
rect 11576 107382 11578 107434
rect 11522 107380 11578 107382
rect 11626 107434 11682 107436
rect 11626 107382 11628 107434
rect 11628 107382 11680 107434
rect 11680 107382 11682 107434
rect 11626 107380 11682 107382
rect 10780 106988 10836 107044
rect 10108 106818 10164 106820
rect 10108 106766 10110 106818
rect 10110 106766 10162 106818
rect 10162 106766 10164 106818
rect 10108 106764 10164 106766
rect 9996 106204 10052 106260
rect 9212 102844 9268 102900
rect 9212 102620 9268 102676
rect 11452 107042 11508 107044
rect 11452 106990 11454 107042
rect 11454 106990 11506 107042
rect 11506 106990 11508 107042
rect 11452 106988 11508 106990
rect 12572 108610 12628 108612
rect 12572 108558 12574 108610
rect 12574 108558 12626 108610
rect 12626 108558 12628 108610
rect 12572 108556 12628 108558
rect 12796 110012 12852 110068
rect 12908 109228 12964 109284
rect 14820 112922 14876 112924
rect 14820 112870 14822 112922
rect 14822 112870 14874 112922
rect 14874 112870 14876 112922
rect 14820 112868 14876 112870
rect 14924 112922 14980 112924
rect 14924 112870 14926 112922
rect 14926 112870 14978 112922
rect 14978 112870 14980 112922
rect 14924 112868 14980 112870
rect 15028 112922 15084 112924
rect 15028 112870 15030 112922
rect 15030 112870 15082 112922
rect 15082 112870 15084 112922
rect 15028 112868 15084 112870
rect 14700 112530 14756 112532
rect 14700 112478 14702 112530
rect 14702 112478 14754 112530
rect 14754 112478 14756 112530
rect 14700 112476 14756 112478
rect 14820 111354 14876 111356
rect 14820 111302 14822 111354
rect 14822 111302 14874 111354
rect 14874 111302 14876 111354
rect 14820 111300 14876 111302
rect 14924 111354 14980 111356
rect 14924 111302 14926 111354
rect 14926 111302 14978 111354
rect 14978 111302 14980 111354
rect 14924 111300 14980 111302
rect 15028 111354 15084 111356
rect 15028 111302 15030 111354
rect 15030 111302 15082 111354
rect 15082 111302 15084 111354
rect 15028 111300 15084 111302
rect 14476 110684 14532 110740
rect 13916 110012 13972 110068
rect 14252 110124 14308 110180
rect 14028 109340 14084 109396
rect 13468 109228 13524 109284
rect 13692 108444 13748 108500
rect 12236 107714 12292 107716
rect 12236 107662 12238 107714
rect 12238 107662 12290 107714
rect 12290 107662 12292 107714
rect 12236 107660 12292 107662
rect 12124 107548 12180 107604
rect 11788 106988 11844 107044
rect 10444 105308 10500 105364
rect 11418 105866 11474 105868
rect 11418 105814 11420 105866
rect 11420 105814 11472 105866
rect 11472 105814 11474 105866
rect 11418 105812 11474 105814
rect 11522 105866 11578 105868
rect 11522 105814 11524 105866
rect 11524 105814 11576 105866
rect 11576 105814 11578 105866
rect 11522 105812 11578 105814
rect 11626 105866 11682 105868
rect 11626 105814 11628 105866
rect 11628 105814 11680 105866
rect 11680 105814 11682 105866
rect 11626 105812 11682 105814
rect 12460 107042 12516 107044
rect 12460 106990 12462 107042
rect 12462 106990 12514 107042
rect 12514 106990 12516 107042
rect 12460 106988 12516 106990
rect 12348 106316 12404 106372
rect 13580 107826 13636 107828
rect 13580 107774 13582 107826
rect 13582 107774 13634 107826
rect 13634 107774 13636 107826
rect 13580 107772 13636 107774
rect 14820 109786 14876 109788
rect 14820 109734 14822 109786
rect 14822 109734 14874 109786
rect 14874 109734 14876 109786
rect 14820 109732 14876 109734
rect 14924 109786 14980 109788
rect 14924 109734 14926 109786
rect 14926 109734 14978 109786
rect 14978 109734 14980 109786
rect 14924 109732 14980 109734
rect 15028 109786 15084 109788
rect 15028 109734 15030 109786
rect 15030 109734 15082 109786
rect 15082 109734 15084 109786
rect 15028 109732 15084 109734
rect 15036 109228 15092 109284
rect 14924 108610 14980 108612
rect 14924 108558 14926 108610
rect 14926 108558 14978 108610
rect 14978 108558 14980 108610
rect 14924 108556 14980 108558
rect 14820 108218 14876 108220
rect 14820 108166 14822 108218
rect 14822 108166 14874 108218
rect 14874 108166 14876 108218
rect 14820 108164 14876 108166
rect 14924 108218 14980 108220
rect 14924 108166 14926 108218
rect 14926 108166 14978 108218
rect 14978 108166 14980 108218
rect 14924 108164 14980 108166
rect 15028 108218 15084 108220
rect 15028 108166 15030 108218
rect 15030 108166 15082 108218
rect 15082 108166 15084 108218
rect 15028 108164 15084 108166
rect 14924 107996 14980 108052
rect 13580 107042 13636 107044
rect 13580 106990 13582 107042
rect 13582 106990 13634 107042
rect 13634 106990 13636 107042
rect 13580 106988 13636 106990
rect 13468 106930 13524 106932
rect 13468 106878 13470 106930
rect 13470 106878 13522 106930
rect 13522 106878 13524 106930
rect 13468 106876 13524 106878
rect 12684 105868 12740 105924
rect 13580 105868 13636 105924
rect 12684 105644 12740 105700
rect 12796 105532 12852 105588
rect 11788 104690 11844 104692
rect 11788 104638 11790 104690
rect 11790 104638 11842 104690
rect 11842 104638 11844 104690
rect 11788 104636 11844 104638
rect 11228 104412 11284 104468
rect 10108 104076 10164 104132
rect 9884 103906 9940 103908
rect 9884 103854 9886 103906
rect 9886 103854 9938 103906
rect 9938 103854 9940 103906
rect 9884 103852 9940 103854
rect 9548 103740 9604 103796
rect 9548 103346 9604 103348
rect 9548 103294 9550 103346
rect 9550 103294 9602 103346
rect 9602 103294 9604 103346
rect 9548 103292 9604 103294
rect 12460 104412 12516 104468
rect 12684 104860 12740 104916
rect 11418 104298 11474 104300
rect 11418 104246 11420 104298
rect 11420 104246 11472 104298
rect 11472 104246 11474 104298
rect 11418 104244 11474 104246
rect 11522 104298 11578 104300
rect 11522 104246 11524 104298
rect 11524 104246 11576 104298
rect 11576 104246 11578 104298
rect 11522 104244 11578 104246
rect 11626 104298 11682 104300
rect 11626 104246 11628 104298
rect 11628 104246 11680 104298
rect 11680 104246 11682 104298
rect 11626 104244 11682 104246
rect 10108 103740 10164 103796
rect 9436 102732 9492 102788
rect 9212 101836 9268 101892
rect 9324 100828 9380 100884
rect 9212 100716 9268 100772
rect 7420 99036 7476 99092
rect 7084 97804 7140 97860
rect 6860 97692 6916 97748
rect 6748 97634 6804 97636
rect 6748 97582 6750 97634
rect 6750 97582 6802 97634
rect 6802 97582 6804 97634
rect 6748 97580 6804 97582
rect 6636 97468 6692 97524
rect 6636 96178 6692 96180
rect 6636 96126 6638 96178
rect 6638 96126 6690 96178
rect 6690 96126 6692 96178
rect 6636 96124 6692 96126
rect 5852 94892 5908 94948
rect 5740 94610 5796 94612
rect 5740 94558 5742 94610
rect 5742 94558 5794 94610
rect 5794 94558 5796 94610
rect 5740 94556 5796 94558
rect 5516 93602 5572 93604
rect 5516 93550 5518 93602
rect 5518 93550 5570 93602
rect 5570 93550 5572 93602
rect 5516 93548 5572 93550
rect 5404 92204 5460 92260
rect 6524 95506 6580 95508
rect 6524 95454 6526 95506
rect 6526 95454 6578 95506
rect 6578 95454 6580 95506
rect 6524 95452 6580 95454
rect 6188 94108 6244 94164
rect 6300 95116 6356 95172
rect 6076 93884 6132 93940
rect 6188 93548 6244 93604
rect 6076 93324 6132 93380
rect 5292 90748 5348 90804
rect 5852 92204 5908 92260
rect 5740 91586 5796 91588
rect 5740 91534 5742 91586
rect 5742 91534 5794 91586
rect 5794 91534 5796 91586
rect 5740 91532 5796 91534
rect 6412 93884 6468 93940
rect 6412 93436 6468 93492
rect 6636 94780 6692 94836
rect 7196 96012 7252 96068
rect 6860 95452 6916 95508
rect 6972 95170 7028 95172
rect 6972 95118 6974 95170
rect 6974 95118 7026 95170
rect 7026 95118 7028 95170
rect 6972 95116 7028 95118
rect 6748 94668 6804 94724
rect 6524 92988 6580 93044
rect 6076 91474 6132 91476
rect 6076 91422 6078 91474
rect 6078 91422 6130 91474
rect 6130 91422 6132 91474
rect 6076 91420 6132 91422
rect 5740 90690 5796 90692
rect 5740 90638 5742 90690
rect 5742 90638 5794 90690
rect 5794 90638 5796 90690
rect 5740 90636 5796 90638
rect 6636 94108 6692 94164
rect 4614 88618 4670 88620
rect 4614 88566 4616 88618
rect 4616 88566 4668 88618
rect 4668 88566 4670 88618
rect 4614 88564 4670 88566
rect 4718 88618 4774 88620
rect 4718 88566 4720 88618
rect 4720 88566 4772 88618
rect 4772 88566 4774 88618
rect 4718 88564 4774 88566
rect 4822 88618 4878 88620
rect 4822 88566 4824 88618
rect 4824 88566 4876 88618
rect 4876 88566 4878 88618
rect 4822 88564 4878 88566
rect 5068 88284 5124 88340
rect 5068 87388 5124 87444
rect 5292 87500 5348 87556
rect 4614 87050 4670 87052
rect 4614 86998 4616 87050
rect 4616 86998 4668 87050
rect 4668 86998 4670 87050
rect 4614 86996 4670 86998
rect 4718 87050 4774 87052
rect 4718 86998 4720 87050
rect 4720 86998 4772 87050
rect 4772 86998 4774 87050
rect 4718 86996 4774 86998
rect 4822 87050 4878 87052
rect 4822 86998 4824 87050
rect 4824 86998 4876 87050
rect 4876 86998 4878 87050
rect 4822 86996 4878 86998
rect 2492 85372 2548 85428
rect 4614 85482 4670 85484
rect 4614 85430 4616 85482
rect 4616 85430 4668 85482
rect 4668 85430 4670 85482
rect 4614 85428 4670 85430
rect 4718 85482 4774 85484
rect 4718 85430 4720 85482
rect 4720 85430 4772 85482
rect 4772 85430 4774 85482
rect 4718 85428 4774 85430
rect 4822 85482 4878 85484
rect 4822 85430 4824 85482
rect 4824 85430 4876 85482
rect 4876 85430 4878 85482
rect 4822 85428 4878 85430
rect 3052 85090 3108 85092
rect 3052 85038 3054 85090
rect 3054 85038 3106 85090
rect 3106 85038 3108 85090
rect 3052 85036 3108 85038
rect 1708 83410 1764 83412
rect 1708 83358 1710 83410
rect 1710 83358 1762 83410
rect 1762 83358 1764 83410
rect 1708 83356 1764 83358
rect 2492 83356 2548 83412
rect 1708 82684 1764 82740
rect 2044 82684 2100 82740
rect 1820 82236 1876 82292
rect 2268 81900 2324 81956
rect 2828 82514 2884 82516
rect 2828 82462 2830 82514
rect 2830 82462 2882 82514
rect 2882 82462 2884 82514
rect 2828 82460 2884 82462
rect 2604 81228 2660 81284
rect 3276 83410 3332 83412
rect 3276 83358 3278 83410
rect 3278 83358 3330 83410
rect 3330 83358 3332 83410
rect 3276 83356 3332 83358
rect 3276 82684 3332 82740
rect 3052 82124 3108 82180
rect 2044 80162 2100 80164
rect 2044 80110 2046 80162
rect 2046 80110 2098 80162
rect 2098 80110 2100 80162
rect 2044 80108 2100 80110
rect 1708 79996 1764 80052
rect 2492 79996 2548 80052
rect 3388 82514 3444 82516
rect 3388 82462 3390 82514
rect 3390 82462 3442 82514
rect 3442 82462 3444 82514
rect 3388 82460 3444 82462
rect 3724 81900 3780 81956
rect 1708 77308 1764 77364
rect 3164 78540 3220 78596
rect 2828 78204 2884 78260
rect 1932 77308 1988 77364
rect 2940 78034 2996 78036
rect 2940 77982 2942 78034
rect 2942 77982 2994 78034
rect 2994 77982 2996 78034
rect 2940 77980 2996 77982
rect 2044 77084 2100 77140
rect 2716 77138 2772 77140
rect 2716 77086 2718 77138
rect 2718 77086 2770 77138
rect 2770 77086 2772 77138
rect 2716 77084 2772 77086
rect 1708 74620 1764 74676
rect 2044 74844 2100 74900
rect 2268 74620 2324 74676
rect 2492 74172 2548 74228
rect 2940 75628 2996 75684
rect 2828 74844 2884 74900
rect 3500 78034 3556 78036
rect 3500 77982 3502 78034
rect 3502 77982 3554 78034
rect 3554 77982 3556 78034
rect 3500 77980 3556 77982
rect 3500 77250 3556 77252
rect 3500 77198 3502 77250
rect 3502 77198 3554 77250
rect 3554 77198 3556 77250
rect 3500 77196 3556 77198
rect 3500 76524 3556 76580
rect 3724 76524 3780 76580
rect 3612 74898 3668 74900
rect 3612 74846 3614 74898
rect 3614 74846 3666 74898
rect 3666 74846 3668 74898
rect 3612 74844 3668 74846
rect 3164 74284 3220 74340
rect 2940 74172 2996 74228
rect 2940 73500 2996 73556
rect 2044 73442 2100 73444
rect 2044 73390 2046 73442
rect 2046 73390 2098 73442
rect 2098 73390 2100 73442
rect 2044 73388 2100 73390
rect 2716 73388 2772 73444
rect 1820 72546 1876 72548
rect 1820 72494 1822 72546
rect 1822 72494 1874 72546
rect 1874 72494 1876 72546
rect 1820 72492 1876 72494
rect 2380 73276 2436 73332
rect 1708 71932 1764 71988
rect 2268 71874 2324 71876
rect 2268 71822 2270 71874
rect 2270 71822 2322 71874
rect 2322 71822 2324 71874
rect 2268 71820 2324 71822
rect 1820 70476 1876 70532
rect 1932 70700 1988 70756
rect 2604 71762 2660 71764
rect 2604 71710 2606 71762
rect 2606 71710 2658 71762
rect 2658 71710 2660 71762
rect 2604 71708 2660 71710
rect 3052 72156 3108 72212
rect 3612 74172 3668 74228
rect 3500 72380 3556 72436
rect 3276 71820 3332 71876
rect 2604 70754 2660 70756
rect 2604 70702 2606 70754
rect 2606 70702 2658 70754
rect 2658 70702 2660 70754
rect 2604 70700 2660 70702
rect 3612 72156 3668 72212
rect 3388 71762 3444 71764
rect 3388 71710 3390 71762
rect 3390 71710 3442 71762
rect 3442 71710 3444 71762
rect 3388 71708 3444 71710
rect 3052 70476 3108 70532
rect 3276 70700 3332 70756
rect 3052 70082 3108 70084
rect 3052 70030 3054 70082
rect 3054 70030 3106 70082
rect 3106 70030 3108 70082
rect 3052 70028 3108 70030
rect 1820 69244 1876 69300
rect 1596 67004 1652 67060
rect 2044 67170 2100 67172
rect 2044 67118 2046 67170
rect 2046 67118 2098 67170
rect 2098 67118 2100 67170
rect 2044 67116 2100 67118
rect 3388 69020 3444 69076
rect 6076 88844 6132 88900
rect 5740 88338 5796 88340
rect 5740 88286 5742 88338
rect 5742 88286 5794 88338
rect 5794 88286 5796 88338
rect 5740 88284 5796 88286
rect 6524 90748 6580 90804
rect 6524 89180 6580 89236
rect 6412 88956 6468 89012
rect 5852 85762 5908 85764
rect 5852 85710 5854 85762
rect 5854 85710 5906 85762
rect 5906 85710 5908 85762
rect 5852 85708 5908 85710
rect 4956 85036 5012 85092
rect 4956 84476 5012 84532
rect 4614 83914 4670 83916
rect 4614 83862 4616 83914
rect 4616 83862 4668 83914
rect 4668 83862 4670 83914
rect 4614 83860 4670 83862
rect 4718 83914 4774 83916
rect 4718 83862 4720 83914
rect 4720 83862 4772 83914
rect 4772 83862 4774 83914
rect 4718 83860 4774 83862
rect 4822 83914 4878 83916
rect 4822 83862 4824 83914
rect 4824 83862 4876 83914
rect 4876 83862 4878 83914
rect 4822 83860 4878 83862
rect 4172 83356 4228 83412
rect 4060 83244 4116 83300
rect 4060 82460 4116 82516
rect 4620 83298 4676 83300
rect 4620 83246 4622 83298
rect 4622 83246 4674 83298
rect 4674 83246 4676 83298
rect 4620 83244 4676 83246
rect 6860 94780 6916 94836
rect 6748 91084 6804 91140
rect 7196 94780 7252 94836
rect 7084 94332 7140 94388
rect 7644 99202 7700 99204
rect 7644 99150 7646 99202
rect 7646 99150 7698 99202
rect 7698 99150 7700 99202
rect 7644 99148 7700 99150
rect 7532 98028 7588 98084
rect 8540 99372 8596 99428
rect 8988 100210 9044 100212
rect 8988 100158 8990 100210
rect 8990 100158 9042 100210
rect 9042 100158 9044 100210
rect 8988 100156 9044 100158
rect 8764 98924 8820 98980
rect 8016 98810 8072 98812
rect 8016 98758 8018 98810
rect 8018 98758 8070 98810
rect 8070 98758 8072 98810
rect 8016 98756 8072 98758
rect 8120 98810 8176 98812
rect 8120 98758 8122 98810
rect 8122 98758 8174 98810
rect 8174 98758 8176 98810
rect 8120 98756 8176 98758
rect 8224 98810 8280 98812
rect 8224 98758 8226 98810
rect 8226 98758 8278 98810
rect 8278 98758 8280 98810
rect 8224 98756 8280 98758
rect 8764 98364 8820 98420
rect 7308 94220 7364 94276
rect 7084 94108 7140 94164
rect 6972 92930 7028 92932
rect 6972 92878 6974 92930
rect 6974 92878 7026 92930
rect 7026 92878 7028 92930
rect 6972 92876 7028 92878
rect 7308 91420 7364 91476
rect 7532 97244 7588 97300
rect 8016 97242 8072 97244
rect 8016 97190 8018 97242
rect 8018 97190 8070 97242
rect 8070 97190 8072 97242
rect 8016 97188 8072 97190
rect 8120 97242 8176 97244
rect 8120 97190 8122 97242
rect 8122 97190 8174 97242
rect 8174 97190 8176 97242
rect 8120 97188 8176 97190
rect 8224 97242 8280 97244
rect 8224 97190 8226 97242
rect 8226 97190 8278 97242
rect 8278 97190 8280 97242
rect 8224 97188 8280 97190
rect 9660 103068 9716 103124
rect 9884 102844 9940 102900
rect 9660 102732 9716 102788
rect 9660 102226 9716 102228
rect 9660 102174 9662 102226
rect 9662 102174 9714 102226
rect 9714 102174 9716 102226
rect 9660 102172 9716 102174
rect 10668 103740 10724 103796
rect 11116 103794 11172 103796
rect 11116 103742 11118 103794
rect 11118 103742 11170 103794
rect 11170 103742 11172 103794
rect 11116 103740 11172 103742
rect 10220 103292 10276 103348
rect 10108 102620 10164 102676
rect 10220 102508 10276 102564
rect 10332 102732 10388 102788
rect 10108 102338 10164 102340
rect 10108 102286 10110 102338
rect 10110 102286 10162 102338
rect 10162 102286 10164 102338
rect 10108 102284 10164 102286
rect 9884 102060 9940 102116
rect 9548 101612 9604 101668
rect 9884 101666 9940 101668
rect 9884 101614 9886 101666
rect 9886 101614 9938 101666
rect 9938 101614 9940 101666
rect 9884 101612 9940 101614
rect 9772 101276 9828 101332
rect 9772 100828 9828 100884
rect 9548 100380 9604 100436
rect 9436 98476 9492 98532
rect 9548 98418 9604 98420
rect 9548 98366 9550 98418
rect 9550 98366 9602 98418
rect 9602 98366 9604 98418
rect 9548 98364 9604 98366
rect 10220 101388 10276 101444
rect 10444 100604 10500 100660
rect 10108 100380 10164 100436
rect 9884 100156 9940 100212
rect 10108 99986 10164 99988
rect 10108 99934 10110 99986
rect 10110 99934 10162 99986
rect 10162 99934 10164 99986
rect 10108 99932 10164 99934
rect 9884 99036 9940 99092
rect 10668 103122 10724 103124
rect 10668 103070 10670 103122
rect 10670 103070 10722 103122
rect 10722 103070 10724 103122
rect 10668 103068 10724 103070
rect 10780 103010 10836 103012
rect 10780 102958 10782 103010
rect 10782 102958 10834 103010
rect 10834 102958 10836 103010
rect 10780 102956 10836 102958
rect 10668 102844 10724 102900
rect 10668 100380 10724 100436
rect 10780 100940 10836 100996
rect 11116 103068 11172 103124
rect 11116 102844 11172 102900
rect 11788 103404 11844 103460
rect 11228 102956 11284 103012
rect 11228 102732 11284 102788
rect 11418 102730 11474 102732
rect 11418 102678 11420 102730
rect 11420 102678 11472 102730
rect 11472 102678 11474 102730
rect 11418 102676 11474 102678
rect 11522 102730 11578 102732
rect 11522 102678 11524 102730
rect 11524 102678 11576 102730
rect 11576 102678 11578 102730
rect 11522 102676 11578 102678
rect 11626 102730 11682 102732
rect 11626 102678 11628 102730
rect 11628 102678 11680 102730
rect 11680 102678 11682 102730
rect 11626 102676 11682 102678
rect 12572 103180 12628 103236
rect 12796 104748 12852 104804
rect 12908 104076 12964 104132
rect 13020 103180 13076 103236
rect 13804 104412 13860 104468
rect 14588 106876 14644 106932
rect 14820 106650 14876 106652
rect 14820 106598 14822 106650
rect 14822 106598 14874 106650
rect 14874 106598 14876 106650
rect 14820 106596 14876 106598
rect 14924 106650 14980 106652
rect 14924 106598 14926 106650
rect 14926 106598 14978 106650
rect 14978 106598 14980 106650
rect 14924 106596 14980 106598
rect 15028 106650 15084 106652
rect 15028 106598 15030 106650
rect 15030 106598 15082 106650
rect 15082 106598 15084 106650
rect 15028 106596 15084 106598
rect 14588 105868 14644 105924
rect 14252 104636 14308 104692
rect 13804 102956 13860 103012
rect 12124 102284 12180 102340
rect 12012 101276 12068 101332
rect 11418 101162 11474 101164
rect 11418 101110 11420 101162
rect 11420 101110 11472 101162
rect 11472 101110 11474 101162
rect 11418 101108 11474 101110
rect 11522 101162 11578 101164
rect 11522 101110 11524 101162
rect 11524 101110 11576 101162
rect 11576 101110 11578 101162
rect 11522 101108 11578 101110
rect 11626 101162 11682 101164
rect 11626 101110 11628 101162
rect 11628 101110 11680 101162
rect 11680 101110 11682 101162
rect 11626 101108 11682 101110
rect 11116 100940 11172 100996
rect 12236 100940 12292 100996
rect 11004 99260 11060 99316
rect 10556 99036 10612 99092
rect 11418 99594 11474 99596
rect 11418 99542 11420 99594
rect 11420 99542 11472 99594
rect 11472 99542 11474 99594
rect 11418 99540 11474 99542
rect 11522 99594 11578 99596
rect 11522 99542 11524 99594
rect 11524 99542 11576 99594
rect 11576 99542 11578 99594
rect 11522 99540 11578 99542
rect 11626 99594 11682 99596
rect 11626 99542 11628 99594
rect 11628 99542 11680 99594
rect 11680 99542 11682 99594
rect 11626 99540 11682 99542
rect 9996 97580 10052 97636
rect 8988 97244 9044 97300
rect 10332 98028 10388 98084
rect 9996 97132 10052 97188
rect 10108 97244 10164 97300
rect 8876 97074 8932 97076
rect 8876 97022 8878 97074
rect 8878 97022 8930 97074
rect 8930 97022 8932 97074
rect 8876 97020 8932 97022
rect 8764 96850 8820 96852
rect 8764 96798 8766 96850
rect 8766 96798 8818 96850
rect 8818 96798 8820 96850
rect 8764 96796 8820 96798
rect 7756 95788 7812 95844
rect 7644 95170 7700 95172
rect 7644 95118 7646 95170
rect 7646 95118 7698 95170
rect 7698 95118 7700 95170
rect 7644 95116 7700 95118
rect 7532 94892 7588 94948
rect 7644 94780 7700 94836
rect 7532 94274 7588 94276
rect 7532 94222 7534 94274
rect 7534 94222 7586 94274
rect 7586 94222 7588 94274
rect 7532 94220 7588 94222
rect 8016 95674 8072 95676
rect 8016 95622 8018 95674
rect 8018 95622 8070 95674
rect 8070 95622 8072 95674
rect 8016 95620 8072 95622
rect 8120 95674 8176 95676
rect 8120 95622 8122 95674
rect 8122 95622 8174 95674
rect 8174 95622 8176 95674
rect 8120 95620 8176 95622
rect 8224 95674 8280 95676
rect 8224 95622 8226 95674
rect 8226 95622 8278 95674
rect 8278 95622 8280 95674
rect 8428 95676 8484 95732
rect 8224 95620 8280 95622
rect 7868 95452 7924 95508
rect 8540 95564 8596 95620
rect 8092 94668 8148 94724
rect 8540 94220 8596 94276
rect 8016 94106 8072 94108
rect 8016 94054 8018 94106
rect 8018 94054 8070 94106
rect 8070 94054 8072 94106
rect 8016 94052 8072 94054
rect 8120 94106 8176 94108
rect 8120 94054 8122 94106
rect 8122 94054 8174 94106
rect 8174 94054 8176 94106
rect 8120 94052 8176 94054
rect 8224 94106 8280 94108
rect 8224 94054 8226 94106
rect 8226 94054 8278 94106
rect 8278 94054 8280 94106
rect 8224 94052 8280 94054
rect 8316 93884 8372 93940
rect 10332 96908 10388 96964
rect 10220 96572 10276 96628
rect 10220 95452 10276 95508
rect 9660 95228 9716 95284
rect 10444 97916 10500 97972
rect 10556 97132 10612 97188
rect 10780 96124 10836 96180
rect 10668 95676 10724 95732
rect 8764 93660 8820 93716
rect 8316 92876 8372 92932
rect 7532 92204 7588 92260
rect 8016 92538 8072 92540
rect 8016 92486 8018 92538
rect 8018 92486 8070 92538
rect 8070 92486 8072 92538
rect 8016 92484 8072 92486
rect 8120 92538 8176 92540
rect 8120 92486 8122 92538
rect 8122 92486 8174 92538
rect 8174 92486 8176 92538
rect 8120 92484 8176 92486
rect 8224 92538 8280 92540
rect 8224 92486 8226 92538
rect 8226 92486 8278 92538
rect 8278 92486 8280 92538
rect 8224 92484 8280 92486
rect 7420 91084 7476 91140
rect 7196 90748 7252 90804
rect 7532 90690 7588 90692
rect 7532 90638 7534 90690
rect 7534 90638 7586 90690
rect 7586 90638 7588 90690
rect 7532 90636 7588 90638
rect 6860 89180 6916 89236
rect 7196 89010 7252 89012
rect 7196 88958 7198 89010
rect 7198 88958 7250 89010
rect 7250 88958 7252 89010
rect 7196 88956 7252 88958
rect 8016 90970 8072 90972
rect 8016 90918 8018 90970
rect 8018 90918 8070 90970
rect 8070 90918 8072 90970
rect 8016 90916 8072 90918
rect 8120 90970 8176 90972
rect 8120 90918 8122 90970
rect 8122 90918 8174 90970
rect 8174 90918 8176 90970
rect 8120 90916 8176 90918
rect 8224 90970 8280 90972
rect 8224 90918 8226 90970
rect 8226 90918 8278 90970
rect 8278 90918 8280 90970
rect 8224 90916 8280 90918
rect 8428 90748 8484 90804
rect 8988 92316 9044 92372
rect 8764 90690 8820 90692
rect 8764 90638 8766 90690
rect 8766 90638 8818 90690
rect 8818 90638 8820 90690
rect 8764 90636 8820 90638
rect 8876 90524 8932 90580
rect 8092 90466 8148 90468
rect 8092 90414 8094 90466
rect 8094 90414 8146 90466
rect 8146 90414 8148 90466
rect 8092 90412 8148 90414
rect 8016 89402 8072 89404
rect 8016 89350 8018 89402
rect 8018 89350 8070 89402
rect 8070 89350 8072 89402
rect 8016 89348 8072 89350
rect 8120 89402 8176 89404
rect 8120 89350 8122 89402
rect 8122 89350 8174 89402
rect 8174 89350 8176 89402
rect 8120 89348 8176 89350
rect 8224 89402 8280 89404
rect 8224 89350 8226 89402
rect 8226 89350 8278 89402
rect 8278 89350 8280 89402
rect 8224 89348 8280 89350
rect 7644 88956 7700 89012
rect 7756 89180 7812 89236
rect 9212 90524 9268 90580
rect 9996 93884 10052 93940
rect 9548 93436 9604 93492
rect 9884 93436 9940 93492
rect 9884 92988 9940 93044
rect 9772 92258 9828 92260
rect 9772 92206 9774 92258
rect 9774 92206 9826 92258
rect 9826 92206 9828 92258
rect 9772 92204 9828 92206
rect 9660 90748 9716 90804
rect 8092 88898 8148 88900
rect 8092 88846 8094 88898
rect 8094 88846 8146 88898
rect 8146 88846 8148 88898
rect 8092 88844 8148 88846
rect 6748 87388 6804 87444
rect 6524 86770 6580 86772
rect 6524 86718 6526 86770
rect 6526 86718 6578 86770
rect 6578 86718 6580 86770
rect 6524 86716 6580 86718
rect 7532 86658 7588 86660
rect 7532 86606 7534 86658
rect 7534 86606 7586 86658
rect 7586 86606 7588 86658
rect 7532 86604 7588 86606
rect 7308 86098 7364 86100
rect 7308 86046 7310 86098
rect 7310 86046 7362 86098
rect 7362 86046 7364 86098
rect 7308 86044 7364 86046
rect 7084 85932 7140 85988
rect 6972 85762 7028 85764
rect 6972 85710 6974 85762
rect 6974 85710 7026 85762
rect 7026 85710 7028 85762
rect 6972 85708 7028 85710
rect 5740 84530 5796 84532
rect 5740 84478 5742 84530
rect 5742 84478 5794 84530
rect 5794 84478 5796 84530
rect 5740 84476 5796 84478
rect 5740 83356 5796 83412
rect 4844 82850 4900 82852
rect 4844 82798 4846 82850
rect 4846 82798 4898 82850
rect 4898 82798 4900 82850
rect 4844 82796 4900 82798
rect 5628 82796 5684 82852
rect 4614 82346 4670 82348
rect 4614 82294 4616 82346
rect 4616 82294 4668 82346
rect 4668 82294 4670 82346
rect 4614 82292 4670 82294
rect 4718 82346 4774 82348
rect 4718 82294 4720 82346
rect 4720 82294 4772 82346
rect 4772 82294 4774 82346
rect 4718 82292 4774 82294
rect 4822 82346 4878 82348
rect 4822 82294 4824 82346
rect 4824 82294 4876 82346
rect 4876 82294 4878 82346
rect 4822 82292 4878 82294
rect 6188 83410 6244 83412
rect 6188 83358 6190 83410
rect 6190 83358 6242 83410
rect 6242 83358 6244 83410
rect 6188 83356 6244 83358
rect 4844 81788 4900 81844
rect 5628 81842 5684 81844
rect 5628 81790 5630 81842
rect 5630 81790 5682 81842
rect 5682 81790 5684 81842
rect 5628 81788 5684 81790
rect 5068 81730 5124 81732
rect 5068 81678 5070 81730
rect 5070 81678 5122 81730
rect 5122 81678 5124 81730
rect 5068 81676 5124 81678
rect 5180 80892 5236 80948
rect 4614 80778 4670 80780
rect 4614 80726 4616 80778
rect 4616 80726 4668 80778
rect 4668 80726 4670 80778
rect 4614 80724 4670 80726
rect 4718 80778 4774 80780
rect 4718 80726 4720 80778
rect 4720 80726 4772 80778
rect 4772 80726 4774 80778
rect 4718 80724 4774 80726
rect 4822 80778 4878 80780
rect 4822 80726 4824 80778
rect 4824 80726 4876 80778
rect 4876 80726 4878 80778
rect 4822 80724 4878 80726
rect 5068 79996 5124 80052
rect 4614 79210 4670 79212
rect 4614 79158 4616 79210
rect 4616 79158 4668 79210
rect 4668 79158 4670 79210
rect 4614 79156 4670 79158
rect 4718 79210 4774 79212
rect 4718 79158 4720 79210
rect 4720 79158 4772 79210
rect 4772 79158 4774 79210
rect 4718 79156 4774 79158
rect 4822 79210 4878 79212
rect 4822 79158 4824 79210
rect 4824 79158 4876 79210
rect 4876 79158 4878 79210
rect 4822 79156 4878 79158
rect 4508 78876 4564 78932
rect 4060 78652 4116 78708
rect 4060 78204 4116 78260
rect 4844 78876 4900 78932
rect 5740 79996 5796 80052
rect 5068 78594 5124 78596
rect 5068 78542 5070 78594
rect 5070 78542 5122 78594
rect 5122 78542 5124 78594
rect 5068 78540 5124 78542
rect 5852 78652 5908 78708
rect 4614 77642 4670 77644
rect 4614 77590 4616 77642
rect 4616 77590 4668 77642
rect 4668 77590 4670 77642
rect 4614 77588 4670 77590
rect 4718 77642 4774 77644
rect 4718 77590 4720 77642
rect 4720 77590 4772 77642
rect 4772 77590 4774 77642
rect 4718 77588 4774 77590
rect 4822 77642 4878 77644
rect 4822 77590 4824 77642
rect 4824 77590 4876 77642
rect 4876 77590 4878 77642
rect 4822 77588 4878 77590
rect 6188 81058 6244 81060
rect 6188 81006 6190 81058
rect 6190 81006 6242 81058
rect 6242 81006 6244 81058
rect 6188 81004 6244 81006
rect 6524 83244 6580 83300
rect 6748 83356 6804 83412
rect 6748 82460 6804 82516
rect 6636 80892 6692 80948
rect 7308 81170 7364 81172
rect 7308 81118 7310 81170
rect 7310 81118 7362 81170
rect 7362 81118 7364 81170
rect 7308 81116 7364 81118
rect 6972 80892 7028 80948
rect 6076 80108 6132 80164
rect 6524 79996 6580 80052
rect 9772 90578 9828 90580
rect 9772 90526 9774 90578
rect 9774 90526 9826 90578
rect 9826 90526 9828 90578
rect 9772 90524 9828 90526
rect 9884 90412 9940 90468
rect 9436 88732 9492 88788
rect 9548 89906 9604 89908
rect 9548 89854 9550 89906
rect 9550 89854 9602 89906
rect 9602 89854 9604 89906
rect 9548 89852 9604 89854
rect 9100 88396 9156 88452
rect 10668 94444 10724 94500
rect 10780 94668 10836 94724
rect 10444 93884 10500 93940
rect 10332 93826 10388 93828
rect 10332 93774 10334 93826
rect 10334 93774 10386 93826
rect 10386 93774 10388 93826
rect 10332 93772 10388 93774
rect 10332 92988 10388 93044
rect 10220 92370 10276 92372
rect 10220 92318 10222 92370
rect 10222 92318 10274 92370
rect 10274 92318 10276 92370
rect 10220 92316 10276 92318
rect 11900 98924 11956 98980
rect 11788 98530 11844 98532
rect 11788 98478 11790 98530
rect 11790 98478 11842 98530
rect 11842 98478 11844 98530
rect 11788 98476 11844 98478
rect 11418 98026 11474 98028
rect 11418 97974 11420 98026
rect 11420 97974 11472 98026
rect 11472 97974 11474 98026
rect 11418 97972 11474 97974
rect 11522 98026 11578 98028
rect 11522 97974 11524 98026
rect 11524 97974 11576 98026
rect 11576 97974 11578 98026
rect 11522 97972 11578 97974
rect 11626 98026 11682 98028
rect 11626 97974 11628 98026
rect 11628 97974 11680 98026
rect 11680 97974 11682 98026
rect 11626 97972 11682 97974
rect 12012 97132 12068 97188
rect 11418 96458 11474 96460
rect 11418 96406 11420 96458
rect 11420 96406 11472 96458
rect 11472 96406 11474 96458
rect 11418 96404 11474 96406
rect 11522 96458 11578 96460
rect 11522 96406 11524 96458
rect 11524 96406 11576 96458
rect 11576 96406 11578 96458
rect 11522 96404 11578 96406
rect 11626 96458 11682 96460
rect 11626 96406 11628 96458
rect 11628 96406 11680 96458
rect 11680 96406 11682 96458
rect 11626 96404 11682 96406
rect 12012 96236 12068 96292
rect 12124 97020 12180 97076
rect 12348 98252 12404 98308
rect 13580 102396 13636 102452
rect 12572 102338 12628 102340
rect 12572 102286 12574 102338
rect 12574 102286 12626 102338
rect 12626 102286 12628 102338
rect 12572 102284 12628 102286
rect 13468 102284 13524 102340
rect 12796 101276 12852 101332
rect 12908 100940 12964 100996
rect 12572 100882 12628 100884
rect 12572 100830 12574 100882
rect 12574 100830 12626 100882
rect 12626 100830 12628 100882
rect 12572 100828 12628 100830
rect 13468 100770 13524 100772
rect 13468 100718 13470 100770
rect 13470 100718 13522 100770
rect 13522 100718 13524 100770
rect 13468 100716 13524 100718
rect 14252 103516 14308 103572
rect 14140 102284 14196 102340
rect 14028 100940 14084 100996
rect 12460 97020 12516 97076
rect 12572 99372 12628 99428
rect 12348 96348 12404 96404
rect 13580 99874 13636 99876
rect 13580 99822 13582 99874
rect 13582 99822 13634 99874
rect 13634 99822 13636 99874
rect 13580 99820 13636 99822
rect 14140 97522 14196 97524
rect 14140 97470 14142 97522
rect 14142 97470 14194 97522
rect 14194 97470 14196 97522
rect 14140 97468 14196 97470
rect 13468 97020 13524 97076
rect 13692 96962 13748 96964
rect 13692 96910 13694 96962
rect 13694 96910 13746 96962
rect 13746 96910 13748 96962
rect 13692 96908 13748 96910
rect 12572 96796 12628 96852
rect 12124 96178 12180 96180
rect 12124 96126 12126 96178
rect 12126 96126 12178 96178
rect 12178 96126 12180 96178
rect 12124 96124 12180 96126
rect 11788 96012 11844 96068
rect 11004 95900 11060 95956
rect 11900 95900 11956 95956
rect 11340 95676 11396 95732
rect 11116 95452 11172 95508
rect 11228 95340 11284 95396
rect 11340 95116 11396 95172
rect 11788 95058 11844 95060
rect 11788 95006 11790 95058
rect 11790 95006 11842 95058
rect 11842 95006 11844 95058
rect 11788 95004 11844 95006
rect 11418 94890 11474 94892
rect 11418 94838 11420 94890
rect 11420 94838 11472 94890
rect 11472 94838 11474 94890
rect 11418 94836 11474 94838
rect 11522 94890 11578 94892
rect 11522 94838 11524 94890
rect 11524 94838 11576 94890
rect 11576 94838 11578 94890
rect 11522 94836 11578 94838
rect 11626 94890 11682 94892
rect 11626 94838 11628 94890
rect 11628 94838 11680 94890
rect 11680 94838 11682 94890
rect 11626 94836 11682 94838
rect 11676 94556 11732 94612
rect 11340 94498 11396 94500
rect 11340 94446 11342 94498
rect 11342 94446 11394 94498
rect 11394 94446 11396 94498
rect 11340 94444 11396 94446
rect 11228 94332 11284 94388
rect 11116 93938 11172 93940
rect 11116 93886 11118 93938
rect 11118 93886 11170 93938
rect 11170 93886 11172 93938
rect 11116 93884 11172 93886
rect 11004 93100 11060 93156
rect 11418 93322 11474 93324
rect 11418 93270 11420 93322
rect 11420 93270 11472 93322
rect 11472 93270 11474 93322
rect 11418 93268 11474 93270
rect 11522 93322 11578 93324
rect 11522 93270 11524 93322
rect 11524 93270 11576 93322
rect 11576 93270 11578 93322
rect 11522 93268 11578 93270
rect 11626 93322 11682 93324
rect 11626 93270 11628 93322
rect 11628 93270 11680 93322
rect 11680 93270 11682 93322
rect 11626 93268 11682 93270
rect 11564 93154 11620 93156
rect 11564 93102 11566 93154
rect 11566 93102 11618 93154
rect 11618 93102 11620 93154
rect 11564 93100 11620 93102
rect 11340 93042 11396 93044
rect 11340 92990 11342 93042
rect 11342 92990 11394 93042
rect 11394 92990 11396 93042
rect 11340 92988 11396 92990
rect 12124 95954 12180 95956
rect 12124 95902 12126 95954
rect 12126 95902 12178 95954
rect 12178 95902 12180 95954
rect 12124 95900 12180 95902
rect 12348 95116 12404 95172
rect 13132 96460 13188 96516
rect 13356 96572 13412 96628
rect 13356 95788 13412 95844
rect 13244 95506 13300 95508
rect 13244 95454 13246 95506
rect 13246 95454 13298 95506
rect 13298 95454 13300 95506
rect 13244 95452 13300 95454
rect 13580 95282 13636 95284
rect 13580 95230 13582 95282
rect 13582 95230 13634 95282
rect 13634 95230 13636 95282
rect 13580 95228 13636 95230
rect 13692 95170 13748 95172
rect 13692 95118 13694 95170
rect 13694 95118 13746 95170
rect 13746 95118 13748 95170
rect 13692 95116 13748 95118
rect 13692 94780 13748 94836
rect 12124 93436 12180 93492
rect 14252 97244 14308 97300
rect 14140 97132 14196 97188
rect 14820 105082 14876 105084
rect 14820 105030 14822 105082
rect 14822 105030 14874 105082
rect 14874 105030 14876 105082
rect 14820 105028 14876 105030
rect 14924 105082 14980 105084
rect 14924 105030 14926 105082
rect 14926 105030 14978 105082
rect 14978 105030 14980 105082
rect 14924 105028 14980 105030
rect 15028 105082 15084 105084
rect 15028 105030 15030 105082
rect 15030 105030 15082 105082
rect 15082 105030 15084 105082
rect 15028 105028 15084 105030
rect 17276 114940 17332 114996
rect 17500 114828 17556 114884
rect 15708 112476 15764 112532
rect 16604 112530 16660 112532
rect 16604 112478 16606 112530
rect 16606 112478 16658 112530
rect 16658 112478 16660 112530
rect 16604 112476 16660 112478
rect 17388 112476 17444 112532
rect 17388 111746 17444 111748
rect 17388 111694 17390 111746
rect 17390 111694 17442 111746
rect 17442 111694 17444 111746
rect 17388 111692 17444 111694
rect 16716 110908 16772 110964
rect 17500 110962 17556 110964
rect 17500 110910 17502 110962
rect 17502 110910 17554 110962
rect 17554 110910 17556 110962
rect 17500 110908 17556 110910
rect 15372 109394 15428 109396
rect 15372 109342 15374 109394
rect 15374 109342 15426 109394
rect 15426 109342 15428 109394
rect 15372 109340 15428 109342
rect 15820 109394 15876 109396
rect 15820 109342 15822 109394
rect 15822 109342 15874 109394
rect 15874 109342 15876 109394
rect 15820 109340 15876 109342
rect 16716 109394 16772 109396
rect 16716 109342 16718 109394
rect 16718 109342 16770 109394
rect 16770 109342 16772 109394
rect 16716 109340 16772 109342
rect 16156 109282 16212 109284
rect 16156 109230 16158 109282
rect 16158 109230 16210 109282
rect 16210 109230 16212 109282
rect 16156 109228 16212 109230
rect 16940 108834 16996 108836
rect 16940 108782 16942 108834
rect 16942 108782 16994 108834
rect 16994 108782 16996 108834
rect 16940 108780 16996 108782
rect 16044 108498 16100 108500
rect 16044 108446 16046 108498
rect 16046 108446 16098 108498
rect 16098 108446 16100 108498
rect 16044 108444 16100 108446
rect 16940 108332 16996 108388
rect 16604 108220 16660 108276
rect 16268 107772 16324 107828
rect 16156 107042 16212 107044
rect 16156 106990 16158 107042
rect 16158 106990 16210 107042
rect 16210 106990 16212 107042
rect 16156 106988 16212 106990
rect 15260 104524 15316 104580
rect 15036 104300 15092 104356
rect 14700 104130 14756 104132
rect 14700 104078 14702 104130
rect 14702 104078 14754 104130
rect 14754 104078 14756 104130
rect 14700 104076 14756 104078
rect 15708 105868 15764 105924
rect 14812 103682 14868 103684
rect 14812 103630 14814 103682
rect 14814 103630 14866 103682
rect 14866 103630 14868 103682
rect 14812 103628 14868 103630
rect 14820 103514 14876 103516
rect 14820 103462 14822 103514
rect 14822 103462 14874 103514
rect 14874 103462 14876 103514
rect 14820 103460 14876 103462
rect 14924 103514 14980 103516
rect 14924 103462 14926 103514
rect 14926 103462 14978 103514
rect 14978 103462 14980 103514
rect 14924 103460 14980 103462
rect 15028 103514 15084 103516
rect 15028 103462 15030 103514
rect 15030 103462 15082 103514
rect 15082 103462 15084 103514
rect 15028 103460 15084 103462
rect 14924 103122 14980 103124
rect 14924 103070 14926 103122
rect 14926 103070 14978 103122
rect 14978 103070 14980 103122
rect 14924 103068 14980 103070
rect 14820 101946 14876 101948
rect 14820 101894 14822 101946
rect 14822 101894 14874 101946
rect 14874 101894 14876 101946
rect 14820 101892 14876 101894
rect 14924 101946 14980 101948
rect 14924 101894 14926 101946
rect 14926 101894 14978 101946
rect 14978 101894 14980 101946
rect 14924 101892 14980 101894
rect 15028 101946 15084 101948
rect 15028 101894 15030 101946
rect 15030 101894 15082 101946
rect 15082 101894 15084 101946
rect 15028 101892 15084 101894
rect 14588 100716 14644 100772
rect 15484 100658 15540 100660
rect 15484 100606 15486 100658
rect 15486 100606 15538 100658
rect 15538 100606 15540 100658
rect 15484 100604 15540 100606
rect 14820 100378 14876 100380
rect 14820 100326 14822 100378
rect 14822 100326 14874 100378
rect 14874 100326 14876 100378
rect 14820 100324 14876 100326
rect 14924 100378 14980 100380
rect 14924 100326 14926 100378
rect 14926 100326 14978 100378
rect 14978 100326 14980 100378
rect 14924 100324 14980 100326
rect 15028 100378 15084 100380
rect 15028 100326 15030 100378
rect 15030 100326 15082 100378
rect 15082 100326 15084 100378
rect 15028 100324 15084 100326
rect 15484 99314 15540 99316
rect 15484 99262 15486 99314
rect 15486 99262 15538 99314
rect 15538 99262 15540 99314
rect 15484 99260 15540 99262
rect 15148 99036 15204 99092
rect 14820 98810 14876 98812
rect 14820 98758 14822 98810
rect 14822 98758 14874 98810
rect 14874 98758 14876 98810
rect 14820 98756 14876 98758
rect 14924 98810 14980 98812
rect 14924 98758 14926 98810
rect 14926 98758 14978 98810
rect 14978 98758 14980 98810
rect 14924 98756 14980 98758
rect 15028 98810 15084 98812
rect 15028 98758 15030 98810
rect 15030 98758 15082 98810
rect 15082 98758 15084 98810
rect 15028 98756 15084 98758
rect 15484 99036 15540 99092
rect 15036 97692 15092 97748
rect 14700 97634 14756 97636
rect 14700 97582 14702 97634
rect 14702 97582 14754 97634
rect 14754 97582 14756 97634
rect 14700 97580 14756 97582
rect 14364 97132 14420 97188
rect 14588 97468 14644 97524
rect 14028 96962 14084 96964
rect 14028 96910 14030 96962
rect 14030 96910 14082 96962
rect 14082 96910 14084 96962
rect 14028 96908 14084 96910
rect 13916 96236 13972 96292
rect 14028 96348 14084 96404
rect 14252 96348 14308 96404
rect 14364 95788 14420 95844
rect 13916 94386 13972 94388
rect 13916 94334 13918 94386
rect 13918 94334 13970 94386
rect 13970 94334 13972 94386
rect 13916 94332 13972 94334
rect 14140 95228 14196 95284
rect 13916 94108 13972 94164
rect 13468 93772 13524 93828
rect 12460 93714 12516 93716
rect 12460 93662 12462 93714
rect 12462 93662 12514 93714
rect 12514 93662 12516 93714
rect 12460 93660 12516 93662
rect 13132 93714 13188 93716
rect 13132 93662 13134 93714
rect 13134 93662 13186 93714
rect 13186 93662 13188 93714
rect 13132 93660 13188 93662
rect 13356 93436 13412 93492
rect 13356 92764 13412 92820
rect 11900 92706 11956 92708
rect 11900 92654 11902 92706
rect 11902 92654 11954 92706
rect 11954 92654 11956 92706
rect 11900 92652 11956 92654
rect 10892 92316 10948 92372
rect 12348 92316 12404 92372
rect 10444 92204 10500 92260
rect 10108 90748 10164 90804
rect 10556 90748 10612 90804
rect 10444 90524 10500 90580
rect 10332 89852 10388 89908
rect 10108 89010 10164 89012
rect 10108 88958 10110 89010
rect 10110 88958 10162 89010
rect 10162 88958 10164 89010
rect 10108 88956 10164 88958
rect 10892 90690 10948 90692
rect 10892 90638 10894 90690
rect 10894 90638 10946 90690
rect 10946 90638 10948 90690
rect 10892 90636 10948 90638
rect 11418 91754 11474 91756
rect 11418 91702 11420 91754
rect 11420 91702 11472 91754
rect 11472 91702 11474 91754
rect 11418 91700 11474 91702
rect 11522 91754 11578 91756
rect 11522 91702 11524 91754
rect 11524 91702 11576 91754
rect 11576 91702 11578 91754
rect 11522 91700 11578 91702
rect 11626 91754 11682 91756
rect 11626 91702 11628 91754
rect 11628 91702 11680 91754
rect 11680 91702 11682 91754
rect 11626 91700 11682 91702
rect 11452 90802 11508 90804
rect 11452 90750 11454 90802
rect 11454 90750 11506 90802
rect 11506 90750 11508 90802
rect 11452 90748 11508 90750
rect 11228 90524 11284 90580
rect 11418 90186 11474 90188
rect 11418 90134 11420 90186
rect 11420 90134 11472 90186
rect 11472 90134 11474 90186
rect 11418 90132 11474 90134
rect 11522 90186 11578 90188
rect 11522 90134 11524 90186
rect 11524 90134 11576 90186
rect 11576 90134 11578 90186
rect 11522 90132 11578 90134
rect 11626 90186 11682 90188
rect 11626 90134 11628 90186
rect 11628 90134 11680 90186
rect 11680 90134 11682 90186
rect 11626 90132 11682 90134
rect 11900 90524 11956 90580
rect 12012 90636 12068 90692
rect 12012 90412 12068 90468
rect 11788 89740 11844 89796
rect 11116 88844 11172 88900
rect 11418 88618 11474 88620
rect 11418 88566 11420 88618
rect 11420 88566 11472 88618
rect 11472 88566 11474 88618
rect 11418 88564 11474 88566
rect 11522 88618 11578 88620
rect 11522 88566 11524 88618
rect 11524 88566 11576 88618
rect 11576 88566 11578 88618
rect 11522 88564 11578 88566
rect 11626 88618 11682 88620
rect 11626 88566 11628 88618
rect 11628 88566 11680 88618
rect 11680 88566 11682 88618
rect 11626 88564 11682 88566
rect 7756 88114 7812 88116
rect 7756 88062 7758 88114
rect 7758 88062 7810 88114
rect 7810 88062 7812 88114
rect 7756 88060 7812 88062
rect 9212 88114 9268 88116
rect 9212 88062 9214 88114
rect 9214 88062 9266 88114
rect 9266 88062 9268 88114
rect 9212 88060 9268 88062
rect 7980 87948 8036 88004
rect 8876 87948 8932 88004
rect 8016 87834 8072 87836
rect 8016 87782 8018 87834
rect 8018 87782 8070 87834
rect 8070 87782 8072 87834
rect 8016 87780 8072 87782
rect 8120 87834 8176 87836
rect 8120 87782 8122 87834
rect 8122 87782 8174 87834
rect 8174 87782 8176 87834
rect 8120 87780 8176 87782
rect 8224 87834 8280 87836
rect 8224 87782 8226 87834
rect 8226 87782 8278 87834
rect 8278 87782 8280 87834
rect 8224 87780 8280 87782
rect 7868 87276 7924 87332
rect 12348 88060 12404 88116
rect 9660 87276 9716 87332
rect 10108 87276 10164 87332
rect 8652 86380 8708 86436
rect 8016 86266 8072 86268
rect 8016 86214 8018 86266
rect 8018 86214 8070 86266
rect 8070 86214 8072 86266
rect 8016 86212 8072 86214
rect 8120 86266 8176 86268
rect 8120 86214 8122 86266
rect 8122 86214 8174 86266
rect 8174 86214 8176 86266
rect 8120 86212 8176 86214
rect 8224 86266 8280 86268
rect 8224 86214 8226 86266
rect 8226 86214 8278 86266
rect 8278 86214 8280 86266
rect 8224 86212 8280 86214
rect 8652 85986 8708 85988
rect 8652 85934 8654 85986
rect 8654 85934 8706 85986
rect 8706 85934 8708 85986
rect 8652 85932 8708 85934
rect 7756 85874 7812 85876
rect 7756 85822 7758 85874
rect 7758 85822 7810 85874
rect 7810 85822 7812 85874
rect 7756 85820 7812 85822
rect 8316 85708 8372 85764
rect 8016 84698 8072 84700
rect 8016 84646 8018 84698
rect 8018 84646 8070 84698
rect 8070 84646 8072 84698
rect 8016 84644 8072 84646
rect 8120 84698 8176 84700
rect 8120 84646 8122 84698
rect 8122 84646 8174 84698
rect 8174 84646 8176 84698
rect 8120 84644 8176 84646
rect 8224 84698 8280 84700
rect 8224 84646 8226 84698
rect 8226 84646 8278 84698
rect 8278 84646 8280 84698
rect 8224 84644 8280 84646
rect 8988 86716 9044 86772
rect 11418 87050 11474 87052
rect 11418 86998 11420 87050
rect 11420 86998 11472 87050
rect 11472 86998 11474 87050
rect 11418 86996 11474 86998
rect 11522 87050 11578 87052
rect 11522 86998 11524 87050
rect 11524 86998 11576 87050
rect 11576 86998 11578 87050
rect 11522 86996 11578 86998
rect 11626 87050 11682 87052
rect 11626 86998 11628 87050
rect 11628 86998 11680 87050
rect 11680 86998 11682 87050
rect 11626 86996 11682 86998
rect 10108 86716 10164 86772
rect 11228 86716 11284 86772
rect 9212 86546 9268 86548
rect 9212 86494 9214 86546
rect 9214 86494 9266 86546
rect 9266 86494 9268 86546
rect 9212 86492 9268 86494
rect 10892 86546 10948 86548
rect 10892 86494 10894 86546
rect 10894 86494 10946 86546
rect 10946 86494 10948 86546
rect 10892 86492 10948 86494
rect 12236 86658 12292 86660
rect 12236 86606 12238 86658
rect 12238 86606 12290 86658
rect 12290 86606 12292 86658
rect 12236 86604 12292 86606
rect 8988 86380 9044 86436
rect 9548 86434 9604 86436
rect 9548 86382 9550 86434
rect 9550 86382 9602 86434
rect 9602 86382 9604 86434
rect 9548 86380 9604 86382
rect 9660 85932 9716 85988
rect 9772 86044 9828 86100
rect 10780 86434 10836 86436
rect 10780 86382 10782 86434
rect 10782 86382 10834 86434
rect 10834 86382 10836 86434
rect 10780 86380 10836 86382
rect 11004 85820 11060 85876
rect 8876 85596 8932 85652
rect 8988 84530 9044 84532
rect 8988 84478 8990 84530
rect 8990 84478 9042 84530
rect 9042 84478 9044 84530
rect 8988 84476 9044 84478
rect 10220 84418 10276 84420
rect 10220 84366 10222 84418
rect 10222 84366 10274 84418
rect 10274 84366 10276 84418
rect 10220 84364 10276 84366
rect 10332 84476 10388 84532
rect 9884 84252 9940 84308
rect 8764 84028 8820 84084
rect 7756 81900 7812 81956
rect 7644 81788 7700 81844
rect 7756 81004 7812 81060
rect 8016 83130 8072 83132
rect 8016 83078 8018 83130
rect 8018 83078 8070 83130
rect 8070 83078 8072 83130
rect 8016 83076 8072 83078
rect 8120 83130 8176 83132
rect 8120 83078 8122 83130
rect 8122 83078 8174 83130
rect 8174 83078 8176 83130
rect 8120 83076 8176 83078
rect 8224 83130 8280 83132
rect 8224 83078 8226 83130
rect 8226 83078 8278 83130
rect 8278 83078 8280 83130
rect 8224 83076 8280 83078
rect 10108 84028 10164 84084
rect 8092 81788 8148 81844
rect 9548 81900 9604 81956
rect 8016 81562 8072 81564
rect 8016 81510 8018 81562
rect 8018 81510 8070 81562
rect 8070 81510 8072 81562
rect 8016 81508 8072 81510
rect 8120 81562 8176 81564
rect 8120 81510 8122 81562
rect 8122 81510 8174 81562
rect 8174 81510 8176 81562
rect 8120 81508 8176 81510
rect 8224 81562 8280 81564
rect 8224 81510 8226 81562
rect 8226 81510 8278 81562
rect 8278 81510 8280 81562
rect 8224 81508 8280 81510
rect 7868 80444 7924 80500
rect 9436 81340 9492 81396
rect 8016 79994 8072 79996
rect 8016 79942 8018 79994
rect 8018 79942 8070 79994
rect 8070 79942 8072 79994
rect 8016 79940 8072 79942
rect 8120 79994 8176 79996
rect 8120 79942 8122 79994
rect 8122 79942 8174 79994
rect 8174 79942 8176 79994
rect 8120 79940 8176 79942
rect 8224 79994 8280 79996
rect 8224 79942 8226 79994
rect 8226 79942 8278 79994
rect 8278 79942 8280 79994
rect 8224 79940 8280 79942
rect 6188 78818 6244 78820
rect 6188 78766 6190 78818
rect 6190 78766 6242 78818
rect 6242 78766 6244 78818
rect 6188 78764 6244 78766
rect 6412 78540 6468 78596
rect 6860 78594 6916 78596
rect 6860 78542 6862 78594
rect 6862 78542 6914 78594
rect 6914 78542 6916 78594
rect 6860 78540 6916 78542
rect 5964 78092 6020 78148
rect 4060 76412 4116 76468
rect 4620 76636 4676 76692
rect 5068 76524 5124 76580
rect 5292 76466 5348 76468
rect 5292 76414 5294 76466
rect 5294 76414 5346 76466
rect 5346 76414 5348 76466
rect 5292 76412 5348 76414
rect 4614 76074 4670 76076
rect 4614 76022 4616 76074
rect 4616 76022 4668 76074
rect 4668 76022 4670 76074
rect 4614 76020 4670 76022
rect 4718 76074 4774 76076
rect 4718 76022 4720 76074
rect 4720 76022 4772 76074
rect 4772 76022 4774 76074
rect 4718 76020 4774 76022
rect 4822 76074 4878 76076
rect 4822 76022 4824 76074
rect 4824 76022 4876 76074
rect 4876 76022 4878 76074
rect 4822 76020 4878 76022
rect 4956 75682 5012 75684
rect 4956 75630 4958 75682
rect 4958 75630 5010 75682
rect 5010 75630 5012 75682
rect 4956 75628 5012 75630
rect 4172 74786 4228 74788
rect 4172 74734 4174 74786
rect 4174 74734 4226 74786
rect 4226 74734 4228 74786
rect 4172 74732 4228 74734
rect 4060 74284 4116 74340
rect 4614 74506 4670 74508
rect 4614 74454 4616 74506
rect 4616 74454 4668 74506
rect 4668 74454 4670 74506
rect 4614 74452 4670 74454
rect 4718 74506 4774 74508
rect 4718 74454 4720 74506
rect 4720 74454 4772 74506
rect 4772 74454 4774 74506
rect 4718 74452 4774 74454
rect 4822 74506 4878 74508
rect 4822 74454 4824 74506
rect 4824 74454 4876 74506
rect 4876 74454 4878 74506
rect 4822 74452 4878 74454
rect 5292 74786 5348 74788
rect 5292 74734 5294 74786
rect 5294 74734 5346 74786
rect 5346 74734 5348 74786
rect 5292 74732 5348 74734
rect 5516 76300 5572 76356
rect 7868 78764 7924 78820
rect 8316 78876 8372 78932
rect 7868 78594 7924 78596
rect 7868 78542 7870 78594
rect 7870 78542 7922 78594
rect 7922 78542 7924 78594
rect 7868 78540 7924 78542
rect 8016 78426 8072 78428
rect 8016 78374 8018 78426
rect 8018 78374 8070 78426
rect 8070 78374 8072 78426
rect 8016 78372 8072 78374
rect 8120 78426 8176 78428
rect 8120 78374 8122 78426
rect 8122 78374 8174 78426
rect 8174 78374 8176 78426
rect 8120 78372 8176 78374
rect 8224 78426 8280 78428
rect 8224 78374 8226 78426
rect 8226 78374 8278 78426
rect 8278 78374 8280 78426
rect 8224 78372 8280 78374
rect 8764 78428 8820 78484
rect 7868 78034 7924 78036
rect 7868 77982 7870 78034
rect 7870 77982 7922 78034
rect 7922 77982 7924 78034
rect 7868 77980 7924 77982
rect 6972 77644 7028 77700
rect 8540 77644 8596 77700
rect 8016 76858 8072 76860
rect 8016 76806 8018 76858
rect 8018 76806 8070 76858
rect 8070 76806 8072 76858
rect 8016 76804 8072 76806
rect 8120 76858 8176 76860
rect 8120 76806 8122 76858
rect 8122 76806 8174 76858
rect 8174 76806 8176 76858
rect 8120 76804 8176 76806
rect 8224 76858 8280 76860
rect 8224 76806 8226 76858
rect 8226 76806 8278 76858
rect 8278 76806 8280 76858
rect 8224 76804 8280 76806
rect 6076 76524 6132 76580
rect 5740 76354 5796 76356
rect 5740 76302 5742 76354
rect 5742 76302 5794 76354
rect 5794 76302 5796 76354
rect 5740 76300 5796 76302
rect 4844 73890 4900 73892
rect 4844 73838 4846 73890
rect 4846 73838 4898 73890
rect 4898 73838 4900 73890
rect 4844 73836 4900 73838
rect 4614 72938 4670 72940
rect 4614 72886 4616 72938
rect 4616 72886 4668 72938
rect 4668 72886 4670 72938
rect 4614 72884 4670 72886
rect 4718 72938 4774 72940
rect 4718 72886 4720 72938
rect 4720 72886 4772 72938
rect 4772 72886 4774 72938
rect 4718 72884 4774 72886
rect 4822 72938 4878 72940
rect 4822 72886 4824 72938
rect 4824 72886 4876 72938
rect 4876 72886 4878 72938
rect 4822 72884 4878 72886
rect 4396 72492 4452 72548
rect 4172 71820 4228 71876
rect 3948 71650 4004 71652
rect 3948 71598 3950 71650
rect 3950 71598 4002 71650
rect 4002 71598 4004 71650
rect 3948 71596 4004 71598
rect 3836 71036 3892 71092
rect 3948 70754 4004 70756
rect 3948 70702 3950 70754
rect 3950 70702 4002 70754
rect 4002 70702 4004 70754
rect 3948 70700 4004 70702
rect 4172 70700 4228 70756
rect 3500 68796 3556 68852
rect 2492 68626 2548 68628
rect 2492 68574 2494 68626
rect 2494 68574 2546 68626
rect 2546 68574 2548 68626
rect 2492 68572 2548 68574
rect 2828 68626 2884 68628
rect 2828 68574 2830 68626
rect 2830 68574 2882 68626
rect 2882 68574 2884 68626
rect 2828 68572 2884 68574
rect 3388 68626 3444 68628
rect 3388 68574 3390 68626
rect 3390 68574 3442 68626
rect 3442 68574 3444 68626
rect 3388 68572 3444 68574
rect 3500 68348 3556 68404
rect 3948 68402 4004 68404
rect 3948 68350 3950 68402
rect 3950 68350 4002 68402
rect 4002 68350 4004 68402
rect 3948 68348 4004 68350
rect 2716 67116 2772 67172
rect 2380 66834 2436 66836
rect 2380 66782 2382 66834
rect 2382 66782 2434 66834
rect 2434 66782 2436 66834
rect 2380 66780 2436 66782
rect 1708 66556 1764 66612
rect 1708 64594 1764 64596
rect 1708 64542 1710 64594
rect 1710 64542 1762 64594
rect 1762 64542 1764 64594
rect 1708 64540 1764 64542
rect 1932 64540 1988 64596
rect 2492 65490 2548 65492
rect 2492 65438 2494 65490
rect 2494 65438 2546 65490
rect 2546 65438 2548 65490
rect 2492 65436 2548 65438
rect 2828 65772 2884 65828
rect 3052 65602 3108 65604
rect 3052 65550 3054 65602
rect 3054 65550 3106 65602
rect 3106 65550 3108 65602
rect 3052 65548 3108 65550
rect 2268 64540 2324 64596
rect 2044 64482 2100 64484
rect 2044 64430 2046 64482
rect 2046 64430 2098 64482
rect 2098 64430 2100 64482
rect 2044 64428 2100 64430
rect 1820 63922 1876 63924
rect 1820 63870 1822 63922
rect 1822 63870 1874 63922
rect 1874 63870 1876 63922
rect 1820 63868 1876 63870
rect 3052 64594 3108 64596
rect 3052 64542 3054 64594
rect 3054 64542 3106 64594
rect 3106 64542 3108 64594
rect 3052 64540 3108 64542
rect 2828 64482 2884 64484
rect 2828 64430 2830 64482
rect 2830 64430 2882 64482
rect 2882 64430 2884 64482
rect 2828 64428 2884 64430
rect 2716 63922 2772 63924
rect 2716 63870 2718 63922
rect 2718 63870 2770 63922
rect 2770 63870 2772 63922
rect 2716 63868 2772 63870
rect 1708 61180 1764 61236
rect 2044 61458 2100 61460
rect 2044 61406 2046 61458
rect 2046 61406 2098 61458
rect 2098 61406 2100 61458
rect 2044 61404 2100 61406
rect 2380 61292 2436 61348
rect 3052 63756 3108 63812
rect 3836 66946 3892 66948
rect 3836 66894 3838 66946
rect 3838 66894 3890 66946
rect 3890 66894 3892 66946
rect 3836 66892 3892 66894
rect 3500 65772 3556 65828
rect 3276 65548 3332 65604
rect 3836 65324 3892 65380
rect 3164 62972 3220 63028
rect 3276 64092 3332 64148
rect 3724 63868 3780 63924
rect 3500 63756 3556 63812
rect 3724 63196 3780 63252
rect 3500 61740 3556 61796
rect 2716 61292 2772 61348
rect 2492 61180 2548 61236
rect 2156 60620 2212 60676
rect 1708 58492 1764 58548
rect 2044 58380 2100 58436
rect 3276 61404 3332 61460
rect 2604 60562 2660 60564
rect 2604 60510 2606 60562
rect 2606 60510 2658 60562
rect 2658 60510 2660 60562
rect 2604 60508 2660 60510
rect 3948 64428 4004 64484
rect 4172 68348 4228 68404
rect 4508 71820 4564 71876
rect 4956 72492 5012 72548
rect 5068 72434 5124 72436
rect 5068 72382 5070 72434
rect 5070 72382 5122 72434
rect 5122 72382 5124 72434
rect 5068 72380 5124 72382
rect 4508 71596 4564 71652
rect 5180 71596 5236 71652
rect 4614 71370 4670 71372
rect 4614 71318 4616 71370
rect 4616 71318 4668 71370
rect 4668 71318 4670 71370
rect 4614 71316 4670 71318
rect 4718 71370 4774 71372
rect 4718 71318 4720 71370
rect 4720 71318 4772 71370
rect 4772 71318 4774 71370
rect 4718 71316 4774 71318
rect 4822 71370 4878 71372
rect 4822 71318 4824 71370
rect 4824 71318 4876 71370
rect 4876 71318 4878 71370
rect 4822 71316 4878 71318
rect 4508 70700 4564 70756
rect 5068 70588 5124 70644
rect 5180 70476 5236 70532
rect 4614 69802 4670 69804
rect 4614 69750 4616 69802
rect 4616 69750 4668 69802
rect 4668 69750 4670 69802
rect 4614 69748 4670 69750
rect 4718 69802 4774 69804
rect 4718 69750 4720 69802
rect 4720 69750 4772 69802
rect 4772 69750 4774 69802
rect 4718 69748 4774 69750
rect 4822 69802 4878 69804
rect 4822 69750 4824 69802
rect 4824 69750 4876 69802
rect 4876 69750 4878 69802
rect 4822 69748 4878 69750
rect 4396 68514 4452 68516
rect 4396 68462 4398 68514
rect 4398 68462 4450 68514
rect 4450 68462 4452 68514
rect 4396 68460 4452 68462
rect 4614 68234 4670 68236
rect 4614 68182 4616 68234
rect 4616 68182 4668 68234
rect 4668 68182 4670 68234
rect 4614 68180 4670 68182
rect 4718 68234 4774 68236
rect 4718 68182 4720 68234
rect 4720 68182 4772 68234
rect 4772 68182 4774 68234
rect 4718 68180 4774 68182
rect 4822 68234 4878 68236
rect 4822 68182 4824 68234
rect 4824 68182 4876 68234
rect 4876 68182 4878 68234
rect 4822 68180 4878 68182
rect 4956 67900 5012 67956
rect 4732 67058 4788 67060
rect 4732 67006 4734 67058
rect 4734 67006 4786 67058
rect 4786 67006 4788 67058
rect 4732 67004 4788 67006
rect 4614 66666 4670 66668
rect 4614 66614 4616 66666
rect 4616 66614 4668 66666
rect 4668 66614 4670 66666
rect 4614 66612 4670 66614
rect 4718 66666 4774 66668
rect 4718 66614 4720 66666
rect 4720 66614 4772 66666
rect 4772 66614 4774 66666
rect 4718 66612 4774 66614
rect 4822 66666 4878 66668
rect 4822 66614 4824 66666
rect 4824 66614 4876 66666
rect 4876 66614 4878 66666
rect 4822 66612 4878 66614
rect 4396 65602 4452 65604
rect 4396 65550 4398 65602
rect 4398 65550 4450 65602
rect 4450 65550 4452 65602
rect 4396 65548 4452 65550
rect 4620 65324 4676 65380
rect 4284 65212 4340 65268
rect 4614 65098 4670 65100
rect 4614 65046 4616 65098
rect 4616 65046 4668 65098
rect 4668 65046 4670 65098
rect 4614 65044 4670 65046
rect 4718 65098 4774 65100
rect 4718 65046 4720 65098
rect 4720 65046 4772 65098
rect 4772 65046 4774 65098
rect 4718 65044 4774 65046
rect 4822 65098 4878 65100
rect 4822 65046 4824 65098
rect 4824 65046 4876 65098
rect 4876 65046 4878 65098
rect 4822 65044 4878 65046
rect 4284 64764 4340 64820
rect 4172 64706 4228 64708
rect 4172 64654 4174 64706
rect 4174 64654 4226 64706
rect 4226 64654 4228 64706
rect 4172 64652 4228 64654
rect 4172 64092 4228 64148
rect 4172 61346 4228 61348
rect 4172 61294 4174 61346
rect 4174 61294 4226 61346
rect 4226 61294 4228 61346
rect 4172 61292 4228 61294
rect 3724 60674 3780 60676
rect 3724 60622 3726 60674
rect 3726 60622 3778 60674
rect 3778 60622 3780 60674
rect 3724 60620 3780 60622
rect 3388 60562 3444 60564
rect 3388 60510 3390 60562
rect 3390 60510 3442 60562
rect 3442 60510 3444 60562
rect 3388 60508 3444 60510
rect 3836 60508 3892 60564
rect 3276 59836 3332 59892
rect 2380 58604 2436 58660
rect 2940 58658 2996 58660
rect 2940 58606 2942 58658
rect 2942 58606 2994 58658
rect 2994 58606 2996 58658
rect 2940 58604 2996 58606
rect 2492 58492 2548 58548
rect 2828 58492 2884 58548
rect 2268 58210 2324 58212
rect 2268 58158 2270 58210
rect 2270 58158 2322 58210
rect 2322 58158 2324 58210
rect 2268 58156 2324 58158
rect 1820 57820 1876 57876
rect 3724 58658 3780 58660
rect 3724 58606 3726 58658
rect 3726 58606 3778 58658
rect 3778 58606 3780 58658
rect 3724 58604 3780 58606
rect 3612 57260 3668 57316
rect 3164 57036 3220 57092
rect 3500 57090 3556 57092
rect 3500 57038 3502 57090
rect 3502 57038 3554 57090
rect 3554 57038 3556 57090
rect 3500 57036 3556 57038
rect 3612 56754 3668 56756
rect 3612 56702 3614 56754
rect 3614 56702 3666 56754
rect 3666 56702 3668 56754
rect 3612 56700 3668 56702
rect 3500 56588 3556 56644
rect 3388 56364 3444 56420
rect 1708 55804 1764 55860
rect 2156 54514 2212 54516
rect 2156 54462 2158 54514
rect 2158 54462 2210 54514
rect 2210 54462 2212 54514
rect 2156 54460 2212 54462
rect 1820 53676 1876 53732
rect 2492 55804 2548 55860
rect 2828 54626 2884 54628
rect 2828 54574 2830 54626
rect 2830 54574 2882 54626
rect 2882 54574 2884 54626
rect 2828 54572 2884 54574
rect 3276 54460 3332 54516
rect 3612 56194 3668 56196
rect 3612 56142 3614 56194
rect 3614 56142 3666 56194
rect 3666 56142 3668 56194
rect 3612 56140 3668 56142
rect 3836 58210 3892 58212
rect 3836 58158 3838 58210
rect 3838 58158 3890 58210
rect 3890 58158 3892 58210
rect 3836 58156 3892 58158
rect 3836 56194 3892 56196
rect 3836 56142 3838 56194
rect 3838 56142 3890 56194
rect 3890 56142 3892 56194
rect 3836 56140 3892 56142
rect 4172 58716 4228 58772
rect 4060 58322 4116 58324
rect 4060 58270 4062 58322
rect 4062 58270 4114 58322
rect 4114 58270 4116 58322
rect 4060 58268 4116 58270
rect 4060 56754 4116 56756
rect 4060 56702 4062 56754
rect 4062 56702 4114 56754
rect 4114 56702 4116 56754
rect 4060 56700 4116 56702
rect 4620 64594 4676 64596
rect 4620 64542 4622 64594
rect 4622 64542 4674 64594
rect 4674 64542 4676 64594
rect 4620 64540 4676 64542
rect 4508 63922 4564 63924
rect 4508 63870 4510 63922
rect 4510 63870 4562 63922
rect 4562 63870 4564 63922
rect 4508 63868 4564 63870
rect 4614 63530 4670 63532
rect 4614 63478 4616 63530
rect 4616 63478 4668 63530
rect 4668 63478 4670 63530
rect 4614 63476 4670 63478
rect 4718 63530 4774 63532
rect 4718 63478 4720 63530
rect 4720 63478 4772 63530
rect 4772 63478 4774 63530
rect 4718 63476 4774 63478
rect 4822 63530 4878 63532
rect 4822 63478 4824 63530
rect 4824 63478 4876 63530
rect 4876 63478 4878 63530
rect 4822 63476 4878 63478
rect 4620 63250 4676 63252
rect 4620 63198 4622 63250
rect 4622 63198 4674 63250
rect 4674 63198 4676 63250
rect 4620 63196 4676 63198
rect 5180 67730 5236 67732
rect 5180 67678 5182 67730
rect 5182 67678 5234 67730
rect 5234 67678 5236 67730
rect 5180 67676 5236 67678
rect 5180 66162 5236 66164
rect 5180 66110 5182 66162
rect 5182 66110 5234 66162
rect 5234 66110 5236 66162
rect 5180 66108 5236 66110
rect 5068 63420 5124 63476
rect 5180 63868 5236 63924
rect 4956 62860 5012 62916
rect 4614 61962 4670 61964
rect 4614 61910 4616 61962
rect 4616 61910 4668 61962
rect 4668 61910 4670 61962
rect 4614 61908 4670 61910
rect 4718 61962 4774 61964
rect 4718 61910 4720 61962
rect 4720 61910 4772 61962
rect 4772 61910 4774 61962
rect 4718 61908 4774 61910
rect 4822 61962 4878 61964
rect 4822 61910 4824 61962
rect 4824 61910 4876 61962
rect 4876 61910 4878 61962
rect 4822 61908 4878 61910
rect 4620 61682 4676 61684
rect 4620 61630 4622 61682
rect 4622 61630 4674 61682
rect 4674 61630 4676 61682
rect 4620 61628 4676 61630
rect 4396 60508 4452 60564
rect 4614 60394 4670 60396
rect 4614 60342 4616 60394
rect 4616 60342 4668 60394
rect 4668 60342 4670 60394
rect 4614 60340 4670 60342
rect 4718 60394 4774 60396
rect 4718 60342 4720 60394
rect 4720 60342 4772 60394
rect 4772 60342 4774 60394
rect 4718 60340 4774 60342
rect 4822 60394 4878 60396
rect 4822 60342 4824 60394
rect 4824 60342 4876 60394
rect 4876 60342 4878 60394
rect 4822 60340 4878 60342
rect 4620 59836 4676 59892
rect 4620 58940 4676 58996
rect 4614 58826 4670 58828
rect 4614 58774 4616 58826
rect 4616 58774 4668 58826
rect 4668 58774 4670 58826
rect 4614 58772 4670 58774
rect 4718 58826 4774 58828
rect 4718 58774 4720 58826
rect 4720 58774 4772 58826
rect 4772 58774 4774 58826
rect 4718 58772 4774 58774
rect 4822 58826 4878 58828
rect 4822 58774 4824 58826
rect 4824 58774 4876 58826
rect 4876 58774 4878 58826
rect 4822 58772 4878 58774
rect 4620 58546 4676 58548
rect 4620 58494 4622 58546
rect 4622 58494 4674 58546
rect 4674 58494 4676 58546
rect 4620 58492 4676 58494
rect 4614 57258 4670 57260
rect 4614 57206 4616 57258
rect 4616 57206 4668 57258
rect 4668 57206 4670 57258
rect 4614 57204 4670 57206
rect 4718 57258 4774 57260
rect 4718 57206 4720 57258
rect 4720 57206 4772 57258
rect 4772 57206 4774 57258
rect 4718 57204 4774 57206
rect 4822 57258 4878 57260
rect 4822 57206 4824 57258
rect 4824 57206 4876 57258
rect 4876 57206 4878 57258
rect 4822 57204 4878 57206
rect 4396 56700 4452 56756
rect 4620 56812 4676 56868
rect 4284 56476 4340 56532
rect 3724 54684 3780 54740
rect 3836 55580 3892 55636
rect 3500 54572 3556 54628
rect 3276 54290 3332 54292
rect 3276 54238 3278 54290
rect 3278 54238 3330 54290
rect 3330 54238 3332 54290
rect 3276 54236 3332 54238
rect 3948 54236 4004 54292
rect 1708 53618 1764 53620
rect 1708 53566 1710 53618
rect 1710 53566 1762 53618
rect 1762 53566 1764 53618
rect 1708 53564 1764 53566
rect 1708 50428 1764 50484
rect 1820 49644 1876 49700
rect 1820 49308 1876 49364
rect 1932 53564 1988 53620
rect 1932 53116 1988 53172
rect 2940 53452 2996 53508
rect 2828 53116 2884 53172
rect 2156 52834 2212 52836
rect 2156 52782 2158 52834
rect 2158 52782 2210 52834
rect 2210 52782 2212 52834
rect 2156 52780 2212 52782
rect 2268 52050 2324 52052
rect 2268 51998 2270 52050
rect 2270 51998 2322 52050
rect 2322 51998 2324 52050
rect 2268 51996 2324 51998
rect 2716 52722 2772 52724
rect 2716 52670 2718 52722
rect 2718 52670 2770 52722
rect 2770 52670 2772 52722
rect 2716 52668 2772 52670
rect 2044 51100 2100 51156
rect 2156 50092 2212 50148
rect 2044 49922 2100 49924
rect 2044 49870 2046 49922
rect 2046 49870 2098 49922
rect 2098 49870 2100 49922
rect 2044 49868 2100 49870
rect 1708 47516 1764 47572
rect 1820 48860 1876 48916
rect 1708 47346 1764 47348
rect 1708 47294 1710 47346
rect 1710 47294 1762 47346
rect 1762 47294 1764 47346
rect 1708 47292 1764 47294
rect 2156 47404 2212 47460
rect 2044 47234 2100 47236
rect 2044 47182 2046 47234
rect 2046 47182 2098 47234
rect 2098 47182 2100 47234
rect 2044 47180 2100 47182
rect 1820 46844 1876 46900
rect 1708 45052 1764 45108
rect 1932 44828 1988 44884
rect 2828 52274 2884 52276
rect 2828 52222 2830 52274
rect 2830 52222 2882 52274
rect 2882 52222 2884 52274
rect 2828 52220 2884 52222
rect 2716 51154 2772 51156
rect 2716 51102 2718 51154
rect 2718 51102 2770 51154
rect 2770 51102 2772 51154
rect 2716 51100 2772 51102
rect 2492 50482 2548 50484
rect 2492 50430 2494 50482
rect 2494 50430 2546 50482
rect 2546 50430 2548 50482
rect 2492 50428 2548 50430
rect 4172 56082 4228 56084
rect 4172 56030 4174 56082
rect 4174 56030 4226 56082
rect 4226 56030 4228 56082
rect 4172 56028 4228 56030
rect 6076 74898 6132 74900
rect 6076 74846 6078 74898
rect 6078 74846 6130 74898
rect 6130 74846 6132 74898
rect 6076 74844 6132 74846
rect 7084 76524 7140 76580
rect 6524 76300 6580 76356
rect 6860 76466 6916 76468
rect 6860 76414 6862 76466
rect 6862 76414 6914 76466
rect 6914 76414 6916 76466
rect 6860 76412 6916 76414
rect 6300 76188 6356 76244
rect 7084 76076 7140 76132
rect 8764 76636 8820 76692
rect 7644 76242 7700 76244
rect 7644 76190 7646 76242
rect 7646 76190 7698 76242
rect 7698 76190 7700 76242
rect 7644 76188 7700 76190
rect 6860 75852 6916 75908
rect 6972 75404 7028 75460
rect 6860 74898 6916 74900
rect 6860 74846 6862 74898
rect 6862 74846 6914 74898
rect 6914 74846 6916 74898
rect 6860 74844 6916 74846
rect 5964 74732 6020 74788
rect 5964 74284 6020 74340
rect 6524 73948 6580 74004
rect 5740 73836 5796 73892
rect 6188 72658 6244 72660
rect 6188 72606 6190 72658
rect 6190 72606 6242 72658
rect 6242 72606 6244 72658
rect 6188 72604 6244 72606
rect 6076 72380 6132 72436
rect 5740 71596 5796 71652
rect 6076 70978 6132 70980
rect 6076 70926 6078 70978
rect 6078 70926 6130 70978
rect 6130 70926 6132 70978
rect 6076 70924 6132 70926
rect 7196 74002 7252 74004
rect 7196 73950 7198 74002
rect 7198 73950 7250 74002
rect 7250 73950 7252 74002
rect 7196 73948 7252 73950
rect 7196 72716 7252 72772
rect 6972 72658 7028 72660
rect 6972 72606 6974 72658
rect 6974 72606 7026 72658
rect 7026 72606 7028 72658
rect 6972 72604 7028 72606
rect 6636 72380 6692 72436
rect 5628 70588 5684 70644
rect 5516 70140 5572 70196
rect 5964 70700 6020 70756
rect 5852 70476 5908 70532
rect 5964 67564 6020 67620
rect 5852 65996 5908 66052
rect 6076 66108 6132 66164
rect 5740 64764 5796 64820
rect 6076 64428 6132 64484
rect 6300 67730 6356 67732
rect 6300 67678 6302 67730
rect 6302 67678 6354 67730
rect 6354 67678 6356 67730
rect 6300 67676 6356 67678
rect 6412 66892 6468 66948
rect 6524 65660 6580 65716
rect 7756 76076 7812 76132
rect 8016 75290 8072 75292
rect 8016 75238 8018 75290
rect 8018 75238 8070 75290
rect 8070 75238 8072 75290
rect 8016 75236 8072 75238
rect 8120 75290 8176 75292
rect 8120 75238 8122 75290
rect 8122 75238 8174 75290
rect 8174 75238 8176 75290
rect 8120 75236 8176 75238
rect 8224 75290 8280 75292
rect 8224 75238 8226 75290
rect 8226 75238 8278 75290
rect 8278 75238 8280 75290
rect 8224 75236 8280 75238
rect 7980 75122 8036 75124
rect 7980 75070 7982 75122
rect 7982 75070 8034 75122
rect 8034 75070 8036 75122
rect 7980 75068 8036 75070
rect 8540 76354 8596 76356
rect 8540 76302 8542 76354
rect 8542 76302 8594 76354
rect 8594 76302 8596 76354
rect 8540 76300 8596 76302
rect 9772 81116 9828 81172
rect 10220 83020 10276 83076
rect 10668 84306 10724 84308
rect 10668 84254 10670 84306
rect 10670 84254 10722 84306
rect 10722 84254 10724 84306
rect 10668 84252 10724 84254
rect 10332 82962 10388 82964
rect 10332 82910 10334 82962
rect 10334 82910 10386 82962
rect 10386 82910 10388 82962
rect 10332 82908 10388 82910
rect 10780 82962 10836 82964
rect 10780 82910 10782 82962
rect 10782 82910 10834 82962
rect 10834 82910 10836 82962
rect 10780 82908 10836 82910
rect 10668 81564 10724 81620
rect 10780 81676 10836 81732
rect 10220 81394 10276 81396
rect 10220 81342 10222 81394
rect 10222 81342 10274 81394
rect 10274 81342 10276 81394
rect 10220 81340 10276 81342
rect 9996 79548 10052 79604
rect 9884 78988 9940 79044
rect 9884 78034 9940 78036
rect 9884 77982 9886 78034
rect 9886 77982 9938 78034
rect 9938 77982 9940 78034
rect 9884 77980 9940 77982
rect 9660 77250 9716 77252
rect 9660 77198 9662 77250
rect 9662 77198 9714 77250
rect 9714 77198 9716 77250
rect 9660 77196 9716 77198
rect 9548 76860 9604 76916
rect 9772 76466 9828 76468
rect 9772 76414 9774 76466
rect 9774 76414 9826 76466
rect 9826 76414 9828 76466
rect 9772 76412 9828 76414
rect 8988 76188 9044 76244
rect 9772 75794 9828 75796
rect 9772 75742 9774 75794
rect 9774 75742 9826 75794
rect 9826 75742 9828 75794
rect 9772 75740 9828 75742
rect 8540 75404 8596 75460
rect 8652 75516 8708 75572
rect 6860 70978 6916 70980
rect 6860 70926 6862 70978
rect 6862 70926 6914 70978
rect 6914 70926 6916 70978
rect 6860 70924 6916 70926
rect 6748 70866 6804 70868
rect 6748 70814 6750 70866
rect 6750 70814 6802 70866
rect 6802 70814 6804 70866
rect 6748 70812 6804 70814
rect 8016 73722 8072 73724
rect 8016 73670 8018 73722
rect 8018 73670 8070 73722
rect 8070 73670 8072 73722
rect 8016 73668 8072 73670
rect 8120 73722 8176 73724
rect 8120 73670 8122 73722
rect 8122 73670 8174 73722
rect 8174 73670 8176 73722
rect 8120 73668 8176 73670
rect 8224 73722 8280 73724
rect 8224 73670 8226 73722
rect 8226 73670 8278 73722
rect 8278 73670 8280 73722
rect 8224 73668 8280 73670
rect 8764 75122 8820 75124
rect 8764 75070 8766 75122
rect 8766 75070 8818 75122
rect 8818 75070 8820 75122
rect 8764 75068 8820 75070
rect 8764 73836 8820 73892
rect 8428 73500 8484 73556
rect 7868 72716 7924 72772
rect 7980 72658 8036 72660
rect 7980 72606 7982 72658
rect 7982 72606 8034 72658
rect 8034 72606 8036 72658
rect 7980 72604 8036 72606
rect 7644 72492 7700 72548
rect 8092 72492 8148 72548
rect 8988 73948 9044 74004
rect 8016 72154 8072 72156
rect 8016 72102 8018 72154
rect 8018 72102 8070 72154
rect 8070 72102 8072 72154
rect 8016 72100 8072 72102
rect 8120 72154 8176 72156
rect 8120 72102 8122 72154
rect 8122 72102 8174 72154
rect 8174 72102 8176 72154
rect 8120 72100 8176 72102
rect 8224 72154 8280 72156
rect 8224 72102 8226 72154
rect 8226 72102 8278 72154
rect 8278 72102 8280 72154
rect 8224 72100 8280 72102
rect 8540 72716 8596 72772
rect 8428 71708 8484 71764
rect 7084 70364 7140 70420
rect 7084 67618 7140 67620
rect 7084 67566 7086 67618
rect 7086 67566 7138 67618
rect 7138 67566 7140 67618
rect 7084 67564 7140 67566
rect 6860 66050 6916 66052
rect 6860 65998 6862 66050
rect 6862 65998 6914 66050
rect 6914 65998 6916 66050
rect 6860 65996 6916 65998
rect 6412 64092 6468 64148
rect 6188 63980 6244 64036
rect 6076 63922 6132 63924
rect 6076 63870 6078 63922
rect 6078 63870 6130 63922
rect 6130 63870 6132 63922
rect 6076 63868 6132 63870
rect 5180 62076 5236 62132
rect 5292 61740 5348 61796
rect 5180 61068 5236 61124
rect 5068 57874 5124 57876
rect 5068 57822 5070 57874
rect 5070 57822 5122 57874
rect 5122 57822 5124 57874
rect 5068 57820 5124 57822
rect 5180 59388 5236 59444
rect 5404 56924 5460 56980
rect 5852 63420 5908 63476
rect 5852 62188 5908 62244
rect 5292 56700 5348 56756
rect 5964 62076 6020 62132
rect 6188 61628 6244 61684
rect 6076 61570 6132 61572
rect 6076 61518 6078 61570
rect 6078 61518 6130 61570
rect 6130 61518 6132 61570
rect 6076 61516 6132 61518
rect 5740 61068 5796 61124
rect 5740 60508 5796 60564
rect 5740 60172 5796 60228
rect 6636 64764 6692 64820
rect 6636 63756 6692 63812
rect 6636 63308 6692 63364
rect 6748 62524 6804 62580
rect 5740 59442 5796 59444
rect 5740 59390 5742 59442
rect 5742 59390 5794 59442
rect 5794 59390 5796 59442
rect 5740 59388 5796 59390
rect 6524 62300 6580 62356
rect 5628 58434 5684 58436
rect 5628 58382 5630 58434
rect 5630 58382 5682 58434
rect 5682 58382 5684 58434
rect 5628 58380 5684 58382
rect 5516 56700 5572 56756
rect 5628 57260 5684 57316
rect 6636 62242 6692 62244
rect 6636 62190 6638 62242
rect 6638 62190 6690 62242
rect 6690 62190 6692 62242
rect 6636 62188 6692 62190
rect 7420 70812 7476 70868
rect 7980 71036 8036 71092
rect 8876 72492 8932 72548
rect 9772 75404 9828 75460
rect 10556 79324 10612 79380
rect 10332 78876 10388 78932
rect 10332 78652 10388 78708
rect 10108 77250 10164 77252
rect 10108 77198 10110 77250
rect 10110 77198 10162 77250
rect 10162 77198 10164 77250
rect 10108 77196 10164 77198
rect 10108 76466 10164 76468
rect 10108 76414 10110 76466
rect 10110 76414 10162 76466
rect 10162 76414 10164 76466
rect 10108 76412 10164 76414
rect 10220 75740 10276 75796
rect 9996 75122 10052 75124
rect 9996 75070 9998 75122
rect 9998 75070 10050 75122
rect 10050 75070 10052 75122
rect 9996 75068 10052 75070
rect 9324 73948 9380 74004
rect 10780 77138 10836 77140
rect 10780 77086 10782 77138
rect 10782 77086 10834 77138
rect 10834 77086 10836 77138
rect 10780 77084 10836 77086
rect 10444 76578 10500 76580
rect 10444 76526 10446 76578
rect 10446 76526 10498 76578
rect 10498 76526 10500 76578
rect 10444 76524 10500 76526
rect 10444 75516 10500 75572
rect 9996 74060 10052 74116
rect 9772 73836 9828 73892
rect 9548 73500 9604 73556
rect 9324 72604 9380 72660
rect 9100 72268 9156 72324
rect 8764 71762 8820 71764
rect 8764 71710 8766 71762
rect 8766 71710 8818 71762
rect 8818 71710 8820 71762
rect 8764 71708 8820 71710
rect 8988 71596 9044 71652
rect 7980 70754 8036 70756
rect 7980 70702 7982 70754
rect 7982 70702 8034 70754
rect 8034 70702 8036 70754
rect 7980 70700 8036 70702
rect 8016 70586 8072 70588
rect 8016 70534 8018 70586
rect 8018 70534 8070 70586
rect 8070 70534 8072 70586
rect 8016 70532 8072 70534
rect 8120 70586 8176 70588
rect 8120 70534 8122 70586
rect 8122 70534 8174 70586
rect 8174 70534 8176 70586
rect 8120 70532 8176 70534
rect 8224 70586 8280 70588
rect 8224 70534 8226 70586
rect 8226 70534 8278 70586
rect 8278 70534 8280 70586
rect 8224 70532 8280 70534
rect 8540 70588 8596 70644
rect 8876 71090 8932 71092
rect 8876 71038 8878 71090
rect 8878 71038 8930 71090
rect 8930 71038 8932 71090
rect 8876 71036 8932 71038
rect 9436 71596 9492 71652
rect 9660 71650 9716 71652
rect 9660 71598 9662 71650
rect 9662 71598 9714 71650
rect 9714 71598 9716 71650
rect 9660 71596 9716 71598
rect 9548 71484 9604 71540
rect 9548 70306 9604 70308
rect 9548 70254 9550 70306
rect 9550 70254 9602 70306
rect 9602 70254 9604 70306
rect 9548 70252 9604 70254
rect 9436 69804 9492 69860
rect 8428 69132 8484 69188
rect 8016 69018 8072 69020
rect 8016 68966 8018 69018
rect 8018 68966 8070 69018
rect 8070 68966 8072 69018
rect 8016 68964 8072 68966
rect 8120 69018 8176 69020
rect 8120 68966 8122 69018
rect 8122 68966 8174 69018
rect 8174 68966 8176 69018
rect 8120 68964 8176 68966
rect 8224 69018 8280 69020
rect 8224 68966 8226 69018
rect 8226 68966 8278 69018
rect 8278 68966 8280 69018
rect 8224 68964 8280 68966
rect 7756 67954 7812 67956
rect 7756 67902 7758 67954
rect 7758 67902 7810 67954
rect 7810 67902 7812 67954
rect 7756 67900 7812 67902
rect 9324 69298 9380 69300
rect 9324 69246 9326 69298
rect 9326 69246 9378 69298
rect 9378 69246 9380 69298
rect 9324 69244 9380 69246
rect 9212 69186 9268 69188
rect 9212 69134 9214 69186
rect 9214 69134 9266 69186
rect 9266 69134 9268 69186
rect 9212 69132 9268 69134
rect 9436 69186 9492 69188
rect 9436 69134 9438 69186
rect 9438 69134 9490 69186
rect 9490 69134 9492 69186
rect 9436 69132 9492 69134
rect 8016 67450 8072 67452
rect 8016 67398 8018 67450
rect 8018 67398 8070 67450
rect 8070 67398 8072 67450
rect 8016 67396 8072 67398
rect 8120 67450 8176 67452
rect 8120 67398 8122 67450
rect 8122 67398 8174 67450
rect 8174 67398 8176 67450
rect 8120 67396 8176 67398
rect 8224 67450 8280 67452
rect 8224 67398 8226 67450
rect 8226 67398 8278 67450
rect 8278 67398 8280 67450
rect 8224 67396 8280 67398
rect 7980 66946 8036 66948
rect 7980 66894 7982 66946
rect 7982 66894 8034 66946
rect 8034 66894 8036 66946
rect 7980 66892 8036 66894
rect 7868 66780 7924 66836
rect 7420 65660 7476 65716
rect 7196 65436 7252 65492
rect 7196 64652 7252 64708
rect 7084 63868 7140 63924
rect 7084 62300 7140 62356
rect 8316 66332 8372 66388
rect 8016 65882 8072 65884
rect 8016 65830 8018 65882
rect 8018 65830 8070 65882
rect 8070 65830 8072 65882
rect 8016 65828 8072 65830
rect 8120 65882 8176 65884
rect 8120 65830 8122 65882
rect 8122 65830 8174 65882
rect 8174 65830 8176 65882
rect 8120 65828 8176 65830
rect 8224 65882 8280 65884
rect 8224 65830 8226 65882
rect 8226 65830 8278 65882
rect 8278 65830 8280 65882
rect 8224 65828 8280 65830
rect 7644 65436 7700 65492
rect 8428 65436 8484 65492
rect 8016 64314 8072 64316
rect 8016 64262 8018 64314
rect 8018 64262 8070 64314
rect 8070 64262 8072 64314
rect 8016 64260 8072 64262
rect 8120 64314 8176 64316
rect 8120 64262 8122 64314
rect 8122 64262 8174 64314
rect 8174 64262 8176 64314
rect 8120 64260 8176 64262
rect 8224 64314 8280 64316
rect 8224 64262 8226 64314
rect 8226 64262 8278 64314
rect 8278 64262 8280 64314
rect 8224 64260 8280 64262
rect 7420 63922 7476 63924
rect 7420 63870 7422 63922
rect 7422 63870 7474 63922
rect 7474 63870 7476 63922
rect 7420 63868 7476 63870
rect 6860 61570 6916 61572
rect 6860 61518 6862 61570
rect 6862 61518 6914 61570
rect 6914 61518 6916 61570
rect 6860 61516 6916 61518
rect 6748 61292 6804 61348
rect 7084 61404 7140 61460
rect 6748 60396 6804 60452
rect 6188 59106 6244 59108
rect 6188 59054 6190 59106
rect 6190 59054 6242 59106
rect 6242 59054 6244 59106
rect 6188 59052 6244 59054
rect 5852 57932 5908 57988
rect 6076 57708 6132 57764
rect 6524 59218 6580 59220
rect 6524 59166 6526 59218
rect 6526 59166 6578 59218
rect 6578 59166 6580 59218
rect 6524 59164 6580 59166
rect 7532 63810 7588 63812
rect 7532 63758 7534 63810
rect 7534 63758 7586 63810
rect 7586 63758 7588 63810
rect 7532 63756 7588 63758
rect 8428 62860 8484 62916
rect 8016 62746 8072 62748
rect 8016 62694 8018 62746
rect 8018 62694 8070 62746
rect 8070 62694 8072 62746
rect 8016 62692 8072 62694
rect 8120 62746 8176 62748
rect 8120 62694 8122 62746
rect 8122 62694 8174 62746
rect 8174 62694 8176 62746
rect 8120 62692 8176 62694
rect 8224 62746 8280 62748
rect 8224 62694 8226 62746
rect 8226 62694 8278 62746
rect 8278 62694 8280 62746
rect 8224 62692 8280 62694
rect 7980 62524 8036 62580
rect 7756 62354 7812 62356
rect 7756 62302 7758 62354
rect 7758 62302 7810 62354
rect 7810 62302 7812 62354
rect 7756 62300 7812 62302
rect 8428 62524 8484 62580
rect 8316 62466 8372 62468
rect 8316 62414 8318 62466
rect 8318 62414 8370 62466
rect 8370 62414 8372 62466
rect 8316 62412 8372 62414
rect 7532 61346 7588 61348
rect 7532 61294 7534 61346
rect 7534 61294 7586 61346
rect 7586 61294 7588 61346
rect 7532 61292 7588 61294
rect 7532 60732 7588 60788
rect 6860 59164 6916 59220
rect 7420 59388 7476 59444
rect 6748 59052 6804 59108
rect 6300 57820 6356 57876
rect 6076 57148 6132 57204
rect 5852 56754 5908 56756
rect 5852 56702 5854 56754
rect 5854 56702 5906 56754
rect 5906 56702 5908 56754
rect 5852 56700 5908 56702
rect 5628 56588 5684 56644
rect 5180 56476 5236 56532
rect 4956 56028 5012 56084
rect 4284 55804 4340 55860
rect 4614 55690 4670 55692
rect 4614 55638 4616 55690
rect 4616 55638 4668 55690
rect 4668 55638 4670 55690
rect 4614 55636 4670 55638
rect 4718 55690 4774 55692
rect 4718 55638 4720 55690
rect 4720 55638 4772 55690
rect 4772 55638 4774 55690
rect 4718 55636 4774 55638
rect 4822 55690 4878 55692
rect 4822 55638 4824 55690
rect 4824 55638 4876 55690
rect 4876 55638 4878 55690
rect 4822 55636 4878 55638
rect 4060 53900 4116 53956
rect 2940 50092 2996 50148
rect 3052 51100 3108 51156
rect 2604 49756 2660 49812
rect 2492 49532 2548 49588
rect 2492 48130 2548 48132
rect 2492 48078 2494 48130
rect 2494 48078 2546 48130
rect 2546 48078 2548 48130
rect 2492 48076 2548 48078
rect 2492 47570 2548 47572
rect 2492 47518 2494 47570
rect 2494 47518 2546 47570
rect 2546 47518 2548 47570
rect 2492 47516 2548 47518
rect 3164 50428 3220 50484
rect 4396 54626 4452 54628
rect 4396 54574 4398 54626
rect 4398 54574 4450 54626
rect 4450 54574 4452 54626
rect 4396 54572 4452 54574
rect 4614 54122 4670 54124
rect 4614 54070 4616 54122
rect 4616 54070 4668 54122
rect 4668 54070 4670 54122
rect 4614 54068 4670 54070
rect 4718 54122 4774 54124
rect 4718 54070 4720 54122
rect 4720 54070 4772 54122
rect 4772 54070 4774 54122
rect 4718 54068 4774 54070
rect 4822 54122 4878 54124
rect 4822 54070 4824 54122
rect 4824 54070 4876 54122
rect 4876 54070 4878 54122
rect 4822 54068 4878 54070
rect 3836 53730 3892 53732
rect 3836 53678 3838 53730
rect 3838 53678 3890 53730
rect 3890 53678 3892 53730
rect 3836 53676 3892 53678
rect 4172 53618 4228 53620
rect 4172 53566 4174 53618
rect 4174 53566 4226 53618
rect 4226 53566 4228 53618
rect 4172 53564 4228 53566
rect 3836 53228 3892 53284
rect 4508 53900 4564 53956
rect 3724 52332 3780 52388
rect 3388 52274 3444 52276
rect 3388 52222 3390 52274
rect 3390 52222 3442 52274
rect 3442 52222 3444 52274
rect 3388 52220 3444 52222
rect 4732 53900 4788 53956
rect 4620 53788 4676 53844
rect 4956 53564 5012 53620
rect 5516 55804 5572 55860
rect 5292 54738 5348 54740
rect 5292 54686 5294 54738
rect 5294 54686 5346 54738
rect 5346 54686 5348 54738
rect 5292 54684 5348 54686
rect 5292 53788 5348 53844
rect 5404 54572 5460 54628
rect 4620 52892 4676 52948
rect 4732 52668 4788 52724
rect 5180 53228 5236 53284
rect 4614 52554 4670 52556
rect 4614 52502 4616 52554
rect 4616 52502 4668 52554
rect 4668 52502 4670 52554
rect 4614 52500 4670 52502
rect 4718 52554 4774 52556
rect 4718 52502 4720 52554
rect 4720 52502 4772 52554
rect 4772 52502 4774 52554
rect 4718 52500 4774 52502
rect 4822 52554 4878 52556
rect 4822 52502 4824 52554
rect 4824 52502 4876 52554
rect 4876 52502 4878 52554
rect 4822 52500 4878 52502
rect 4284 52220 4340 52276
rect 3724 52162 3780 52164
rect 3724 52110 3726 52162
rect 3726 52110 3778 52162
rect 3778 52110 3780 52162
rect 3724 52108 3780 52110
rect 3612 51378 3668 51380
rect 3612 51326 3614 51378
rect 3614 51326 3666 51378
rect 3666 51326 3668 51378
rect 3612 51324 3668 51326
rect 3836 51154 3892 51156
rect 3836 51102 3838 51154
rect 3838 51102 3890 51154
rect 3890 51102 3892 51154
rect 3836 51100 3892 51102
rect 3276 49980 3332 50036
rect 3164 49810 3220 49812
rect 3164 49758 3166 49810
rect 3166 49758 3218 49810
rect 3218 49758 3220 49810
rect 3164 49756 3220 49758
rect 2940 48300 2996 48356
rect 3052 48076 3108 48132
rect 4060 50764 4116 50820
rect 4732 52332 4788 52388
rect 4508 51996 4564 52052
rect 4396 51938 4452 51940
rect 4396 51886 4398 51938
rect 4398 51886 4450 51938
rect 4450 51886 4452 51938
rect 4396 51884 4452 51886
rect 5068 53004 5124 53060
rect 6412 56924 6468 56980
rect 6188 56476 6244 56532
rect 5628 53730 5684 53732
rect 5628 53678 5630 53730
rect 5630 53678 5682 53730
rect 5682 53678 5684 53730
rect 5628 53676 5684 53678
rect 5852 53788 5908 53844
rect 5740 53004 5796 53060
rect 5740 52668 5796 52724
rect 6076 54572 6132 54628
rect 6188 54402 6244 54404
rect 6188 54350 6190 54402
rect 6190 54350 6242 54402
rect 6242 54350 6244 54402
rect 6188 54348 6244 54350
rect 6300 53788 6356 53844
rect 6300 53564 6356 53620
rect 6300 53228 6356 53284
rect 5628 51996 5684 52052
rect 4732 51602 4788 51604
rect 4732 51550 4734 51602
rect 4734 51550 4786 51602
rect 4786 51550 4788 51602
rect 4732 51548 4788 51550
rect 4614 50986 4670 50988
rect 4614 50934 4616 50986
rect 4616 50934 4668 50986
rect 4668 50934 4670 50986
rect 4614 50932 4670 50934
rect 4718 50986 4774 50988
rect 4718 50934 4720 50986
rect 4720 50934 4772 50986
rect 4772 50934 4774 50986
rect 4718 50932 4774 50934
rect 4822 50986 4878 50988
rect 4822 50934 4824 50986
rect 4824 50934 4876 50986
rect 4876 50934 4878 50986
rect 4822 50932 4878 50934
rect 4620 50764 4676 50820
rect 4284 49980 4340 50036
rect 3612 49026 3668 49028
rect 3612 48974 3614 49026
rect 3614 48974 3666 49026
rect 3666 48974 3668 49026
rect 3612 48972 3668 48974
rect 3612 48748 3668 48804
rect 3164 47628 3220 47684
rect 3500 47682 3556 47684
rect 3500 47630 3502 47682
rect 3502 47630 3554 47682
rect 3554 47630 3556 47682
rect 3500 47628 3556 47630
rect 2604 47292 2660 47348
rect 3164 47458 3220 47460
rect 3164 47406 3166 47458
rect 3166 47406 3218 47458
rect 3218 47406 3220 47458
rect 3164 47404 3220 47406
rect 3500 47292 3556 47348
rect 2380 45724 2436 45780
rect 2380 45276 2436 45332
rect 1820 43708 1876 43764
rect 1708 42364 1764 42420
rect 1708 39676 1764 39732
rect 3612 46732 3668 46788
rect 3164 46562 3220 46564
rect 3164 46510 3166 46562
rect 3166 46510 3218 46562
rect 3218 46510 3220 46562
rect 3164 46508 3220 46510
rect 3612 46396 3668 46452
rect 2828 45276 2884 45332
rect 3612 45164 3668 45220
rect 2828 45106 2884 45108
rect 2828 45054 2830 45106
rect 2830 45054 2882 45106
rect 2882 45054 2884 45106
rect 2828 45052 2884 45054
rect 2828 44828 2884 44884
rect 2828 44380 2884 44436
rect 2492 44156 2548 44212
rect 2156 43762 2212 43764
rect 2156 43710 2158 43762
rect 2158 43710 2210 43762
rect 2210 43710 2212 43762
rect 2156 43708 2212 43710
rect 2380 43708 2436 43764
rect 2492 43650 2548 43652
rect 2492 43598 2494 43650
rect 2494 43598 2546 43650
rect 2546 43598 2548 43650
rect 2492 43596 2548 43598
rect 3052 44098 3108 44100
rect 3052 44046 3054 44098
rect 3054 44046 3106 44098
rect 3106 44046 3108 44098
rect 3052 44044 3108 44046
rect 2044 40962 2100 40964
rect 2044 40910 2046 40962
rect 2046 40910 2098 40962
rect 2098 40910 2100 40962
rect 2044 40908 2100 40910
rect 2044 40348 2100 40404
rect 2044 39788 2100 39844
rect 1820 39004 1876 39060
rect 1708 36988 1764 37044
rect 2044 36258 2100 36260
rect 2044 36206 2046 36258
rect 2046 36206 2098 36258
rect 2098 36206 2100 36258
rect 2044 36204 2100 36206
rect 1932 35196 1988 35252
rect 1708 34300 1764 34356
rect 2044 33292 2100 33348
rect 2380 40796 2436 40852
rect 2492 40460 2548 40516
rect 3164 43596 3220 43652
rect 2716 41970 2772 41972
rect 2716 41918 2718 41970
rect 2718 41918 2770 41970
rect 2770 41918 2772 41970
rect 2716 41916 2772 41918
rect 3052 43484 3108 43540
rect 3388 44994 3444 44996
rect 3388 44942 3390 44994
rect 3390 44942 3442 44994
rect 3442 44942 3444 44994
rect 3388 44940 3444 44942
rect 5180 51490 5236 51492
rect 5180 51438 5182 51490
rect 5182 51438 5234 51490
rect 5234 51438 5236 51490
rect 5180 51436 5236 51438
rect 5852 52274 5908 52276
rect 5852 52222 5854 52274
rect 5854 52222 5906 52274
rect 5906 52222 5908 52274
rect 5852 52220 5908 52222
rect 6636 57820 6692 57876
rect 6636 55916 6692 55972
rect 6860 56866 6916 56868
rect 6860 56814 6862 56866
rect 6862 56814 6914 56866
rect 6914 56814 6916 56866
rect 6860 56812 6916 56814
rect 6748 56140 6804 56196
rect 8016 61178 8072 61180
rect 8016 61126 8018 61178
rect 8018 61126 8070 61178
rect 8070 61126 8072 61178
rect 8016 61124 8072 61126
rect 8120 61178 8176 61180
rect 8120 61126 8122 61178
rect 8122 61126 8174 61178
rect 8174 61126 8176 61178
rect 8120 61124 8176 61126
rect 8224 61178 8280 61180
rect 8224 61126 8226 61178
rect 8226 61126 8278 61178
rect 8278 61126 8280 61178
rect 8224 61124 8280 61126
rect 8316 60786 8372 60788
rect 8316 60734 8318 60786
rect 8318 60734 8370 60786
rect 8370 60734 8372 60786
rect 8316 60732 8372 60734
rect 7868 60060 7924 60116
rect 8428 60172 8484 60228
rect 7756 59218 7812 59220
rect 7756 59166 7758 59218
rect 7758 59166 7810 59218
rect 7810 59166 7812 59218
rect 7756 59164 7812 59166
rect 7532 58156 7588 58212
rect 7756 58492 7812 58548
rect 7084 57874 7140 57876
rect 7084 57822 7086 57874
rect 7086 57822 7138 57874
rect 7138 57822 7140 57874
rect 7084 57820 7140 57822
rect 7532 57260 7588 57316
rect 7532 56754 7588 56756
rect 7532 56702 7534 56754
rect 7534 56702 7586 56754
rect 7586 56702 7588 56754
rect 7532 56700 7588 56702
rect 7420 55970 7476 55972
rect 7420 55918 7422 55970
rect 7422 55918 7474 55970
rect 7474 55918 7476 55970
rect 7420 55916 7476 55918
rect 7756 55356 7812 55412
rect 6636 53788 6692 53844
rect 6748 53564 6804 53620
rect 6748 52444 6804 52500
rect 7084 52274 7140 52276
rect 7084 52222 7086 52274
rect 7086 52222 7138 52274
rect 7138 52222 7140 52274
rect 7084 52220 7140 52222
rect 6188 52050 6244 52052
rect 6188 51998 6190 52050
rect 6190 51998 6242 52050
rect 6242 51998 6244 52050
rect 6188 51996 6244 51998
rect 5964 51548 6020 51604
rect 5404 51212 5460 51268
rect 5180 50706 5236 50708
rect 5180 50654 5182 50706
rect 5182 50654 5234 50706
rect 5234 50654 5236 50706
rect 5180 50652 5236 50654
rect 4620 49532 4676 49588
rect 4614 49418 4670 49420
rect 4614 49366 4616 49418
rect 4616 49366 4668 49418
rect 4668 49366 4670 49418
rect 4614 49364 4670 49366
rect 4718 49418 4774 49420
rect 4718 49366 4720 49418
rect 4720 49366 4772 49418
rect 4772 49366 4774 49418
rect 4718 49364 4774 49366
rect 4822 49418 4878 49420
rect 4822 49366 4824 49418
rect 4824 49366 4876 49418
rect 4876 49366 4878 49418
rect 4822 49364 4878 49366
rect 4396 49196 4452 49252
rect 3948 49026 4004 49028
rect 3948 48974 3950 49026
rect 3950 48974 4002 49026
rect 4002 48974 4004 49026
rect 3948 48972 4004 48974
rect 5068 49196 5124 49252
rect 3724 44716 3780 44772
rect 3836 48524 3892 48580
rect 4172 48802 4228 48804
rect 4172 48750 4174 48802
rect 4174 48750 4226 48802
rect 4226 48750 4228 48802
rect 4172 48748 4228 48750
rect 4060 47628 4116 47684
rect 4172 48412 4228 48468
rect 3836 44604 3892 44660
rect 3948 47516 4004 47572
rect 4060 46898 4116 46900
rect 4060 46846 4062 46898
rect 4062 46846 4114 46898
rect 4114 46846 4116 46898
rect 4060 46844 4116 46846
rect 4060 45388 4116 45444
rect 4284 47292 4340 47348
rect 4396 48972 4452 49028
rect 3948 44492 4004 44548
rect 4284 46396 4340 46452
rect 3724 44434 3780 44436
rect 3724 44382 3726 44434
rect 3726 44382 3778 44434
rect 3778 44382 3780 44434
rect 3724 44380 3780 44382
rect 3388 44210 3444 44212
rect 3388 44158 3390 44210
rect 3390 44158 3442 44210
rect 3442 44158 3444 44210
rect 3388 44156 3444 44158
rect 3836 44098 3892 44100
rect 3836 44046 3838 44098
rect 3838 44046 3890 44098
rect 3890 44046 3892 44098
rect 3836 44044 3892 44046
rect 3836 43372 3892 43428
rect 3724 41970 3780 41972
rect 3724 41918 3726 41970
rect 3726 41918 3778 41970
rect 3778 41918 3780 41970
rect 3724 41916 3780 41918
rect 3388 41692 3444 41748
rect 3052 40908 3108 40964
rect 3500 41244 3556 41300
rect 3836 41132 3892 41188
rect 2940 40572 2996 40628
rect 3164 40796 3220 40852
rect 3500 40796 3556 40852
rect 2828 40348 2884 40404
rect 3612 40402 3668 40404
rect 3612 40350 3614 40402
rect 3614 40350 3666 40402
rect 3666 40350 3668 40402
rect 3612 40348 3668 40350
rect 3724 40178 3780 40180
rect 3724 40126 3726 40178
rect 3726 40126 3778 40178
rect 3778 40126 3780 40178
rect 3724 40124 3780 40126
rect 4620 48748 4676 48804
rect 4620 47964 4676 48020
rect 4956 48300 5012 48356
rect 4614 47850 4670 47852
rect 4614 47798 4616 47850
rect 4616 47798 4668 47850
rect 4668 47798 4670 47850
rect 4614 47796 4670 47798
rect 4718 47850 4774 47852
rect 4718 47798 4720 47850
rect 4720 47798 4772 47850
rect 4772 47798 4774 47850
rect 4718 47796 4774 47798
rect 4822 47850 4878 47852
rect 4822 47798 4824 47850
rect 4824 47798 4876 47850
rect 4876 47798 4878 47850
rect 4956 47852 5012 47908
rect 4822 47796 4878 47798
rect 4732 47570 4788 47572
rect 4732 47518 4734 47570
rect 4734 47518 4786 47570
rect 4786 47518 4788 47570
rect 4732 47516 4788 47518
rect 4508 47404 4564 47460
rect 4844 47012 4900 47068
rect 4956 47404 5012 47460
rect 4508 46562 4564 46564
rect 4508 46510 4510 46562
rect 4510 46510 4562 46562
rect 4562 46510 4564 46562
rect 4508 46508 4564 46510
rect 5068 47180 5124 47236
rect 5292 49084 5348 49140
rect 5964 51266 6020 51268
rect 5964 51214 5966 51266
rect 5966 51214 6018 51266
rect 6018 51214 6020 51266
rect 5964 51212 6020 51214
rect 6188 51212 6244 51268
rect 6412 51100 6468 51156
rect 5628 50988 5684 51044
rect 5964 50876 6020 50932
rect 5628 49868 5684 49924
rect 5628 49138 5684 49140
rect 5628 49086 5630 49138
rect 5630 49086 5682 49138
rect 5682 49086 5684 49138
rect 5628 49084 5684 49086
rect 5740 48802 5796 48804
rect 5740 48750 5742 48802
rect 5742 48750 5794 48802
rect 5794 48750 5796 48802
rect 5740 48748 5796 48750
rect 5852 48524 5908 48580
rect 5852 48354 5908 48356
rect 5852 48302 5854 48354
rect 5854 48302 5906 48354
rect 5906 48302 5908 48354
rect 5852 48300 5908 48302
rect 5516 47628 5572 47684
rect 5180 46732 5236 46788
rect 5404 46620 5460 46676
rect 5516 46844 5572 46900
rect 4844 46396 4900 46452
rect 4614 46282 4670 46284
rect 4614 46230 4616 46282
rect 4616 46230 4668 46282
rect 4668 46230 4670 46282
rect 4614 46228 4670 46230
rect 4718 46282 4774 46284
rect 4718 46230 4720 46282
rect 4720 46230 4772 46282
rect 4772 46230 4774 46282
rect 4718 46228 4774 46230
rect 4822 46282 4878 46284
rect 4822 46230 4824 46282
rect 4824 46230 4876 46282
rect 4876 46230 4878 46282
rect 4822 46228 4878 46230
rect 5180 45666 5236 45668
rect 5180 45614 5182 45666
rect 5182 45614 5234 45666
rect 5234 45614 5236 45666
rect 5180 45612 5236 45614
rect 5180 45388 5236 45444
rect 4620 45164 4676 45220
rect 4844 44994 4900 44996
rect 4844 44942 4846 44994
rect 4846 44942 4898 44994
rect 4898 44942 4900 44994
rect 4844 44940 4900 44942
rect 4614 44714 4670 44716
rect 4614 44662 4616 44714
rect 4616 44662 4668 44714
rect 4668 44662 4670 44714
rect 4614 44660 4670 44662
rect 4718 44714 4774 44716
rect 4718 44662 4720 44714
rect 4720 44662 4772 44714
rect 4772 44662 4774 44714
rect 4718 44660 4774 44662
rect 4822 44714 4878 44716
rect 4822 44662 4824 44714
rect 4824 44662 4876 44714
rect 4876 44662 4878 44714
rect 4822 44660 4878 44662
rect 4172 43596 4228 43652
rect 4396 43484 4452 43540
rect 5180 44098 5236 44100
rect 5180 44046 5182 44098
rect 5182 44046 5234 44098
rect 5234 44046 5236 44098
rect 5180 44044 5236 44046
rect 4614 43146 4670 43148
rect 4614 43094 4616 43146
rect 4616 43094 4668 43146
rect 4668 43094 4670 43146
rect 4614 43092 4670 43094
rect 4718 43146 4774 43148
rect 4718 43094 4720 43146
rect 4720 43094 4772 43146
rect 4772 43094 4774 43146
rect 4718 43092 4774 43094
rect 4822 43146 4878 43148
rect 4822 43094 4824 43146
rect 4824 43094 4876 43146
rect 4876 43094 4878 43146
rect 4822 43092 4878 43094
rect 4956 42812 5012 42868
rect 4620 42588 4676 42644
rect 4172 41970 4228 41972
rect 4172 41918 4174 41970
rect 4174 41918 4226 41970
rect 4226 41918 4228 41970
rect 4172 41916 4228 41918
rect 4844 42028 4900 42084
rect 5740 47180 5796 47236
rect 5852 47068 5908 47124
rect 5852 46844 5908 46900
rect 5740 45330 5796 45332
rect 5740 45278 5742 45330
rect 5742 45278 5794 45330
rect 5794 45278 5796 45330
rect 5740 45276 5796 45278
rect 6188 50594 6244 50596
rect 6188 50542 6190 50594
rect 6190 50542 6242 50594
rect 6242 50542 6244 50594
rect 6188 50540 6244 50542
rect 7308 53788 7364 53844
rect 7644 53452 7700 53508
rect 7644 52556 7700 52612
rect 7532 52332 7588 52388
rect 7196 51100 7252 51156
rect 7756 51602 7812 51604
rect 7756 51550 7758 51602
rect 7758 51550 7810 51602
rect 7810 51550 7812 51602
rect 7756 51548 7812 51550
rect 8016 59610 8072 59612
rect 8016 59558 8018 59610
rect 8018 59558 8070 59610
rect 8070 59558 8072 59610
rect 8016 59556 8072 59558
rect 8120 59610 8176 59612
rect 8120 59558 8122 59610
rect 8122 59558 8174 59610
rect 8174 59558 8176 59610
rect 8120 59556 8176 59558
rect 8224 59610 8280 59612
rect 8224 59558 8226 59610
rect 8226 59558 8278 59610
rect 8278 59558 8280 59610
rect 8224 59556 8280 59558
rect 8016 58042 8072 58044
rect 8016 57990 8018 58042
rect 8018 57990 8070 58042
rect 8070 57990 8072 58042
rect 8016 57988 8072 57990
rect 8120 58042 8176 58044
rect 8120 57990 8122 58042
rect 8122 57990 8174 58042
rect 8174 57990 8176 58042
rect 8120 57988 8176 57990
rect 8224 58042 8280 58044
rect 8224 57990 8226 58042
rect 8226 57990 8278 58042
rect 8278 57990 8280 58042
rect 8224 57988 8280 57990
rect 8540 60114 8596 60116
rect 8540 60062 8542 60114
rect 8542 60062 8594 60114
rect 8594 60062 8596 60114
rect 8540 60060 8596 60062
rect 8540 59388 8596 59444
rect 8876 66780 8932 66836
rect 8988 66444 9044 66500
rect 8988 64818 9044 64820
rect 8988 64766 8990 64818
rect 8990 64766 9042 64818
rect 9042 64766 9044 64818
rect 8988 64764 9044 64766
rect 9772 70588 9828 70644
rect 9772 70418 9828 70420
rect 9772 70366 9774 70418
rect 9774 70366 9826 70418
rect 9826 70366 9828 70418
rect 9772 70364 9828 70366
rect 9660 67788 9716 67844
rect 9660 67618 9716 67620
rect 9660 67566 9662 67618
rect 9662 67566 9714 67618
rect 9714 67566 9716 67618
rect 9660 67564 9716 67566
rect 9660 66946 9716 66948
rect 9660 66894 9662 66946
rect 9662 66894 9714 66946
rect 9714 66894 9716 66946
rect 9660 66892 9716 66894
rect 9548 66444 9604 66500
rect 10108 72604 10164 72660
rect 9996 72268 10052 72324
rect 10108 71932 10164 71988
rect 12012 85596 12068 85652
rect 11418 85482 11474 85484
rect 11418 85430 11420 85482
rect 11420 85430 11472 85482
rect 11472 85430 11474 85482
rect 11418 85428 11474 85430
rect 11522 85482 11578 85484
rect 11522 85430 11524 85482
rect 11524 85430 11576 85482
rect 11576 85430 11578 85482
rect 11522 85428 11578 85430
rect 11626 85482 11682 85484
rect 11626 85430 11628 85482
rect 11628 85430 11680 85482
rect 11680 85430 11682 85482
rect 11626 85428 11682 85430
rect 11452 84364 11508 84420
rect 11116 84306 11172 84308
rect 11116 84254 11118 84306
rect 11118 84254 11170 84306
rect 11170 84254 11172 84306
rect 11116 84252 11172 84254
rect 11418 83914 11474 83916
rect 11418 83862 11420 83914
rect 11420 83862 11472 83914
rect 11472 83862 11474 83914
rect 11418 83860 11474 83862
rect 11522 83914 11578 83916
rect 11522 83862 11524 83914
rect 11524 83862 11576 83914
rect 11576 83862 11578 83914
rect 11522 83860 11578 83862
rect 11626 83914 11682 83916
rect 11626 83862 11628 83914
rect 11628 83862 11680 83914
rect 11680 83862 11682 83914
rect 11626 83860 11682 83862
rect 11564 83244 11620 83300
rect 11228 83020 11284 83076
rect 11116 82962 11172 82964
rect 11116 82910 11118 82962
rect 11118 82910 11170 82962
rect 11170 82910 11172 82962
rect 11116 82908 11172 82910
rect 11418 82346 11474 82348
rect 11418 82294 11420 82346
rect 11420 82294 11472 82346
rect 11472 82294 11474 82346
rect 11418 82292 11474 82294
rect 11522 82346 11578 82348
rect 11522 82294 11524 82346
rect 11524 82294 11576 82346
rect 11576 82294 11578 82346
rect 11522 82292 11578 82294
rect 11626 82346 11682 82348
rect 11626 82294 11628 82346
rect 11628 82294 11680 82346
rect 11680 82294 11682 82346
rect 11626 82292 11682 82294
rect 11004 81564 11060 81620
rect 11564 81730 11620 81732
rect 11564 81678 11566 81730
rect 11566 81678 11618 81730
rect 11618 81678 11620 81730
rect 11564 81676 11620 81678
rect 12124 82460 12180 82516
rect 11564 81340 11620 81396
rect 11340 81228 11396 81284
rect 11116 80946 11172 80948
rect 11116 80894 11118 80946
rect 11118 80894 11170 80946
rect 11170 80894 11172 80946
rect 11116 80892 11172 80894
rect 11418 80778 11474 80780
rect 11418 80726 11420 80778
rect 11420 80726 11472 80778
rect 11472 80726 11474 80778
rect 11418 80724 11474 80726
rect 11522 80778 11578 80780
rect 11522 80726 11524 80778
rect 11524 80726 11576 80778
rect 11576 80726 11578 80778
rect 11522 80724 11578 80726
rect 11626 80778 11682 80780
rect 11626 80726 11628 80778
rect 11628 80726 11680 80778
rect 11680 80726 11682 80778
rect 11626 80724 11682 80726
rect 11676 79602 11732 79604
rect 11676 79550 11678 79602
rect 11678 79550 11730 79602
rect 11730 79550 11732 79602
rect 11676 79548 11732 79550
rect 12012 79548 12068 79604
rect 12012 79324 12068 79380
rect 11418 79210 11474 79212
rect 11418 79158 11420 79210
rect 11420 79158 11472 79210
rect 11472 79158 11474 79210
rect 11418 79156 11474 79158
rect 11522 79210 11578 79212
rect 11522 79158 11524 79210
rect 11524 79158 11576 79210
rect 11576 79158 11578 79210
rect 11522 79156 11578 79158
rect 11626 79210 11682 79212
rect 11626 79158 11628 79210
rect 11628 79158 11680 79210
rect 11680 79158 11682 79210
rect 11626 79156 11682 79158
rect 11004 78876 11060 78932
rect 11004 78652 11060 78708
rect 11418 77642 11474 77644
rect 11418 77590 11420 77642
rect 11420 77590 11472 77642
rect 11472 77590 11474 77642
rect 11418 77588 11474 77590
rect 11522 77642 11578 77644
rect 11522 77590 11524 77642
rect 11524 77590 11576 77642
rect 11576 77590 11578 77642
rect 11522 77588 11578 77590
rect 11626 77642 11682 77644
rect 11626 77590 11628 77642
rect 11628 77590 11680 77642
rect 11680 77590 11682 77642
rect 11626 77588 11682 77590
rect 11228 76972 11284 77028
rect 11116 76690 11172 76692
rect 11116 76638 11118 76690
rect 11118 76638 11170 76690
rect 11170 76638 11172 76690
rect 11116 76636 11172 76638
rect 11900 77084 11956 77140
rect 11788 76466 11844 76468
rect 11788 76414 11790 76466
rect 11790 76414 11842 76466
rect 11842 76414 11844 76466
rect 11788 76412 11844 76414
rect 11004 76242 11060 76244
rect 11004 76190 11006 76242
rect 11006 76190 11058 76242
rect 11058 76190 11060 76242
rect 11004 76188 11060 76190
rect 11418 76074 11474 76076
rect 11418 76022 11420 76074
rect 11420 76022 11472 76074
rect 11472 76022 11474 76074
rect 11418 76020 11474 76022
rect 11522 76074 11578 76076
rect 11522 76022 11524 76074
rect 11524 76022 11576 76074
rect 11576 76022 11578 76074
rect 11522 76020 11578 76022
rect 11626 76074 11682 76076
rect 11626 76022 11628 76074
rect 11628 76022 11680 76074
rect 11680 76022 11682 76074
rect 11626 76020 11682 76022
rect 11004 75516 11060 75572
rect 11228 75122 11284 75124
rect 11228 75070 11230 75122
rect 11230 75070 11282 75122
rect 11282 75070 11284 75122
rect 11228 75068 11284 75070
rect 11452 74898 11508 74900
rect 11452 74846 11454 74898
rect 11454 74846 11506 74898
rect 11506 74846 11508 74898
rect 11452 74844 11508 74846
rect 10444 72156 10500 72212
rect 10556 71986 10612 71988
rect 10556 71934 10558 71986
rect 10558 71934 10610 71986
rect 10610 71934 10612 71986
rect 10556 71932 10612 71934
rect 9996 70364 10052 70420
rect 10892 73500 10948 73556
rect 10668 71148 10724 71204
rect 10780 71762 10836 71764
rect 10780 71710 10782 71762
rect 10782 71710 10834 71762
rect 10834 71710 10836 71762
rect 10780 71708 10836 71710
rect 10444 70924 10500 70980
rect 10780 70700 10836 70756
rect 10444 70588 10500 70644
rect 10220 70418 10276 70420
rect 10220 70366 10222 70418
rect 10222 70366 10274 70418
rect 10274 70366 10276 70418
rect 10220 70364 10276 70366
rect 10668 70364 10724 70420
rect 9996 69132 10052 69188
rect 10444 69186 10500 69188
rect 10444 69134 10446 69186
rect 10446 69134 10498 69186
rect 10498 69134 10500 69186
rect 10444 69132 10500 69134
rect 10668 67730 10724 67732
rect 10668 67678 10670 67730
rect 10670 67678 10722 67730
rect 10722 67678 10724 67730
rect 10668 67676 10724 67678
rect 9212 64316 9268 64372
rect 8876 63810 8932 63812
rect 8876 63758 8878 63810
rect 8878 63758 8930 63810
rect 8930 63758 8932 63810
rect 8876 63756 8932 63758
rect 8988 63868 9044 63924
rect 8764 62748 8820 62804
rect 8764 62300 8820 62356
rect 8988 60732 9044 60788
rect 8988 60172 9044 60228
rect 9100 59276 9156 59332
rect 8876 58268 8932 58324
rect 9100 58380 9156 58436
rect 8988 57932 9044 57988
rect 8540 57874 8596 57876
rect 8540 57822 8542 57874
rect 8542 57822 8594 57874
rect 8594 57822 8596 57874
rect 8540 57820 8596 57822
rect 8428 56700 8484 56756
rect 8016 56474 8072 56476
rect 8016 56422 8018 56474
rect 8018 56422 8070 56474
rect 8070 56422 8072 56474
rect 8016 56420 8072 56422
rect 8120 56474 8176 56476
rect 8120 56422 8122 56474
rect 8122 56422 8174 56474
rect 8174 56422 8176 56474
rect 8120 56420 8176 56422
rect 8224 56474 8280 56476
rect 8224 56422 8226 56474
rect 8226 56422 8278 56474
rect 8278 56422 8280 56474
rect 8224 56420 8280 56422
rect 8652 56364 8708 56420
rect 8988 56252 9044 56308
rect 8092 55804 8148 55860
rect 7980 55410 8036 55412
rect 7980 55358 7982 55410
rect 7982 55358 8034 55410
rect 8034 55358 8036 55410
rect 7980 55356 8036 55358
rect 8876 56194 8932 56196
rect 8876 56142 8878 56194
rect 8878 56142 8930 56194
rect 8930 56142 8932 56194
rect 8876 56140 8932 56142
rect 8652 55356 8708 55412
rect 8016 54906 8072 54908
rect 8016 54854 8018 54906
rect 8018 54854 8070 54906
rect 8070 54854 8072 54906
rect 8016 54852 8072 54854
rect 8120 54906 8176 54908
rect 8120 54854 8122 54906
rect 8122 54854 8174 54906
rect 8174 54854 8176 54906
rect 8120 54852 8176 54854
rect 8224 54906 8280 54908
rect 8224 54854 8226 54906
rect 8226 54854 8278 54906
rect 8278 54854 8280 54906
rect 8224 54852 8280 54854
rect 8204 54124 8260 54180
rect 8540 54236 8596 54292
rect 8016 53338 8072 53340
rect 8016 53286 8018 53338
rect 8018 53286 8070 53338
rect 8070 53286 8072 53338
rect 8016 53284 8072 53286
rect 8120 53338 8176 53340
rect 8120 53286 8122 53338
rect 8122 53286 8174 53338
rect 8174 53286 8176 53338
rect 8120 53284 8176 53286
rect 8224 53338 8280 53340
rect 8224 53286 8226 53338
rect 8226 53286 8278 53338
rect 8278 53286 8280 53338
rect 8224 53284 8280 53286
rect 8092 52444 8148 52500
rect 8428 52220 8484 52276
rect 8540 53842 8596 53844
rect 8540 53790 8542 53842
rect 8542 53790 8594 53842
rect 8594 53790 8596 53842
rect 8540 53788 8596 53790
rect 8428 51996 8484 52052
rect 8016 51770 8072 51772
rect 8016 51718 8018 51770
rect 8018 51718 8070 51770
rect 8070 51718 8072 51770
rect 8016 51716 8072 51718
rect 8120 51770 8176 51772
rect 8120 51718 8122 51770
rect 8122 51718 8174 51770
rect 8174 51718 8176 51770
rect 8120 51716 8176 51718
rect 8224 51770 8280 51772
rect 8224 51718 8226 51770
rect 8226 51718 8278 51770
rect 8278 51718 8280 51770
rect 8224 51716 8280 51718
rect 9212 58322 9268 58324
rect 9212 58270 9214 58322
rect 9214 58270 9266 58322
rect 9266 58270 9268 58322
rect 9212 58268 9268 58270
rect 9212 54796 9268 54852
rect 8988 53676 9044 53732
rect 9100 54012 9156 54068
rect 8764 53564 8820 53620
rect 8652 53340 8708 53396
rect 9100 53228 9156 53284
rect 9212 53004 9268 53060
rect 9212 52668 9268 52724
rect 8988 51772 9044 51828
rect 8764 51660 8820 51716
rect 8988 51436 9044 51492
rect 8764 51378 8820 51380
rect 8764 51326 8766 51378
rect 8766 51326 8818 51378
rect 8818 51326 8820 51378
rect 8764 51324 8820 51326
rect 8204 51266 8260 51268
rect 8204 51214 8206 51266
rect 8206 51214 8258 51266
rect 8258 51214 8260 51266
rect 8204 51212 8260 51214
rect 7868 50988 7924 51044
rect 8652 50988 8708 51044
rect 6860 50652 6916 50708
rect 6748 50428 6804 50484
rect 6300 49980 6356 50036
rect 6188 49532 6244 49588
rect 6524 49756 6580 49812
rect 6412 48748 6468 48804
rect 6300 46562 6356 46564
rect 6300 46510 6302 46562
rect 6302 46510 6354 46562
rect 6354 46510 6356 46562
rect 6300 46508 6356 46510
rect 6524 48524 6580 48580
rect 6748 50204 6804 50260
rect 6412 46172 6468 46228
rect 6412 45778 6468 45780
rect 6412 45726 6414 45778
rect 6414 45726 6466 45778
rect 6466 45726 6468 45778
rect 6412 45724 6468 45726
rect 6188 45500 6244 45556
rect 6524 45612 6580 45668
rect 6076 45388 6132 45444
rect 5964 45052 6020 45108
rect 6300 44940 6356 44996
rect 6188 44546 6244 44548
rect 6188 44494 6190 44546
rect 6190 44494 6242 44546
rect 6242 44494 6244 44546
rect 6188 44492 6244 44494
rect 5068 41916 5124 41972
rect 4614 41578 4670 41580
rect 4614 41526 4616 41578
rect 4616 41526 4668 41578
rect 4668 41526 4670 41578
rect 4614 41524 4670 41526
rect 4718 41578 4774 41580
rect 4718 41526 4720 41578
rect 4720 41526 4772 41578
rect 4772 41526 4774 41578
rect 4718 41524 4774 41526
rect 4822 41578 4878 41580
rect 4822 41526 4824 41578
rect 4824 41526 4876 41578
rect 4876 41526 4878 41578
rect 4822 41524 4878 41526
rect 5628 44210 5684 44212
rect 5628 44158 5630 44210
rect 5630 44158 5682 44210
rect 5682 44158 5684 44210
rect 5628 44156 5684 44158
rect 4956 41244 5012 41300
rect 4284 40572 4340 40628
rect 4396 40962 4452 40964
rect 4396 40910 4398 40962
rect 4398 40910 4450 40962
rect 4450 40910 4452 40962
rect 4396 40908 4452 40910
rect 3164 40012 3220 40068
rect 2268 39058 2324 39060
rect 2268 39006 2270 39058
rect 2270 39006 2322 39058
rect 2322 39006 2324 39058
rect 2268 39004 2324 39006
rect 3500 39004 3556 39060
rect 3612 38892 3668 38948
rect 2380 38274 2436 38276
rect 2380 38222 2382 38274
rect 2382 38222 2434 38274
rect 2434 38222 2436 38274
rect 2380 38220 2436 38222
rect 2380 38050 2436 38052
rect 2380 37998 2382 38050
rect 2382 37998 2434 38050
rect 2434 37998 2436 38050
rect 2380 37996 2436 37998
rect 3388 38050 3444 38052
rect 3388 37998 3390 38050
rect 3390 37998 3442 38050
rect 3442 37998 3444 38050
rect 3388 37996 3444 37998
rect 2492 36988 2548 37044
rect 2940 37938 2996 37940
rect 2940 37886 2942 37938
rect 2942 37886 2994 37938
rect 2994 37886 2996 37938
rect 2940 37884 2996 37886
rect 3276 36652 3332 36708
rect 2940 35026 2996 35028
rect 2940 34974 2942 35026
rect 2942 34974 2994 35026
rect 2994 34974 2996 35026
rect 2940 34972 2996 34974
rect 2380 33516 2436 33572
rect 2156 31836 2212 31892
rect 1708 31666 1764 31668
rect 1708 31614 1710 31666
rect 1710 31614 1762 31666
rect 1762 31614 1764 31666
rect 1708 31612 1764 31614
rect 2044 31724 2100 31780
rect 1708 28924 1764 28980
rect 1708 28588 1764 28644
rect 2604 33458 2660 33460
rect 2604 33406 2606 33458
rect 2606 33406 2658 33458
rect 2658 33406 2660 33458
rect 2604 33404 2660 33406
rect 3500 34914 3556 34916
rect 3500 34862 3502 34914
rect 3502 34862 3554 34914
rect 3554 34862 3556 34914
rect 3500 34860 3556 34862
rect 2716 33292 2772 33348
rect 3388 33516 3444 33572
rect 2604 32786 2660 32788
rect 2604 32734 2606 32786
rect 2606 32734 2658 32786
rect 2658 32734 2660 32786
rect 2604 32732 2660 32734
rect 3052 32786 3108 32788
rect 3052 32734 3054 32786
rect 3054 32734 3106 32786
rect 3106 32734 3108 32786
rect 3052 32732 3108 32734
rect 3500 33458 3556 33460
rect 3500 33406 3502 33458
rect 3502 33406 3554 33458
rect 3554 33406 3556 33458
rect 3500 33404 3556 33406
rect 3388 33346 3444 33348
rect 3388 33294 3390 33346
rect 3390 33294 3442 33346
rect 3442 33294 3444 33346
rect 3388 33292 3444 33294
rect 3388 31948 3444 32004
rect 2828 31778 2884 31780
rect 2828 31726 2830 31778
rect 2830 31726 2882 31778
rect 2882 31726 2884 31778
rect 2828 31724 2884 31726
rect 1820 28028 1876 28084
rect 2492 29314 2548 29316
rect 2492 29262 2494 29314
rect 2494 29262 2546 29314
rect 2546 29262 2548 29314
rect 2492 29260 2548 29262
rect 2156 27804 2212 27860
rect 2716 28754 2772 28756
rect 2716 28702 2718 28754
rect 2718 28702 2770 28754
rect 2770 28702 2772 28754
rect 2716 28700 2772 28702
rect 2604 28588 2660 28644
rect 3164 29260 3220 29316
rect 4060 39788 4116 39844
rect 3948 38892 4004 38948
rect 3948 37996 4004 38052
rect 3724 36428 3780 36484
rect 3836 37826 3892 37828
rect 3836 37774 3838 37826
rect 3838 37774 3890 37826
rect 3890 37774 3892 37826
rect 3836 37772 3892 37774
rect 4172 37996 4228 38052
rect 3948 36594 4004 36596
rect 3948 36542 3950 36594
rect 3950 36542 4002 36594
rect 4002 36542 4004 36594
rect 3948 36540 4004 36542
rect 4060 37100 4116 37156
rect 3948 36204 4004 36260
rect 3836 35980 3892 36036
rect 3836 34300 3892 34356
rect 3724 32732 3780 32788
rect 3612 29986 3668 29988
rect 3612 29934 3614 29986
rect 3614 29934 3666 29986
rect 3666 29934 3668 29986
rect 3612 29932 3668 29934
rect 3612 29538 3668 29540
rect 3612 29486 3614 29538
rect 3614 29486 3666 29538
rect 3666 29486 3668 29538
rect 3612 29484 3668 29486
rect 2940 28642 2996 28644
rect 2940 28590 2942 28642
rect 2942 28590 2994 28642
rect 2994 28590 2996 28642
rect 2940 28588 2996 28590
rect 3500 28754 3556 28756
rect 3500 28702 3502 28754
rect 3502 28702 3554 28754
rect 3554 28702 3556 28754
rect 3500 28700 3556 28702
rect 2940 28028 2996 28084
rect 2828 27132 2884 27188
rect 1708 26796 1764 26852
rect 1708 26236 1764 26292
rect 1932 26348 1988 26404
rect 1820 23548 1876 23604
rect 1708 23324 1764 23380
rect 2044 25452 2100 25508
rect 2940 26796 2996 26852
rect 4060 35196 4116 35252
rect 3948 32450 4004 32452
rect 3948 32398 3950 32450
rect 3950 32398 4002 32450
rect 4002 32398 4004 32450
rect 3948 32396 4004 32398
rect 4060 31836 4116 31892
rect 4172 31164 4228 31220
rect 3948 30156 4004 30212
rect 4396 39900 4452 39956
rect 4614 40010 4670 40012
rect 4614 39958 4616 40010
rect 4616 39958 4668 40010
rect 4668 39958 4670 40010
rect 4614 39956 4670 39958
rect 4718 40010 4774 40012
rect 4718 39958 4720 40010
rect 4720 39958 4772 40010
rect 4772 39958 4774 40010
rect 4718 39956 4774 39958
rect 4822 40010 4878 40012
rect 4822 39958 4824 40010
rect 4824 39958 4876 40010
rect 4876 39958 4878 40010
rect 4822 39956 4878 39958
rect 4396 39676 4452 39732
rect 4620 39004 4676 39060
rect 4614 38442 4670 38444
rect 4614 38390 4616 38442
rect 4616 38390 4668 38442
rect 4668 38390 4670 38442
rect 4614 38388 4670 38390
rect 4718 38442 4774 38444
rect 4718 38390 4720 38442
rect 4720 38390 4772 38442
rect 4772 38390 4774 38442
rect 4718 38388 4774 38390
rect 4822 38442 4878 38444
rect 4822 38390 4824 38442
rect 4824 38390 4876 38442
rect 4876 38390 4878 38442
rect 4822 38388 4878 38390
rect 4396 37772 4452 37828
rect 4396 37324 4452 37380
rect 5068 39730 5124 39732
rect 5068 39678 5070 39730
rect 5070 39678 5122 39730
rect 5122 39678 5124 39730
rect 5068 39676 5124 39678
rect 5180 39228 5236 39284
rect 5068 38946 5124 38948
rect 5068 38894 5070 38946
rect 5070 38894 5122 38946
rect 5122 38894 5124 38946
rect 5068 38892 5124 38894
rect 5292 38892 5348 38948
rect 4956 37324 5012 37380
rect 5068 37154 5124 37156
rect 5068 37102 5070 37154
rect 5070 37102 5122 37154
rect 5122 37102 5124 37154
rect 5068 37100 5124 37102
rect 4732 36988 4788 37044
rect 4614 36874 4670 36876
rect 4614 36822 4616 36874
rect 4616 36822 4668 36874
rect 4668 36822 4670 36874
rect 4614 36820 4670 36822
rect 4718 36874 4774 36876
rect 4718 36822 4720 36874
rect 4720 36822 4772 36874
rect 4772 36822 4774 36874
rect 4718 36820 4774 36822
rect 4822 36874 4878 36876
rect 4822 36822 4824 36874
rect 4824 36822 4876 36874
rect 4876 36822 4878 36874
rect 4822 36820 4878 36822
rect 4396 36258 4452 36260
rect 4396 36206 4398 36258
rect 4398 36206 4450 36258
rect 4450 36206 4452 36258
rect 4396 36204 4452 36206
rect 4732 36482 4788 36484
rect 4732 36430 4734 36482
rect 4734 36430 4786 36482
rect 4786 36430 4788 36482
rect 4732 36428 4788 36430
rect 5068 36428 5124 36484
rect 5180 36540 5236 36596
rect 4956 36370 5012 36372
rect 4956 36318 4958 36370
rect 4958 36318 5010 36370
rect 5010 36318 5012 36370
rect 4956 36316 5012 36318
rect 4956 36092 5012 36148
rect 4844 35810 4900 35812
rect 4844 35758 4846 35810
rect 4846 35758 4898 35810
rect 4898 35758 4900 35810
rect 4844 35756 4900 35758
rect 4614 35306 4670 35308
rect 4614 35254 4616 35306
rect 4616 35254 4668 35306
rect 4668 35254 4670 35306
rect 4614 35252 4670 35254
rect 4718 35306 4774 35308
rect 4718 35254 4720 35306
rect 4720 35254 4772 35306
rect 4772 35254 4774 35306
rect 4718 35252 4774 35254
rect 4822 35306 4878 35308
rect 4822 35254 4824 35306
rect 4824 35254 4876 35306
rect 4876 35254 4878 35306
rect 4822 35252 4878 35254
rect 4844 35084 4900 35140
rect 4620 34860 4676 34916
rect 4614 33738 4670 33740
rect 4614 33686 4616 33738
rect 4616 33686 4668 33738
rect 4668 33686 4670 33738
rect 4614 33684 4670 33686
rect 4718 33738 4774 33740
rect 4718 33686 4720 33738
rect 4720 33686 4772 33738
rect 4772 33686 4774 33738
rect 4718 33684 4774 33686
rect 4822 33738 4878 33740
rect 4822 33686 4824 33738
rect 4824 33686 4876 33738
rect 4876 33686 4878 33738
rect 4822 33684 4878 33686
rect 4844 33404 4900 33460
rect 4396 33122 4452 33124
rect 4396 33070 4398 33122
rect 4398 33070 4450 33122
rect 4450 33070 4452 33122
rect 4396 33068 4452 33070
rect 5180 33516 5236 33572
rect 5180 33292 5236 33348
rect 4844 32396 4900 32452
rect 4614 32170 4670 32172
rect 4614 32118 4616 32170
rect 4616 32118 4668 32170
rect 4668 32118 4670 32170
rect 4614 32116 4670 32118
rect 4718 32170 4774 32172
rect 4718 32118 4720 32170
rect 4720 32118 4772 32170
rect 4772 32118 4774 32170
rect 4718 32116 4774 32118
rect 4822 32170 4878 32172
rect 4822 32118 4824 32170
rect 4824 32118 4876 32170
rect 4876 32118 4878 32170
rect 4822 32116 4878 32118
rect 4620 31948 4676 32004
rect 4732 31778 4788 31780
rect 4732 31726 4734 31778
rect 4734 31726 4786 31778
rect 4786 31726 4788 31778
rect 4732 31724 4788 31726
rect 5180 31500 5236 31556
rect 5068 31276 5124 31332
rect 4614 30602 4670 30604
rect 4614 30550 4616 30602
rect 4616 30550 4668 30602
rect 4668 30550 4670 30602
rect 4614 30548 4670 30550
rect 4718 30602 4774 30604
rect 4718 30550 4720 30602
rect 4720 30550 4772 30602
rect 4772 30550 4774 30602
rect 4718 30548 4774 30550
rect 4822 30602 4878 30604
rect 4822 30550 4824 30602
rect 4824 30550 4876 30602
rect 4876 30550 4878 30602
rect 4822 30548 4878 30550
rect 4732 30434 4788 30436
rect 4732 30382 4734 30434
rect 4734 30382 4786 30434
rect 4786 30382 4788 30434
rect 4732 30380 4788 30382
rect 3948 29820 4004 29876
rect 3388 26402 3444 26404
rect 3388 26350 3390 26402
rect 3390 26350 3442 26402
rect 3442 26350 3444 26402
rect 3388 26348 3444 26350
rect 4396 29986 4452 29988
rect 4396 29934 4398 29986
rect 4398 29934 4450 29986
rect 4450 29934 4452 29986
rect 4396 29932 4452 29934
rect 5180 30268 5236 30324
rect 5068 30210 5124 30212
rect 5068 30158 5070 30210
rect 5070 30158 5122 30210
rect 5122 30158 5124 30210
rect 5068 30156 5124 30158
rect 4732 29820 4788 29876
rect 5180 29932 5236 29988
rect 4284 29372 4340 29428
rect 4284 28754 4340 28756
rect 4284 28702 4286 28754
rect 4286 28702 4338 28754
rect 4338 28702 4340 28754
rect 4284 28700 4340 28702
rect 4172 28642 4228 28644
rect 4172 28590 4174 28642
rect 4174 28590 4226 28642
rect 4226 28590 4228 28642
rect 4172 28588 4228 28590
rect 3612 27132 3668 27188
rect 4284 28476 4340 28532
rect 3276 25564 3332 25620
rect 2716 25452 2772 25508
rect 2268 25340 2324 25396
rect 2044 23378 2100 23380
rect 2044 23326 2046 23378
rect 2046 23326 2098 23378
rect 2098 23326 2100 23378
rect 2044 23324 2100 23326
rect 1820 22092 1876 22148
rect 1820 20914 1876 20916
rect 1820 20862 1822 20914
rect 1822 20862 1874 20914
rect 1874 20862 1876 20914
rect 1820 20860 1876 20862
rect 2044 20748 2100 20804
rect 1708 18172 1764 18228
rect 2940 24722 2996 24724
rect 2940 24670 2942 24722
rect 2942 24670 2994 24722
rect 2994 24670 2996 24722
rect 2940 24668 2996 24670
rect 3500 25506 3556 25508
rect 3500 25454 3502 25506
rect 3502 25454 3554 25506
rect 3554 25454 3556 25506
rect 3500 25452 3556 25454
rect 3612 24834 3668 24836
rect 3612 24782 3614 24834
rect 3614 24782 3666 24834
rect 3666 24782 3668 24834
rect 3612 24780 3668 24782
rect 3500 24722 3556 24724
rect 3500 24670 3502 24722
rect 3502 24670 3554 24722
rect 3554 24670 3556 24722
rect 3500 24668 3556 24670
rect 3836 27186 3892 27188
rect 3836 27134 3838 27186
rect 3838 27134 3890 27186
rect 3890 27134 3892 27186
rect 3836 27132 3892 27134
rect 4284 26348 4340 26404
rect 4060 25506 4116 25508
rect 4060 25454 4062 25506
rect 4062 25454 4114 25506
rect 4114 25454 4116 25506
rect 4060 25452 4116 25454
rect 4614 29034 4670 29036
rect 4614 28982 4616 29034
rect 4616 28982 4668 29034
rect 4668 28982 4670 29034
rect 4614 28980 4670 28982
rect 4718 29034 4774 29036
rect 4718 28982 4720 29034
rect 4720 28982 4772 29034
rect 4772 28982 4774 29034
rect 4718 28980 4774 28982
rect 4822 29034 4878 29036
rect 4822 28982 4824 29034
rect 4824 28982 4876 29034
rect 4876 28982 4878 29034
rect 4822 28980 4878 28982
rect 4620 28700 4676 28756
rect 5068 28082 5124 28084
rect 5068 28030 5070 28082
rect 5070 28030 5122 28082
rect 5122 28030 5124 28082
rect 5068 28028 5124 28030
rect 4614 27466 4670 27468
rect 4614 27414 4616 27466
rect 4616 27414 4668 27466
rect 4668 27414 4670 27466
rect 4614 27412 4670 27414
rect 4718 27466 4774 27468
rect 4718 27414 4720 27466
rect 4720 27414 4772 27466
rect 4772 27414 4774 27466
rect 4718 27412 4774 27414
rect 4822 27466 4878 27468
rect 4822 27414 4824 27466
rect 4824 27414 4876 27466
rect 4876 27414 4878 27466
rect 4822 27412 4878 27414
rect 5068 27186 5124 27188
rect 5068 27134 5070 27186
rect 5070 27134 5122 27186
rect 5122 27134 5124 27186
rect 5068 27132 5124 27134
rect 5852 44210 5908 44212
rect 5852 44158 5854 44210
rect 5854 44158 5906 44210
rect 5906 44158 5908 44210
rect 5852 44156 5908 44158
rect 5740 42028 5796 42084
rect 5628 41244 5684 41300
rect 5516 40572 5572 40628
rect 5516 40012 5572 40068
rect 5628 39788 5684 39844
rect 5628 39228 5684 39284
rect 6860 49138 6916 49140
rect 6860 49086 6862 49138
rect 6862 49086 6914 49138
rect 6914 49086 6916 49138
rect 6860 49084 6916 49086
rect 6972 48972 7028 49028
rect 7084 49756 7140 49812
rect 6860 48300 6916 48356
rect 6748 47292 6804 47348
rect 6860 46508 6916 46564
rect 6748 45612 6804 45668
rect 7084 47852 7140 47908
rect 7084 47068 7140 47124
rect 7084 46060 7140 46116
rect 6972 45388 7028 45444
rect 6636 45276 6692 45332
rect 7308 50594 7364 50596
rect 7308 50542 7310 50594
rect 7310 50542 7362 50594
rect 7362 50542 7364 50594
rect 7308 50540 7364 50542
rect 7868 50540 7924 50596
rect 7532 50428 7588 50484
rect 8016 50202 8072 50204
rect 8016 50150 8018 50202
rect 8018 50150 8070 50202
rect 8070 50150 8072 50202
rect 8016 50148 8072 50150
rect 8120 50202 8176 50204
rect 8120 50150 8122 50202
rect 8122 50150 8174 50202
rect 8174 50150 8176 50202
rect 8120 50148 8176 50150
rect 8224 50202 8280 50204
rect 8224 50150 8226 50202
rect 8226 50150 8278 50202
rect 8278 50150 8280 50202
rect 8224 50148 8280 50150
rect 8428 50204 8484 50260
rect 8204 49868 8260 49924
rect 7868 49196 7924 49252
rect 8652 49810 8708 49812
rect 8652 49758 8654 49810
rect 8654 49758 8706 49810
rect 8706 49758 8708 49810
rect 8652 49756 8708 49758
rect 8764 50204 8820 50260
rect 8428 49084 8484 49140
rect 7308 48972 7364 49028
rect 8016 48634 8072 48636
rect 8016 48582 8018 48634
rect 8018 48582 8070 48634
rect 8070 48582 8072 48634
rect 8016 48580 8072 48582
rect 8120 48634 8176 48636
rect 8120 48582 8122 48634
rect 8122 48582 8174 48634
rect 8174 48582 8176 48634
rect 8120 48580 8176 48582
rect 8224 48634 8280 48636
rect 8224 48582 8226 48634
rect 8226 48582 8278 48634
rect 8278 48582 8280 48634
rect 8224 48580 8280 48582
rect 8652 49196 8708 49252
rect 7532 48466 7588 48468
rect 7532 48414 7534 48466
rect 7534 48414 7586 48466
rect 7586 48414 7588 48466
rect 7532 48412 7588 48414
rect 8316 48242 8372 48244
rect 8316 48190 8318 48242
rect 8318 48190 8370 48242
rect 8370 48190 8372 48242
rect 8316 48188 8372 48190
rect 8540 48300 8596 48356
rect 7420 48076 7476 48132
rect 8428 48130 8484 48132
rect 8428 48078 8430 48130
rect 8430 48078 8482 48130
rect 8482 48078 8484 48130
rect 8428 48076 8484 48078
rect 8204 47628 8260 47684
rect 8016 47066 8072 47068
rect 8016 47014 8018 47066
rect 8018 47014 8070 47066
rect 8070 47014 8072 47066
rect 8016 47012 8072 47014
rect 8120 47066 8176 47068
rect 8120 47014 8122 47066
rect 8122 47014 8174 47066
rect 8174 47014 8176 47066
rect 8120 47012 8176 47014
rect 8224 47066 8280 47068
rect 8224 47014 8226 47066
rect 8226 47014 8278 47066
rect 8278 47014 8280 47066
rect 8224 47012 8280 47014
rect 7308 46060 7364 46116
rect 7980 45890 8036 45892
rect 7980 45838 7982 45890
rect 7982 45838 8034 45890
rect 8034 45838 8036 45890
rect 7980 45836 8036 45838
rect 8204 45836 8260 45892
rect 8204 45612 8260 45668
rect 8428 45724 8484 45780
rect 7756 45500 7812 45556
rect 8016 45498 8072 45500
rect 7196 45388 7252 45444
rect 8016 45446 8018 45498
rect 8018 45446 8070 45498
rect 8070 45446 8072 45498
rect 8016 45444 8072 45446
rect 8120 45498 8176 45500
rect 8120 45446 8122 45498
rect 8122 45446 8174 45498
rect 8174 45446 8176 45498
rect 8120 45444 8176 45446
rect 8224 45498 8280 45500
rect 8224 45446 8226 45498
rect 8226 45446 8278 45498
rect 8278 45446 8280 45498
rect 8428 45500 8484 45556
rect 8224 45444 8280 45446
rect 7084 45276 7140 45332
rect 8428 45276 8484 45332
rect 7196 44994 7252 44996
rect 7196 44942 7198 44994
rect 7198 44942 7250 44994
rect 7250 44942 7252 44994
rect 7196 44940 7252 44942
rect 7532 44940 7588 44996
rect 6748 44828 6804 44884
rect 6748 44604 6804 44660
rect 7532 44604 7588 44660
rect 6300 44156 6356 44212
rect 6188 44044 6244 44100
rect 6076 42866 6132 42868
rect 6076 42814 6078 42866
rect 6078 42814 6130 42866
rect 6130 42814 6132 42866
rect 6076 42812 6132 42814
rect 6412 43484 6468 43540
rect 6524 41132 6580 41188
rect 6300 41074 6356 41076
rect 6300 41022 6302 41074
rect 6302 41022 6354 41074
rect 6354 41022 6356 41074
rect 6300 41020 6356 41022
rect 6524 40460 6580 40516
rect 6412 39676 6468 39732
rect 6076 38892 6132 38948
rect 5516 37212 5572 37268
rect 5740 38444 5796 38500
rect 5404 33292 5460 33348
rect 5404 31500 5460 31556
rect 4956 26290 5012 26292
rect 4956 26238 4958 26290
rect 4958 26238 5010 26290
rect 5010 26238 5012 26290
rect 4956 26236 5012 26238
rect 4614 25898 4670 25900
rect 4614 25846 4616 25898
rect 4616 25846 4668 25898
rect 4668 25846 4670 25898
rect 4614 25844 4670 25846
rect 4718 25898 4774 25900
rect 4718 25846 4720 25898
rect 4720 25846 4772 25898
rect 4772 25846 4774 25898
rect 4718 25844 4774 25846
rect 4822 25898 4878 25900
rect 4822 25846 4824 25898
rect 4824 25846 4876 25898
rect 4876 25846 4878 25898
rect 4822 25844 4878 25846
rect 5068 25618 5124 25620
rect 5068 25566 5070 25618
rect 5070 25566 5122 25618
rect 5122 25566 5124 25618
rect 5068 25564 5124 25566
rect 4620 25394 4676 25396
rect 4620 25342 4622 25394
rect 4622 25342 4674 25394
rect 4674 25342 4676 25394
rect 4620 25340 4676 25342
rect 5628 36540 5684 36596
rect 5628 35756 5684 35812
rect 6412 37490 6468 37492
rect 6412 37438 6414 37490
rect 6414 37438 6466 37490
rect 6466 37438 6468 37490
rect 6412 37436 6468 37438
rect 5852 37212 5908 37268
rect 5964 37154 6020 37156
rect 5964 37102 5966 37154
rect 5966 37102 6018 37154
rect 6018 37102 6020 37154
rect 5964 37100 6020 37102
rect 5964 36482 6020 36484
rect 5964 36430 5966 36482
rect 5966 36430 6018 36482
rect 6018 36430 6020 36482
rect 5964 36428 6020 36430
rect 6412 36204 6468 36260
rect 5516 30828 5572 30884
rect 6860 44492 6916 44548
rect 6748 44322 6804 44324
rect 6748 44270 6750 44322
rect 6750 44270 6802 44322
rect 6802 44270 6804 44322
rect 6748 44268 6804 44270
rect 7308 44268 7364 44324
rect 6748 43932 6804 43988
rect 7196 42924 7252 42980
rect 6972 42476 7028 42532
rect 6860 41804 6916 41860
rect 7196 41020 7252 41076
rect 7644 44268 7700 44324
rect 7868 44492 7924 44548
rect 7980 44994 8036 44996
rect 7980 44942 7982 44994
rect 7982 44942 8034 44994
rect 8034 44942 8036 44994
rect 7980 44940 8036 44942
rect 7980 44380 8036 44436
rect 8652 44940 8708 44996
rect 7868 44210 7924 44212
rect 7868 44158 7870 44210
rect 7870 44158 7922 44210
rect 7922 44158 7924 44210
rect 7868 44156 7924 44158
rect 7756 42700 7812 42756
rect 7532 41692 7588 41748
rect 7308 40796 7364 40852
rect 7644 41186 7700 41188
rect 7644 41134 7646 41186
rect 7646 41134 7698 41186
rect 7698 41134 7700 41186
rect 7644 41132 7700 41134
rect 7196 40012 7252 40068
rect 7756 40684 7812 40740
rect 8016 43930 8072 43932
rect 8016 43878 8018 43930
rect 8018 43878 8070 43930
rect 8070 43878 8072 43930
rect 8016 43876 8072 43878
rect 8120 43930 8176 43932
rect 8120 43878 8122 43930
rect 8122 43878 8174 43930
rect 8174 43878 8176 43930
rect 8120 43876 8176 43878
rect 8224 43930 8280 43932
rect 8224 43878 8226 43930
rect 8226 43878 8278 43930
rect 8278 43878 8280 43930
rect 8224 43876 8280 43878
rect 9100 51212 9156 51268
rect 9100 48860 9156 48916
rect 9212 48076 9268 48132
rect 9212 47852 9268 47908
rect 9100 47628 9156 47684
rect 8988 46562 9044 46564
rect 8988 46510 8990 46562
rect 8990 46510 9042 46562
rect 9042 46510 9044 46562
rect 8988 46508 9044 46510
rect 9212 45836 9268 45892
rect 9212 45388 9268 45444
rect 9100 45106 9156 45108
rect 9100 45054 9102 45106
rect 9102 45054 9154 45106
rect 9154 45054 9156 45106
rect 9100 45052 9156 45054
rect 8988 44940 9044 44996
rect 8876 44380 8932 44436
rect 8652 44044 8708 44100
rect 8540 43484 8596 43540
rect 8652 43820 8708 43876
rect 8540 42924 8596 42980
rect 8016 42362 8072 42364
rect 8016 42310 8018 42362
rect 8018 42310 8070 42362
rect 8070 42310 8072 42362
rect 8016 42308 8072 42310
rect 8120 42362 8176 42364
rect 8120 42310 8122 42362
rect 8122 42310 8174 42362
rect 8174 42310 8176 42362
rect 8120 42308 8176 42310
rect 8224 42362 8280 42364
rect 8224 42310 8226 42362
rect 8226 42310 8278 42362
rect 8278 42310 8280 42362
rect 8224 42308 8280 42310
rect 8316 42140 8372 42196
rect 8092 41970 8148 41972
rect 8092 41918 8094 41970
rect 8094 41918 8146 41970
rect 8146 41918 8148 41970
rect 8092 41916 8148 41918
rect 8092 41132 8148 41188
rect 8016 40794 8072 40796
rect 8016 40742 8018 40794
rect 8018 40742 8070 40794
rect 8070 40742 8072 40794
rect 8016 40740 8072 40742
rect 8120 40794 8176 40796
rect 8120 40742 8122 40794
rect 8122 40742 8174 40794
rect 8174 40742 8176 40794
rect 8120 40740 8176 40742
rect 8224 40794 8280 40796
rect 8224 40742 8226 40794
rect 8226 40742 8278 40794
rect 8278 40742 8280 40794
rect 8224 40740 8280 40742
rect 7756 40460 7812 40516
rect 8204 40514 8260 40516
rect 8204 40462 8206 40514
rect 8206 40462 8258 40514
rect 8258 40462 8260 40514
rect 8204 40460 8260 40462
rect 7756 40012 7812 40068
rect 7756 38892 7812 38948
rect 7644 38780 7700 38836
rect 6748 38332 6804 38388
rect 7420 38332 7476 38388
rect 7196 37660 7252 37716
rect 6972 36876 7028 36932
rect 6860 36706 6916 36708
rect 6860 36654 6862 36706
rect 6862 36654 6914 36706
rect 6914 36654 6916 36706
rect 6860 36652 6916 36654
rect 6748 36316 6804 36372
rect 6748 36092 6804 36148
rect 6524 33740 6580 33796
rect 5964 33628 6020 33684
rect 6300 32396 6356 32452
rect 5852 31276 5908 31332
rect 5628 30940 5684 30996
rect 5852 30268 5908 30324
rect 5740 30156 5796 30212
rect 5516 29932 5572 29988
rect 5628 29484 5684 29540
rect 6300 31218 6356 31220
rect 6300 31166 6302 31218
rect 6302 31166 6354 31218
rect 6354 31166 6356 31218
rect 6300 31164 6356 31166
rect 6748 33404 6804 33460
rect 7420 37436 7476 37492
rect 7532 37772 7588 37828
rect 7532 37378 7588 37380
rect 7532 37326 7534 37378
rect 7534 37326 7586 37378
rect 7586 37326 7588 37378
rect 7532 37324 7588 37326
rect 7420 37212 7476 37268
rect 7084 34972 7140 35028
rect 7196 34354 7252 34356
rect 7196 34302 7198 34354
rect 7198 34302 7250 34354
rect 7250 34302 7252 34354
rect 7196 34300 7252 34302
rect 7084 33628 7140 33684
rect 7532 34018 7588 34020
rect 7532 33966 7534 34018
rect 7534 33966 7586 34018
rect 7586 33966 7588 34018
rect 7532 33964 7588 33966
rect 6972 32620 7028 32676
rect 7196 31612 7252 31668
rect 7196 31164 7252 31220
rect 6412 30828 6468 30884
rect 6188 30098 6244 30100
rect 6188 30046 6190 30098
rect 6190 30046 6242 30098
rect 6242 30046 6244 30098
rect 6188 30044 6244 30046
rect 5964 28028 6020 28084
rect 5852 27804 5908 27860
rect 5628 27186 5684 27188
rect 5628 27134 5630 27186
rect 5630 27134 5682 27186
rect 5682 27134 5684 27186
rect 5628 27132 5684 27134
rect 5852 27020 5908 27076
rect 5740 25340 5796 25396
rect 3164 23378 3220 23380
rect 3164 23326 3166 23378
rect 3166 23326 3218 23378
rect 3218 23326 3220 23378
rect 3164 23324 3220 23326
rect 4508 24892 4564 24948
rect 2716 21980 2772 22036
rect 2380 21196 2436 21252
rect 4060 24722 4116 24724
rect 4060 24670 4062 24722
rect 4062 24670 4114 24722
rect 4114 24670 4116 24722
rect 4060 24668 4116 24670
rect 4956 24892 5012 24948
rect 4614 24330 4670 24332
rect 4614 24278 4616 24330
rect 4616 24278 4668 24330
rect 4668 24278 4670 24330
rect 4614 24276 4670 24278
rect 4718 24330 4774 24332
rect 4718 24278 4720 24330
rect 4720 24278 4772 24330
rect 4772 24278 4774 24330
rect 4718 24276 4774 24278
rect 4822 24330 4878 24332
rect 4822 24278 4824 24330
rect 4824 24278 4876 24330
rect 4876 24278 4878 24330
rect 4822 24276 4878 24278
rect 4060 24108 4116 24164
rect 4620 24108 4676 24164
rect 5740 24892 5796 24948
rect 4956 23548 5012 23604
rect 4620 23378 4676 23380
rect 4620 23326 4622 23378
rect 4622 23326 4674 23378
rect 4674 23326 4676 23378
rect 4620 23324 4676 23326
rect 3276 22204 3332 22260
rect 3052 21196 3108 21252
rect 1820 15538 1876 15540
rect 1820 15486 1822 15538
rect 1822 15486 1874 15538
rect 1874 15486 1876 15538
rect 1820 15484 1876 15486
rect 1708 12796 1764 12852
rect 1820 10780 1876 10836
rect 2716 20802 2772 20804
rect 2716 20750 2718 20802
rect 2718 20750 2770 20802
rect 2770 20750 2772 20802
rect 2716 20748 2772 20750
rect 2716 19964 2772 20020
rect 3500 21980 3556 22036
rect 4508 23154 4564 23156
rect 4508 23102 4510 23154
rect 4510 23102 4562 23154
rect 4562 23102 4564 23154
rect 4508 23100 4564 23102
rect 4614 22762 4670 22764
rect 4614 22710 4616 22762
rect 4616 22710 4668 22762
rect 4668 22710 4670 22762
rect 4614 22708 4670 22710
rect 4718 22762 4774 22764
rect 4718 22710 4720 22762
rect 4720 22710 4772 22762
rect 4772 22710 4774 22762
rect 4718 22708 4774 22710
rect 4822 22762 4878 22764
rect 4822 22710 4824 22762
rect 4824 22710 4876 22762
rect 4876 22710 4878 22762
rect 4822 22708 4878 22710
rect 3836 22540 3892 22596
rect 4620 22540 4676 22596
rect 3724 22204 3780 22260
rect 4396 22092 4452 22148
rect 3612 21196 3668 21252
rect 4614 21194 4670 21196
rect 4614 21142 4616 21194
rect 4616 21142 4668 21194
rect 4668 21142 4670 21194
rect 4614 21140 4670 21142
rect 4718 21194 4774 21196
rect 4718 21142 4720 21194
rect 4720 21142 4772 21194
rect 4772 21142 4774 21194
rect 4718 21140 4774 21142
rect 4822 21194 4878 21196
rect 4822 21142 4824 21194
rect 4824 21142 4876 21194
rect 4876 21142 4878 21194
rect 4822 21140 4878 21142
rect 3052 20300 3108 20356
rect 3388 20300 3444 20356
rect 3276 20130 3332 20132
rect 3276 20078 3278 20130
rect 3278 20078 3330 20130
rect 3330 20078 3332 20130
rect 3276 20076 3332 20078
rect 3500 20076 3556 20132
rect 2604 18508 2660 18564
rect 2492 18172 2548 18228
rect 2044 17612 2100 17668
rect 2044 15148 2100 15204
rect 2044 14924 2100 14980
rect 2604 15148 2660 15204
rect 3948 20018 4004 20020
rect 3948 19966 3950 20018
rect 3950 19966 4002 20018
rect 4002 19966 4004 20018
rect 3948 19964 4004 19966
rect 3836 19852 3892 19908
rect 5068 20860 5124 20916
rect 4396 20076 4452 20132
rect 4956 19906 5012 19908
rect 4956 19854 4958 19906
rect 4958 19854 5010 19906
rect 5010 19854 5012 19906
rect 4956 19852 5012 19854
rect 4508 19794 4564 19796
rect 4508 19742 4510 19794
rect 4510 19742 4562 19794
rect 4562 19742 4564 19794
rect 4508 19740 4564 19742
rect 4614 19626 4670 19628
rect 4614 19574 4616 19626
rect 4616 19574 4668 19626
rect 4668 19574 4670 19626
rect 4614 19572 4670 19574
rect 4718 19626 4774 19628
rect 4718 19574 4720 19626
rect 4720 19574 4772 19626
rect 4772 19574 4774 19626
rect 4718 19572 4774 19574
rect 4822 19626 4878 19628
rect 4822 19574 4824 19626
rect 4824 19574 4876 19626
rect 4876 19574 4878 19626
rect 4822 19572 4878 19574
rect 3836 18508 3892 18564
rect 3724 18450 3780 18452
rect 3724 18398 3726 18450
rect 3726 18398 3778 18450
rect 3778 18398 3780 18450
rect 3724 18396 3780 18398
rect 2940 17612 2996 17668
rect 3052 17388 3108 17444
rect 4396 18396 4452 18452
rect 4172 17666 4228 17668
rect 4172 17614 4174 17666
rect 4174 17614 4226 17666
rect 4226 17614 4228 17666
rect 4172 17612 4228 17614
rect 3388 17442 3444 17444
rect 3388 17390 3390 17442
rect 3390 17390 3442 17442
rect 3442 17390 3444 17442
rect 3388 17388 3444 17390
rect 4956 18284 5012 18340
rect 4614 18058 4670 18060
rect 4614 18006 4616 18058
rect 4616 18006 4668 18058
rect 4668 18006 4670 18058
rect 4614 18004 4670 18006
rect 4718 18058 4774 18060
rect 4718 18006 4720 18058
rect 4720 18006 4772 18058
rect 4772 18006 4774 18058
rect 4718 18004 4774 18006
rect 4822 18058 4878 18060
rect 4822 18006 4824 18058
rect 4824 18006 4876 18058
rect 4876 18006 4878 18058
rect 4822 18004 4878 18006
rect 4614 16490 4670 16492
rect 4614 16438 4616 16490
rect 4616 16438 4668 16490
rect 4668 16438 4670 16490
rect 4614 16436 4670 16438
rect 4718 16490 4774 16492
rect 4718 16438 4720 16490
rect 4720 16438 4772 16490
rect 4772 16438 4774 16490
rect 4718 16436 4774 16438
rect 4822 16490 4878 16492
rect 4822 16438 4824 16490
rect 4824 16438 4876 16490
rect 4876 16438 4878 16490
rect 4822 16436 4878 16438
rect 2268 14700 2324 14756
rect 2380 14924 2436 14980
rect 2044 11340 2100 11396
rect 2268 13970 2324 13972
rect 2268 13918 2270 13970
rect 2270 13918 2322 13970
rect 2322 13918 2324 13970
rect 2268 13916 2324 13918
rect 2716 14924 2772 14980
rect 3500 15148 3556 15204
rect 3836 15148 3892 15204
rect 2492 14476 2548 14532
rect 2492 13804 2548 13860
rect 2828 14418 2884 14420
rect 2828 14366 2830 14418
rect 2830 14366 2882 14418
rect 2882 14366 2884 14418
rect 2828 14364 2884 14366
rect 3276 14364 3332 14420
rect 2716 13858 2772 13860
rect 2716 13806 2718 13858
rect 2718 13806 2770 13858
rect 2770 13806 2772 13858
rect 2716 13804 2772 13806
rect 3388 13916 3444 13972
rect 3612 13804 3668 13860
rect 2380 12348 2436 12404
rect 2716 12124 2772 12180
rect 2044 11170 2100 11172
rect 2044 11118 2046 11170
rect 2046 11118 2098 11170
rect 2098 11118 2100 11170
rect 2044 11116 2100 11118
rect 2268 10892 2324 10948
rect 2156 10780 2212 10836
rect 1932 9100 1988 9156
rect 2044 10220 2100 10276
rect 2156 8316 2212 8372
rect 2380 10220 2436 10276
rect 2604 10892 2660 10948
rect 2380 9154 2436 9156
rect 2380 9102 2382 9154
rect 2382 9102 2434 9154
rect 2434 9102 2436 9154
rect 2380 9100 2436 9102
rect 3052 12178 3108 12180
rect 3052 12126 3054 12178
rect 3054 12126 3106 12178
rect 3106 12126 3108 12178
rect 3052 12124 3108 12126
rect 3388 13634 3444 13636
rect 3388 13582 3390 13634
rect 3390 13582 3442 13634
rect 3442 13582 3444 13634
rect 3388 13580 3444 13582
rect 2828 11282 2884 11284
rect 2828 11230 2830 11282
rect 2830 11230 2882 11282
rect 2882 11230 2884 11282
rect 2828 11228 2884 11230
rect 2716 10108 2772 10164
rect 2604 8428 2660 8484
rect 3500 11340 3556 11396
rect 3388 10220 3444 10276
rect 2828 8316 2884 8372
rect 3164 8316 3220 8372
rect 3724 8316 3780 8372
rect 2940 7644 2996 7700
rect 2828 7532 2884 7588
rect 1708 7474 1764 7476
rect 1708 7422 1710 7474
rect 1710 7422 1762 7474
rect 1762 7422 1764 7474
rect 1708 7420 1764 7422
rect 2492 7420 2548 7476
rect 4172 13468 4228 13524
rect 4060 12402 4116 12404
rect 4060 12350 4062 12402
rect 4062 12350 4114 12402
rect 4114 12350 4116 12402
rect 4060 12348 4116 12350
rect 3948 11618 4004 11620
rect 3948 11566 3950 11618
rect 3950 11566 4002 11618
rect 4002 11566 4004 11618
rect 3948 11564 4004 11566
rect 4614 14922 4670 14924
rect 4614 14870 4616 14922
rect 4616 14870 4668 14922
rect 4668 14870 4670 14922
rect 4614 14868 4670 14870
rect 4718 14922 4774 14924
rect 4718 14870 4720 14922
rect 4720 14870 4772 14922
rect 4772 14870 4774 14922
rect 4718 14868 4774 14870
rect 4822 14922 4878 14924
rect 4822 14870 4824 14922
rect 4824 14870 4876 14922
rect 4876 14870 4878 14922
rect 4822 14868 4878 14870
rect 4620 14418 4676 14420
rect 4620 14366 4622 14418
rect 4622 14366 4674 14418
rect 4674 14366 4676 14418
rect 4620 14364 4676 14366
rect 5180 17724 5236 17780
rect 4956 14364 5012 14420
rect 5180 16828 5236 16884
rect 6636 30882 6692 30884
rect 6636 30830 6638 30882
rect 6638 30830 6690 30882
rect 6690 30830 6692 30882
rect 6636 30828 6692 30830
rect 6748 30268 6804 30324
rect 8428 40236 8484 40292
rect 8016 39226 8072 39228
rect 8016 39174 8018 39226
rect 8018 39174 8070 39226
rect 8070 39174 8072 39226
rect 8016 39172 8072 39174
rect 8120 39226 8176 39228
rect 8120 39174 8122 39226
rect 8122 39174 8174 39226
rect 8174 39174 8176 39226
rect 8120 39172 8176 39174
rect 8224 39226 8280 39228
rect 8224 39174 8226 39226
rect 8226 39174 8278 39226
rect 8278 39174 8280 39226
rect 8224 39172 8280 39174
rect 8540 40348 8596 40404
rect 8540 38892 8596 38948
rect 8428 38108 8484 38164
rect 8016 37658 8072 37660
rect 8016 37606 8018 37658
rect 8018 37606 8070 37658
rect 8070 37606 8072 37658
rect 8016 37604 8072 37606
rect 8120 37658 8176 37660
rect 8120 37606 8122 37658
rect 8122 37606 8174 37658
rect 8174 37606 8176 37658
rect 8120 37604 8176 37606
rect 8224 37658 8280 37660
rect 8224 37606 8226 37658
rect 8226 37606 8278 37658
rect 8278 37606 8280 37658
rect 8224 37604 8280 37606
rect 7980 37212 8036 37268
rect 8204 37490 8260 37492
rect 8204 37438 8206 37490
rect 8206 37438 8258 37490
rect 8258 37438 8260 37490
rect 8204 37436 8260 37438
rect 8316 37266 8372 37268
rect 8316 37214 8318 37266
rect 8318 37214 8370 37266
rect 8370 37214 8372 37266
rect 8316 37212 8372 37214
rect 8204 36988 8260 37044
rect 8204 36764 8260 36820
rect 8764 37436 8820 37492
rect 8652 37324 8708 37380
rect 8016 36090 8072 36092
rect 8016 36038 8018 36090
rect 8018 36038 8070 36090
rect 8070 36038 8072 36090
rect 8016 36036 8072 36038
rect 8120 36090 8176 36092
rect 8120 36038 8122 36090
rect 8122 36038 8174 36090
rect 8174 36038 8176 36090
rect 8120 36036 8176 36038
rect 8224 36090 8280 36092
rect 8224 36038 8226 36090
rect 8226 36038 8278 36090
rect 8278 36038 8280 36090
rect 8224 36036 8280 36038
rect 8988 40402 9044 40404
rect 8988 40350 8990 40402
rect 8990 40350 9042 40402
rect 9042 40350 9044 40402
rect 8988 40348 9044 40350
rect 9436 64764 9492 64820
rect 11116 72604 11172 72660
rect 11004 71874 11060 71876
rect 11004 71822 11006 71874
rect 11006 71822 11058 71874
rect 11058 71822 11060 71874
rect 11004 71820 11060 71822
rect 11418 74506 11474 74508
rect 11418 74454 11420 74506
rect 11420 74454 11472 74506
rect 11472 74454 11474 74506
rect 11418 74452 11474 74454
rect 11522 74506 11578 74508
rect 11522 74454 11524 74506
rect 11524 74454 11576 74506
rect 11576 74454 11578 74506
rect 11522 74452 11578 74454
rect 11626 74506 11682 74508
rect 11626 74454 11628 74506
rect 11628 74454 11680 74506
rect 11680 74454 11682 74506
rect 11626 74452 11682 74454
rect 11900 74844 11956 74900
rect 11788 74396 11844 74452
rect 11900 74508 11956 74564
rect 11788 74172 11844 74228
rect 11676 74002 11732 74004
rect 11676 73950 11678 74002
rect 11678 73950 11730 74002
rect 11730 73950 11732 74002
rect 11676 73948 11732 73950
rect 11418 72938 11474 72940
rect 11418 72886 11420 72938
rect 11420 72886 11472 72938
rect 11472 72886 11474 72938
rect 11418 72884 11474 72886
rect 11522 72938 11578 72940
rect 11522 72886 11524 72938
rect 11524 72886 11576 72938
rect 11576 72886 11578 72938
rect 11522 72884 11578 72886
rect 11626 72938 11682 72940
rect 11626 72886 11628 72938
rect 11628 72886 11680 72938
rect 11680 72886 11682 72938
rect 11626 72884 11682 72886
rect 11228 72156 11284 72212
rect 11676 72044 11732 72100
rect 11788 71932 11844 71988
rect 11564 71874 11620 71876
rect 11564 71822 11566 71874
rect 11566 71822 11618 71874
rect 11618 71822 11620 71874
rect 11564 71820 11620 71822
rect 11418 71370 11474 71372
rect 11418 71318 11420 71370
rect 11420 71318 11472 71370
rect 11472 71318 11474 71370
rect 11418 71316 11474 71318
rect 11522 71370 11578 71372
rect 11522 71318 11524 71370
rect 11524 71318 11576 71370
rect 11576 71318 11578 71370
rect 11522 71316 11578 71318
rect 11626 71370 11682 71372
rect 11626 71318 11628 71370
rect 11628 71318 11680 71370
rect 11680 71318 11682 71370
rect 11626 71316 11682 71318
rect 11228 70978 11284 70980
rect 11228 70926 11230 70978
rect 11230 70926 11282 70978
rect 11282 70926 11284 70978
rect 11228 70924 11284 70926
rect 11340 70418 11396 70420
rect 11340 70366 11342 70418
rect 11342 70366 11394 70418
rect 11394 70366 11396 70418
rect 11340 70364 11396 70366
rect 11788 70588 11844 70644
rect 10892 70252 10948 70308
rect 11418 69802 11474 69804
rect 11418 69750 11420 69802
rect 11420 69750 11472 69802
rect 11472 69750 11474 69802
rect 11418 69748 11474 69750
rect 11522 69802 11578 69804
rect 11522 69750 11524 69802
rect 11524 69750 11576 69802
rect 11576 69750 11578 69802
rect 11522 69748 11578 69750
rect 11626 69802 11682 69804
rect 11626 69750 11628 69802
rect 11628 69750 11680 69802
rect 11680 69750 11682 69802
rect 11626 69748 11682 69750
rect 12796 92316 12852 92372
rect 12684 91532 12740 91588
rect 13692 93660 13748 93716
rect 14028 93436 14084 93492
rect 13804 93212 13860 93268
rect 13580 92204 13636 92260
rect 12908 91420 12964 91476
rect 12684 90578 12740 90580
rect 12684 90526 12686 90578
rect 12686 90526 12738 90578
rect 12738 90526 12740 90578
rect 12684 90524 12740 90526
rect 13580 91420 13636 91476
rect 13692 91250 13748 91252
rect 13692 91198 13694 91250
rect 13694 91198 13746 91250
rect 13746 91198 13748 91250
rect 13692 91196 13748 91198
rect 13468 90748 13524 90804
rect 13356 90524 13412 90580
rect 12908 89964 12964 90020
rect 14028 92428 14084 92484
rect 14820 97242 14876 97244
rect 14820 97190 14822 97242
rect 14822 97190 14874 97242
rect 14874 97190 14876 97242
rect 14820 97188 14876 97190
rect 14924 97242 14980 97244
rect 14924 97190 14926 97242
rect 14926 97190 14978 97242
rect 14978 97190 14980 97242
rect 14924 97188 14980 97190
rect 15028 97242 15084 97244
rect 15028 97190 15030 97242
rect 15030 97190 15082 97242
rect 15082 97190 15084 97242
rect 15028 97188 15084 97190
rect 15148 96572 15204 96628
rect 14700 96178 14756 96180
rect 14700 96126 14702 96178
rect 14702 96126 14754 96178
rect 14754 96126 14756 96178
rect 14700 96124 14756 96126
rect 15596 97580 15652 97636
rect 16828 107772 16884 107828
rect 16492 106034 16548 106036
rect 16492 105982 16494 106034
rect 16494 105982 16546 106034
rect 16546 105982 16548 106034
rect 16492 105980 16548 105982
rect 15820 104300 15876 104356
rect 16044 104188 16100 104244
rect 15932 98140 15988 98196
rect 15932 97634 15988 97636
rect 15932 97582 15934 97634
rect 15934 97582 15986 97634
rect 15986 97582 15988 97634
rect 15932 97580 15988 97582
rect 15596 96460 15652 96516
rect 15820 96460 15876 96516
rect 15372 96348 15428 96404
rect 14812 95900 14868 95956
rect 15596 96236 15652 96292
rect 15260 95788 15316 95844
rect 14820 95674 14876 95676
rect 14820 95622 14822 95674
rect 14822 95622 14874 95674
rect 14874 95622 14876 95674
rect 14820 95620 14876 95622
rect 14924 95674 14980 95676
rect 14924 95622 14926 95674
rect 14926 95622 14978 95674
rect 14978 95622 14980 95674
rect 14924 95620 14980 95622
rect 15028 95674 15084 95676
rect 15028 95622 15030 95674
rect 15030 95622 15082 95674
rect 15082 95622 15084 95674
rect 15028 95620 15084 95622
rect 14812 95452 14868 95508
rect 14364 95004 14420 95060
rect 14364 94108 14420 94164
rect 14252 93714 14308 93716
rect 14252 93662 14254 93714
rect 14254 93662 14306 93714
rect 14306 93662 14308 93714
rect 14252 93660 14308 93662
rect 14700 94444 14756 94500
rect 15820 95842 15876 95844
rect 15820 95790 15822 95842
rect 15822 95790 15874 95842
rect 15874 95790 15876 95842
rect 15820 95788 15876 95790
rect 15932 95676 15988 95732
rect 15596 95282 15652 95284
rect 15596 95230 15598 95282
rect 15598 95230 15650 95282
rect 15650 95230 15652 95282
rect 15596 95228 15652 95230
rect 15372 95116 15428 95172
rect 15932 95004 15988 95060
rect 17500 108108 17556 108164
rect 17388 105980 17444 106036
rect 17164 103964 17220 104020
rect 16492 103180 16548 103236
rect 16828 103852 16884 103908
rect 18222 116842 18278 116844
rect 18222 116790 18224 116842
rect 18224 116790 18276 116842
rect 18276 116790 18278 116842
rect 18222 116788 18278 116790
rect 18326 116842 18382 116844
rect 18326 116790 18328 116842
rect 18328 116790 18380 116842
rect 18380 116790 18382 116842
rect 18326 116788 18382 116790
rect 18430 116842 18486 116844
rect 18430 116790 18432 116842
rect 18432 116790 18484 116842
rect 18484 116790 18486 116842
rect 18430 116788 18486 116790
rect 17724 116450 17780 116452
rect 17724 116398 17726 116450
rect 17726 116398 17778 116450
rect 17778 116398 17780 116450
rect 17724 116396 17780 116398
rect 18396 116396 18452 116452
rect 18222 115274 18278 115276
rect 18222 115222 18224 115274
rect 18224 115222 18276 115274
rect 18276 115222 18278 115274
rect 18222 115220 18278 115222
rect 18326 115274 18382 115276
rect 18326 115222 18328 115274
rect 18328 115222 18380 115274
rect 18380 115222 18382 115274
rect 18326 115220 18382 115222
rect 18430 115274 18486 115276
rect 18430 115222 18432 115274
rect 18432 115222 18484 115274
rect 18484 115222 18486 115274
rect 18430 115220 18486 115222
rect 18620 114940 18676 114996
rect 18060 114882 18116 114884
rect 18060 114830 18062 114882
rect 18062 114830 18114 114882
rect 18114 114830 18116 114882
rect 18060 114828 18116 114830
rect 20076 114828 20132 114884
rect 20076 114268 20132 114324
rect 18222 113706 18278 113708
rect 18222 113654 18224 113706
rect 18224 113654 18276 113706
rect 18276 113654 18278 113706
rect 18222 113652 18278 113654
rect 18326 113706 18382 113708
rect 18326 113654 18328 113706
rect 18328 113654 18380 113706
rect 18380 113654 18382 113706
rect 18326 113652 18382 113654
rect 18430 113706 18486 113708
rect 18430 113654 18432 113706
rect 18432 113654 18484 113706
rect 18484 113654 18486 113706
rect 18430 113652 18486 113654
rect 18620 113314 18676 113316
rect 18620 113262 18622 113314
rect 18622 113262 18674 113314
rect 18674 113262 18676 113314
rect 18620 113260 18676 113262
rect 18222 112138 18278 112140
rect 18222 112086 18224 112138
rect 18224 112086 18276 112138
rect 18276 112086 18278 112138
rect 18222 112084 18278 112086
rect 18326 112138 18382 112140
rect 18326 112086 18328 112138
rect 18328 112086 18380 112138
rect 18380 112086 18382 112138
rect 18326 112084 18382 112086
rect 18430 112138 18486 112140
rect 18430 112086 18432 112138
rect 18432 112086 18484 112138
rect 18484 112086 18486 112138
rect 18430 112084 18486 112086
rect 18172 111692 18228 111748
rect 18222 110570 18278 110572
rect 18222 110518 18224 110570
rect 18224 110518 18276 110570
rect 18276 110518 18278 110570
rect 18222 110516 18278 110518
rect 18326 110570 18382 110572
rect 18326 110518 18328 110570
rect 18328 110518 18380 110570
rect 18380 110518 18382 110570
rect 18326 110516 18382 110518
rect 18430 110570 18486 110572
rect 18430 110518 18432 110570
rect 18432 110518 18484 110570
rect 18484 110518 18486 110570
rect 18430 110516 18486 110518
rect 19180 113260 19236 113316
rect 20076 113260 20132 113316
rect 19292 112476 19348 112532
rect 19964 112530 20020 112532
rect 19964 112478 19966 112530
rect 19966 112478 20018 112530
rect 20018 112478 20020 112530
rect 19964 112476 20020 112478
rect 18956 111746 19012 111748
rect 18956 111694 18958 111746
rect 18958 111694 19010 111746
rect 19010 111694 19012 111746
rect 18956 111692 19012 111694
rect 20076 110962 20132 110964
rect 20076 110910 20078 110962
rect 20078 110910 20130 110962
rect 20130 110910 20132 110962
rect 20076 110908 20132 110910
rect 18222 109002 18278 109004
rect 18222 108950 18224 109002
rect 18224 108950 18276 109002
rect 18276 108950 18278 109002
rect 18222 108948 18278 108950
rect 18326 109002 18382 109004
rect 18326 108950 18328 109002
rect 18328 108950 18380 109002
rect 18380 108950 18382 109002
rect 18326 108948 18382 108950
rect 18430 109002 18486 109004
rect 18430 108950 18432 109002
rect 18432 108950 18484 109002
rect 18484 108950 18486 109002
rect 18430 108948 18486 108950
rect 17724 106988 17780 107044
rect 17724 106818 17780 106820
rect 17724 106766 17726 106818
rect 17726 106766 17778 106818
rect 17778 106766 17780 106818
rect 17724 106764 17780 106766
rect 17612 105532 17668 105588
rect 17500 103794 17556 103796
rect 17500 103742 17502 103794
rect 17502 103742 17554 103794
rect 17554 103742 17556 103794
rect 17500 103740 17556 103742
rect 16716 99148 16772 99204
rect 16492 97244 16548 97300
rect 16380 97132 16436 97188
rect 16380 96796 16436 96852
rect 16268 96236 16324 96292
rect 17612 102396 17668 102452
rect 17500 100716 17556 100772
rect 17388 98924 17444 98980
rect 17388 97692 17444 97748
rect 16604 96012 16660 96068
rect 16716 97020 16772 97076
rect 16940 97020 16996 97076
rect 16716 96178 16772 96180
rect 16716 96126 16718 96178
rect 16718 96126 16770 96178
rect 16770 96126 16772 96178
rect 16716 96124 16772 96126
rect 16716 95676 16772 95732
rect 16268 95452 16324 95508
rect 16828 95506 16884 95508
rect 16828 95454 16830 95506
rect 16830 95454 16882 95506
rect 16882 95454 16884 95506
rect 16828 95452 16884 95454
rect 16380 95282 16436 95284
rect 16380 95230 16382 95282
rect 16382 95230 16434 95282
rect 16434 95230 16436 95282
rect 16380 95228 16436 95230
rect 14924 94780 14980 94836
rect 15036 94444 15092 94500
rect 14588 93884 14644 93940
rect 14924 94220 14980 94276
rect 14820 94106 14876 94108
rect 14820 94054 14822 94106
rect 14822 94054 14874 94106
rect 14874 94054 14876 94106
rect 14820 94052 14876 94054
rect 14924 94106 14980 94108
rect 14924 94054 14926 94106
rect 14926 94054 14978 94106
rect 14978 94054 14980 94106
rect 14924 94052 14980 94054
rect 15028 94106 15084 94108
rect 15028 94054 15030 94106
rect 15030 94054 15082 94106
rect 15082 94054 15084 94106
rect 15028 94052 15084 94054
rect 15260 93996 15316 94052
rect 14476 93212 14532 93268
rect 14364 92818 14420 92820
rect 14364 92766 14366 92818
rect 14366 92766 14418 92818
rect 14418 92766 14420 92818
rect 14364 92764 14420 92766
rect 14364 91980 14420 92036
rect 14588 92204 14644 92260
rect 14252 91532 14308 91588
rect 14588 91532 14644 91588
rect 14820 92538 14876 92540
rect 14820 92486 14822 92538
rect 14822 92486 14874 92538
rect 14874 92486 14876 92538
rect 14820 92484 14876 92486
rect 14924 92538 14980 92540
rect 14924 92486 14926 92538
rect 14926 92486 14978 92538
rect 14978 92486 14980 92538
rect 14924 92484 14980 92486
rect 15028 92538 15084 92540
rect 15028 92486 15030 92538
rect 15030 92486 15082 92538
rect 15082 92486 15084 92538
rect 15028 92484 15084 92486
rect 15932 94444 15988 94500
rect 16156 94498 16212 94500
rect 16156 94446 16158 94498
rect 16158 94446 16210 94498
rect 16210 94446 16212 94498
rect 16156 94444 16212 94446
rect 15932 93772 15988 93828
rect 16044 94220 16100 94276
rect 16492 95004 16548 95060
rect 16380 93996 16436 94052
rect 15932 93436 15988 93492
rect 15596 93212 15652 93268
rect 16156 92988 16212 93044
rect 15932 92818 15988 92820
rect 15932 92766 15934 92818
rect 15934 92766 15986 92818
rect 15986 92766 15988 92818
rect 15932 92764 15988 92766
rect 15596 92092 15652 92148
rect 15372 91420 15428 91476
rect 15484 91980 15540 92036
rect 15484 91362 15540 91364
rect 15484 91310 15486 91362
rect 15486 91310 15538 91362
rect 15538 91310 15540 91362
rect 15484 91308 15540 91310
rect 14700 91084 14756 91140
rect 14820 90970 14876 90972
rect 14820 90918 14822 90970
rect 14822 90918 14874 90970
rect 14874 90918 14876 90970
rect 14820 90916 14876 90918
rect 14924 90970 14980 90972
rect 14924 90918 14926 90970
rect 14926 90918 14978 90970
rect 14978 90918 14980 90970
rect 14924 90916 14980 90918
rect 15028 90970 15084 90972
rect 15028 90918 15030 90970
rect 15030 90918 15082 90970
rect 15082 90918 15084 90970
rect 15028 90916 15084 90918
rect 15484 90748 15540 90804
rect 13468 89964 13524 90020
rect 13580 89852 13636 89908
rect 12684 89740 12740 89796
rect 14924 90690 14980 90692
rect 14924 90638 14926 90690
rect 14926 90638 14978 90690
rect 14978 90638 14980 90690
rect 14924 90636 14980 90638
rect 15148 90578 15204 90580
rect 15148 90526 15150 90578
rect 15150 90526 15202 90578
rect 15202 90526 15204 90578
rect 15148 90524 15204 90526
rect 15372 90412 15428 90468
rect 14588 89852 14644 89908
rect 13804 89794 13860 89796
rect 13804 89742 13806 89794
rect 13806 89742 13858 89794
rect 13858 89742 13860 89794
rect 13804 89740 13860 89742
rect 13692 89516 13748 89572
rect 13356 88898 13412 88900
rect 13356 88846 13358 88898
rect 13358 88846 13410 88898
rect 13410 88846 13412 88898
rect 13356 88844 13412 88846
rect 12908 88172 12964 88228
rect 13244 88060 13300 88116
rect 13020 87500 13076 87556
rect 13468 88226 13524 88228
rect 13468 88174 13470 88226
rect 13470 88174 13522 88226
rect 13522 88174 13524 88226
rect 13468 88172 13524 88174
rect 13244 87164 13300 87220
rect 13580 85932 13636 85988
rect 12796 84978 12852 84980
rect 12796 84926 12798 84978
rect 12798 84926 12850 84978
rect 12850 84926 12852 84978
rect 12796 84924 12852 84926
rect 12572 83298 12628 83300
rect 12572 83246 12574 83298
rect 12574 83246 12626 83298
rect 12626 83246 12628 83298
rect 12572 83244 12628 83246
rect 12796 83298 12852 83300
rect 12796 83246 12798 83298
rect 12798 83246 12850 83298
rect 12850 83246 12852 83298
rect 12796 83244 12852 83246
rect 12908 82908 12964 82964
rect 15036 89906 15092 89908
rect 15036 89854 15038 89906
rect 15038 89854 15090 89906
rect 15090 89854 15092 89906
rect 15036 89852 15092 89854
rect 14028 89682 14084 89684
rect 14028 89630 14030 89682
rect 14030 89630 14082 89682
rect 14082 89630 14084 89682
rect 14028 89628 14084 89630
rect 13804 88844 13860 88900
rect 14028 88396 14084 88452
rect 13804 87554 13860 87556
rect 13804 87502 13806 87554
rect 13806 87502 13858 87554
rect 13858 87502 13860 87554
rect 13804 87500 13860 87502
rect 13916 87330 13972 87332
rect 13916 87278 13918 87330
rect 13918 87278 13970 87330
rect 13970 87278 13972 87330
rect 13916 87276 13972 87278
rect 14252 87276 14308 87332
rect 13692 85820 13748 85876
rect 13468 83244 13524 83300
rect 16380 93660 16436 93716
rect 16380 92764 16436 92820
rect 16492 93436 16548 93492
rect 16156 92428 16212 92484
rect 15932 91980 15988 92036
rect 16268 91532 16324 91588
rect 15708 91196 15764 91252
rect 16940 92818 16996 92820
rect 16940 92766 16942 92818
rect 16942 92766 16994 92818
rect 16994 92766 16996 92818
rect 16940 92764 16996 92766
rect 16828 92540 16884 92596
rect 16828 91308 16884 91364
rect 14812 89516 14868 89572
rect 15260 89628 15316 89684
rect 14820 89402 14876 89404
rect 14820 89350 14822 89402
rect 14822 89350 14874 89402
rect 14874 89350 14876 89402
rect 14820 89348 14876 89350
rect 14924 89402 14980 89404
rect 14924 89350 14926 89402
rect 14926 89350 14978 89402
rect 14978 89350 14980 89402
rect 14924 89348 14980 89350
rect 15028 89402 15084 89404
rect 15028 89350 15030 89402
rect 15030 89350 15082 89402
rect 15082 89350 15084 89402
rect 15028 89348 15084 89350
rect 14700 88956 14756 89012
rect 15148 88732 15204 88788
rect 14820 87834 14876 87836
rect 14820 87782 14822 87834
rect 14822 87782 14874 87834
rect 14874 87782 14876 87834
rect 14820 87780 14876 87782
rect 14924 87834 14980 87836
rect 14924 87782 14926 87834
rect 14926 87782 14978 87834
rect 14978 87782 14980 87834
rect 14924 87780 14980 87782
rect 15028 87834 15084 87836
rect 15028 87782 15030 87834
rect 15030 87782 15082 87834
rect 15082 87782 15084 87834
rect 15028 87780 15084 87782
rect 14700 87612 14756 87668
rect 15036 87500 15092 87556
rect 15708 89964 15764 90020
rect 15372 88844 15428 88900
rect 15036 87164 15092 87220
rect 15036 86716 15092 86772
rect 14028 84924 14084 84980
rect 13804 84252 13860 84308
rect 14364 84364 14420 84420
rect 12684 79548 12740 79604
rect 12460 78988 12516 79044
rect 12236 78876 12292 78932
rect 12124 76300 12180 76356
rect 12124 75628 12180 75684
rect 12124 74396 12180 74452
rect 13132 79324 13188 79380
rect 13020 78764 13076 78820
rect 13244 78876 13300 78932
rect 13020 78594 13076 78596
rect 13020 78542 13022 78594
rect 13022 78542 13074 78594
rect 13074 78542 13076 78594
rect 13020 78540 13076 78542
rect 13020 77084 13076 77140
rect 12348 75122 12404 75124
rect 12348 75070 12350 75122
rect 12350 75070 12402 75122
rect 12402 75070 12404 75122
rect 12348 75068 12404 75070
rect 12796 76860 12852 76916
rect 12796 76188 12852 76244
rect 12572 74956 12628 75012
rect 12460 74844 12516 74900
rect 12348 74396 12404 74452
rect 12796 74508 12852 74564
rect 13132 76860 13188 76916
rect 13692 81676 13748 81732
rect 13468 78428 13524 78484
rect 13580 78204 13636 78260
rect 13244 76524 13300 76580
rect 13692 78818 13748 78820
rect 13692 78766 13694 78818
rect 13694 78766 13746 78818
rect 13746 78766 13748 78818
rect 13692 78764 13748 78766
rect 13916 81676 13972 81732
rect 14028 81564 14084 81620
rect 13916 78876 13972 78932
rect 13692 77868 13748 77924
rect 13468 77196 13524 77252
rect 13580 76972 13636 77028
rect 13468 75740 13524 75796
rect 13580 75404 13636 75460
rect 13580 75010 13636 75012
rect 13580 74958 13582 75010
rect 13582 74958 13634 75010
rect 13634 74958 13636 75010
rect 13580 74956 13636 74958
rect 13244 74898 13300 74900
rect 13244 74846 13246 74898
rect 13246 74846 13298 74898
rect 13298 74846 13300 74898
rect 13244 74844 13300 74846
rect 13916 76972 13972 77028
rect 14140 81004 14196 81060
rect 14252 80892 14308 80948
rect 14476 83522 14532 83524
rect 14476 83470 14478 83522
rect 14478 83470 14530 83522
rect 14530 83470 14532 83522
rect 14476 83468 14532 83470
rect 15036 86434 15092 86436
rect 15036 86382 15038 86434
rect 15038 86382 15090 86434
rect 15090 86382 15092 86434
rect 15036 86380 15092 86382
rect 14476 81730 14532 81732
rect 14476 81678 14478 81730
rect 14478 81678 14530 81730
rect 14530 81678 14532 81730
rect 14476 81676 14532 81678
rect 14364 80556 14420 80612
rect 14820 86266 14876 86268
rect 14820 86214 14822 86266
rect 14822 86214 14874 86266
rect 14874 86214 14876 86266
rect 14820 86212 14876 86214
rect 14924 86266 14980 86268
rect 14924 86214 14926 86266
rect 14926 86214 14978 86266
rect 14978 86214 14980 86266
rect 14924 86212 14980 86214
rect 15028 86266 15084 86268
rect 15028 86214 15030 86266
rect 15030 86214 15082 86266
rect 15082 86214 15084 86266
rect 15028 86212 15084 86214
rect 15708 89122 15764 89124
rect 15708 89070 15710 89122
rect 15710 89070 15762 89122
rect 15762 89070 15764 89122
rect 15708 89068 15764 89070
rect 15820 89180 15876 89236
rect 16380 90412 16436 90468
rect 16604 90466 16660 90468
rect 16604 90414 16606 90466
rect 16606 90414 16658 90466
rect 16658 90414 16660 90466
rect 16604 90412 16660 90414
rect 16828 89964 16884 90020
rect 17500 97020 17556 97076
rect 17500 96796 17556 96852
rect 17276 95452 17332 95508
rect 17164 94274 17220 94276
rect 17164 94222 17166 94274
rect 17166 94222 17218 94274
rect 17218 94222 17220 94274
rect 17164 94220 17220 94222
rect 17948 108780 18004 108836
rect 18172 108498 18228 108500
rect 18172 108446 18174 108498
rect 18174 108446 18226 108498
rect 18226 108446 18228 108498
rect 18172 108444 18228 108446
rect 18508 108220 18564 108276
rect 18222 107434 18278 107436
rect 18222 107382 18224 107434
rect 18224 107382 18276 107434
rect 18276 107382 18278 107434
rect 18222 107380 18278 107382
rect 18326 107434 18382 107436
rect 18326 107382 18328 107434
rect 18328 107382 18380 107434
rect 18380 107382 18382 107434
rect 18326 107380 18382 107382
rect 18430 107434 18486 107436
rect 18430 107382 18432 107434
rect 18432 107382 18484 107434
rect 18484 107382 18486 107434
rect 18430 107380 18486 107382
rect 18222 105866 18278 105868
rect 18222 105814 18224 105866
rect 18224 105814 18276 105866
rect 18276 105814 18278 105866
rect 18222 105812 18278 105814
rect 18326 105866 18382 105868
rect 18326 105814 18328 105866
rect 18328 105814 18380 105866
rect 18380 105814 18382 105866
rect 18326 105812 18382 105814
rect 18430 105866 18486 105868
rect 18430 105814 18432 105866
rect 18432 105814 18484 105866
rect 18484 105814 18486 105866
rect 18430 105812 18486 105814
rect 19516 109394 19572 109396
rect 19516 109342 19518 109394
rect 19518 109342 19570 109394
rect 19570 109342 19572 109394
rect 19516 109340 19572 109342
rect 18732 109228 18788 109284
rect 19180 108498 19236 108500
rect 19180 108446 19182 108498
rect 19182 108446 19234 108498
rect 19234 108446 19236 108498
rect 19180 108444 19236 108446
rect 19068 108386 19124 108388
rect 19068 108334 19070 108386
rect 19070 108334 19122 108386
rect 19122 108334 19124 108386
rect 19068 108332 19124 108334
rect 18620 104860 18676 104916
rect 18956 107436 19012 107492
rect 19852 107436 19908 107492
rect 20412 109228 20468 109284
rect 20188 108332 20244 108388
rect 19180 106764 19236 106820
rect 19964 106988 20020 107044
rect 18956 106204 19012 106260
rect 17948 104076 18004 104132
rect 18508 104636 18564 104692
rect 18222 104298 18278 104300
rect 18222 104246 18224 104298
rect 18224 104246 18276 104298
rect 18276 104246 18278 104298
rect 18222 104244 18278 104246
rect 18326 104298 18382 104300
rect 18326 104246 18328 104298
rect 18328 104246 18380 104298
rect 18380 104246 18382 104298
rect 18326 104244 18382 104246
rect 18430 104298 18486 104300
rect 18430 104246 18432 104298
rect 18432 104246 18484 104298
rect 18484 104246 18486 104298
rect 18430 104244 18486 104246
rect 18396 104076 18452 104132
rect 17836 102284 17892 102340
rect 17948 100828 18004 100884
rect 18222 102730 18278 102732
rect 18222 102678 18224 102730
rect 18224 102678 18276 102730
rect 18276 102678 18278 102730
rect 18222 102676 18278 102678
rect 18326 102730 18382 102732
rect 18326 102678 18328 102730
rect 18328 102678 18380 102730
rect 18380 102678 18382 102730
rect 18326 102676 18382 102678
rect 18430 102730 18486 102732
rect 18430 102678 18432 102730
rect 18432 102678 18484 102730
rect 18484 102678 18486 102730
rect 18430 102676 18486 102678
rect 18844 102396 18900 102452
rect 20524 108332 20580 108388
rect 20748 107826 20804 107828
rect 20748 107774 20750 107826
rect 20750 107774 20802 107826
rect 20802 107774 20804 107826
rect 20748 107772 20804 107774
rect 21624 117626 21680 117628
rect 21624 117574 21626 117626
rect 21626 117574 21678 117626
rect 21678 117574 21680 117626
rect 21624 117572 21680 117574
rect 21728 117626 21784 117628
rect 21728 117574 21730 117626
rect 21730 117574 21782 117626
rect 21782 117574 21784 117626
rect 21728 117572 21784 117574
rect 21832 117626 21888 117628
rect 21832 117574 21834 117626
rect 21834 117574 21886 117626
rect 21886 117574 21888 117626
rect 21832 117572 21888 117574
rect 21624 116058 21680 116060
rect 21624 116006 21626 116058
rect 21626 116006 21678 116058
rect 21678 116006 21680 116058
rect 21624 116004 21680 116006
rect 21728 116058 21784 116060
rect 21728 116006 21730 116058
rect 21730 116006 21782 116058
rect 21782 116006 21784 116058
rect 21728 116004 21784 116006
rect 21832 116058 21888 116060
rect 21832 116006 21834 116058
rect 21834 116006 21886 116058
rect 21886 116006 21888 116058
rect 21832 116004 21888 116006
rect 22652 114604 22708 114660
rect 21624 114490 21680 114492
rect 21624 114438 21626 114490
rect 21626 114438 21678 114490
rect 21678 114438 21680 114490
rect 21624 114436 21680 114438
rect 21728 114490 21784 114492
rect 21728 114438 21730 114490
rect 21730 114438 21782 114490
rect 21782 114438 21784 114490
rect 21728 114436 21784 114438
rect 21832 114490 21888 114492
rect 21832 114438 21834 114490
rect 21834 114438 21886 114490
rect 21886 114438 21888 114490
rect 21832 114436 21888 114438
rect 21420 114268 21476 114324
rect 22876 114380 22932 114436
rect 25026 118410 25082 118412
rect 25026 118358 25028 118410
rect 25028 118358 25080 118410
rect 25080 118358 25082 118410
rect 25026 118356 25082 118358
rect 25130 118410 25186 118412
rect 25130 118358 25132 118410
rect 25132 118358 25184 118410
rect 25184 118358 25186 118410
rect 25130 118356 25186 118358
rect 25234 118410 25290 118412
rect 25234 118358 25236 118410
rect 25236 118358 25288 118410
rect 25288 118358 25290 118410
rect 25234 118356 25290 118358
rect 24668 117180 24724 117236
rect 25340 117234 25396 117236
rect 25340 117182 25342 117234
rect 25342 117182 25394 117234
rect 25394 117182 25396 117234
rect 25340 117180 25396 117182
rect 24108 114658 24164 114660
rect 24108 114606 24110 114658
rect 24110 114606 24162 114658
rect 24162 114606 24164 114658
rect 24108 114604 24164 114606
rect 24108 114380 24164 114436
rect 21624 112922 21680 112924
rect 21624 112870 21626 112922
rect 21626 112870 21678 112922
rect 21678 112870 21680 112922
rect 21624 112868 21680 112870
rect 21728 112922 21784 112924
rect 21728 112870 21730 112922
rect 21730 112870 21782 112922
rect 21782 112870 21784 112922
rect 21728 112868 21784 112870
rect 21832 112922 21888 112924
rect 21832 112870 21834 112922
rect 21834 112870 21886 112922
rect 21886 112870 21888 112922
rect 21832 112868 21888 112870
rect 21624 111354 21680 111356
rect 21624 111302 21626 111354
rect 21626 111302 21678 111354
rect 21678 111302 21680 111354
rect 21624 111300 21680 111302
rect 21728 111354 21784 111356
rect 21728 111302 21730 111354
rect 21730 111302 21782 111354
rect 21782 111302 21784 111354
rect 21728 111300 21784 111302
rect 21832 111354 21888 111356
rect 21832 111302 21834 111354
rect 21834 111302 21886 111354
rect 21886 111302 21888 111354
rect 21832 111300 21888 111302
rect 21420 110908 21476 110964
rect 21624 109786 21680 109788
rect 21624 109734 21626 109786
rect 21626 109734 21678 109786
rect 21678 109734 21680 109786
rect 21624 109732 21680 109734
rect 21728 109786 21784 109788
rect 21728 109734 21730 109786
rect 21730 109734 21782 109786
rect 21782 109734 21784 109786
rect 21728 109732 21784 109734
rect 21832 109786 21888 109788
rect 21832 109734 21834 109786
rect 21834 109734 21886 109786
rect 21886 109734 21888 109786
rect 21832 109732 21888 109734
rect 21420 108498 21476 108500
rect 21420 108446 21422 108498
rect 21422 108446 21474 108498
rect 21474 108446 21476 108498
rect 21420 108444 21476 108446
rect 21868 108386 21924 108388
rect 21868 108334 21870 108386
rect 21870 108334 21922 108386
rect 21922 108334 21924 108386
rect 21868 108332 21924 108334
rect 22204 108332 22260 108388
rect 22316 108668 22372 108724
rect 21624 108218 21680 108220
rect 21624 108166 21626 108218
rect 21626 108166 21678 108218
rect 21678 108166 21680 108218
rect 21624 108164 21680 108166
rect 21728 108218 21784 108220
rect 21728 108166 21730 108218
rect 21730 108166 21782 108218
rect 21782 108166 21784 108218
rect 21728 108164 21784 108166
rect 21832 108218 21888 108220
rect 21832 108166 21834 108218
rect 21834 108166 21886 108218
rect 21886 108166 21888 108218
rect 21832 108164 21888 108166
rect 21644 107548 21700 107604
rect 23436 111692 23492 111748
rect 23212 108668 23268 108724
rect 22428 107548 22484 107604
rect 23100 108610 23156 108612
rect 23100 108558 23102 108610
rect 23102 108558 23154 108610
rect 23154 108558 23156 108610
rect 23100 108556 23156 108558
rect 21624 106650 21680 106652
rect 21624 106598 21626 106650
rect 21626 106598 21678 106650
rect 21678 106598 21680 106650
rect 21624 106596 21680 106598
rect 21728 106650 21784 106652
rect 21728 106598 21730 106650
rect 21730 106598 21782 106650
rect 21782 106598 21784 106650
rect 21728 106596 21784 106598
rect 21832 106650 21888 106652
rect 21832 106598 21834 106650
rect 21834 106598 21886 106650
rect 21886 106598 21888 106650
rect 21832 106596 21888 106598
rect 20188 105532 20244 105588
rect 21308 106482 21364 106484
rect 21308 106430 21310 106482
rect 21310 106430 21362 106482
rect 21362 106430 21364 106482
rect 21308 106428 21364 106430
rect 22316 106428 22372 106484
rect 22204 106258 22260 106260
rect 22204 106206 22206 106258
rect 22206 106206 22258 106258
rect 22258 106206 22260 106258
rect 22204 106204 22260 106206
rect 20636 105644 20692 105700
rect 22540 106092 22596 106148
rect 23324 106146 23380 106148
rect 23324 106094 23326 106146
rect 23326 106094 23378 106146
rect 23378 106094 23380 106146
rect 23324 106092 23380 106094
rect 20300 105308 20356 105364
rect 19068 104802 19124 104804
rect 19068 104750 19070 104802
rect 19070 104750 19122 104802
rect 19122 104750 19124 104802
rect 19068 104748 19124 104750
rect 20300 104748 20356 104804
rect 18844 101276 18900 101332
rect 19740 102226 19796 102228
rect 19740 102174 19742 102226
rect 19742 102174 19794 102226
rect 19794 102174 19796 102226
rect 19740 102172 19796 102174
rect 18222 101162 18278 101164
rect 18222 101110 18224 101162
rect 18224 101110 18276 101162
rect 18276 101110 18278 101162
rect 18222 101108 18278 101110
rect 18326 101162 18382 101164
rect 18326 101110 18328 101162
rect 18328 101110 18380 101162
rect 18380 101110 18382 101162
rect 18326 101108 18382 101110
rect 18430 101162 18486 101164
rect 18430 101110 18432 101162
rect 18432 101110 18484 101162
rect 18484 101110 18486 101162
rect 18430 101108 18486 101110
rect 18284 100940 18340 100996
rect 18732 100828 18788 100884
rect 18222 99594 18278 99596
rect 18222 99542 18224 99594
rect 18224 99542 18276 99594
rect 18276 99542 18278 99594
rect 18222 99540 18278 99542
rect 18326 99594 18382 99596
rect 18326 99542 18328 99594
rect 18328 99542 18380 99594
rect 18380 99542 18382 99594
rect 18326 99540 18382 99542
rect 18430 99594 18486 99596
rect 18430 99542 18432 99594
rect 18432 99542 18484 99594
rect 18484 99542 18486 99594
rect 18430 99540 18486 99542
rect 18060 99036 18116 99092
rect 18172 99372 18228 99428
rect 17836 98924 17892 98980
rect 17948 98700 18004 98756
rect 19404 100940 19460 100996
rect 18844 99484 18900 99540
rect 19180 99202 19236 99204
rect 19180 99150 19182 99202
rect 19182 99150 19234 99202
rect 19234 99150 19236 99202
rect 19180 99148 19236 99150
rect 19740 99148 19796 99204
rect 20636 102956 20692 103012
rect 20188 102508 20244 102564
rect 21308 105362 21364 105364
rect 21308 105310 21310 105362
rect 21310 105310 21362 105362
rect 21362 105310 21364 105362
rect 21308 105308 21364 105310
rect 22204 105586 22260 105588
rect 22204 105534 22206 105586
rect 22206 105534 22258 105586
rect 22258 105534 22260 105586
rect 22204 105532 22260 105534
rect 21624 105082 21680 105084
rect 21624 105030 21626 105082
rect 21626 105030 21678 105082
rect 21678 105030 21680 105082
rect 21624 105028 21680 105030
rect 21728 105082 21784 105084
rect 21728 105030 21730 105082
rect 21730 105030 21782 105082
rect 21782 105030 21784 105082
rect 21728 105028 21784 105030
rect 21832 105082 21888 105084
rect 21832 105030 21834 105082
rect 21834 105030 21886 105082
rect 21886 105030 21888 105082
rect 21832 105028 21888 105030
rect 21624 103514 21680 103516
rect 21624 103462 21626 103514
rect 21626 103462 21678 103514
rect 21678 103462 21680 103514
rect 21624 103460 21680 103462
rect 21728 103514 21784 103516
rect 21728 103462 21730 103514
rect 21730 103462 21782 103514
rect 21782 103462 21784 103514
rect 21728 103460 21784 103462
rect 21832 103514 21888 103516
rect 21832 103462 21834 103514
rect 21834 103462 21886 103514
rect 21886 103462 21888 103514
rect 21832 103460 21888 103462
rect 22316 104300 22372 104356
rect 23212 105308 23268 105364
rect 23436 104188 23492 104244
rect 23324 103346 23380 103348
rect 23324 103294 23326 103346
rect 23326 103294 23378 103346
rect 23378 103294 23380 103346
rect 23324 103292 23380 103294
rect 24108 113314 24164 113316
rect 24108 113262 24110 113314
rect 24110 113262 24162 113314
rect 24162 113262 24164 113314
rect 24108 113260 24164 113262
rect 24108 111746 24164 111748
rect 24108 111694 24110 111746
rect 24110 111694 24162 111746
rect 24162 111694 24164 111746
rect 24108 111692 24164 111694
rect 23996 108332 24052 108388
rect 23772 106146 23828 106148
rect 23772 106094 23774 106146
rect 23774 106094 23826 106146
rect 23826 106094 23828 106146
rect 23772 106092 23828 106094
rect 23884 105362 23940 105364
rect 23884 105310 23886 105362
rect 23886 105310 23938 105362
rect 23938 105310 23940 105362
rect 23884 105308 23940 105310
rect 23660 104300 23716 104356
rect 23772 104188 23828 104244
rect 22428 103180 22484 103236
rect 21756 102508 21812 102564
rect 22540 103068 22596 103124
rect 22988 103010 23044 103012
rect 22988 102958 22990 103010
rect 22990 102958 23042 103010
rect 23042 102958 23044 103010
rect 22988 102956 23044 102958
rect 23660 102956 23716 103012
rect 20076 100770 20132 100772
rect 20076 100718 20078 100770
rect 20078 100718 20130 100770
rect 20130 100718 20132 100770
rect 20076 100716 20132 100718
rect 19964 99372 20020 99428
rect 19292 99036 19348 99092
rect 17948 98530 18004 98532
rect 17948 98478 17950 98530
rect 17950 98478 18002 98530
rect 18002 98478 18004 98530
rect 17948 98476 18004 98478
rect 18284 98418 18340 98420
rect 18284 98366 18286 98418
rect 18286 98366 18338 98418
rect 18338 98366 18340 98418
rect 18284 98364 18340 98366
rect 18620 98140 18676 98196
rect 19180 98588 19236 98644
rect 18222 98026 18278 98028
rect 18222 97974 18224 98026
rect 18224 97974 18276 98026
rect 18276 97974 18278 98026
rect 18222 97972 18278 97974
rect 18326 98026 18382 98028
rect 18326 97974 18328 98026
rect 18328 97974 18380 98026
rect 18380 97974 18382 98026
rect 18326 97972 18382 97974
rect 18430 98026 18486 98028
rect 18430 97974 18432 98026
rect 18432 97974 18484 98026
rect 18484 97974 18486 98026
rect 18430 97972 18486 97974
rect 18508 97580 18564 97636
rect 18172 97468 18228 97524
rect 17948 97132 18004 97188
rect 18396 97020 18452 97076
rect 18732 97244 18788 97300
rect 17948 96796 18004 96852
rect 19516 98978 19572 98980
rect 19516 98926 19518 98978
rect 19518 98926 19570 98978
rect 19570 98926 19572 98978
rect 19516 98924 19572 98926
rect 20076 98978 20132 98980
rect 20076 98926 20078 98978
rect 20078 98926 20130 98978
rect 20130 98926 20132 98978
rect 20076 98924 20132 98926
rect 20188 98418 20244 98420
rect 20188 98366 20190 98418
rect 20190 98366 20242 98418
rect 20242 98366 20244 98418
rect 20188 98364 20244 98366
rect 18956 97522 19012 97524
rect 18956 97470 18958 97522
rect 18958 97470 19010 97522
rect 19010 97470 19012 97522
rect 18956 97468 19012 97470
rect 18844 97020 18900 97076
rect 17836 96738 17892 96740
rect 17836 96686 17838 96738
rect 17838 96686 17890 96738
rect 17890 96686 17892 96738
rect 17836 96684 17892 96686
rect 18222 96458 18278 96460
rect 18222 96406 18224 96458
rect 18224 96406 18276 96458
rect 18276 96406 18278 96458
rect 18222 96404 18278 96406
rect 18326 96458 18382 96460
rect 18326 96406 18328 96458
rect 18328 96406 18380 96458
rect 18380 96406 18382 96458
rect 18326 96404 18382 96406
rect 18430 96458 18486 96460
rect 18430 96406 18432 96458
rect 18432 96406 18484 96458
rect 18484 96406 18486 96458
rect 18430 96404 18486 96406
rect 17724 96012 17780 96068
rect 17612 95282 17668 95284
rect 17612 95230 17614 95282
rect 17614 95230 17666 95282
rect 17666 95230 17668 95282
rect 17612 95228 17668 95230
rect 17388 95116 17444 95172
rect 17500 94892 17556 94948
rect 17164 92652 17220 92708
rect 17276 92876 17332 92932
rect 17052 89852 17108 89908
rect 17164 92428 17220 92484
rect 16156 88956 16212 89012
rect 16380 89516 16436 89572
rect 16716 89292 16772 89348
rect 15484 88060 15540 88116
rect 15372 86828 15428 86884
rect 15484 87612 15540 87668
rect 16044 88172 16100 88228
rect 16828 89010 16884 89012
rect 16828 88958 16830 89010
rect 16830 88958 16882 89010
rect 16882 88958 16884 89010
rect 16828 88956 16884 88958
rect 17500 93996 17556 94052
rect 17612 93714 17668 93716
rect 17612 93662 17614 93714
rect 17614 93662 17666 93714
rect 17666 93662 17668 93714
rect 17612 93660 17668 93662
rect 17612 93212 17668 93268
rect 18396 95004 18452 95060
rect 18222 94890 18278 94892
rect 18222 94838 18224 94890
rect 18224 94838 18276 94890
rect 18276 94838 18278 94890
rect 18222 94836 18278 94838
rect 18326 94890 18382 94892
rect 18326 94838 18328 94890
rect 18328 94838 18380 94890
rect 18380 94838 18382 94890
rect 18326 94836 18382 94838
rect 18430 94890 18486 94892
rect 18430 94838 18432 94890
rect 18432 94838 18484 94890
rect 18484 94838 18486 94890
rect 18430 94836 18486 94838
rect 18396 94668 18452 94724
rect 18172 94444 18228 94500
rect 18060 94386 18116 94388
rect 18060 94334 18062 94386
rect 18062 94334 18114 94386
rect 18114 94334 18116 94386
rect 18060 94332 18116 94334
rect 18620 94108 18676 94164
rect 19068 96738 19124 96740
rect 19068 96686 19070 96738
rect 19070 96686 19122 96738
rect 19122 96686 19124 96738
rect 19068 96684 19124 96686
rect 18844 95954 18900 95956
rect 18844 95902 18846 95954
rect 18846 95902 18898 95954
rect 18898 95902 18900 95954
rect 18844 95900 18900 95902
rect 18844 95452 18900 95508
rect 18060 93548 18116 93604
rect 18508 93436 18564 93492
rect 18060 93212 18116 93268
rect 18222 93322 18278 93324
rect 18222 93270 18224 93322
rect 18224 93270 18276 93322
rect 18276 93270 18278 93322
rect 18222 93268 18278 93270
rect 18326 93322 18382 93324
rect 18326 93270 18328 93322
rect 18328 93270 18380 93322
rect 18380 93270 18382 93322
rect 18326 93268 18382 93270
rect 18430 93322 18486 93324
rect 18430 93270 18432 93322
rect 18432 93270 18484 93322
rect 18484 93270 18486 93322
rect 18430 93268 18486 93270
rect 17836 92316 17892 92372
rect 17948 92764 18004 92820
rect 17500 92146 17556 92148
rect 17500 92094 17502 92146
rect 17502 92094 17554 92146
rect 17554 92094 17556 92146
rect 17500 92092 17556 92094
rect 17836 91532 17892 91588
rect 18620 92764 18676 92820
rect 19068 95116 19124 95172
rect 18508 92370 18564 92372
rect 18508 92318 18510 92370
rect 18510 92318 18562 92370
rect 18562 92318 18564 92370
rect 18508 92316 18564 92318
rect 18222 91754 18278 91756
rect 18222 91702 18224 91754
rect 18224 91702 18276 91754
rect 18276 91702 18278 91754
rect 18222 91700 18278 91702
rect 18326 91754 18382 91756
rect 18326 91702 18328 91754
rect 18328 91702 18380 91754
rect 18380 91702 18382 91754
rect 18326 91700 18382 91702
rect 18430 91754 18486 91756
rect 18430 91702 18432 91754
rect 18432 91702 18484 91754
rect 18484 91702 18486 91754
rect 18430 91700 18486 91702
rect 19404 97692 19460 97748
rect 19068 94498 19124 94500
rect 19068 94446 19070 94498
rect 19070 94446 19122 94498
rect 19122 94446 19124 94498
rect 19068 94444 19124 94446
rect 19180 94386 19236 94388
rect 19180 94334 19182 94386
rect 19182 94334 19234 94386
rect 19234 94334 19236 94386
rect 19180 94332 19236 94334
rect 19068 93548 19124 93604
rect 18956 92876 19012 92932
rect 18844 91980 18900 92036
rect 18956 91756 19012 91812
rect 18956 91196 19012 91252
rect 18172 90524 18228 90580
rect 17388 89964 17444 90020
rect 17948 90466 18004 90468
rect 17948 90414 17950 90466
rect 17950 90414 18002 90466
rect 18002 90414 18004 90466
rect 17948 90412 18004 90414
rect 18844 90524 18900 90580
rect 17724 89794 17780 89796
rect 17724 89742 17726 89794
rect 17726 89742 17778 89794
rect 17778 89742 17780 89794
rect 17724 89740 17780 89742
rect 17612 89628 17668 89684
rect 18222 90186 18278 90188
rect 18222 90134 18224 90186
rect 18224 90134 18276 90186
rect 18276 90134 18278 90186
rect 18222 90132 18278 90134
rect 18326 90186 18382 90188
rect 18326 90134 18328 90186
rect 18328 90134 18380 90186
rect 18380 90134 18382 90186
rect 18326 90132 18382 90134
rect 18430 90186 18486 90188
rect 18430 90134 18432 90186
rect 18432 90134 18484 90186
rect 18484 90134 18486 90186
rect 18430 90132 18486 90134
rect 18508 89964 18564 90020
rect 17948 89628 18004 89684
rect 18060 89570 18116 89572
rect 18060 89518 18062 89570
rect 18062 89518 18114 89570
rect 18114 89518 18116 89570
rect 18060 89516 18116 89518
rect 17500 89292 17556 89348
rect 18396 89628 18452 89684
rect 18284 89180 18340 89236
rect 17948 89068 18004 89124
rect 16604 88172 16660 88228
rect 16716 88060 16772 88116
rect 16604 87666 16660 87668
rect 16604 87614 16606 87666
rect 16606 87614 16658 87666
rect 16658 87614 16660 87666
rect 16604 87612 16660 87614
rect 15036 85820 15092 85876
rect 14820 84698 14876 84700
rect 14820 84646 14822 84698
rect 14822 84646 14874 84698
rect 14874 84646 14876 84698
rect 14820 84644 14876 84646
rect 14924 84698 14980 84700
rect 14924 84646 14926 84698
rect 14926 84646 14978 84698
rect 14978 84646 14980 84698
rect 14924 84644 14980 84646
rect 15028 84698 15084 84700
rect 15028 84646 15030 84698
rect 15030 84646 15082 84698
rect 15082 84646 15084 84698
rect 15028 84644 15084 84646
rect 14812 84364 14868 84420
rect 14924 83522 14980 83524
rect 14924 83470 14926 83522
rect 14926 83470 14978 83522
rect 14978 83470 14980 83522
rect 14924 83468 14980 83470
rect 14820 83130 14876 83132
rect 14820 83078 14822 83130
rect 14822 83078 14874 83130
rect 14874 83078 14876 83130
rect 14820 83076 14876 83078
rect 14924 83130 14980 83132
rect 14924 83078 14926 83130
rect 14926 83078 14978 83130
rect 14978 83078 14980 83130
rect 14924 83076 14980 83078
rect 15028 83130 15084 83132
rect 15028 83078 15030 83130
rect 15030 83078 15082 83130
rect 15082 83078 15084 83130
rect 15028 83076 15084 83078
rect 14812 81676 14868 81732
rect 14820 81562 14876 81564
rect 14820 81510 14822 81562
rect 14822 81510 14874 81562
rect 14874 81510 14876 81562
rect 14820 81508 14876 81510
rect 14924 81562 14980 81564
rect 14924 81510 14926 81562
rect 14926 81510 14978 81562
rect 14978 81510 14980 81562
rect 14924 81508 14980 81510
rect 15028 81562 15084 81564
rect 15028 81510 15030 81562
rect 15030 81510 15082 81562
rect 15082 81510 15084 81562
rect 15028 81508 15084 81510
rect 14820 79994 14876 79996
rect 14820 79942 14822 79994
rect 14822 79942 14874 79994
rect 14874 79942 14876 79994
rect 14820 79940 14876 79942
rect 14924 79994 14980 79996
rect 14924 79942 14926 79994
rect 14926 79942 14978 79994
rect 14978 79942 14980 79994
rect 14924 79940 14980 79942
rect 15028 79994 15084 79996
rect 15028 79942 15030 79994
rect 15030 79942 15082 79994
rect 15082 79942 15084 79994
rect 15028 79940 15084 79942
rect 15260 83692 15316 83748
rect 15484 86268 15540 86324
rect 15932 85986 15988 85988
rect 15932 85934 15934 85986
rect 15934 85934 15986 85986
rect 15986 85934 15988 85986
rect 15932 85932 15988 85934
rect 15484 85260 15540 85316
rect 16156 84924 16212 84980
rect 15484 84364 15540 84420
rect 16492 86828 16548 86884
rect 16828 85708 16884 85764
rect 16716 85650 16772 85652
rect 16716 85598 16718 85650
rect 16718 85598 16770 85650
rect 16770 85598 16772 85650
rect 16716 85596 16772 85598
rect 16380 85260 16436 85316
rect 16604 85036 16660 85092
rect 16268 84252 16324 84308
rect 15932 83692 15988 83748
rect 15596 83634 15652 83636
rect 15596 83582 15598 83634
rect 15598 83582 15650 83634
rect 15650 83582 15652 83634
rect 15596 83580 15652 83582
rect 15372 82908 15428 82964
rect 15708 83468 15764 83524
rect 15932 82908 15988 82964
rect 15596 82738 15652 82740
rect 15596 82686 15598 82738
rect 15598 82686 15650 82738
rect 15650 82686 15652 82738
rect 15596 82684 15652 82686
rect 15820 82348 15876 82404
rect 14812 79714 14868 79716
rect 14812 79662 14814 79714
rect 14814 79662 14866 79714
rect 14866 79662 14868 79714
rect 14812 79660 14868 79662
rect 14924 79602 14980 79604
rect 14924 79550 14926 79602
rect 14926 79550 14978 79602
rect 14978 79550 14980 79602
rect 14924 79548 14980 79550
rect 14700 79100 14756 79156
rect 14252 78428 14308 78484
rect 14820 78426 14876 78428
rect 14820 78374 14822 78426
rect 14822 78374 14874 78426
rect 14874 78374 14876 78426
rect 14820 78372 14876 78374
rect 14924 78426 14980 78428
rect 14924 78374 14926 78426
rect 14926 78374 14978 78426
rect 14978 78374 14980 78426
rect 14924 78372 14980 78374
rect 15028 78426 15084 78428
rect 15028 78374 15030 78426
rect 15030 78374 15082 78426
rect 15082 78374 15084 78426
rect 15028 78372 15084 78374
rect 14700 78204 14756 78260
rect 14364 78092 14420 78148
rect 15036 77250 15092 77252
rect 15036 77198 15038 77250
rect 15038 77198 15090 77250
rect 15090 77198 15092 77250
rect 15036 77196 15092 77198
rect 14820 76858 14876 76860
rect 14820 76806 14822 76858
rect 14822 76806 14874 76858
rect 14874 76806 14876 76858
rect 14820 76804 14876 76806
rect 14924 76858 14980 76860
rect 14924 76806 14926 76858
rect 14926 76806 14978 76858
rect 14978 76806 14980 76858
rect 14924 76804 14980 76806
rect 15028 76858 15084 76860
rect 15028 76806 15030 76858
rect 15030 76806 15082 76858
rect 15082 76806 15084 76858
rect 15028 76804 15084 76806
rect 14028 76466 14084 76468
rect 14028 76414 14030 76466
rect 14030 76414 14082 76466
rect 14082 76414 14084 76466
rect 14028 76412 14084 76414
rect 16604 83580 16660 83636
rect 16828 83244 16884 83300
rect 16044 82684 16100 82740
rect 16716 82738 16772 82740
rect 16716 82686 16718 82738
rect 16718 82686 16770 82738
rect 16770 82686 16772 82738
rect 16716 82684 16772 82686
rect 16380 82012 16436 82068
rect 15596 78204 15652 78260
rect 15260 75964 15316 76020
rect 14820 75290 14876 75292
rect 14820 75238 14822 75290
rect 14822 75238 14874 75290
rect 14874 75238 14876 75290
rect 14820 75236 14876 75238
rect 14924 75290 14980 75292
rect 14924 75238 14926 75290
rect 14926 75238 14978 75290
rect 14978 75238 14980 75290
rect 14924 75236 14980 75238
rect 15028 75290 15084 75292
rect 15028 75238 15030 75290
rect 15030 75238 15082 75290
rect 15082 75238 15084 75290
rect 15028 75236 15084 75238
rect 15596 75292 15652 75348
rect 15148 75122 15204 75124
rect 15148 75070 15150 75122
rect 15150 75070 15202 75122
rect 15202 75070 15204 75122
rect 15148 75068 15204 75070
rect 12572 74060 12628 74116
rect 12236 72828 12292 72884
rect 12236 72156 12292 72212
rect 11900 70082 11956 70084
rect 11900 70030 11902 70082
rect 11902 70030 11954 70082
rect 11954 70030 11956 70082
rect 11900 70028 11956 70030
rect 11788 69186 11844 69188
rect 11788 69134 11790 69186
rect 11790 69134 11842 69186
rect 11842 69134 11844 69186
rect 11788 69132 11844 69134
rect 12012 68684 12068 68740
rect 11418 68234 11474 68236
rect 11418 68182 11420 68234
rect 11420 68182 11472 68234
rect 11472 68182 11474 68234
rect 11418 68180 11474 68182
rect 11522 68234 11578 68236
rect 11522 68182 11524 68234
rect 11524 68182 11576 68234
rect 11576 68182 11578 68234
rect 11522 68180 11578 68182
rect 11626 68234 11682 68236
rect 11626 68182 11628 68234
rect 11628 68182 11680 68234
rect 11680 68182 11682 68234
rect 11626 68180 11682 68182
rect 11676 67842 11732 67844
rect 11676 67790 11678 67842
rect 11678 67790 11730 67842
rect 11730 67790 11732 67842
rect 11676 67788 11732 67790
rect 11452 67618 11508 67620
rect 11452 67566 11454 67618
rect 11454 67566 11506 67618
rect 11506 67566 11508 67618
rect 11452 67564 11508 67566
rect 10780 67004 10836 67060
rect 10332 64540 10388 64596
rect 9884 64482 9940 64484
rect 9884 64430 9886 64482
rect 9886 64430 9938 64482
rect 9938 64430 9940 64482
rect 9884 64428 9940 64430
rect 9660 63868 9716 63924
rect 10108 63922 10164 63924
rect 10108 63870 10110 63922
rect 10110 63870 10162 63922
rect 10162 63870 10164 63922
rect 10108 63868 10164 63870
rect 9996 63756 10052 63812
rect 9660 63698 9716 63700
rect 9660 63646 9662 63698
rect 9662 63646 9714 63698
rect 9714 63646 9716 63698
rect 9660 63644 9716 63646
rect 9660 63250 9716 63252
rect 9660 63198 9662 63250
rect 9662 63198 9714 63250
rect 9714 63198 9716 63250
rect 9660 63196 9716 63198
rect 10220 63196 10276 63252
rect 10108 62636 10164 62692
rect 9996 62524 10052 62580
rect 10444 64428 10500 64484
rect 9996 61516 10052 61572
rect 9660 60956 9716 61012
rect 9772 60674 9828 60676
rect 9772 60622 9774 60674
rect 9774 60622 9826 60674
rect 9826 60622 9828 60674
rect 9772 60620 9828 60622
rect 9884 59442 9940 59444
rect 9884 59390 9886 59442
rect 9886 59390 9938 59442
rect 9938 59390 9940 59442
rect 9884 59388 9940 59390
rect 9660 59164 9716 59220
rect 9548 58268 9604 58324
rect 10332 61010 10388 61012
rect 10332 60958 10334 61010
rect 10334 60958 10386 61010
rect 10386 60958 10388 61010
rect 10332 60956 10388 60958
rect 10332 60786 10388 60788
rect 10332 60734 10334 60786
rect 10334 60734 10386 60786
rect 10386 60734 10388 60786
rect 10332 60732 10388 60734
rect 10108 60620 10164 60676
rect 9660 58044 9716 58100
rect 11564 67058 11620 67060
rect 11564 67006 11566 67058
rect 11566 67006 11618 67058
rect 11618 67006 11620 67058
rect 11564 67004 11620 67006
rect 11004 66946 11060 66948
rect 11004 66894 11006 66946
rect 11006 66894 11058 66946
rect 11058 66894 11060 66946
rect 11004 66892 11060 66894
rect 11418 66666 11474 66668
rect 11418 66614 11420 66666
rect 11420 66614 11472 66666
rect 11472 66614 11474 66666
rect 11418 66612 11474 66614
rect 11522 66666 11578 66668
rect 11522 66614 11524 66666
rect 11524 66614 11576 66666
rect 11576 66614 11578 66666
rect 11522 66612 11578 66614
rect 11626 66666 11682 66668
rect 11626 66614 11628 66666
rect 11628 66614 11680 66666
rect 11680 66614 11682 66666
rect 11626 66612 11682 66614
rect 11418 65098 11474 65100
rect 11418 65046 11420 65098
rect 11420 65046 11472 65098
rect 11472 65046 11474 65098
rect 11418 65044 11474 65046
rect 11522 65098 11578 65100
rect 11522 65046 11524 65098
rect 11524 65046 11576 65098
rect 11576 65046 11578 65098
rect 11522 65044 11578 65046
rect 11626 65098 11682 65100
rect 11626 65046 11628 65098
rect 11628 65046 11680 65098
rect 11680 65046 11682 65098
rect 11626 65044 11682 65046
rect 11228 64594 11284 64596
rect 11228 64542 11230 64594
rect 11230 64542 11282 64594
rect 11282 64542 11284 64594
rect 11228 64540 11284 64542
rect 10556 61628 10612 61684
rect 11418 63530 11474 63532
rect 11418 63478 11420 63530
rect 11420 63478 11472 63530
rect 11472 63478 11474 63530
rect 11418 63476 11474 63478
rect 11522 63530 11578 63532
rect 11522 63478 11524 63530
rect 11524 63478 11576 63530
rect 11576 63478 11578 63530
rect 11522 63476 11578 63478
rect 11626 63530 11682 63532
rect 11626 63478 11628 63530
rect 11628 63478 11680 63530
rect 11680 63478 11682 63530
rect 11626 63476 11682 63478
rect 12012 66892 12068 66948
rect 12012 63868 12068 63924
rect 11564 63196 11620 63252
rect 11228 62748 11284 62804
rect 11788 63138 11844 63140
rect 11788 63086 11790 63138
rect 11790 63086 11842 63138
rect 11842 63086 11844 63138
rect 11788 63084 11844 63086
rect 11004 62578 11060 62580
rect 11004 62526 11006 62578
rect 11006 62526 11058 62578
rect 11058 62526 11060 62578
rect 11004 62524 11060 62526
rect 11418 61962 11474 61964
rect 11418 61910 11420 61962
rect 11420 61910 11472 61962
rect 11472 61910 11474 61962
rect 11418 61908 11474 61910
rect 11522 61962 11578 61964
rect 11522 61910 11524 61962
rect 11524 61910 11576 61962
rect 11576 61910 11578 61962
rect 11522 61908 11578 61910
rect 11626 61962 11682 61964
rect 11626 61910 11628 61962
rect 11628 61910 11680 61962
rect 11680 61910 11682 61962
rect 11626 61908 11682 61910
rect 11788 61292 11844 61348
rect 10444 60508 10500 60564
rect 10780 60508 10836 60564
rect 10444 59778 10500 59780
rect 10444 59726 10446 59778
rect 10446 59726 10498 59778
rect 10498 59726 10500 59778
rect 10444 59724 10500 59726
rect 10444 59276 10500 59332
rect 9660 56588 9716 56644
rect 9772 56476 9828 56532
rect 9548 56140 9604 56196
rect 9436 55410 9492 55412
rect 9436 55358 9438 55410
rect 9438 55358 9490 55410
rect 9490 55358 9492 55410
rect 9436 55356 9492 55358
rect 10108 57820 10164 57876
rect 10444 58828 10500 58884
rect 10556 58546 10612 58548
rect 10556 58494 10558 58546
rect 10558 58494 10610 58546
rect 10610 58494 10612 58546
rect 10556 58492 10612 58494
rect 11452 60898 11508 60900
rect 11452 60846 11454 60898
rect 11454 60846 11506 60898
rect 11506 60846 11508 60898
rect 11452 60844 11508 60846
rect 11228 60396 11284 60452
rect 11418 60394 11474 60396
rect 11418 60342 11420 60394
rect 11420 60342 11472 60394
rect 11472 60342 11474 60394
rect 11418 60340 11474 60342
rect 11522 60394 11578 60396
rect 11522 60342 11524 60394
rect 11524 60342 11576 60394
rect 11576 60342 11578 60394
rect 11522 60340 11578 60342
rect 11626 60394 11682 60396
rect 11626 60342 11628 60394
rect 11628 60342 11680 60394
rect 11680 60342 11682 60394
rect 11626 60340 11682 60342
rect 12460 70754 12516 70756
rect 12460 70702 12462 70754
rect 12462 70702 12514 70754
rect 12514 70702 12516 70754
rect 12460 70700 12516 70702
rect 13132 73836 13188 73892
rect 12684 72828 12740 72884
rect 12908 72658 12964 72660
rect 12908 72606 12910 72658
rect 12910 72606 12962 72658
rect 12962 72606 12964 72658
rect 12908 72604 12964 72606
rect 12684 70082 12740 70084
rect 12684 70030 12686 70082
rect 12686 70030 12738 70082
rect 12738 70030 12740 70082
rect 12684 70028 12740 70030
rect 12796 72268 12852 72324
rect 12908 71986 12964 71988
rect 12908 71934 12910 71986
rect 12910 71934 12962 71986
rect 12962 71934 12964 71986
rect 12908 71932 12964 71934
rect 13020 71148 13076 71204
rect 12908 70588 12964 70644
rect 14028 74898 14084 74900
rect 14028 74846 14030 74898
rect 14030 74846 14082 74898
rect 14082 74846 14084 74898
rect 14028 74844 14084 74846
rect 13804 74172 13860 74228
rect 14028 74620 14084 74676
rect 14588 74898 14644 74900
rect 14588 74846 14590 74898
rect 14590 74846 14642 74898
rect 14642 74846 14644 74898
rect 14588 74844 14644 74846
rect 15036 74898 15092 74900
rect 15036 74846 15038 74898
rect 15038 74846 15090 74898
rect 15090 74846 15092 74898
rect 15036 74844 15092 74846
rect 14924 74732 14980 74788
rect 14252 74508 14308 74564
rect 13692 73948 13748 74004
rect 14028 73442 14084 73444
rect 14028 73390 14030 73442
rect 14030 73390 14082 73442
rect 14082 73390 14084 73442
rect 14028 73388 14084 73390
rect 13804 73330 13860 73332
rect 13804 73278 13806 73330
rect 13806 73278 13858 73330
rect 13858 73278 13860 73330
rect 13804 73276 13860 73278
rect 14252 73276 14308 73332
rect 13692 73164 13748 73220
rect 14028 72716 14084 72772
rect 13580 72546 13636 72548
rect 13580 72494 13582 72546
rect 13582 72494 13634 72546
rect 13634 72494 13636 72546
rect 13580 72492 13636 72494
rect 14140 72268 14196 72324
rect 15708 74060 15764 74116
rect 14588 73890 14644 73892
rect 14588 73838 14590 73890
rect 14590 73838 14642 73890
rect 14642 73838 14644 73890
rect 14588 73836 14644 73838
rect 15372 73836 15428 73892
rect 14820 73722 14876 73724
rect 14820 73670 14822 73722
rect 14822 73670 14874 73722
rect 14874 73670 14876 73722
rect 14820 73668 14876 73670
rect 14924 73722 14980 73724
rect 14924 73670 14926 73722
rect 14926 73670 14978 73722
rect 14978 73670 14980 73722
rect 14924 73668 14980 73670
rect 15028 73722 15084 73724
rect 15028 73670 15030 73722
rect 15030 73670 15082 73722
rect 15082 73670 15084 73722
rect 15028 73668 15084 73670
rect 14700 73388 14756 73444
rect 15260 73388 15316 73444
rect 14588 72492 14644 72548
rect 15148 73218 15204 73220
rect 15148 73166 15150 73218
rect 15150 73166 15202 73218
rect 15202 73166 15204 73218
rect 15148 73164 15204 73166
rect 15148 72380 15204 72436
rect 14252 72044 14308 72100
rect 13468 71538 13524 71540
rect 13468 71486 13470 71538
rect 13470 71486 13522 71538
rect 13522 71486 13524 71538
rect 13468 71484 13524 71486
rect 13916 71538 13972 71540
rect 13916 71486 13918 71538
rect 13918 71486 13970 71538
rect 13970 71486 13972 71538
rect 13916 71484 13972 71486
rect 14364 71986 14420 71988
rect 14364 71934 14366 71986
rect 14366 71934 14418 71986
rect 14418 71934 14420 71986
rect 14364 71932 14420 71934
rect 14820 72154 14876 72156
rect 14820 72102 14822 72154
rect 14822 72102 14874 72154
rect 14874 72102 14876 72154
rect 14820 72100 14876 72102
rect 14924 72154 14980 72156
rect 14924 72102 14926 72154
rect 14926 72102 14978 72154
rect 14978 72102 14980 72154
rect 14924 72100 14980 72102
rect 15028 72154 15084 72156
rect 15028 72102 15030 72154
rect 15030 72102 15082 72154
rect 15082 72102 15084 72154
rect 15028 72100 15084 72102
rect 14252 71484 14308 71540
rect 13468 71148 13524 71204
rect 13244 71036 13300 71092
rect 12908 70194 12964 70196
rect 12908 70142 12910 70194
rect 12910 70142 12962 70194
rect 12962 70142 12964 70194
rect 12908 70140 12964 70142
rect 12236 68684 12292 68740
rect 12684 69634 12740 69636
rect 12684 69582 12686 69634
rect 12686 69582 12738 69634
rect 12738 69582 12740 69634
rect 12684 69580 12740 69582
rect 12460 67788 12516 67844
rect 12908 67954 12964 67956
rect 12908 67902 12910 67954
rect 12910 67902 12962 67954
rect 12962 67902 12964 67954
rect 12908 67900 12964 67902
rect 12460 67618 12516 67620
rect 12460 67566 12462 67618
rect 12462 67566 12514 67618
rect 12514 67566 12516 67618
rect 12460 67564 12516 67566
rect 12460 67340 12516 67396
rect 12460 65660 12516 65716
rect 12572 67058 12628 67060
rect 12572 67006 12574 67058
rect 12574 67006 12626 67058
rect 12626 67006 12628 67058
rect 12572 67004 12628 67006
rect 13132 69804 13188 69860
rect 13580 70588 13636 70644
rect 13692 70924 13748 70980
rect 13356 70140 13412 70196
rect 13468 70028 13524 70084
rect 13468 69468 13524 69524
rect 13244 69356 13300 69412
rect 13916 70924 13972 70980
rect 13804 70812 13860 70868
rect 14140 70812 14196 70868
rect 14028 70700 14084 70756
rect 14028 70140 14084 70196
rect 14140 70588 14196 70644
rect 14028 69410 14084 69412
rect 14028 69358 14030 69410
rect 14030 69358 14082 69410
rect 14082 69358 14084 69410
rect 14028 69356 14084 69358
rect 12796 66834 12852 66836
rect 12796 66782 12798 66834
rect 12798 66782 12850 66834
rect 12850 66782 12852 66834
rect 12796 66780 12852 66782
rect 13468 68348 13524 68404
rect 13468 67954 13524 67956
rect 13468 67902 13470 67954
rect 13470 67902 13522 67954
rect 13522 67902 13524 67954
rect 13468 67900 13524 67902
rect 13916 69186 13972 69188
rect 13916 69134 13918 69186
rect 13918 69134 13970 69186
rect 13970 69134 13972 69186
rect 13916 69132 13972 69134
rect 13692 68236 13748 68292
rect 12908 66386 12964 66388
rect 12908 66334 12910 66386
rect 12910 66334 12962 66386
rect 12962 66334 12964 66386
rect 12908 66332 12964 66334
rect 12684 65436 12740 65492
rect 12236 63084 12292 63140
rect 12460 63138 12516 63140
rect 12460 63086 12462 63138
rect 12462 63086 12514 63138
rect 12514 63086 12516 63138
rect 12460 63084 12516 63086
rect 12236 62524 12292 62580
rect 12460 62748 12516 62804
rect 12684 63868 12740 63924
rect 12684 62914 12740 62916
rect 12684 62862 12686 62914
rect 12686 62862 12738 62914
rect 12738 62862 12740 62914
rect 12684 62860 12740 62862
rect 12124 61740 12180 61796
rect 12684 62300 12740 62356
rect 12124 61458 12180 61460
rect 12124 61406 12126 61458
rect 12126 61406 12178 61458
rect 12178 61406 12180 61458
rect 12124 61404 12180 61406
rect 12348 61740 12404 61796
rect 13132 65378 13188 65380
rect 13132 65326 13134 65378
rect 13134 65326 13186 65378
rect 13186 65326 13188 65378
rect 13132 65324 13188 65326
rect 13132 64204 13188 64260
rect 13020 63084 13076 63140
rect 13020 62578 13076 62580
rect 13020 62526 13022 62578
rect 13022 62526 13074 62578
rect 13074 62526 13076 62578
rect 13020 62524 13076 62526
rect 12348 61292 12404 61348
rect 12684 61346 12740 61348
rect 12684 61294 12686 61346
rect 12686 61294 12738 61346
rect 12738 61294 12740 61346
rect 12684 61292 12740 61294
rect 11900 60002 11956 60004
rect 11900 59950 11902 60002
rect 11902 59950 11954 60002
rect 11954 59950 11956 60002
rect 11900 59948 11956 59950
rect 11900 58940 11956 58996
rect 11418 58826 11474 58828
rect 11418 58774 11420 58826
rect 11420 58774 11472 58826
rect 11472 58774 11474 58826
rect 11418 58772 11474 58774
rect 11522 58826 11578 58828
rect 11522 58774 11524 58826
rect 11524 58774 11576 58826
rect 11576 58774 11578 58826
rect 11522 58772 11578 58774
rect 11626 58826 11682 58828
rect 11626 58774 11628 58826
rect 11628 58774 11680 58826
rect 11680 58774 11682 58826
rect 11626 58772 11682 58774
rect 11788 58658 11844 58660
rect 11788 58606 11790 58658
rect 11790 58606 11842 58658
rect 11842 58606 11844 58658
rect 11788 58604 11844 58606
rect 10892 58380 10948 58436
rect 10556 58268 10612 58324
rect 11340 58322 11396 58324
rect 11340 58270 11342 58322
rect 11342 58270 11394 58322
rect 11394 58270 11396 58322
rect 11340 58268 11396 58270
rect 11004 58210 11060 58212
rect 11004 58158 11006 58210
rect 11006 58158 11058 58210
rect 11058 58158 11060 58210
rect 11004 58156 11060 58158
rect 10332 57484 10388 57540
rect 10108 56476 10164 56532
rect 10220 56588 10276 56644
rect 10332 56140 10388 56196
rect 10668 57650 10724 57652
rect 10668 57598 10670 57650
rect 10670 57598 10722 57650
rect 10722 57598 10724 57650
rect 10668 57596 10724 57598
rect 9772 55916 9828 55972
rect 9660 55132 9716 55188
rect 10332 55970 10388 55972
rect 10332 55918 10334 55970
rect 10334 55918 10386 55970
rect 10386 55918 10388 55970
rect 10332 55916 10388 55918
rect 10108 55804 10164 55860
rect 9996 54908 10052 54964
rect 10444 55804 10500 55860
rect 9660 53788 9716 53844
rect 10780 56978 10836 56980
rect 10780 56926 10782 56978
rect 10782 56926 10834 56978
rect 10834 56926 10836 56978
rect 10780 56924 10836 56926
rect 11340 57596 11396 57652
rect 11116 57538 11172 57540
rect 11116 57486 11118 57538
rect 11118 57486 11170 57538
rect 11170 57486 11172 57538
rect 11116 57484 11172 57486
rect 10892 56252 10948 56308
rect 10892 55858 10948 55860
rect 10892 55806 10894 55858
rect 10894 55806 10946 55858
rect 10946 55806 10948 55858
rect 10892 55804 10948 55806
rect 10668 55074 10724 55076
rect 10668 55022 10670 55074
rect 10670 55022 10722 55074
rect 10722 55022 10724 55074
rect 10668 55020 10724 55022
rect 10556 54796 10612 54852
rect 9548 53116 9604 53172
rect 9996 53564 10052 53620
rect 10220 53842 10276 53844
rect 10220 53790 10222 53842
rect 10222 53790 10274 53842
rect 10274 53790 10276 53842
rect 10220 53788 10276 53790
rect 9884 52220 9940 52276
rect 10220 53004 10276 53060
rect 10556 54124 10612 54180
rect 10108 52332 10164 52388
rect 9436 51772 9492 51828
rect 9548 51660 9604 51716
rect 10444 53676 10500 53732
rect 10780 53452 10836 53508
rect 10556 52892 10612 52948
rect 10332 52274 10388 52276
rect 10332 52222 10334 52274
rect 10334 52222 10386 52274
rect 10386 52222 10388 52274
rect 10332 52220 10388 52222
rect 9996 51324 10052 51380
rect 10332 50204 10388 50260
rect 10108 49810 10164 49812
rect 10108 49758 10110 49810
rect 10110 49758 10162 49810
rect 10162 49758 10164 49810
rect 10108 49756 10164 49758
rect 9772 49532 9828 49588
rect 9436 48412 9492 48468
rect 9660 48130 9716 48132
rect 9660 48078 9662 48130
rect 9662 48078 9714 48130
rect 9714 48078 9716 48130
rect 9660 48076 9716 48078
rect 9548 47852 9604 47908
rect 9548 47404 9604 47460
rect 9996 48636 10052 48692
rect 9996 48466 10052 48468
rect 9996 48414 9998 48466
rect 9998 48414 10050 48466
rect 10050 48414 10052 48466
rect 9996 48412 10052 48414
rect 9996 47964 10052 48020
rect 10668 52668 10724 52724
rect 10892 52668 10948 52724
rect 11418 57258 11474 57260
rect 11418 57206 11420 57258
rect 11420 57206 11472 57258
rect 11472 57206 11474 57258
rect 11418 57204 11474 57206
rect 11522 57258 11578 57260
rect 11522 57206 11524 57258
rect 11524 57206 11576 57258
rect 11576 57206 11578 57258
rect 11522 57204 11578 57206
rect 11626 57258 11682 57260
rect 11626 57206 11628 57258
rect 11628 57206 11680 57258
rect 11680 57206 11682 57258
rect 11626 57204 11682 57206
rect 12012 58044 12068 58100
rect 11900 57484 11956 57540
rect 12012 56924 12068 56980
rect 11900 56588 11956 56644
rect 11228 56194 11284 56196
rect 11228 56142 11230 56194
rect 11230 56142 11282 56194
rect 11282 56142 11284 56194
rect 11228 56140 11284 56142
rect 11452 56140 11508 56196
rect 11452 55804 11508 55860
rect 12348 60732 12404 60788
rect 12236 57932 12292 57988
rect 12236 57148 12292 57204
rect 12236 56476 12292 56532
rect 11418 55690 11474 55692
rect 11418 55638 11420 55690
rect 11420 55638 11472 55690
rect 11472 55638 11474 55690
rect 11418 55636 11474 55638
rect 11522 55690 11578 55692
rect 11522 55638 11524 55690
rect 11524 55638 11576 55690
rect 11576 55638 11578 55690
rect 11522 55636 11578 55638
rect 11626 55690 11682 55692
rect 11626 55638 11628 55690
rect 11628 55638 11680 55690
rect 11680 55638 11682 55690
rect 11626 55636 11682 55638
rect 11340 55468 11396 55524
rect 11564 55186 11620 55188
rect 11564 55134 11566 55186
rect 11566 55134 11618 55186
rect 11618 55134 11620 55186
rect 11564 55132 11620 55134
rect 12012 55186 12068 55188
rect 12012 55134 12014 55186
rect 12014 55134 12066 55186
rect 12066 55134 12068 55186
rect 12012 55132 12068 55134
rect 12012 54908 12068 54964
rect 11418 54122 11474 54124
rect 11418 54070 11420 54122
rect 11420 54070 11472 54122
rect 11472 54070 11474 54122
rect 11418 54068 11474 54070
rect 11522 54122 11578 54124
rect 11522 54070 11524 54122
rect 11524 54070 11576 54122
rect 11576 54070 11578 54122
rect 11522 54068 11578 54070
rect 11626 54122 11682 54124
rect 11626 54070 11628 54122
rect 11628 54070 11680 54122
rect 11680 54070 11682 54122
rect 11626 54068 11682 54070
rect 11900 54012 11956 54068
rect 11116 53788 11172 53844
rect 11788 53842 11844 53844
rect 11788 53790 11790 53842
rect 11790 53790 11842 53842
rect 11842 53790 11844 53842
rect 11788 53788 11844 53790
rect 11228 53676 11284 53732
rect 11116 53004 11172 53060
rect 12908 60620 12964 60676
rect 12572 58604 12628 58660
rect 12572 58322 12628 58324
rect 12572 58270 12574 58322
rect 12574 58270 12626 58322
rect 12626 58270 12628 58322
rect 12572 58268 12628 58270
rect 12908 60284 12964 60340
rect 12908 58940 12964 58996
rect 13020 58492 13076 58548
rect 13132 61292 13188 61348
rect 12460 57932 12516 57988
rect 13132 57708 13188 57764
rect 12460 56924 12516 56980
rect 12684 57148 12740 57204
rect 12572 56082 12628 56084
rect 12572 56030 12574 56082
rect 12574 56030 12626 56082
rect 12626 56030 12628 56082
rect 12572 56028 12628 56030
rect 11788 53452 11844 53508
rect 11788 53228 11844 53284
rect 11004 52386 11060 52388
rect 11004 52334 11006 52386
rect 11006 52334 11058 52386
rect 11058 52334 11060 52386
rect 11004 52332 11060 52334
rect 10556 52220 10612 52276
rect 10668 51436 10724 51492
rect 10556 50652 10612 50708
rect 10668 49980 10724 50036
rect 11228 52556 11284 52612
rect 11418 52554 11474 52556
rect 11418 52502 11420 52554
rect 11420 52502 11472 52554
rect 11472 52502 11474 52554
rect 11418 52500 11474 52502
rect 11522 52554 11578 52556
rect 11522 52502 11524 52554
rect 11524 52502 11576 52554
rect 11576 52502 11578 52554
rect 11522 52500 11578 52502
rect 11626 52554 11682 52556
rect 11626 52502 11628 52554
rect 11628 52502 11680 52554
rect 11680 52502 11682 52554
rect 11626 52500 11682 52502
rect 12012 53452 12068 53508
rect 12124 53340 12180 53396
rect 12124 53058 12180 53060
rect 12124 53006 12126 53058
rect 12126 53006 12178 53058
rect 12178 53006 12180 53058
rect 12124 53004 12180 53006
rect 11116 51548 11172 51604
rect 11676 51100 11732 51156
rect 11418 50986 11474 50988
rect 11418 50934 11420 50986
rect 11420 50934 11472 50986
rect 11472 50934 11474 50986
rect 11418 50932 11474 50934
rect 11522 50986 11578 50988
rect 11522 50934 11524 50986
rect 11524 50934 11576 50986
rect 11576 50934 11578 50986
rect 11522 50932 11578 50934
rect 11626 50986 11682 50988
rect 11626 50934 11628 50986
rect 11628 50934 11680 50986
rect 11680 50934 11682 50986
rect 11626 50932 11682 50934
rect 12124 52162 12180 52164
rect 12124 52110 12126 52162
rect 12126 52110 12178 52162
rect 12178 52110 12180 52162
rect 12124 52108 12180 52110
rect 12012 51100 12068 51156
rect 10556 48802 10612 48804
rect 10556 48750 10558 48802
rect 10558 48750 10610 48802
rect 10610 48750 10612 48802
rect 10556 48748 10612 48750
rect 10444 48412 10500 48468
rect 11004 49698 11060 49700
rect 11004 49646 11006 49698
rect 11006 49646 11058 49698
rect 11058 49646 11060 49698
rect 11004 49644 11060 49646
rect 10780 49532 10836 49588
rect 12572 55410 12628 55412
rect 12572 55358 12574 55410
rect 12574 55358 12626 55410
rect 12626 55358 12628 55410
rect 12572 55356 12628 55358
rect 12796 57036 12852 57092
rect 12908 56476 12964 56532
rect 14028 68626 14084 68628
rect 14028 68574 14030 68626
rect 14030 68574 14082 68626
rect 14082 68574 14084 68626
rect 14028 68572 14084 68574
rect 13916 67564 13972 67620
rect 14476 71148 14532 71204
rect 15036 71932 15092 71988
rect 14924 71484 14980 71540
rect 15260 72268 15316 72324
rect 15596 73500 15652 73556
rect 15372 72156 15428 72212
rect 14924 70924 14980 70980
rect 15484 73052 15540 73108
rect 15596 72828 15652 72884
rect 16604 81116 16660 81172
rect 16492 80946 16548 80948
rect 16492 80894 16494 80946
rect 16494 80894 16546 80946
rect 16546 80894 16548 80946
rect 16492 80892 16548 80894
rect 16940 82012 16996 82068
rect 17052 87836 17108 87892
rect 17276 87276 17332 87332
rect 18396 88844 18452 88900
rect 18620 89234 18676 89236
rect 18620 89182 18622 89234
rect 18622 89182 18674 89234
rect 18674 89182 18676 89234
rect 18620 89180 18676 89182
rect 19852 97468 19908 97524
rect 19516 97132 19572 97188
rect 19964 97804 20020 97860
rect 20076 97634 20132 97636
rect 20076 97582 20078 97634
rect 20078 97582 20130 97634
rect 20130 97582 20132 97634
rect 20076 97580 20132 97582
rect 20188 96962 20244 96964
rect 20188 96910 20190 96962
rect 20190 96910 20242 96962
rect 20242 96910 20244 96962
rect 20188 96908 20244 96910
rect 19852 96684 19908 96740
rect 19740 96236 19796 96292
rect 19628 95900 19684 95956
rect 19516 94668 19572 94724
rect 20188 96572 20244 96628
rect 19740 94668 19796 94724
rect 19852 95788 19908 95844
rect 19180 92876 19236 92932
rect 19404 92428 19460 92484
rect 19292 91980 19348 92036
rect 19180 91868 19236 91924
rect 19404 90802 19460 90804
rect 19404 90750 19406 90802
rect 19406 90750 19458 90802
rect 19458 90750 19460 90802
rect 19404 90748 19460 90750
rect 18956 88732 19012 88788
rect 18222 88618 18278 88620
rect 18222 88566 18224 88618
rect 18224 88566 18276 88618
rect 18276 88566 18278 88618
rect 18222 88564 18278 88566
rect 18326 88618 18382 88620
rect 18326 88566 18328 88618
rect 18328 88566 18380 88618
rect 18380 88566 18382 88618
rect 18326 88564 18382 88566
rect 18430 88618 18486 88620
rect 18430 88566 18432 88618
rect 18432 88566 18484 88618
rect 18484 88566 18486 88618
rect 18430 88564 18486 88566
rect 17276 85932 17332 85988
rect 17052 85596 17108 85652
rect 17724 88114 17780 88116
rect 17724 88062 17726 88114
rect 17726 88062 17778 88114
rect 17778 88062 17780 88114
rect 17724 88060 17780 88062
rect 18060 88114 18116 88116
rect 18060 88062 18062 88114
rect 18062 88062 18114 88114
rect 18114 88062 18116 88114
rect 18060 88060 18116 88062
rect 18508 88114 18564 88116
rect 18508 88062 18510 88114
rect 18510 88062 18562 88114
rect 18562 88062 18564 88114
rect 18508 88060 18564 88062
rect 17612 87948 17668 88004
rect 17500 87666 17556 87668
rect 17500 87614 17502 87666
rect 17502 87614 17554 87666
rect 17554 87614 17556 87666
rect 17500 87612 17556 87614
rect 18620 87836 18676 87892
rect 17836 87330 17892 87332
rect 17836 87278 17838 87330
rect 17838 87278 17890 87330
rect 17890 87278 17892 87330
rect 17836 87276 17892 87278
rect 17948 86828 18004 86884
rect 18222 87050 18278 87052
rect 18222 86998 18224 87050
rect 18224 86998 18276 87050
rect 18276 86998 18278 87050
rect 18222 86996 18278 86998
rect 18326 87050 18382 87052
rect 18326 86998 18328 87050
rect 18328 86998 18380 87050
rect 18380 86998 18382 87050
rect 18326 86996 18382 86998
rect 18430 87050 18486 87052
rect 18430 86998 18432 87050
rect 18432 86998 18484 87050
rect 18484 86998 18486 87050
rect 18430 86996 18486 86998
rect 18620 86604 18676 86660
rect 18844 87724 18900 87780
rect 18956 86882 19012 86884
rect 18956 86830 18958 86882
rect 18958 86830 19010 86882
rect 19010 86830 19012 86882
rect 18956 86828 19012 86830
rect 19292 88956 19348 89012
rect 19740 94332 19796 94388
rect 19628 92316 19684 92372
rect 19740 94108 19796 94164
rect 20076 95954 20132 95956
rect 20076 95902 20078 95954
rect 20078 95902 20130 95954
rect 20130 95902 20132 95954
rect 20076 95900 20132 95902
rect 20076 95676 20132 95732
rect 19852 92876 19908 92932
rect 19740 92428 19796 92484
rect 19628 91196 19684 91252
rect 19964 90802 20020 90804
rect 19964 90750 19966 90802
rect 19966 90750 20018 90802
rect 20018 90750 20020 90802
rect 19964 90748 20020 90750
rect 20300 93548 20356 93604
rect 20972 102284 21028 102340
rect 20636 99484 20692 99540
rect 20748 99036 20804 99092
rect 20524 96626 20580 96628
rect 20524 96574 20526 96626
rect 20526 96574 20578 96626
rect 20578 96574 20580 96626
rect 20524 96572 20580 96574
rect 20636 96124 20692 96180
rect 20636 95954 20692 95956
rect 20636 95902 20638 95954
rect 20638 95902 20690 95954
rect 20690 95902 20692 95954
rect 20636 95900 20692 95902
rect 20524 95506 20580 95508
rect 20524 95454 20526 95506
rect 20526 95454 20578 95506
rect 20578 95454 20580 95506
rect 20524 95452 20580 95454
rect 20860 97580 20916 97636
rect 20860 96012 20916 96068
rect 20748 93884 20804 93940
rect 22764 102450 22820 102452
rect 22764 102398 22766 102450
rect 22766 102398 22818 102450
rect 22818 102398 22820 102450
rect 22764 102396 22820 102398
rect 21868 102338 21924 102340
rect 21868 102286 21870 102338
rect 21870 102286 21922 102338
rect 21922 102286 21924 102338
rect 21868 102284 21924 102286
rect 21308 101500 21364 101556
rect 21084 99148 21140 99204
rect 21624 101946 21680 101948
rect 21624 101894 21626 101946
rect 21626 101894 21678 101946
rect 21678 101894 21680 101946
rect 21624 101892 21680 101894
rect 21728 101946 21784 101948
rect 21728 101894 21730 101946
rect 21730 101894 21782 101946
rect 21782 101894 21784 101946
rect 21728 101892 21784 101894
rect 21832 101946 21888 101948
rect 21832 101894 21834 101946
rect 21834 101894 21886 101946
rect 21886 101894 21888 101946
rect 21832 101892 21888 101894
rect 21868 100716 21924 100772
rect 21420 100604 21476 100660
rect 21624 100378 21680 100380
rect 21624 100326 21626 100378
rect 21626 100326 21678 100378
rect 21678 100326 21680 100378
rect 21624 100324 21680 100326
rect 21728 100378 21784 100380
rect 21728 100326 21730 100378
rect 21730 100326 21782 100378
rect 21782 100326 21784 100378
rect 21728 100324 21784 100326
rect 21832 100378 21888 100380
rect 21832 100326 21834 100378
rect 21834 100326 21886 100378
rect 21886 100326 21888 100378
rect 21832 100324 21888 100326
rect 22316 99932 22372 99988
rect 21196 98530 21252 98532
rect 21196 98478 21198 98530
rect 21198 98478 21250 98530
rect 21250 98478 21252 98530
rect 21196 98476 21252 98478
rect 21756 99202 21812 99204
rect 21756 99150 21758 99202
rect 21758 99150 21810 99202
rect 21810 99150 21812 99202
rect 21756 99148 21812 99150
rect 21980 99036 22036 99092
rect 21624 98810 21680 98812
rect 21624 98758 21626 98810
rect 21626 98758 21678 98810
rect 21678 98758 21680 98810
rect 21624 98756 21680 98758
rect 21728 98810 21784 98812
rect 21728 98758 21730 98810
rect 21730 98758 21782 98810
rect 21782 98758 21784 98810
rect 21728 98756 21784 98758
rect 21832 98810 21888 98812
rect 21832 98758 21834 98810
rect 21834 98758 21886 98810
rect 21886 98758 21888 98810
rect 21832 98756 21888 98758
rect 21868 98642 21924 98644
rect 21868 98590 21870 98642
rect 21870 98590 21922 98642
rect 21922 98590 21924 98642
rect 21868 98588 21924 98590
rect 21868 98194 21924 98196
rect 21868 98142 21870 98194
rect 21870 98142 21922 98194
rect 21922 98142 21924 98194
rect 21868 98140 21924 98142
rect 22764 98924 22820 98980
rect 21980 97804 22036 97860
rect 21420 97522 21476 97524
rect 21420 97470 21422 97522
rect 21422 97470 21474 97522
rect 21474 97470 21476 97522
rect 21420 97468 21476 97470
rect 21624 97242 21680 97244
rect 21624 97190 21626 97242
rect 21626 97190 21678 97242
rect 21678 97190 21680 97242
rect 21624 97188 21680 97190
rect 21728 97242 21784 97244
rect 21728 97190 21730 97242
rect 21730 97190 21782 97242
rect 21782 97190 21784 97242
rect 21728 97188 21784 97190
rect 21832 97242 21888 97244
rect 21832 97190 21834 97242
rect 21834 97190 21886 97242
rect 21886 97190 21888 97242
rect 21832 97188 21888 97190
rect 21308 96796 21364 96852
rect 22204 98476 22260 98532
rect 22540 97746 22596 97748
rect 22540 97694 22542 97746
rect 22542 97694 22594 97746
rect 22594 97694 22596 97746
rect 22540 97692 22596 97694
rect 22204 97580 22260 97636
rect 22092 96850 22148 96852
rect 22092 96798 22094 96850
rect 22094 96798 22146 96850
rect 22146 96798 22148 96850
rect 22092 96796 22148 96798
rect 22876 97522 22932 97524
rect 22876 97470 22878 97522
rect 22878 97470 22930 97522
rect 22930 97470 22932 97522
rect 22876 97468 22932 97470
rect 21084 95788 21140 95844
rect 22316 95900 22372 95956
rect 21644 95788 21700 95844
rect 21624 95674 21680 95676
rect 21624 95622 21626 95674
rect 21626 95622 21678 95674
rect 21678 95622 21680 95674
rect 21624 95620 21680 95622
rect 21728 95674 21784 95676
rect 21728 95622 21730 95674
rect 21730 95622 21782 95674
rect 21782 95622 21784 95674
rect 21728 95620 21784 95622
rect 21832 95674 21888 95676
rect 21832 95622 21834 95674
rect 21834 95622 21886 95674
rect 21886 95622 21888 95674
rect 21832 95620 21888 95622
rect 20972 94556 21028 94612
rect 20524 93714 20580 93716
rect 20524 93662 20526 93714
rect 20526 93662 20578 93714
rect 20578 93662 20580 93714
rect 20524 93660 20580 93662
rect 20188 92706 20244 92708
rect 20188 92654 20190 92706
rect 20190 92654 20242 92706
rect 20242 92654 20244 92706
rect 20188 92652 20244 92654
rect 20636 92652 20692 92708
rect 20300 92258 20356 92260
rect 20300 92206 20302 92258
rect 20302 92206 20354 92258
rect 20354 92206 20356 92258
rect 20300 92204 20356 92206
rect 20748 92428 20804 92484
rect 20300 91196 20356 91252
rect 19740 90578 19796 90580
rect 19740 90526 19742 90578
rect 19742 90526 19794 90578
rect 19794 90526 19796 90578
rect 19740 90524 19796 90526
rect 20188 90300 20244 90356
rect 19964 89682 20020 89684
rect 19964 89630 19966 89682
rect 19966 89630 20018 89682
rect 20018 89630 20020 89682
rect 19964 89628 20020 89630
rect 19628 89292 19684 89348
rect 19628 88732 19684 88788
rect 19292 88226 19348 88228
rect 19292 88174 19294 88226
rect 19294 88174 19346 88226
rect 19346 88174 19348 88226
rect 19292 88172 19348 88174
rect 19180 88114 19236 88116
rect 19180 88062 19182 88114
rect 19182 88062 19234 88114
rect 19234 88062 19236 88114
rect 19180 88060 19236 88062
rect 19404 87612 19460 87668
rect 19180 86658 19236 86660
rect 19180 86606 19182 86658
rect 19182 86606 19234 86658
rect 19234 86606 19236 86658
rect 19180 86604 19236 86606
rect 18172 85708 18228 85764
rect 18732 85820 18788 85876
rect 18222 85482 18278 85484
rect 18222 85430 18224 85482
rect 18224 85430 18276 85482
rect 18276 85430 18278 85482
rect 18222 85428 18278 85430
rect 18326 85482 18382 85484
rect 18326 85430 18328 85482
rect 18328 85430 18380 85482
rect 18380 85430 18382 85482
rect 18326 85428 18382 85430
rect 18430 85482 18486 85484
rect 18430 85430 18432 85482
rect 18432 85430 18484 85482
rect 18484 85430 18486 85482
rect 18430 85428 18486 85430
rect 17052 84364 17108 84420
rect 15932 75292 15988 75348
rect 16044 74620 16100 74676
rect 16604 79548 16660 79604
rect 16492 76466 16548 76468
rect 16492 76414 16494 76466
rect 16494 76414 16546 76466
rect 16546 76414 16548 76466
rect 16492 76412 16548 76414
rect 16380 75068 16436 75124
rect 16492 74620 16548 74676
rect 15820 73388 15876 73444
rect 15820 73164 15876 73220
rect 16268 72604 16324 72660
rect 15932 72380 15988 72436
rect 15596 72268 15652 72324
rect 16380 72546 16436 72548
rect 16380 72494 16382 72546
rect 16382 72494 16434 72546
rect 16434 72494 16436 72546
rect 16380 72492 16436 72494
rect 16380 72044 16436 72100
rect 15484 71708 15540 71764
rect 15708 71762 15764 71764
rect 15708 71710 15710 71762
rect 15710 71710 15762 71762
rect 15762 71710 15764 71762
rect 15708 71708 15764 71710
rect 16492 71932 16548 71988
rect 15372 71484 15428 71540
rect 16156 71484 16212 71540
rect 15484 70812 15540 70868
rect 14028 67340 14084 67396
rect 13580 66444 13636 66500
rect 13468 66274 13524 66276
rect 13468 66222 13470 66274
rect 13470 66222 13522 66274
rect 13522 66222 13524 66274
rect 13468 66220 13524 66222
rect 13804 66220 13860 66276
rect 14252 66274 14308 66276
rect 14252 66222 14254 66274
rect 14254 66222 14306 66274
rect 14306 66222 14308 66274
rect 14252 66220 14308 66222
rect 13692 65996 13748 66052
rect 13468 65602 13524 65604
rect 13468 65550 13470 65602
rect 13470 65550 13522 65602
rect 13522 65550 13524 65602
rect 13468 65548 13524 65550
rect 13804 65324 13860 65380
rect 14588 70476 14644 70532
rect 14820 70586 14876 70588
rect 14820 70534 14822 70586
rect 14822 70534 14874 70586
rect 14874 70534 14876 70586
rect 14820 70532 14876 70534
rect 14924 70586 14980 70588
rect 14924 70534 14926 70586
rect 14926 70534 14978 70586
rect 14978 70534 14980 70586
rect 14924 70532 14980 70534
rect 15028 70586 15084 70588
rect 15028 70534 15030 70586
rect 15030 70534 15082 70586
rect 15082 70534 15084 70586
rect 15028 70532 15084 70534
rect 15148 70140 15204 70196
rect 15036 70028 15092 70084
rect 16044 70924 16100 70980
rect 15596 70588 15652 70644
rect 15484 69916 15540 69972
rect 15036 69468 15092 69524
rect 14812 69410 14868 69412
rect 14812 69358 14814 69410
rect 14814 69358 14866 69410
rect 14866 69358 14868 69410
rect 14812 69356 14868 69358
rect 15260 69298 15316 69300
rect 15260 69246 15262 69298
rect 15262 69246 15314 69298
rect 15314 69246 15316 69298
rect 15260 69244 15316 69246
rect 14700 69132 14756 69188
rect 14820 69018 14876 69020
rect 14820 68966 14822 69018
rect 14822 68966 14874 69018
rect 14874 68966 14876 69018
rect 14820 68964 14876 68966
rect 14924 69018 14980 69020
rect 14924 68966 14926 69018
rect 14926 68966 14978 69018
rect 14978 68966 14980 69018
rect 14924 68964 14980 68966
rect 15028 69018 15084 69020
rect 15028 68966 15030 69018
rect 15030 68966 15082 69018
rect 15082 68966 15084 69018
rect 15028 68964 15084 68966
rect 15820 69916 15876 69972
rect 16380 70924 16436 70980
rect 16492 71596 16548 71652
rect 15932 69468 15988 69524
rect 15596 69132 15652 69188
rect 16156 69244 16212 69300
rect 15596 68908 15652 68964
rect 14588 68572 14644 68628
rect 15820 68684 15876 68740
rect 14476 68236 14532 68292
rect 14820 67450 14876 67452
rect 14820 67398 14822 67450
rect 14822 67398 14874 67450
rect 14874 67398 14876 67450
rect 14820 67396 14876 67398
rect 14924 67450 14980 67452
rect 14924 67398 14926 67450
rect 14926 67398 14978 67450
rect 14978 67398 14980 67450
rect 14924 67396 14980 67398
rect 15028 67450 15084 67452
rect 15028 67398 15030 67450
rect 15030 67398 15082 67450
rect 15082 67398 15084 67450
rect 15028 67396 15084 67398
rect 16268 69132 16324 69188
rect 16044 68572 16100 68628
rect 15484 66834 15540 66836
rect 15484 66782 15486 66834
rect 15486 66782 15538 66834
rect 15538 66782 15540 66834
rect 15484 66780 15540 66782
rect 15260 66332 15316 66388
rect 14476 65772 14532 65828
rect 14820 65882 14876 65884
rect 14820 65830 14822 65882
rect 14822 65830 14874 65882
rect 14874 65830 14876 65882
rect 14820 65828 14876 65830
rect 14924 65882 14980 65884
rect 14924 65830 14926 65882
rect 14926 65830 14978 65882
rect 14978 65830 14980 65882
rect 14924 65828 14980 65830
rect 15028 65882 15084 65884
rect 15028 65830 15030 65882
rect 15030 65830 15082 65882
rect 15082 65830 15084 65882
rect 15028 65828 15084 65830
rect 16492 67340 16548 67396
rect 14476 65602 14532 65604
rect 14476 65550 14478 65602
rect 14478 65550 14530 65602
rect 14530 65550 14532 65602
rect 14476 65548 14532 65550
rect 14364 65436 14420 65492
rect 16380 66834 16436 66836
rect 16380 66782 16382 66834
rect 16382 66782 16434 66834
rect 16434 66782 16436 66834
rect 16380 66780 16436 66782
rect 14028 65324 14084 65380
rect 15484 65436 15540 65492
rect 14812 65324 14868 65380
rect 15596 64764 15652 64820
rect 14252 64482 14308 64484
rect 14252 64430 14254 64482
rect 14254 64430 14306 64482
rect 14306 64430 14308 64482
rect 14252 64428 14308 64430
rect 14820 64314 14876 64316
rect 14820 64262 14822 64314
rect 14822 64262 14874 64314
rect 14874 64262 14876 64314
rect 14820 64260 14876 64262
rect 14924 64314 14980 64316
rect 14924 64262 14926 64314
rect 14926 64262 14978 64314
rect 14978 64262 14980 64314
rect 14924 64260 14980 64262
rect 15028 64314 15084 64316
rect 15028 64262 15030 64314
rect 15030 64262 15082 64314
rect 15082 64262 15084 64314
rect 15028 64260 15084 64262
rect 13356 63868 13412 63924
rect 13916 63644 13972 63700
rect 13468 63138 13524 63140
rect 13468 63086 13470 63138
rect 13470 63086 13522 63138
rect 13522 63086 13524 63138
rect 13468 63084 13524 63086
rect 14924 63532 14980 63588
rect 14476 63308 14532 63364
rect 13916 63084 13972 63140
rect 15484 63308 15540 63364
rect 15820 63420 15876 63476
rect 14028 62914 14084 62916
rect 14028 62862 14030 62914
rect 14030 62862 14082 62914
rect 14082 62862 14084 62914
rect 14028 62860 14084 62862
rect 13916 62636 13972 62692
rect 14820 62746 14876 62748
rect 14820 62694 14822 62746
rect 14822 62694 14874 62746
rect 14874 62694 14876 62746
rect 14820 62692 14876 62694
rect 14924 62746 14980 62748
rect 14924 62694 14926 62746
rect 14926 62694 14978 62746
rect 14978 62694 14980 62746
rect 14924 62692 14980 62694
rect 15028 62746 15084 62748
rect 15028 62694 15030 62746
rect 15030 62694 15082 62746
rect 15082 62694 15084 62746
rect 15028 62692 15084 62694
rect 14364 62354 14420 62356
rect 14364 62302 14366 62354
rect 14366 62302 14418 62354
rect 14418 62302 14420 62354
rect 14364 62300 14420 62302
rect 13580 61740 13636 61796
rect 14364 61852 14420 61908
rect 13916 61458 13972 61460
rect 13916 61406 13918 61458
rect 13918 61406 13970 61458
rect 13970 61406 13972 61458
rect 13916 61404 13972 61406
rect 13804 60732 13860 60788
rect 14140 61292 14196 61348
rect 14028 60732 14084 60788
rect 13692 60172 13748 60228
rect 13356 58940 13412 58996
rect 15372 62354 15428 62356
rect 15372 62302 15374 62354
rect 15374 62302 15426 62354
rect 15426 62302 15428 62354
rect 15372 62300 15428 62302
rect 14924 61570 14980 61572
rect 14924 61518 14926 61570
rect 14926 61518 14978 61570
rect 14978 61518 14980 61570
rect 14924 61516 14980 61518
rect 15260 61570 15316 61572
rect 15260 61518 15262 61570
rect 15262 61518 15314 61570
rect 15314 61518 15316 61570
rect 15260 61516 15316 61518
rect 14820 61178 14876 61180
rect 14820 61126 14822 61178
rect 14822 61126 14874 61178
rect 14874 61126 14876 61178
rect 14820 61124 14876 61126
rect 14924 61178 14980 61180
rect 14924 61126 14926 61178
rect 14926 61126 14978 61178
rect 14978 61126 14980 61178
rect 14924 61124 14980 61126
rect 15028 61178 15084 61180
rect 15028 61126 15030 61178
rect 15030 61126 15082 61178
rect 15082 61126 15084 61178
rect 15028 61124 15084 61126
rect 14252 60396 14308 60452
rect 14364 60732 14420 60788
rect 14252 60060 14308 60116
rect 13916 59836 13972 59892
rect 13804 59724 13860 59780
rect 14028 59778 14084 59780
rect 14028 59726 14030 59778
rect 14030 59726 14082 59778
rect 14082 59726 14084 59778
rect 14028 59724 14084 59726
rect 14364 59948 14420 60004
rect 13580 58716 13636 58772
rect 13468 57874 13524 57876
rect 13468 57822 13470 57874
rect 13470 57822 13522 57874
rect 13522 57822 13524 57874
rect 13468 57820 13524 57822
rect 13580 57372 13636 57428
rect 13804 58492 13860 58548
rect 14028 58322 14084 58324
rect 14028 58270 14030 58322
rect 14030 58270 14082 58322
rect 14082 58270 14084 58322
rect 14028 58268 14084 58270
rect 13244 56140 13300 56196
rect 12908 56082 12964 56084
rect 12908 56030 12910 56082
rect 12910 56030 12962 56082
rect 12962 56030 12964 56082
rect 12908 56028 12964 56030
rect 12796 55468 12852 55524
rect 12908 55692 12964 55748
rect 12796 54626 12852 54628
rect 12796 54574 12798 54626
rect 12798 54574 12850 54626
rect 12850 54574 12852 54626
rect 12796 54572 12852 54574
rect 12348 54012 12404 54068
rect 12348 53564 12404 53620
rect 12348 52556 12404 52612
rect 11452 49980 11508 50036
rect 11900 49980 11956 50036
rect 11228 49810 11284 49812
rect 11228 49758 11230 49810
rect 11230 49758 11282 49810
rect 11282 49758 11284 49810
rect 11228 49756 11284 49758
rect 11900 49756 11956 49812
rect 11418 49418 11474 49420
rect 11418 49366 11420 49418
rect 11420 49366 11472 49418
rect 11472 49366 11474 49418
rect 11418 49364 11474 49366
rect 11522 49418 11578 49420
rect 11522 49366 11524 49418
rect 11524 49366 11576 49418
rect 11576 49366 11578 49418
rect 11522 49364 11578 49366
rect 11626 49418 11682 49420
rect 11626 49366 11628 49418
rect 11628 49366 11680 49418
rect 11680 49366 11682 49418
rect 11626 49364 11682 49366
rect 10780 49308 10836 49364
rect 11340 49196 11396 49252
rect 11116 49084 11172 49140
rect 11004 48860 11060 48916
rect 10892 48188 10948 48244
rect 10780 48130 10836 48132
rect 10780 48078 10782 48130
rect 10782 48078 10834 48130
rect 10834 48078 10836 48130
rect 10780 48076 10836 48078
rect 10108 47852 10164 47908
rect 10332 47740 10388 47796
rect 10220 47628 10276 47684
rect 10556 47740 10612 47796
rect 10108 47292 10164 47348
rect 9996 47012 10052 47068
rect 10444 47346 10500 47348
rect 10444 47294 10446 47346
rect 10446 47294 10498 47346
rect 10498 47294 10500 47346
rect 10444 47292 10500 47294
rect 10780 47292 10836 47348
rect 10668 47180 10724 47236
rect 10332 47068 10388 47124
rect 10108 46508 10164 46564
rect 10556 47068 10612 47124
rect 9436 45890 9492 45892
rect 9436 45838 9438 45890
rect 9438 45838 9490 45890
rect 9490 45838 9492 45890
rect 9436 45836 9492 45838
rect 9436 45500 9492 45556
rect 9772 45388 9828 45444
rect 10332 46508 10388 46564
rect 10444 45612 10500 45668
rect 9548 45218 9604 45220
rect 9548 45166 9550 45218
rect 9550 45166 9602 45218
rect 9602 45166 9604 45218
rect 9548 45164 9604 45166
rect 9436 44546 9492 44548
rect 9436 44494 9438 44546
rect 9438 44494 9490 44546
rect 9490 44494 9492 44546
rect 9436 44492 9492 44494
rect 9100 38162 9156 38164
rect 9100 38110 9102 38162
rect 9102 38110 9154 38162
rect 9154 38110 9156 38162
rect 9100 38108 9156 38110
rect 7868 35644 7924 35700
rect 7756 34802 7812 34804
rect 7756 34750 7758 34802
rect 7758 34750 7810 34802
rect 7810 34750 7812 34802
rect 7756 34748 7812 34750
rect 8540 35922 8596 35924
rect 8540 35870 8542 35922
rect 8542 35870 8594 35922
rect 8594 35870 8596 35922
rect 8540 35868 8596 35870
rect 8764 35756 8820 35812
rect 8652 35026 8708 35028
rect 8652 34974 8654 35026
rect 8654 34974 8706 35026
rect 8706 34974 8708 35026
rect 8652 34972 8708 34974
rect 8016 34522 8072 34524
rect 8016 34470 8018 34522
rect 8018 34470 8070 34522
rect 8070 34470 8072 34522
rect 8016 34468 8072 34470
rect 8120 34522 8176 34524
rect 8120 34470 8122 34522
rect 8122 34470 8174 34522
rect 8174 34470 8176 34522
rect 8120 34468 8176 34470
rect 8224 34522 8280 34524
rect 8224 34470 8226 34522
rect 8226 34470 8278 34522
rect 8278 34470 8280 34522
rect 8224 34468 8280 34470
rect 8652 34802 8708 34804
rect 8652 34750 8654 34802
rect 8654 34750 8706 34802
rect 8706 34750 8708 34802
rect 8652 34748 8708 34750
rect 8428 34300 8484 34356
rect 7868 34130 7924 34132
rect 7868 34078 7870 34130
rect 7870 34078 7922 34130
rect 7922 34078 7924 34130
rect 7868 34076 7924 34078
rect 8092 34130 8148 34132
rect 8092 34078 8094 34130
rect 8094 34078 8146 34130
rect 8146 34078 8148 34130
rect 8092 34076 8148 34078
rect 7644 31276 7700 31332
rect 7756 33628 7812 33684
rect 7644 31052 7700 31108
rect 7532 30994 7588 30996
rect 7532 30942 7534 30994
rect 7534 30942 7586 30994
rect 7586 30942 7588 30994
rect 7532 30940 7588 30942
rect 6860 29820 6916 29876
rect 7308 30268 7364 30324
rect 7196 29820 7252 29876
rect 7084 29484 7140 29540
rect 6860 28754 6916 28756
rect 6860 28702 6862 28754
rect 6862 28702 6914 28754
rect 6914 28702 6916 28754
rect 6860 28700 6916 28702
rect 7644 30322 7700 30324
rect 7644 30270 7646 30322
rect 7646 30270 7698 30322
rect 7698 30270 7700 30322
rect 7644 30268 7700 30270
rect 8316 33964 8372 34020
rect 8428 33852 8484 33908
rect 8540 33628 8596 33684
rect 8652 33740 8708 33796
rect 8204 33404 8260 33460
rect 8016 32954 8072 32956
rect 8016 32902 8018 32954
rect 8018 32902 8070 32954
rect 8070 32902 8072 32954
rect 8016 32900 8072 32902
rect 8120 32954 8176 32956
rect 8120 32902 8122 32954
rect 8122 32902 8174 32954
rect 8174 32902 8176 32954
rect 8120 32900 8176 32902
rect 8224 32954 8280 32956
rect 8224 32902 8226 32954
rect 8226 32902 8278 32954
rect 8278 32902 8280 32954
rect 8224 32900 8280 32902
rect 8988 34748 9044 34804
rect 9100 34412 9156 34468
rect 8988 33852 9044 33908
rect 9100 34076 9156 34132
rect 8764 32732 8820 32788
rect 8764 32450 8820 32452
rect 8764 32398 8766 32450
rect 8766 32398 8818 32450
rect 8818 32398 8820 32450
rect 8764 32396 8820 32398
rect 8764 32172 8820 32228
rect 8016 31386 8072 31388
rect 8016 31334 8018 31386
rect 8018 31334 8070 31386
rect 8070 31334 8072 31386
rect 8016 31332 8072 31334
rect 8120 31386 8176 31388
rect 8120 31334 8122 31386
rect 8122 31334 8174 31386
rect 8174 31334 8176 31386
rect 8120 31332 8176 31334
rect 8224 31386 8280 31388
rect 8224 31334 8226 31386
rect 8226 31334 8278 31386
rect 8278 31334 8280 31386
rect 8224 31332 8280 31334
rect 7980 31052 8036 31108
rect 8428 30994 8484 30996
rect 8428 30942 8430 30994
rect 8430 30942 8482 30994
rect 8482 30942 8484 30994
rect 8428 30940 8484 30942
rect 8092 30882 8148 30884
rect 8092 30830 8094 30882
rect 8094 30830 8146 30882
rect 8146 30830 8148 30882
rect 8092 30828 8148 30830
rect 7868 30492 7924 30548
rect 8092 30380 8148 30436
rect 8428 30380 8484 30436
rect 6412 27186 6468 27188
rect 6412 27134 6414 27186
rect 6414 27134 6466 27186
rect 6466 27134 6468 27186
rect 6412 27132 6468 27134
rect 6860 27244 6916 27300
rect 6748 27074 6804 27076
rect 6748 27022 6750 27074
rect 6750 27022 6802 27074
rect 6802 27022 6804 27074
rect 6748 27020 6804 27022
rect 6188 26348 6244 26404
rect 7308 27132 7364 27188
rect 6412 25564 6468 25620
rect 6636 25452 6692 25508
rect 6076 24892 6132 24948
rect 5516 22540 5572 22596
rect 6636 23266 6692 23268
rect 6636 23214 6638 23266
rect 6638 23214 6690 23266
rect 6690 23214 6692 23266
rect 6636 23212 6692 23214
rect 6300 22988 6356 23044
rect 6188 20690 6244 20692
rect 6188 20638 6190 20690
rect 6190 20638 6242 20690
rect 6242 20638 6244 20690
rect 6188 20636 6244 20638
rect 6860 21308 6916 21364
rect 7196 25228 7252 25284
rect 8316 29932 8372 29988
rect 8016 29818 8072 29820
rect 8016 29766 8018 29818
rect 8018 29766 8070 29818
rect 8070 29766 8072 29818
rect 8016 29764 8072 29766
rect 8120 29818 8176 29820
rect 8120 29766 8122 29818
rect 8122 29766 8174 29818
rect 8174 29766 8176 29818
rect 8120 29764 8176 29766
rect 8224 29818 8280 29820
rect 8224 29766 8226 29818
rect 8226 29766 8278 29818
rect 8278 29766 8280 29818
rect 8540 29820 8596 29876
rect 8224 29764 8280 29766
rect 8540 29036 8596 29092
rect 7756 28700 7812 28756
rect 8016 28250 8072 28252
rect 8016 28198 8018 28250
rect 8018 28198 8070 28250
rect 8070 28198 8072 28250
rect 8016 28196 8072 28198
rect 8120 28250 8176 28252
rect 8120 28198 8122 28250
rect 8122 28198 8174 28250
rect 8174 28198 8176 28250
rect 8120 28196 8176 28198
rect 8224 28250 8280 28252
rect 8224 28198 8226 28250
rect 8226 28198 8278 28250
rect 8278 28198 8280 28250
rect 8224 28196 8280 28198
rect 7756 27186 7812 27188
rect 7756 27134 7758 27186
rect 7758 27134 7810 27186
rect 7810 27134 7812 27186
rect 7756 27132 7812 27134
rect 8092 27804 8148 27860
rect 8316 27132 8372 27188
rect 7196 22988 7252 23044
rect 7308 22930 7364 22932
rect 7308 22878 7310 22930
rect 7310 22878 7362 22930
rect 7362 22878 7364 22930
rect 7308 22876 7364 22878
rect 7196 21084 7252 21140
rect 6636 20188 6692 20244
rect 5404 20130 5460 20132
rect 5404 20078 5406 20130
rect 5406 20078 5458 20130
rect 5458 20078 5460 20130
rect 5404 20076 5460 20078
rect 7084 20690 7140 20692
rect 7084 20638 7086 20690
rect 7086 20638 7138 20690
rect 7138 20638 7140 20690
rect 7084 20636 7140 20638
rect 6412 19292 6468 19348
rect 8016 26682 8072 26684
rect 8016 26630 8018 26682
rect 8018 26630 8070 26682
rect 8070 26630 8072 26682
rect 8016 26628 8072 26630
rect 8120 26682 8176 26684
rect 8120 26630 8122 26682
rect 8122 26630 8174 26682
rect 8174 26630 8176 26682
rect 8120 26628 8176 26630
rect 8224 26682 8280 26684
rect 8224 26630 8226 26682
rect 8226 26630 8278 26682
rect 8278 26630 8280 26682
rect 8224 26628 8280 26630
rect 8016 25114 8072 25116
rect 8016 25062 8018 25114
rect 8018 25062 8070 25114
rect 8070 25062 8072 25114
rect 8016 25060 8072 25062
rect 8120 25114 8176 25116
rect 8120 25062 8122 25114
rect 8122 25062 8174 25114
rect 8174 25062 8176 25114
rect 8120 25060 8176 25062
rect 8224 25114 8280 25116
rect 8224 25062 8226 25114
rect 8226 25062 8278 25114
rect 8278 25062 8280 25114
rect 8224 25060 8280 25062
rect 7756 24946 7812 24948
rect 7756 24894 7758 24946
rect 7758 24894 7810 24946
rect 7810 24894 7812 24946
rect 7756 24892 7812 24894
rect 8016 23546 8072 23548
rect 8016 23494 8018 23546
rect 8018 23494 8070 23546
rect 8070 23494 8072 23546
rect 8016 23492 8072 23494
rect 8120 23546 8176 23548
rect 8120 23494 8122 23546
rect 8122 23494 8174 23546
rect 8174 23494 8176 23546
rect 8120 23492 8176 23494
rect 8224 23546 8280 23548
rect 8224 23494 8226 23546
rect 8226 23494 8278 23546
rect 8278 23494 8280 23546
rect 8224 23492 8280 23494
rect 7532 23266 7588 23268
rect 7532 23214 7534 23266
rect 7534 23214 7586 23266
rect 7586 23214 7588 23266
rect 7532 23212 7588 23214
rect 7420 20972 7476 21028
rect 8316 22876 8372 22932
rect 8204 22540 8260 22596
rect 7308 20690 7364 20692
rect 7308 20638 7310 20690
rect 7310 20638 7362 20690
rect 7362 20638 7364 20690
rect 7308 20636 7364 20638
rect 8016 21978 8072 21980
rect 8016 21926 8018 21978
rect 8018 21926 8070 21978
rect 8070 21926 8072 21978
rect 8016 21924 8072 21926
rect 8120 21978 8176 21980
rect 8120 21926 8122 21978
rect 8122 21926 8174 21978
rect 8174 21926 8176 21978
rect 8120 21924 8176 21926
rect 8224 21978 8280 21980
rect 8224 21926 8226 21978
rect 8226 21926 8278 21978
rect 8278 21926 8280 21978
rect 8224 21924 8280 21926
rect 8540 27356 8596 27412
rect 9100 30940 9156 30996
rect 8876 30882 8932 30884
rect 8876 30830 8878 30882
rect 8878 30830 8930 30882
rect 8930 30830 8932 30882
rect 8876 30828 8932 30830
rect 9324 42924 9380 42980
rect 9324 36988 9380 37044
rect 8988 30044 9044 30100
rect 8988 29820 9044 29876
rect 8988 27858 9044 27860
rect 8988 27806 8990 27858
rect 8990 27806 9042 27858
rect 9042 27806 9044 27858
rect 8988 27804 9044 27806
rect 8876 27692 8932 27748
rect 9324 30098 9380 30100
rect 9324 30046 9326 30098
rect 9326 30046 9378 30098
rect 9378 30046 9380 30098
rect 9324 30044 9380 30046
rect 9212 27580 9268 27636
rect 9212 27244 9268 27300
rect 8988 25228 9044 25284
rect 8652 23436 8708 23492
rect 8652 22540 8708 22596
rect 7980 21644 8036 21700
rect 8428 21698 8484 21700
rect 8428 21646 8430 21698
rect 8430 21646 8482 21698
rect 8482 21646 8484 21698
rect 8428 21644 8484 21646
rect 8316 21362 8372 21364
rect 8316 21310 8318 21362
rect 8318 21310 8370 21362
rect 8370 21310 8372 21362
rect 8316 21308 8372 21310
rect 8204 20914 8260 20916
rect 8204 20862 8206 20914
rect 8206 20862 8258 20914
rect 8258 20862 8260 20914
rect 8204 20860 8260 20862
rect 7756 20690 7812 20692
rect 7756 20638 7758 20690
rect 7758 20638 7810 20690
rect 7810 20638 7812 20690
rect 7756 20636 7812 20638
rect 8016 20410 8072 20412
rect 8016 20358 8018 20410
rect 8018 20358 8070 20410
rect 8070 20358 8072 20410
rect 8016 20356 8072 20358
rect 8120 20410 8176 20412
rect 8120 20358 8122 20410
rect 8122 20358 8174 20410
rect 8174 20358 8176 20410
rect 8120 20356 8176 20358
rect 8224 20410 8280 20412
rect 8224 20358 8226 20410
rect 8226 20358 8278 20410
rect 8278 20358 8280 20410
rect 8224 20356 8280 20358
rect 7196 19292 7252 19348
rect 6076 19234 6132 19236
rect 6076 19182 6078 19234
rect 6078 19182 6130 19234
rect 6130 19182 6132 19234
rect 6076 19180 6132 19182
rect 5964 18956 6020 19012
rect 5740 17724 5796 17780
rect 6636 19234 6692 19236
rect 6636 19182 6638 19234
rect 6638 19182 6690 19234
rect 6690 19182 6692 19234
rect 6636 19180 6692 19182
rect 6524 19010 6580 19012
rect 6524 18958 6526 19010
rect 6526 18958 6578 19010
rect 6578 18958 6580 19010
rect 6524 18956 6580 18958
rect 6636 18508 6692 18564
rect 6636 17724 6692 17780
rect 6076 16882 6132 16884
rect 6076 16830 6078 16882
rect 6078 16830 6130 16882
rect 6130 16830 6132 16882
rect 6076 16828 6132 16830
rect 5628 16770 5684 16772
rect 5628 16718 5630 16770
rect 5630 16718 5682 16770
rect 5682 16718 5684 16770
rect 5628 16716 5684 16718
rect 6076 15372 6132 15428
rect 6188 15260 6244 15316
rect 5628 15202 5684 15204
rect 5628 15150 5630 15202
rect 5630 15150 5682 15202
rect 5682 15150 5684 15202
rect 5628 15148 5684 15150
rect 5068 14588 5124 14644
rect 4284 12124 4340 12180
rect 4956 13580 5012 13636
rect 4614 13354 4670 13356
rect 4614 13302 4616 13354
rect 4616 13302 4668 13354
rect 4668 13302 4670 13354
rect 4614 13300 4670 13302
rect 4718 13354 4774 13356
rect 4718 13302 4720 13354
rect 4720 13302 4772 13354
rect 4772 13302 4774 13354
rect 4718 13300 4774 13302
rect 4822 13354 4878 13356
rect 4822 13302 4824 13354
rect 4824 13302 4876 13354
rect 4876 13302 4878 13354
rect 4822 13300 4878 13302
rect 5516 14588 5572 14644
rect 5964 14418 6020 14420
rect 5964 14366 5966 14418
rect 5966 14366 6018 14418
rect 6018 14366 6020 14418
rect 5964 14364 6020 14366
rect 5852 14252 5908 14308
rect 5516 13020 5572 13076
rect 4614 11786 4670 11788
rect 4614 11734 4616 11786
rect 4616 11734 4668 11786
rect 4668 11734 4670 11786
rect 4614 11732 4670 11734
rect 4718 11786 4774 11788
rect 4718 11734 4720 11786
rect 4720 11734 4772 11786
rect 4772 11734 4774 11786
rect 4718 11732 4774 11734
rect 4822 11786 4878 11788
rect 4822 11734 4824 11786
rect 4824 11734 4876 11786
rect 4876 11734 4878 11786
rect 4822 11732 4878 11734
rect 4508 11340 4564 11396
rect 4284 11116 4340 11172
rect 4956 11282 5012 11284
rect 4956 11230 4958 11282
rect 4958 11230 5010 11282
rect 5010 11230 5012 11282
rect 4956 11228 5012 11230
rect 3948 9100 4004 9156
rect 3388 6524 3444 6580
rect 2044 6300 2100 6356
rect 1708 4732 1764 4788
rect 2492 4732 2548 4788
rect 5068 10780 5124 10836
rect 4614 10218 4670 10220
rect 4614 10166 4616 10218
rect 4616 10166 4668 10218
rect 4668 10166 4670 10218
rect 4614 10164 4670 10166
rect 4718 10218 4774 10220
rect 4718 10166 4720 10218
rect 4720 10166 4772 10218
rect 4772 10166 4774 10218
rect 4718 10164 4774 10166
rect 4822 10218 4878 10220
rect 4822 10166 4824 10218
rect 4824 10166 4876 10218
rect 4876 10166 4878 10218
rect 4822 10164 4878 10166
rect 5068 10108 5124 10164
rect 5180 11228 5236 11284
rect 4844 9996 4900 10052
rect 4508 9884 4564 9940
rect 5964 13468 6020 13524
rect 5964 12348 6020 12404
rect 5852 11340 5908 11396
rect 6188 12850 6244 12852
rect 6188 12798 6190 12850
rect 6190 12798 6242 12850
rect 6242 12798 6244 12850
rect 6188 12796 6244 12798
rect 6524 15538 6580 15540
rect 6524 15486 6526 15538
rect 6526 15486 6578 15538
rect 6578 15486 6580 15538
rect 6524 15484 6580 15486
rect 6412 11676 6468 11732
rect 6748 16716 6804 16772
rect 8652 20802 8708 20804
rect 8652 20750 8654 20802
rect 8654 20750 8706 20802
rect 8706 20750 8708 20802
rect 8652 20748 8708 20750
rect 9100 24668 9156 24724
rect 9212 23660 9268 23716
rect 9660 44716 9716 44772
rect 9772 44156 9828 44212
rect 9660 43426 9716 43428
rect 9660 43374 9662 43426
rect 9662 43374 9714 43426
rect 9714 43374 9716 43426
rect 9660 43372 9716 43374
rect 9660 43148 9716 43204
rect 9660 42924 9716 42980
rect 9548 42252 9604 42308
rect 9548 41692 9604 41748
rect 9548 40290 9604 40292
rect 9548 40238 9550 40290
rect 9550 40238 9602 40290
rect 9602 40238 9604 40290
rect 9548 40236 9604 40238
rect 9548 40012 9604 40068
rect 9548 39116 9604 39172
rect 10108 44940 10164 44996
rect 11228 48412 11284 48468
rect 11788 49026 11844 49028
rect 11788 48974 11790 49026
rect 11790 48974 11842 49026
rect 11842 48974 11844 49026
rect 11788 48972 11844 48974
rect 11788 48636 11844 48692
rect 11418 47850 11474 47852
rect 11418 47798 11420 47850
rect 11420 47798 11472 47850
rect 11472 47798 11474 47850
rect 11418 47796 11474 47798
rect 11522 47850 11578 47852
rect 11522 47798 11524 47850
rect 11524 47798 11576 47850
rect 11576 47798 11578 47850
rect 11522 47796 11578 47798
rect 11626 47850 11682 47852
rect 11626 47798 11628 47850
rect 11628 47798 11680 47850
rect 11680 47798 11682 47850
rect 11626 47796 11682 47798
rect 11452 47628 11508 47684
rect 10892 46956 10948 47012
rect 11340 47292 11396 47348
rect 10892 46732 10948 46788
rect 10668 44492 10724 44548
rect 10780 44828 10836 44884
rect 12236 50316 12292 50372
rect 13132 54348 13188 54404
rect 12908 53842 12964 53844
rect 12908 53790 12910 53842
rect 12910 53790 12962 53842
rect 12962 53790 12964 53842
rect 12908 53788 12964 53790
rect 13132 53676 13188 53732
rect 14476 58828 14532 58884
rect 14364 58268 14420 58324
rect 14476 58604 14532 58660
rect 14924 60508 14980 60564
rect 14820 59610 14876 59612
rect 14820 59558 14822 59610
rect 14822 59558 14874 59610
rect 14874 59558 14876 59610
rect 14820 59556 14876 59558
rect 14924 59610 14980 59612
rect 14924 59558 14926 59610
rect 14926 59558 14978 59610
rect 14978 59558 14980 59610
rect 14924 59556 14980 59558
rect 15028 59610 15084 59612
rect 15028 59558 15030 59610
rect 15030 59558 15082 59610
rect 15082 59558 15084 59610
rect 15028 59556 15084 59558
rect 14812 59388 14868 59444
rect 14700 59276 14756 59332
rect 13916 57036 13972 57092
rect 14364 58044 14420 58100
rect 13580 56978 13636 56980
rect 13580 56926 13582 56978
rect 13582 56926 13634 56978
rect 13634 56926 13636 56978
rect 13580 56924 13636 56926
rect 13804 56924 13860 56980
rect 13692 56476 13748 56532
rect 13692 56082 13748 56084
rect 13692 56030 13694 56082
rect 13694 56030 13746 56082
rect 13746 56030 13748 56082
rect 13692 56028 13748 56030
rect 13468 55356 13524 55412
rect 12684 53340 12740 53396
rect 13580 55244 13636 55300
rect 13580 54236 13636 54292
rect 13916 56364 13972 56420
rect 13916 55804 13972 55860
rect 14364 57260 14420 57316
rect 14588 58380 14644 58436
rect 14588 57372 14644 57428
rect 14588 56978 14644 56980
rect 14588 56926 14590 56978
rect 14590 56926 14642 56978
rect 14642 56926 14644 56978
rect 14588 56924 14644 56926
rect 15036 59164 15092 59220
rect 15036 58604 15092 58660
rect 15148 58380 15204 58436
rect 15260 60508 15316 60564
rect 15372 60284 15428 60340
rect 15596 62300 15652 62356
rect 16380 66386 16436 66388
rect 16380 66334 16382 66386
rect 16382 66334 16434 66386
rect 16434 66334 16436 66386
rect 16380 66332 16436 66334
rect 16380 65996 16436 66052
rect 16828 78316 16884 78372
rect 16940 81676 16996 81732
rect 16828 75794 16884 75796
rect 16828 75742 16830 75794
rect 16830 75742 16882 75794
rect 16882 75742 16884 75794
rect 16828 75740 16884 75742
rect 16828 74898 16884 74900
rect 16828 74846 16830 74898
rect 16830 74846 16882 74898
rect 16882 74846 16884 74898
rect 16828 74844 16884 74846
rect 16716 72604 16772 72660
rect 16716 72156 16772 72212
rect 16716 71148 16772 71204
rect 16828 70978 16884 70980
rect 16828 70926 16830 70978
rect 16830 70926 16882 70978
rect 16882 70926 16884 70978
rect 16828 70924 16884 70926
rect 16716 70700 16772 70756
rect 16716 69468 16772 69524
rect 17612 84306 17668 84308
rect 17612 84254 17614 84306
rect 17614 84254 17666 84306
rect 17666 84254 17668 84306
rect 17612 84252 17668 84254
rect 17052 80556 17108 80612
rect 17612 83298 17668 83300
rect 17612 83246 17614 83298
rect 17614 83246 17666 83298
rect 17666 83246 17668 83298
rect 17612 83244 17668 83246
rect 17500 82962 17556 82964
rect 17500 82910 17502 82962
rect 17502 82910 17554 82962
rect 17554 82910 17556 82962
rect 17500 82908 17556 82910
rect 17164 80892 17220 80948
rect 16940 69356 16996 69412
rect 17276 82348 17332 82404
rect 16828 69298 16884 69300
rect 16828 69246 16830 69298
rect 16830 69246 16882 69298
rect 16882 69246 16884 69298
rect 16828 69244 16884 69246
rect 16716 68796 16772 68852
rect 16940 68348 16996 68404
rect 16492 63980 16548 64036
rect 16604 64428 16660 64484
rect 16268 63420 16324 63476
rect 16380 63308 16436 63364
rect 16044 62300 16100 62356
rect 16268 62860 16324 62916
rect 15820 62076 15876 62132
rect 15596 61740 15652 61796
rect 15484 60172 15540 60228
rect 15820 60956 15876 61012
rect 16156 61180 16212 61236
rect 16268 61404 16324 61460
rect 16380 60620 16436 60676
rect 16268 60284 16324 60340
rect 15484 58716 15540 58772
rect 15596 58828 15652 58884
rect 14820 58042 14876 58044
rect 14820 57990 14822 58042
rect 14822 57990 14874 58042
rect 14874 57990 14876 58042
rect 14820 57988 14876 57990
rect 14924 58042 14980 58044
rect 14924 57990 14926 58042
rect 14926 57990 14978 58042
rect 14978 57990 14980 58042
rect 14924 57988 14980 57990
rect 15028 58042 15084 58044
rect 15028 57990 15030 58042
rect 15030 57990 15082 58042
rect 15082 57990 15084 58042
rect 15028 57988 15084 57990
rect 15260 57932 15316 57988
rect 15484 57148 15540 57204
rect 15372 56812 15428 56868
rect 15036 56700 15092 56756
rect 14820 56474 14876 56476
rect 14820 56422 14822 56474
rect 14822 56422 14874 56474
rect 14874 56422 14876 56474
rect 14820 56420 14876 56422
rect 14924 56474 14980 56476
rect 14924 56422 14926 56474
rect 14926 56422 14978 56474
rect 14978 56422 14980 56474
rect 14924 56420 14980 56422
rect 15028 56474 15084 56476
rect 15028 56422 15030 56474
rect 15030 56422 15082 56474
rect 15082 56422 15084 56474
rect 15028 56420 15084 56422
rect 15036 56194 15092 56196
rect 15036 56142 15038 56194
rect 15038 56142 15090 56194
rect 15090 56142 15092 56194
rect 15036 56140 15092 56142
rect 14140 55692 14196 55748
rect 14028 55132 14084 55188
rect 12572 53228 12628 53284
rect 12572 52444 12628 52500
rect 12572 50876 12628 50932
rect 12796 52556 12852 52612
rect 12460 50428 12516 50484
rect 12236 49084 12292 49140
rect 12348 49026 12404 49028
rect 12348 48974 12350 49026
rect 12350 48974 12402 49026
rect 12402 48974 12404 49026
rect 12348 48972 12404 48974
rect 12572 48914 12628 48916
rect 12572 48862 12574 48914
rect 12574 48862 12626 48914
rect 12626 48862 12628 48914
rect 12572 48860 12628 48862
rect 12236 48748 12292 48804
rect 12796 48860 12852 48916
rect 11788 47068 11844 47124
rect 12012 47404 12068 47460
rect 12236 47404 12292 47460
rect 12012 47234 12068 47236
rect 12012 47182 12014 47234
rect 12014 47182 12066 47234
rect 12066 47182 12068 47234
rect 12012 47180 12068 47182
rect 11452 46508 11508 46564
rect 11418 46282 11474 46284
rect 11418 46230 11420 46282
rect 11420 46230 11472 46282
rect 11472 46230 11474 46282
rect 11418 46228 11474 46230
rect 11522 46282 11578 46284
rect 11522 46230 11524 46282
rect 11524 46230 11576 46282
rect 11576 46230 11578 46282
rect 11522 46228 11578 46230
rect 11626 46282 11682 46284
rect 11626 46230 11628 46282
rect 11628 46230 11680 46282
rect 11680 46230 11682 46282
rect 11626 46228 11682 46230
rect 11116 45778 11172 45780
rect 11116 45726 11118 45778
rect 11118 45726 11170 45778
rect 11170 45726 11172 45778
rect 11116 45724 11172 45726
rect 11676 45778 11732 45780
rect 11676 45726 11678 45778
rect 11678 45726 11730 45778
rect 11730 45726 11732 45778
rect 11676 45724 11732 45726
rect 11452 45500 11508 45556
rect 10780 44380 10836 44436
rect 10556 43820 10612 43876
rect 10332 43036 10388 43092
rect 11004 43820 11060 43876
rect 11004 43650 11060 43652
rect 11004 43598 11006 43650
rect 11006 43598 11058 43650
rect 11058 43598 11060 43650
rect 11004 43596 11060 43598
rect 10892 43148 10948 43204
rect 9996 42252 10052 42308
rect 9884 42140 9940 42196
rect 9884 41858 9940 41860
rect 9884 41806 9886 41858
rect 9886 41806 9938 41858
rect 9938 41806 9940 41858
rect 9884 41804 9940 41806
rect 10780 42588 10836 42644
rect 10444 42476 10500 42532
rect 10444 41916 10500 41972
rect 10780 41804 10836 41860
rect 9996 41244 10052 41300
rect 10556 41298 10612 41300
rect 10556 41246 10558 41298
rect 10558 41246 10610 41298
rect 10610 41246 10612 41298
rect 10556 41244 10612 41246
rect 10332 40796 10388 40852
rect 11004 42530 11060 42532
rect 11004 42478 11006 42530
rect 11006 42478 11058 42530
rect 11058 42478 11060 42530
rect 11004 42476 11060 42478
rect 11418 44714 11474 44716
rect 11418 44662 11420 44714
rect 11420 44662 11472 44714
rect 11472 44662 11474 44714
rect 11418 44660 11474 44662
rect 11522 44714 11578 44716
rect 11522 44662 11524 44714
rect 11524 44662 11576 44714
rect 11576 44662 11578 44714
rect 11522 44660 11578 44662
rect 11626 44714 11682 44716
rect 11626 44662 11628 44714
rect 11628 44662 11680 44714
rect 11680 44662 11682 44714
rect 11626 44660 11682 44662
rect 12684 48466 12740 48468
rect 12684 48414 12686 48466
rect 12686 48414 12738 48466
rect 12738 48414 12740 48466
rect 12684 48412 12740 48414
rect 13692 52892 13748 52948
rect 13580 52556 13636 52612
rect 13692 52668 13748 52724
rect 13356 52332 13412 52388
rect 13244 50876 13300 50932
rect 13132 50652 13188 50708
rect 13020 50482 13076 50484
rect 13020 50430 13022 50482
rect 13022 50430 13074 50482
rect 13074 50430 13076 50482
rect 13020 50428 13076 50430
rect 13020 48748 13076 48804
rect 12460 47628 12516 47684
rect 12460 45948 12516 46004
rect 11900 45836 11956 45892
rect 12236 45778 12292 45780
rect 12236 45726 12238 45778
rect 12238 45726 12290 45778
rect 12290 45726 12292 45778
rect 12236 45724 12292 45726
rect 12124 45666 12180 45668
rect 12124 45614 12126 45666
rect 12126 45614 12178 45666
rect 12178 45614 12180 45666
rect 12124 45612 12180 45614
rect 12348 45164 12404 45220
rect 12124 44716 12180 44772
rect 11340 44380 11396 44436
rect 11340 43538 11396 43540
rect 11340 43486 11342 43538
rect 11342 43486 11394 43538
rect 11394 43486 11396 43538
rect 11340 43484 11396 43486
rect 10892 41244 10948 41300
rect 11676 44268 11732 44324
rect 11788 43484 11844 43540
rect 10780 40796 10836 40852
rect 10892 40684 10948 40740
rect 10108 40012 10164 40068
rect 9996 39116 10052 39172
rect 10668 39788 10724 39844
rect 10892 39116 10948 39172
rect 11418 43146 11474 43148
rect 11418 43094 11420 43146
rect 11420 43094 11472 43146
rect 11472 43094 11474 43146
rect 11418 43092 11474 43094
rect 11522 43146 11578 43148
rect 11522 43094 11524 43146
rect 11524 43094 11576 43146
rect 11576 43094 11578 43146
rect 11522 43092 11578 43094
rect 11626 43146 11682 43148
rect 11626 43094 11628 43146
rect 11628 43094 11680 43146
rect 11680 43094 11682 43146
rect 11626 43092 11682 43094
rect 11564 42530 11620 42532
rect 11564 42478 11566 42530
rect 11566 42478 11618 42530
rect 11618 42478 11620 42530
rect 11564 42476 11620 42478
rect 11228 42194 11284 42196
rect 11228 42142 11230 42194
rect 11230 42142 11282 42194
rect 11282 42142 11284 42194
rect 11228 42140 11284 42142
rect 11676 42082 11732 42084
rect 11676 42030 11678 42082
rect 11678 42030 11730 42082
rect 11730 42030 11732 42082
rect 11676 42028 11732 42030
rect 11418 41578 11474 41580
rect 11418 41526 11420 41578
rect 11420 41526 11472 41578
rect 11472 41526 11474 41578
rect 11418 41524 11474 41526
rect 11522 41578 11578 41580
rect 11522 41526 11524 41578
rect 11524 41526 11576 41578
rect 11576 41526 11578 41578
rect 11522 41524 11578 41526
rect 11626 41578 11682 41580
rect 11626 41526 11628 41578
rect 11628 41526 11680 41578
rect 11680 41526 11682 41578
rect 11626 41524 11682 41526
rect 11788 41298 11844 41300
rect 11788 41246 11790 41298
rect 11790 41246 11842 41298
rect 11842 41246 11844 41298
rect 11788 41244 11844 41246
rect 11228 40796 11284 40852
rect 11564 40684 11620 40740
rect 11228 40572 11284 40628
rect 11116 40514 11172 40516
rect 11116 40462 11118 40514
rect 11118 40462 11170 40514
rect 11170 40462 11172 40514
rect 11116 40460 11172 40462
rect 11788 40402 11844 40404
rect 11788 40350 11790 40402
rect 11790 40350 11842 40402
rect 11842 40350 11844 40402
rect 11788 40348 11844 40350
rect 11418 40010 11474 40012
rect 11418 39958 11420 40010
rect 11420 39958 11472 40010
rect 11472 39958 11474 40010
rect 11418 39956 11474 39958
rect 11522 40010 11578 40012
rect 11522 39958 11524 40010
rect 11524 39958 11576 40010
rect 11576 39958 11578 40010
rect 11522 39956 11578 39958
rect 11626 40010 11682 40012
rect 11626 39958 11628 40010
rect 11628 39958 11680 40010
rect 11680 39958 11682 40010
rect 11788 40012 11844 40068
rect 11626 39956 11682 39958
rect 11676 39788 11732 39844
rect 9660 38220 9716 38276
rect 10108 38108 10164 38164
rect 10780 38050 10836 38052
rect 10780 37998 10782 38050
rect 10782 37998 10834 38050
rect 10834 37998 10836 38050
rect 10780 37996 10836 37998
rect 10332 37548 10388 37604
rect 9660 37490 9716 37492
rect 9660 37438 9662 37490
rect 9662 37438 9714 37490
rect 9714 37438 9716 37490
rect 9660 37436 9716 37438
rect 10108 37378 10164 37380
rect 10108 37326 10110 37378
rect 10110 37326 10162 37378
rect 10162 37326 10164 37378
rect 10108 37324 10164 37326
rect 9996 37266 10052 37268
rect 9996 37214 9998 37266
rect 9998 37214 10050 37266
rect 10050 37214 10052 37266
rect 9996 37212 10052 37214
rect 9996 36316 10052 36372
rect 10108 35922 10164 35924
rect 10108 35870 10110 35922
rect 10110 35870 10162 35922
rect 10162 35870 10164 35922
rect 10108 35868 10164 35870
rect 9660 35810 9716 35812
rect 9660 35758 9662 35810
rect 9662 35758 9714 35810
rect 9714 35758 9716 35810
rect 9660 35756 9716 35758
rect 10444 36876 10500 36932
rect 10332 35532 10388 35588
rect 9772 34802 9828 34804
rect 9772 34750 9774 34802
rect 9774 34750 9826 34802
rect 9826 34750 9828 34802
rect 9772 34748 9828 34750
rect 10108 34914 10164 34916
rect 10108 34862 10110 34914
rect 10110 34862 10162 34914
rect 10162 34862 10164 34914
rect 10108 34860 10164 34862
rect 10444 34860 10500 34916
rect 10556 36764 10612 36820
rect 10108 34524 10164 34580
rect 9548 33740 9604 33796
rect 9772 34130 9828 34132
rect 9772 34078 9774 34130
rect 9774 34078 9826 34130
rect 9826 34078 9828 34130
rect 9772 34076 9828 34078
rect 9884 33180 9940 33236
rect 9996 33964 10052 34020
rect 9772 31948 9828 32004
rect 9548 30940 9604 30996
rect 9548 30268 9604 30324
rect 10108 33852 10164 33908
rect 10780 35586 10836 35588
rect 10780 35534 10782 35586
rect 10782 35534 10834 35586
rect 10834 35534 10836 35586
rect 10780 35532 10836 35534
rect 10780 34972 10836 35028
rect 10668 34524 10724 34580
rect 10332 33852 10388 33908
rect 10556 33852 10612 33908
rect 10668 33516 10724 33572
rect 9996 32172 10052 32228
rect 10444 33346 10500 33348
rect 10444 33294 10446 33346
rect 10446 33294 10498 33346
rect 10498 33294 10500 33346
rect 10444 33292 10500 33294
rect 10556 33234 10612 33236
rect 10556 33182 10558 33234
rect 10558 33182 10610 33234
rect 10610 33182 10612 33234
rect 10556 33180 10612 33182
rect 9772 31778 9828 31780
rect 9772 31726 9774 31778
rect 9774 31726 9826 31778
rect 9826 31726 9828 31778
rect 9772 31724 9828 31726
rect 11676 38722 11732 38724
rect 11676 38670 11678 38722
rect 11678 38670 11730 38722
rect 11730 38670 11732 38722
rect 11676 38668 11732 38670
rect 11788 38556 11844 38612
rect 11228 38444 11284 38500
rect 11004 37378 11060 37380
rect 11004 37326 11006 37378
rect 11006 37326 11058 37378
rect 11058 37326 11060 37378
rect 11004 37324 11060 37326
rect 11004 36876 11060 36932
rect 11004 35196 11060 35252
rect 11418 38442 11474 38444
rect 11418 38390 11420 38442
rect 11420 38390 11472 38442
rect 11472 38390 11474 38442
rect 11418 38388 11474 38390
rect 11522 38442 11578 38444
rect 11522 38390 11524 38442
rect 11524 38390 11576 38442
rect 11576 38390 11578 38442
rect 11522 38388 11578 38390
rect 11626 38442 11682 38444
rect 11626 38390 11628 38442
rect 11628 38390 11680 38442
rect 11680 38390 11682 38442
rect 11626 38388 11682 38390
rect 11228 38108 11284 38164
rect 11228 37548 11284 37604
rect 11564 37212 11620 37268
rect 11452 37100 11508 37156
rect 11418 36874 11474 36876
rect 11418 36822 11420 36874
rect 11420 36822 11472 36874
rect 11472 36822 11474 36874
rect 11418 36820 11474 36822
rect 11522 36874 11578 36876
rect 11522 36822 11524 36874
rect 11524 36822 11576 36874
rect 11576 36822 11578 36874
rect 11522 36820 11578 36822
rect 11626 36874 11682 36876
rect 11626 36822 11628 36874
rect 11628 36822 11680 36874
rect 11680 36822 11682 36874
rect 11626 36820 11682 36822
rect 11228 35532 11284 35588
rect 11676 35586 11732 35588
rect 11676 35534 11678 35586
rect 11678 35534 11730 35586
rect 11730 35534 11732 35586
rect 11676 35532 11732 35534
rect 11418 35306 11474 35308
rect 11418 35254 11420 35306
rect 11420 35254 11472 35306
rect 11472 35254 11474 35306
rect 11418 35252 11474 35254
rect 11522 35306 11578 35308
rect 11522 35254 11524 35306
rect 11524 35254 11576 35306
rect 11576 35254 11578 35306
rect 11522 35252 11578 35254
rect 11626 35306 11682 35308
rect 11626 35254 11628 35306
rect 11628 35254 11680 35306
rect 11680 35254 11682 35306
rect 11626 35252 11682 35254
rect 11676 35138 11732 35140
rect 11676 35086 11678 35138
rect 11678 35086 11730 35138
rect 11730 35086 11732 35138
rect 11676 35084 11732 35086
rect 11340 34914 11396 34916
rect 11340 34862 11342 34914
rect 11342 34862 11394 34914
rect 11394 34862 11396 34914
rect 11340 34860 11396 34862
rect 11116 34300 11172 34356
rect 11788 34748 11844 34804
rect 11788 34300 11844 34356
rect 11116 34130 11172 34132
rect 11116 34078 11118 34130
rect 11118 34078 11170 34130
rect 11170 34078 11172 34130
rect 11116 34076 11172 34078
rect 11228 33852 11284 33908
rect 11116 33346 11172 33348
rect 11116 33294 11118 33346
rect 11118 33294 11170 33346
rect 11170 33294 11172 33346
rect 11116 33292 11172 33294
rect 10892 32844 10948 32900
rect 11004 32786 11060 32788
rect 11004 32734 11006 32786
rect 11006 32734 11058 32786
rect 11058 32734 11060 32786
rect 11004 32732 11060 32734
rect 10780 32060 10836 32116
rect 10668 31948 10724 32004
rect 9884 31388 9940 31444
rect 9884 30044 9940 30100
rect 9660 29932 9716 29988
rect 9660 29314 9716 29316
rect 9660 29262 9662 29314
rect 9662 29262 9714 29314
rect 9714 29262 9716 29314
rect 9660 29260 9716 29262
rect 9660 27746 9716 27748
rect 9660 27694 9662 27746
rect 9662 27694 9714 27746
rect 9714 27694 9716 27746
rect 9660 27692 9716 27694
rect 9548 27356 9604 27412
rect 9660 27074 9716 27076
rect 9660 27022 9662 27074
rect 9662 27022 9714 27074
rect 9714 27022 9716 27074
rect 9660 27020 9716 27022
rect 9548 26066 9604 26068
rect 9548 26014 9550 26066
rect 9550 26014 9602 26066
rect 9602 26014 9604 26066
rect 9548 26012 9604 26014
rect 9660 25228 9716 25284
rect 9884 28140 9940 28196
rect 10220 31388 10276 31444
rect 10332 31836 10388 31892
rect 10556 30268 10612 30324
rect 10332 30210 10388 30212
rect 10332 30158 10334 30210
rect 10334 30158 10386 30210
rect 10386 30158 10388 30210
rect 10332 30156 10388 30158
rect 11418 33738 11474 33740
rect 11418 33686 11420 33738
rect 11420 33686 11472 33738
rect 11472 33686 11474 33738
rect 11418 33684 11474 33686
rect 11522 33738 11578 33740
rect 11522 33686 11524 33738
rect 11524 33686 11576 33738
rect 11576 33686 11578 33738
rect 11522 33684 11578 33686
rect 11626 33738 11682 33740
rect 11626 33686 11628 33738
rect 11628 33686 11680 33738
rect 11680 33686 11682 33738
rect 11626 33684 11682 33686
rect 12236 44322 12292 44324
rect 12236 44270 12238 44322
rect 12238 44270 12290 44322
rect 12290 44270 12292 44322
rect 12236 44268 12292 44270
rect 12012 44210 12068 44212
rect 12012 44158 12014 44210
rect 12014 44158 12066 44210
rect 12066 44158 12068 44210
rect 12012 44156 12068 44158
rect 12124 42924 12180 42980
rect 12012 42476 12068 42532
rect 12572 44380 12628 44436
rect 12460 44044 12516 44100
rect 12908 47234 12964 47236
rect 12908 47182 12910 47234
rect 12910 47182 12962 47234
rect 12962 47182 12964 47234
rect 12908 47180 12964 47182
rect 12796 45948 12852 46004
rect 12908 45052 12964 45108
rect 13132 48412 13188 48468
rect 13244 46732 13300 46788
rect 13244 45164 13300 45220
rect 12908 44268 12964 44324
rect 12684 42812 12740 42868
rect 12460 42364 12516 42420
rect 12124 41916 12180 41972
rect 12348 41970 12404 41972
rect 12348 41918 12350 41970
rect 12350 41918 12402 41970
rect 12402 41918 12404 41970
rect 12348 41916 12404 41918
rect 12236 41804 12292 41860
rect 12012 41244 12068 41300
rect 12236 41244 12292 41300
rect 12236 40796 12292 40852
rect 12460 40348 12516 40404
rect 12236 40290 12292 40292
rect 12236 40238 12238 40290
rect 12238 40238 12290 40290
rect 12290 40238 12292 40290
rect 12236 40236 12292 40238
rect 12348 40012 12404 40068
rect 12348 38834 12404 38836
rect 12348 38782 12350 38834
rect 12350 38782 12402 38834
rect 12402 38782 12404 38834
rect 12348 38780 12404 38782
rect 12236 38220 12292 38276
rect 12348 37884 12404 37940
rect 12796 44156 12852 44212
rect 13020 41858 13076 41860
rect 13020 41806 13022 41858
rect 13022 41806 13074 41858
rect 13074 41806 13076 41858
rect 13020 41804 13076 41806
rect 13020 41020 13076 41076
rect 12908 40572 12964 40628
rect 12796 40460 12852 40516
rect 12796 38332 12852 38388
rect 12684 37996 12740 38052
rect 12236 37548 12292 37604
rect 12124 36594 12180 36596
rect 12124 36542 12126 36594
rect 12126 36542 12178 36594
rect 12178 36542 12180 36594
rect 12124 36540 12180 36542
rect 12124 36316 12180 36372
rect 12796 36988 12852 37044
rect 12908 36876 12964 36932
rect 12684 36428 12740 36484
rect 12796 36764 12852 36820
rect 12572 36316 12628 36372
rect 12572 35980 12628 36036
rect 12348 34860 12404 34916
rect 12572 35532 12628 35588
rect 12124 34354 12180 34356
rect 12124 34302 12126 34354
rect 12126 34302 12178 34354
rect 12178 34302 12180 34354
rect 12124 34300 12180 34302
rect 12460 34018 12516 34020
rect 12460 33966 12462 34018
rect 12462 33966 12514 34018
rect 12514 33966 12516 34018
rect 12460 33964 12516 33966
rect 12348 33852 12404 33908
rect 12012 33516 12068 33572
rect 12012 33346 12068 33348
rect 12012 33294 12014 33346
rect 12014 33294 12066 33346
rect 12066 33294 12068 33346
rect 12012 33292 12068 33294
rect 11340 33122 11396 33124
rect 11340 33070 11342 33122
rect 11342 33070 11394 33122
rect 11394 33070 11396 33122
rect 11340 33068 11396 33070
rect 11452 32786 11508 32788
rect 11452 32734 11454 32786
rect 11454 32734 11506 32786
rect 11506 32734 11508 32786
rect 11452 32732 11508 32734
rect 11676 32284 11732 32340
rect 11004 31554 11060 31556
rect 11004 31502 11006 31554
rect 11006 31502 11058 31554
rect 11058 31502 11060 31554
rect 11004 31500 11060 31502
rect 10668 30156 10724 30212
rect 10444 30044 10500 30100
rect 10220 29932 10276 29988
rect 10892 30098 10948 30100
rect 10892 30046 10894 30098
rect 10894 30046 10946 30098
rect 10946 30046 10948 30098
rect 10892 30044 10948 30046
rect 10780 29986 10836 29988
rect 10780 29934 10782 29986
rect 10782 29934 10834 29986
rect 10834 29934 10836 29986
rect 10780 29932 10836 29934
rect 10556 29484 10612 29540
rect 10332 28140 10388 28196
rect 10444 28700 10500 28756
rect 10220 27970 10276 27972
rect 10220 27918 10222 27970
rect 10222 27918 10274 27970
rect 10274 27918 10276 27970
rect 10220 27916 10276 27918
rect 11418 32170 11474 32172
rect 11228 32060 11284 32116
rect 11418 32118 11420 32170
rect 11420 32118 11472 32170
rect 11472 32118 11474 32170
rect 11418 32116 11474 32118
rect 11522 32170 11578 32172
rect 11522 32118 11524 32170
rect 11524 32118 11576 32170
rect 11576 32118 11578 32170
rect 11522 32116 11578 32118
rect 11626 32170 11682 32172
rect 11626 32118 11628 32170
rect 11628 32118 11680 32170
rect 11680 32118 11682 32170
rect 11626 32116 11682 32118
rect 11564 31778 11620 31780
rect 11564 31726 11566 31778
rect 11566 31726 11618 31778
rect 11618 31726 11620 31778
rect 11564 31724 11620 31726
rect 11340 31500 11396 31556
rect 11418 30602 11474 30604
rect 11418 30550 11420 30602
rect 11420 30550 11472 30602
rect 11472 30550 11474 30602
rect 11418 30548 11474 30550
rect 11522 30602 11578 30604
rect 11522 30550 11524 30602
rect 11524 30550 11576 30602
rect 11576 30550 11578 30602
rect 11522 30548 11578 30550
rect 11626 30602 11682 30604
rect 11626 30550 11628 30602
rect 11628 30550 11680 30602
rect 11680 30550 11682 30602
rect 11626 30548 11682 30550
rect 11452 30322 11508 30324
rect 11452 30270 11454 30322
rect 11454 30270 11506 30322
rect 11506 30270 11508 30322
rect 11452 30268 11508 30270
rect 10892 29426 10948 29428
rect 10892 29374 10894 29426
rect 10894 29374 10946 29426
rect 10946 29374 10948 29426
rect 10892 29372 10948 29374
rect 12908 35756 12964 35812
rect 12684 34972 12740 35028
rect 12796 33852 12852 33908
rect 12012 32844 12068 32900
rect 12348 32956 12404 33012
rect 12684 33180 12740 33236
rect 12796 32844 12852 32900
rect 12124 32060 12180 32116
rect 12124 31612 12180 31668
rect 12572 31666 12628 31668
rect 12572 31614 12574 31666
rect 12574 31614 12626 31666
rect 12626 31614 12628 31666
rect 12572 31612 12628 31614
rect 12908 32060 12964 32116
rect 12012 30210 12068 30212
rect 12012 30158 12014 30210
rect 12014 30158 12066 30210
rect 12066 30158 12068 30210
rect 12012 30156 12068 30158
rect 11900 30044 11956 30100
rect 12908 30940 12964 30996
rect 12572 30322 12628 30324
rect 12572 30270 12574 30322
rect 12574 30270 12626 30322
rect 12626 30270 12628 30322
rect 12572 30268 12628 30270
rect 12796 30156 12852 30212
rect 12684 29932 12740 29988
rect 12348 29650 12404 29652
rect 12348 29598 12350 29650
rect 12350 29598 12402 29650
rect 12402 29598 12404 29650
rect 12348 29596 12404 29598
rect 11116 29148 11172 29204
rect 12012 29148 12068 29204
rect 11418 29034 11474 29036
rect 11418 28982 11420 29034
rect 11420 28982 11472 29034
rect 11472 28982 11474 29034
rect 11418 28980 11474 28982
rect 11522 29034 11578 29036
rect 11522 28982 11524 29034
rect 11524 28982 11576 29034
rect 11576 28982 11578 29034
rect 11522 28980 11578 28982
rect 11626 29034 11682 29036
rect 11626 28982 11628 29034
rect 11628 28982 11680 29034
rect 11680 28982 11682 29034
rect 11626 28980 11682 28982
rect 11116 28700 11172 28756
rect 10780 28140 10836 28196
rect 10780 27970 10836 27972
rect 10780 27918 10782 27970
rect 10782 27918 10834 27970
rect 10834 27918 10836 27970
rect 10780 27916 10836 27918
rect 11788 28700 11844 28756
rect 12460 28812 12516 28868
rect 11564 28082 11620 28084
rect 11564 28030 11566 28082
rect 11566 28030 11618 28082
rect 11618 28030 11620 28082
rect 11564 28028 11620 28030
rect 11004 27580 11060 27636
rect 10556 27356 10612 27412
rect 9772 24668 9828 24724
rect 9772 24332 9828 24388
rect 8876 22540 8932 22596
rect 8876 20188 8932 20244
rect 9100 20972 9156 21028
rect 9100 19852 9156 19908
rect 7756 19234 7812 19236
rect 7756 19182 7758 19234
rect 7758 19182 7810 19234
rect 7810 19182 7812 19234
rect 7756 19180 7812 19182
rect 6972 18956 7028 19012
rect 7644 19010 7700 19012
rect 7644 18958 7646 19010
rect 7646 18958 7698 19010
rect 7698 18958 7700 19010
rect 7644 18956 7700 18958
rect 8540 19180 8596 19236
rect 8016 18842 8072 18844
rect 8016 18790 8018 18842
rect 8018 18790 8070 18842
rect 8070 18790 8072 18842
rect 8016 18788 8072 18790
rect 8120 18842 8176 18844
rect 8120 18790 8122 18842
rect 8122 18790 8174 18842
rect 8174 18790 8176 18842
rect 8120 18788 8176 18790
rect 8224 18842 8280 18844
rect 8224 18790 8226 18842
rect 8226 18790 8278 18842
rect 8278 18790 8280 18842
rect 8224 18788 8280 18790
rect 7532 18396 7588 18452
rect 7420 17052 7476 17108
rect 7868 18060 7924 18116
rect 7196 16940 7252 16996
rect 6860 15148 6916 15204
rect 7084 15372 7140 15428
rect 7420 15426 7476 15428
rect 7420 15374 7422 15426
rect 7422 15374 7474 15426
rect 7474 15374 7476 15426
rect 7420 15372 7476 15374
rect 7420 15148 7476 15204
rect 6972 13356 7028 13412
rect 7308 14418 7364 14420
rect 7308 14366 7310 14418
rect 7310 14366 7362 14418
rect 7362 14366 7364 14418
rect 7308 14364 7364 14366
rect 7084 12850 7140 12852
rect 7084 12798 7086 12850
rect 7086 12798 7138 12850
rect 7138 12798 7140 12850
rect 7084 12796 7140 12798
rect 7420 12738 7476 12740
rect 7420 12686 7422 12738
rect 7422 12686 7474 12738
rect 7474 12686 7476 12738
rect 7420 12684 7476 12686
rect 7308 12066 7364 12068
rect 7308 12014 7310 12066
rect 7310 12014 7362 12066
rect 7362 12014 7364 12066
rect 7308 12012 7364 12014
rect 6076 11340 6132 11396
rect 6748 11452 6804 11508
rect 8540 18450 8596 18452
rect 8540 18398 8542 18450
rect 8542 18398 8594 18450
rect 8594 18398 8596 18450
rect 8540 18396 8596 18398
rect 8540 18060 8596 18116
rect 9100 18284 9156 18340
rect 8988 17778 9044 17780
rect 8988 17726 8990 17778
rect 8990 17726 9042 17778
rect 9042 17726 9044 17778
rect 8988 17724 9044 17726
rect 8428 17388 8484 17444
rect 8016 17274 8072 17276
rect 8016 17222 8018 17274
rect 8018 17222 8070 17274
rect 8070 17222 8072 17274
rect 8016 17220 8072 17222
rect 8120 17274 8176 17276
rect 8120 17222 8122 17274
rect 8122 17222 8174 17274
rect 8174 17222 8176 17274
rect 8120 17220 8176 17222
rect 8224 17274 8280 17276
rect 8224 17222 8226 17274
rect 8226 17222 8278 17274
rect 8278 17222 8280 17274
rect 8224 17220 8280 17222
rect 8204 17052 8260 17108
rect 7756 16994 7812 16996
rect 7756 16942 7758 16994
rect 7758 16942 7810 16994
rect 7810 16942 7812 16994
rect 7756 16940 7812 16942
rect 9212 18060 9268 18116
rect 9324 23436 9380 23492
rect 8016 15706 8072 15708
rect 8016 15654 8018 15706
rect 8018 15654 8070 15706
rect 8070 15654 8072 15706
rect 8016 15652 8072 15654
rect 8120 15706 8176 15708
rect 8120 15654 8122 15706
rect 8122 15654 8174 15706
rect 8174 15654 8176 15706
rect 8120 15652 8176 15654
rect 8224 15706 8280 15708
rect 8224 15654 8226 15706
rect 8226 15654 8278 15706
rect 8278 15654 8280 15706
rect 8224 15652 8280 15654
rect 7756 15538 7812 15540
rect 7756 15486 7758 15538
rect 7758 15486 7810 15538
rect 7810 15486 7812 15538
rect 7756 15484 7812 15486
rect 8540 15484 8596 15540
rect 7868 15260 7924 15316
rect 7980 15148 8036 15204
rect 9436 20860 9492 20916
rect 9436 20690 9492 20692
rect 9436 20638 9438 20690
rect 9438 20638 9490 20690
rect 9490 20638 9492 20690
rect 9436 20636 9492 20638
rect 9436 17442 9492 17444
rect 9436 17390 9438 17442
rect 9438 17390 9490 17442
rect 9490 17390 9492 17442
rect 9436 17388 9492 17390
rect 9660 22540 9716 22596
rect 10108 24108 10164 24164
rect 10332 26012 10388 26068
rect 10444 25282 10500 25284
rect 10444 25230 10446 25282
rect 10446 25230 10498 25282
rect 10498 25230 10500 25282
rect 10444 25228 10500 25230
rect 10444 24332 10500 24388
rect 10108 22540 10164 22596
rect 9660 21756 9716 21812
rect 9884 21644 9940 21700
rect 10220 20860 10276 20916
rect 9772 20802 9828 20804
rect 9772 20750 9774 20802
rect 9774 20750 9826 20802
rect 9826 20750 9828 20802
rect 9772 20748 9828 20750
rect 9772 20524 9828 20580
rect 9660 18396 9716 18452
rect 10444 21420 10500 21476
rect 10780 26290 10836 26292
rect 10780 26238 10782 26290
rect 10782 26238 10834 26290
rect 10834 26238 10836 26290
rect 10780 26236 10836 26238
rect 10780 25900 10836 25956
rect 10780 24108 10836 24164
rect 10668 23826 10724 23828
rect 10668 23774 10670 23826
rect 10670 23774 10722 23826
rect 10722 23774 10724 23826
rect 10668 23772 10724 23774
rect 11340 27580 11396 27636
rect 11418 27466 11474 27468
rect 11418 27414 11420 27466
rect 11420 27414 11472 27466
rect 11472 27414 11474 27466
rect 11418 27412 11474 27414
rect 11522 27466 11578 27468
rect 11522 27414 11524 27466
rect 11524 27414 11576 27466
rect 11576 27414 11578 27466
rect 11522 27412 11578 27414
rect 11626 27466 11682 27468
rect 11626 27414 11628 27466
rect 11628 27414 11680 27466
rect 11680 27414 11682 27466
rect 11626 27412 11682 27414
rect 10556 21084 10612 21140
rect 11116 26236 11172 26292
rect 10780 20972 10836 21028
rect 10556 20690 10612 20692
rect 10556 20638 10558 20690
rect 10558 20638 10610 20690
rect 10610 20638 10612 20690
rect 10556 20636 10612 20638
rect 9996 20188 10052 20244
rect 10668 20578 10724 20580
rect 10668 20526 10670 20578
rect 10670 20526 10722 20578
rect 10722 20526 10724 20578
rect 10668 20524 10724 20526
rect 10556 20188 10612 20244
rect 10108 18508 10164 18564
rect 10332 18284 10388 18340
rect 10220 17388 10276 17444
rect 9772 16268 9828 16324
rect 8540 14364 8596 14420
rect 8016 14138 8072 14140
rect 8016 14086 8018 14138
rect 8018 14086 8070 14138
rect 8070 14086 8072 14138
rect 8016 14084 8072 14086
rect 8120 14138 8176 14140
rect 8120 14086 8122 14138
rect 8122 14086 8174 14138
rect 8174 14086 8176 14138
rect 8120 14084 8176 14086
rect 8224 14138 8280 14140
rect 8224 14086 8226 14138
rect 8226 14086 8278 14138
rect 8278 14086 8280 14138
rect 8224 14084 8280 14086
rect 8316 13804 8372 13860
rect 8092 13746 8148 13748
rect 8092 13694 8094 13746
rect 8094 13694 8146 13746
rect 8146 13694 8148 13746
rect 8092 13692 8148 13694
rect 7644 13356 7700 13412
rect 8652 13356 8708 13412
rect 8764 14588 8820 14644
rect 9884 14700 9940 14756
rect 10444 17836 10500 17892
rect 10332 17106 10388 17108
rect 10332 17054 10334 17106
rect 10334 17054 10386 17106
rect 10386 17054 10388 17106
rect 10332 17052 10388 17054
rect 10220 16828 10276 16884
rect 8092 13074 8148 13076
rect 8092 13022 8094 13074
rect 8094 13022 8146 13074
rect 8146 13022 8148 13074
rect 8092 13020 8148 13022
rect 8540 12738 8596 12740
rect 8540 12686 8542 12738
rect 8542 12686 8594 12738
rect 8594 12686 8596 12738
rect 8540 12684 8596 12686
rect 8016 12570 8072 12572
rect 8016 12518 8018 12570
rect 8018 12518 8070 12570
rect 8070 12518 8072 12570
rect 8016 12516 8072 12518
rect 8120 12570 8176 12572
rect 8120 12518 8122 12570
rect 8122 12518 8174 12570
rect 8174 12518 8176 12570
rect 8120 12516 8176 12518
rect 8224 12570 8280 12572
rect 8224 12518 8226 12570
rect 8226 12518 8278 12570
rect 8278 12518 8280 12570
rect 8224 12516 8280 12518
rect 9884 13916 9940 13972
rect 10220 16044 10276 16100
rect 9996 13580 10052 13636
rect 10780 19964 10836 20020
rect 10780 18508 10836 18564
rect 11004 22540 11060 22596
rect 11004 21026 11060 21028
rect 11004 20974 11006 21026
rect 11006 20974 11058 21026
rect 11058 20974 11060 21026
rect 11004 20972 11060 20974
rect 11418 25898 11474 25900
rect 11418 25846 11420 25898
rect 11420 25846 11472 25898
rect 11472 25846 11474 25898
rect 11418 25844 11474 25846
rect 11522 25898 11578 25900
rect 11522 25846 11524 25898
rect 11524 25846 11576 25898
rect 11576 25846 11578 25898
rect 11522 25844 11578 25846
rect 11626 25898 11682 25900
rect 11626 25846 11628 25898
rect 11628 25846 11680 25898
rect 11680 25846 11682 25898
rect 11626 25844 11682 25846
rect 12572 28140 12628 28196
rect 12460 28028 12516 28084
rect 12348 27580 12404 27636
rect 12908 29986 12964 29988
rect 12908 29934 12910 29986
rect 12910 29934 12962 29986
rect 12962 29934 12964 29986
rect 12908 29932 12964 29934
rect 12908 28754 12964 28756
rect 12908 28702 12910 28754
rect 12910 28702 12962 28754
rect 12962 28702 12964 28754
rect 12908 28700 12964 28702
rect 12796 27468 12852 27524
rect 12908 27020 12964 27076
rect 11788 24892 11844 24948
rect 11900 25228 11956 25284
rect 11418 24330 11474 24332
rect 11418 24278 11420 24330
rect 11420 24278 11472 24330
rect 11472 24278 11474 24330
rect 11418 24276 11474 24278
rect 11522 24330 11578 24332
rect 11522 24278 11524 24330
rect 11524 24278 11576 24330
rect 11576 24278 11578 24330
rect 11522 24276 11578 24278
rect 11626 24330 11682 24332
rect 11626 24278 11628 24330
rect 11628 24278 11680 24330
rect 11680 24278 11682 24330
rect 11626 24276 11682 24278
rect 11564 23996 11620 24052
rect 11228 23938 11284 23940
rect 11228 23886 11230 23938
rect 11230 23886 11282 23938
rect 11282 23886 11284 23938
rect 11228 23884 11284 23886
rect 12012 23884 12068 23940
rect 11676 23826 11732 23828
rect 11676 23774 11678 23826
rect 11678 23774 11730 23826
rect 11730 23774 11732 23826
rect 11676 23772 11732 23774
rect 11564 23660 11620 23716
rect 12124 26178 12180 26180
rect 12124 26126 12126 26178
rect 12126 26126 12178 26178
rect 12178 26126 12180 26178
rect 12124 26124 12180 26126
rect 11418 22762 11474 22764
rect 11418 22710 11420 22762
rect 11420 22710 11472 22762
rect 11472 22710 11474 22762
rect 11418 22708 11474 22710
rect 11522 22762 11578 22764
rect 11522 22710 11524 22762
rect 11524 22710 11576 22762
rect 11576 22710 11578 22762
rect 11522 22708 11578 22710
rect 11626 22762 11682 22764
rect 11626 22710 11628 22762
rect 11628 22710 11680 22762
rect 11680 22710 11682 22762
rect 11626 22708 11682 22710
rect 11788 22316 11844 22372
rect 11900 22876 11956 22932
rect 11418 21194 11474 21196
rect 11418 21142 11420 21194
rect 11420 21142 11472 21194
rect 11472 21142 11474 21194
rect 11418 21140 11474 21142
rect 11522 21194 11578 21196
rect 11522 21142 11524 21194
rect 11524 21142 11576 21194
rect 11576 21142 11578 21194
rect 11522 21140 11578 21142
rect 11626 21194 11682 21196
rect 11626 21142 11628 21194
rect 11628 21142 11680 21194
rect 11680 21142 11682 21194
rect 11626 21140 11682 21142
rect 11676 21026 11732 21028
rect 11676 20974 11678 21026
rect 11678 20974 11730 21026
rect 11730 20974 11732 21026
rect 11676 20972 11732 20974
rect 11340 20860 11396 20916
rect 11788 20748 11844 20804
rect 11452 20242 11508 20244
rect 11452 20190 11454 20242
rect 11454 20190 11506 20242
rect 11506 20190 11508 20242
rect 11452 20188 11508 20190
rect 12012 22540 12068 22596
rect 11418 19626 11474 19628
rect 11418 19574 11420 19626
rect 11420 19574 11472 19626
rect 11472 19574 11474 19626
rect 11418 19572 11474 19574
rect 11522 19626 11578 19628
rect 11522 19574 11524 19626
rect 11524 19574 11576 19626
rect 11576 19574 11578 19626
rect 11522 19572 11578 19574
rect 11626 19626 11682 19628
rect 11626 19574 11628 19626
rect 11628 19574 11680 19626
rect 11680 19574 11682 19626
rect 11626 19572 11682 19574
rect 11564 18450 11620 18452
rect 11564 18398 11566 18450
rect 11566 18398 11618 18450
rect 11618 18398 11620 18450
rect 11564 18396 11620 18398
rect 11418 18058 11474 18060
rect 11418 18006 11420 18058
rect 11420 18006 11472 18058
rect 11472 18006 11474 18058
rect 11418 18004 11474 18006
rect 11522 18058 11578 18060
rect 11522 18006 11524 18058
rect 11524 18006 11576 18058
rect 11576 18006 11578 18058
rect 11522 18004 11578 18006
rect 11626 18058 11682 18060
rect 11626 18006 11628 18058
rect 11628 18006 11680 18058
rect 11680 18006 11682 18058
rect 11626 18004 11682 18006
rect 11228 17836 11284 17892
rect 11676 17666 11732 17668
rect 11676 17614 11678 17666
rect 11678 17614 11730 17666
rect 11730 17614 11732 17666
rect 11676 17612 11732 17614
rect 10780 16882 10836 16884
rect 10780 16830 10782 16882
rect 10782 16830 10834 16882
rect 10834 16830 10836 16882
rect 10780 16828 10836 16830
rect 11116 15820 11172 15876
rect 10444 13804 10500 13860
rect 9772 13468 9828 13524
rect 9548 13356 9604 13412
rect 9324 12738 9380 12740
rect 9324 12686 9326 12738
rect 9326 12686 9378 12738
rect 9378 12686 9380 12738
rect 9324 12684 9380 12686
rect 9884 13356 9940 13412
rect 7868 11506 7924 11508
rect 7868 11454 7870 11506
rect 7870 11454 7922 11506
rect 7922 11454 7924 11506
rect 7868 11452 7924 11454
rect 6300 11282 6356 11284
rect 6300 11230 6302 11282
rect 6302 11230 6354 11282
rect 6354 11230 6356 11282
rect 6300 11228 6356 11230
rect 6300 10332 6356 10388
rect 4614 8650 4670 8652
rect 4614 8598 4616 8650
rect 4616 8598 4668 8650
rect 4668 8598 4670 8650
rect 4614 8596 4670 8598
rect 4718 8650 4774 8652
rect 4718 8598 4720 8650
rect 4720 8598 4772 8650
rect 4772 8598 4774 8650
rect 4718 8596 4774 8598
rect 4822 8650 4878 8652
rect 4822 8598 4824 8650
rect 4824 8598 4876 8650
rect 4876 8598 4878 8650
rect 4822 8596 4878 8598
rect 4732 8316 4788 8372
rect 5068 7980 5124 8036
rect 5516 8428 5572 8484
rect 5180 7868 5236 7924
rect 5404 7980 5460 8036
rect 5068 7698 5124 7700
rect 5068 7646 5070 7698
rect 5070 7646 5122 7698
rect 5122 7646 5124 7698
rect 5068 7644 5124 7646
rect 4614 7082 4670 7084
rect 4614 7030 4616 7082
rect 4616 7030 4668 7082
rect 4668 7030 4670 7082
rect 4614 7028 4670 7030
rect 4718 7082 4774 7084
rect 4718 7030 4720 7082
rect 4720 7030 4772 7082
rect 4772 7030 4774 7082
rect 4718 7028 4774 7030
rect 4822 7082 4878 7084
rect 4822 7030 4824 7082
rect 4824 7030 4876 7082
rect 4876 7030 4878 7082
rect 4822 7028 4878 7030
rect 4732 6690 4788 6692
rect 4732 6638 4734 6690
rect 4734 6638 4786 6690
rect 4786 6638 4788 6690
rect 4732 6636 4788 6638
rect 6076 7868 6132 7924
rect 5516 7586 5572 7588
rect 5516 7534 5518 7586
rect 5518 7534 5570 7586
rect 5570 7534 5572 7586
rect 5516 7532 5572 7534
rect 6636 11116 6692 11172
rect 6748 10556 6804 10612
rect 9548 12236 9604 12292
rect 10108 12850 10164 12852
rect 10108 12798 10110 12850
rect 10110 12798 10162 12850
rect 10162 12798 10164 12850
rect 10108 12796 10164 12798
rect 11676 17106 11732 17108
rect 11676 17054 11678 17106
rect 11678 17054 11730 17106
rect 11730 17054 11732 17106
rect 11676 17052 11732 17054
rect 11418 16490 11474 16492
rect 11418 16438 11420 16490
rect 11420 16438 11472 16490
rect 11472 16438 11474 16490
rect 11418 16436 11474 16438
rect 11522 16490 11578 16492
rect 11522 16438 11524 16490
rect 11524 16438 11576 16490
rect 11576 16438 11578 16490
rect 11522 16436 11578 16438
rect 11626 16490 11682 16492
rect 11626 16438 11628 16490
rect 11628 16438 11680 16490
rect 11680 16438 11682 16490
rect 11626 16436 11682 16438
rect 11228 15708 11284 15764
rect 11418 14922 11474 14924
rect 11418 14870 11420 14922
rect 11420 14870 11472 14922
rect 11472 14870 11474 14922
rect 11418 14868 11474 14870
rect 11522 14922 11578 14924
rect 11522 14870 11524 14922
rect 11524 14870 11576 14922
rect 11576 14870 11578 14922
rect 11522 14868 11578 14870
rect 11626 14922 11682 14924
rect 11626 14870 11628 14922
rect 11628 14870 11680 14922
rect 11680 14870 11682 14922
rect 11626 14868 11682 14870
rect 11564 13970 11620 13972
rect 11564 13918 11566 13970
rect 11566 13918 11618 13970
rect 11618 13918 11620 13970
rect 11564 13916 11620 13918
rect 10780 13746 10836 13748
rect 10780 13694 10782 13746
rect 10782 13694 10834 13746
rect 10834 13694 10836 13746
rect 10780 13692 10836 13694
rect 10332 13020 10388 13076
rect 9884 12738 9940 12740
rect 9884 12686 9886 12738
rect 9886 12686 9938 12738
rect 9938 12686 9940 12738
rect 9884 12684 9940 12686
rect 8988 12178 9044 12180
rect 8988 12126 8990 12178
rect 8990 12126 9042 12178
rect 9042 12126 9044 12178
rect 8988 12124 9044 12126
rect 8540 12066 8596 12068
rect 8540 12014 8542 12066
rect 8542 12014 8594 12066
rect 8594 12014 8596 12066
rect 8540 12012 8596 12014
rect 7756 10722 7812 10724
rect 7756 10670 7758 10722
rect 7758 10670 7810 10722
rect 7810 10670 7812 10722
rect 7756 10668 7812 10670
rect 6636 9884 6692 9940
rect 7644 10386 7700 10388
rect 7644 10334 7646 10386
rect 7646 10334 7698 10386
rect 7698 10334 7700 10386
rect 7644 10332 7700 10334
rect 8016 11002 8072 11004
rect 8016 10950 8018 11002
rect 8018 10950 8070 11002
rect 8070 10950 8072 11002
rect 8016 10948 8072 10950
rect 8120 11002 8176 11004
rect 8120 10950 8122 11002
rect 8122 10950 8174 11002
rect 8174 10950 8176 11002
rect 8120 10948 8176 10950
rect 8224 11002 8280 11004
rect 8224 10950 8226 11002
rect 8226 10950 8278 11002
rect 8278 10950 8280 11002
rect 8224 10948 8280 10950
rect 9772 12178 9828 12180
rect 9772 12126 9774 12178
rect 9774 12126 9826 12178
rect 9826 12126 9828 12178
rect 9772 12124 9828 12126
rect 8764 11564 8820 11620
rect 10556 12290 10612 12292
rect 10556 12238 10558 12290
rect 10558 12238 10610 12290
rect 10610 12238 10612 12290
rect 10556 12236 10612 12238
rect 9884 11452 9940 11508
rect 10108 11452 10164 11508
rect 8764 10668 8820 10724
rect 8092 10610 8148 10612
rect 8092 10558 8094 10610
rect 8094 10558 8146 10610
rect 8146 10558 8148 10610
rect 8092 10556 8148 10558
rect 9212 11228 9268 11284
rect 8016 9434 8072 9436
rect 8016 9382 8018 9434
rect 8018 9382 8070 9434
rect 8070 9382 8072 9434
rect 8016 9380 8072 9382
rect 8120 9434 8176 9436
rect 8120 9382 8122 9434
rect 8122 9382 8174 9434
rect 8174 9382 8176 9434
rect 8120 9380 8176 9382
rect 8224 9434 8280 9436
rect 8224 9382 8226 9434
rect 8226 9382 8278 9434
rect 8278 9382 8280 9434
rect 8224 9380 8280 9382
rect 10668 11228 10724 11284
rect 10108 11116 10164 11172
rect 10444 11004 10500 11060
rect 9884 10834 9940 10836
rect 9884 10782 9886 10834
rect 9886 10782 9938 10834
rect 9938 10782 9940 10834
rect 9884 10780 9940 10782
rect 10892 13468 10948 13524
rect 11418 13354 11474 13356
rect 11418 13302 11420 13354
rect 11420 13302 11472 13354
rect 11472 13302 11474 13354
rect 11418 13300 11474 13302
rect 11522 13354 11578 13356
rect 11522 13302 11524 13354
rect 11524 13302 11576 13354
rect 11576 13302 11578 13354
rect 11522 13300 11578 13302
rect 11626 13354 11682 13356
rect 11626 13302 11628 13354
rect 11628 13302 11680 13354
rect 11680 13302 11682 13354
rect 11626 13300 11682 13302
rect 11340 13074 11396 13076
rect 11340 13022 11342 13074
rect 11342 13022 11394 13074
rect 11394 13022 11396 13074
rect 11340 13020 11396 13022
rect 13244 41132 13300 41188
rect 13468 50652 13524 50708
rect 13580 51100 13636 51156
rect 13580 50594 13636 50596
rect 13580 50542 13582 50594
rect 13582 50542 13634 50594
rect 13634 50542 13636 50594
rect 13580 50540 13636 50542
rect 13468 50204 13524 50260
rect 13916 50988 13972 51044
rect 14140 54348 14196 54404
rect 14140 52274 14196 52276
rect 14140 52222 14142 52274
rect 14142 52222 14194 52274
rect 14194 52222 14196 52274
rect 14140 52220 14196 52222
rect 13468 49420 13524 49476
rect 13468 45276 13524 45332
rect 13468 45106 13524 45108
rect 13468 45054 13470 45106
rect 13470 45054 13522 45106
rect 13522 45054 13524 45106
rect 13468 45052 13524 45054
rect 13468 44604 13524 44660
rect 14476 55244 14532 55300
rect 14364 55020 14420 55076
rect 14364 53506 14420 53508
rect 14364 53454 14366 53506
rect 14366 53454 14418 53506
rect 14418 53454 14420 53506
rect 14364 53452 14420 53454
rect 14028 49868 14084 49924
rect 14140 49420 14196 49476
rect 14252 50540 14308 50596
rect 13916 49026 13972 49028
rect 13916 48974 13918 49026
rect 13918 48974 13970 49026
rect 13970 48974 13972 49026
rect 13916 48972 13972 48974
rect 13804 48860 13860 48916
rect 13804 47964 13860 48020
rect 15820 58940 15876 58996
rect 15932 58716 15988 58772
rect 15484 56082 15540 56084
rect 15484 56030 15486 56082
rect 15486 56030 15538 56082
rect 15538 56030 15540 56082
rect 15484 56028 15540 56030
rect 15932 56812 15988 56868
rect 15372 55132 15428 55188
rect 14820 54906 14876 54908
rect 14820 54854 14822 54906
rect 14822 54854 14874 54906
rect 14874 54854 14876 54906
rect 14820 54852 14876 54854
rect 14924 54906 14980 54908
rect 14924 54854 14926 54906
rect 14926 54854 14978 54906
rect 14978 54854 14980 54906
rect 14924 54852 14980 54854
rect 15028 54906 15084 54908
rect 15028 54854 15030 54906
rect 15030 54854 15082 54906
rect 15082 54854 15084 54906
rect 15028 54852 15084 54854
rect 15932 55244 15988 55300
rect 14924 53676 14980 53732
rect 14700 53452 14756 53508
rect 15036 53564 15092 53620
rect 14924 53452 14980 53508
rect 14820 53338 14876 53340
rect 14820 53286 14822 53338
rect 14822 53286 14874 53338
rect 14874 53286 14876 53338
rect 14820 53284 14876 53286
rect 14924 53338 14980 53340
rect 14924 53286 14926 53338
rect 14926 53286 14978 53338
rect 14978 53286 14980 53338
rect 14924 53284 14980 53286
rect 15028 53338 15084 53340
rect 15028 53286 15030 53338
rect 15030 53286 15082 53338
rect 15082 53286 15084 53338
rect 15028 53284 15084 53286
rect 15036 53004 15092 53060
rect 14812 52556 14868 52612
rect 15260 53004 15316 53060
rect 15372 53564 15428 53620
rect 14140 49026 14196 49028
rect 14140 48974 14142 49026
rect 14142 48974 14194 49026
rect 14194 48974 14196 49026
rect 14140 48972 14196 48974
rect 14028 48748 14084 48804
rect 14140 48354 14196 48356
rect 14140 48302 14142 48354
rect 14142 48302 14194 48354
rect 14194 48302 14196 48354
rect 14140 48300 14196 48302
rect 14140 48076 14196 48132
rect 14140 47458 14196 47460
rect 14140 47406 14142 47458
rect 14142 47406 14194 47458
rect 14194 47406 14196 47458
rect 14140 47404 14196 47406
rect 14028 47068 14084 47124
rect 13804 45836 13860 45892
rect 14364 48636 14420 48692
rect 14476 48860 14532 48916
rect 14364 47346 14420 47348
rect 14364 47294 14366 47346
rect 14366 47294 14418 47346
rect 14418 47294 14420 47346
rect 14364 47292 14420 47294
rect 14364 47068 14420 47124
rect 13692 45276 13748 45332
rect 13692 44940 13748 44996
rect 13580 44492 13636 44548
rect 13692 44380 13748 44436
rect 13468 44156 13524 44212
rect 13692 43932 13748 43988
rect 15372 52892 15428 52948
rect 15148 52108 15204 52164
rect 14820 51770 14876 51772
rect 14820 51718 14822 51770
rect 14822 51718 14874 51770
rect 14874 51718 14876 51770
rect 14820 51716 14876 51718
rect 14924 51770 14980 51772
rect 14924 51718 14926 51770
rect 14926 51718 14978 51770
rect 14978 51718 14980 51770
rect 14924 51716 14980 51718
rect 15028 51770 15084 51772
rect 15028 51718 15030 51770
rect 15030 51718 15082 51770
rect 15082 51718 15084 51770
rect 15028 51716 15084 51718
rect 14812 50764 14868 50820
rect 15148 50764 15204 50820
rect 15036 50482 15092 50484
rect 15036 50430 15038 50482
rect 15038 50430 15090 50482
rect 15090 50430 15092 50482
rect 15036 50428 15092 50430
rect 14820 50202 14876 50204
rect 14820 50150 14822 50202
rect 14822 50150 14874 50202
rect 14874 50150 14876 50202
rect 14820 50148 14876 50150
rect 14924 50202 14980 50204
rect 14924 50150 14926 50202
rect 14926 50150 14978 50202
rect 14978 50150 14980 50202
rect 14924 50148 14980 50150
rect 15028 50202 15084 50204
rect 15028 50150 15030 50202
rect 15030 50150 15082 50202
rect 15082 50150 15084 50202
rect 15028 50148 15084 50150
rect 15260 50092 15316 50148
rect 15372 50988 15428 51044
rect 15596 53228 15652 53284
rect 15708 53058 15764 53060
rect 15708 53006 15710 53058
rect 15710 53006 15762 53058
rect 15762 53006 15764 53058
rect 15708 53004 15764 53006
rect 15932 53004 15988 53060
rect 15596 51324 15652 51380
rect 15932 50764 15988 50820
rect 15932 50092 15988 50148
rect 15596 49980 15652 50036
rect 15484 49532 15540 49588
rect 15372 49138 15428 49140
rect 15372 49086 15374 49138
rect 15374 49086 15426 49138
rect 15426 49086 15428 49138
rect 15372 49084 15428 49086
rect 15148 48972 15204 49028
rect 14820 48634 14876 48636
rect 14820 48582 14822 48634
rect 14822 48582 14874 48634
rect 14874 48582 14876 48634
rect 14820 48580 14876 48582
rect 14924 48634 14980 48636
rect 14924 48582 14926 48634
rect 14926 48582 14978 48634
rect 14978 48582 14980 48634
rect 14924 48580 14980 48582
rect 15028 48634 15084 48636
rect 15028 48582 15030 48634
rect 15030 48582 15082 48634
rect 15082 48582 15084 48634
rect 15028 48580 15084 48582
rect 15036 48412 15092 48468
rect 15148 48188 15204 48244
rect 14700 47964 14756 48020
rect 14700 47180 14756 47236
rect 14820 47066 14876 47068
rect 14820 47014 14822 47066
rect 14822 47014 14874 47066
rect 14874 47014 14876 47066
rect 14820 47012 14876 47014
rect 14924 47066 14980 47068
rect 14924 47014 14926 47066
rect 14926 47014 14978 47066
rect 14978 47014 14980 47066
rect 14924 47012 14980 47014
rect 15028 47066 15084 47068
rect 15028 47014 15030 47066
rect 15030 47014 15082 47066
rect 15082 47014 15084 47066
rect 15028 47012 15084 47014
rect 15036 46732 15092 46788
rect 15260 47628 15316 47684
rect 14700 45836 14756 45892
rect 14700 45666 14756 45668
rect 14700 45614 14702 45666
rect 14702 45614 14754 45666
rect 14754 45614 14756 45666
rect 14700 45612 14756 45614
rect 14820 45498 14876 45500
rect 14820 45446 14822 45498
rect 14822 45446 14874 45498
rect 14874 45446 14876 45498
rect 14820 45444 14876 45446
rect 14924 45498 14980 45500
rect 14924 45446 14926 45498
rect 14926 45446 14978 45498
rect 14978 45446 14980 45498
rect 14924 45444 14980 45446
rect 15028 45498 15084 45500
rect 15028 45446 15030 45498
rect 15030 45446 15082 45498
rect 15082 45446 15084 45498
rect 15028 45444 15084 45446
rect 14588 45276 14644 45332
rect 14924 45276 14980 45332
rect 14812 44716 14868 44772
rect 14588 44492 14644 44548
rect 13916 44380 13972 44436
rect 13916 44098 13972 44100
rect 13916 44046 13918 44098
rect 13918 44046 13970 44098
rect 13970 44046 13972 44098
rect 13916 44044 13972 44046
rect 13804 43372 13860 43428
rect 13916 43708 13972 43764
rect 13804 42812 13860 42868
rect 13580 41804 13636 41860
rect 13468 40572 13524 40628
rect 15484 46620 15540 46676
rect 15932 48412 15988 48468
rect 16156 59724 16212 59780
rect 16156 59388 16212 59444
rect 16604 61516 16660 61572
rect 16604 60508 16660 60564
rect 16828 66162 16884 66164
rect 16828 66110 16830 66162
rect 16830 66110 16882 66162
rect 16882 66110 16884 66162
rect 16828 66108 16884 66110
rect 17724 81676 17780 81732
rect 18620 85090 18676 85092
rect 18620 85038 18622 85090
rect 18622 85038 18674 85090
rect 18674 85038 18676 85090
rect 18620 85036 18676 85038
rect 18732 84028 18788 84084
rect 18222 83914 18278 83916
rect 18222 83862 18224 83914
rect 18224 83862 18276 83914
rect 18276 83862 18278 83914
rect 18222 83860 18278 83862
rect 18326 83914 18382 83916
rect 18326 83862 18328 83914
rect 18328 83862 18380 83914
rect 18380 83862 18382 83914
rect 18326 83860 18382 83862
rect 18430 83914 18486 83916
rect 18430 83862 18432 83914
rect 18432 83862 18484 83914
rect 18484 83862 18486 83914
rect 18430 83860 18486 83862
rect 18620 83916 18676 83972
rect 18396 83468 18452 83524
rect 19404 85874 19460 85876
rect 19404 85822 19406 85874
rect 19406 85822 19458 85874
rect 19458 85822 19460 85874
rect 19404 85820 19460 85822
rect 19068 85708 19124 85764
rect 19964 88844 20020 88900
rect 20076 88338 20132 88340
rect 20076 88286 20078 88338
rect 20078 88286 20130 88338
rect 20130 88286 20132 88338
rect 20076 88284 20132 88286
rect 21868 94386 21924 94388
rect 21868 94334 21870 94386
rect 21870 94334 21922 94386
rect 21922 94334 21924 94386
rect 21868 94332 21924 94334
rect 21308 93772 21364 93828
rect 21756 94220 21812 94276
rect 21624 94106 21680 94108
rect 21624 94054 21626 94106
rect 21626 94054 21678 94106
rect 21678 94054 21680 94106
rect 21624 94052 21680 94054
rect 21728 94106 21784 94108
rect 21728 94054 21730 94106
rect 21730 94054 21782 94106
rect 21782 94054 21784 94106
rect 21728 94052 21784 94054
rect 21832 94106 21888 94108
rect 21832 94054 21834 94106
rect 21834 94054 21886 94106
rect 21886 94054 21888 94106
rect 21832 94052 21888 94054
rect 21644 93884 21700 93940
rect 21980 93884 22036 93940
rect 21756 93772 21812 93828
rect 22428 93884 22484 93940
rect 21532 92764 21588 92820
rect 21624 92538 21680 92540
rect 21624 92486 21626 92538
rect 21626 92486 21678 92538
rect 21678 92486 21680 92538
rect 21624 92484 21680 92486
rect 21728 92538 21784 92540
rect 21728 92486 21730 92538
rect 21730 92486 21782 92538
rect 21782 92486 21784 92538
rect 21728 92484 21784 92486
rect 21832 92538 21888 92540
rect 21832 92486 21834 92538
rect 21834 92486 21886 92538
rect 21886 92486 21888 92538
rect 21832 92484 21888 92486
rect 21196 92204 21252 92260
rect 22092 92204 22148 92260
rect 21980 91308 22036 91364
rect 22540 92764 22596 92820
rect 22316 92258 22372 92260
rect 22316 92206 22318 92258
rect 22318 92206 22370 92258
rect 22370 92206 22372 92258
rect 22316 92204 22372 92206
rect 22428 92092 22484 92148
rect 22316 91362 22372 91364
rect 22316 91310 22318 91362
rect 22318 91310 22370 91362
rect 22370 91310 22372 91362
rect 22316 91308 22372 91310
rect 21624 90970 21680 90972
rect 21624 90918 21626 90970
rect 21626 90918 21678 90970
rect 21678 90918 21680 90970
rect 21624 90916 21680 90918
rect 21728 90970 21784 90972
rect 21728 90918 21730 90970
rect 21730 90918 21782 90970
rect 21782 90918 21784 90970
rect 21728 90916 21784 90918
rect 21832 90970 21888 90972
rect 21832 90918 21834 90970
rect 21834 90918 21886 90970
rect 21886 90918 21888 90970
rect 21832 90916 21888 90918
rect 22876 92146 22932 92148
rect 22876 92094 22878 92146
rect 22878 92094 22930 92146
rect 22930 92094 22932 92146
rect 22876 92092 22932 92094
rect 22652 91980 22708 92036
rect 23212 102338 23268 102340
rect 23212 102286 23214 102338
rect 23214 102286 23266 102338
rect 23266 102286 23268 102338
rect 23212 102284 23268 102286
rect 23996 104076 24052 104132
rect 25026 116842 25082 116844
rect 25026 116790 25028 116842
rect 25028 116790 25080 116842
rect 25080 116790 25082 116842
rect 25026 116788 25082 116790
rect 25130 116842 25186 116844
rect 25130 116790 25132 116842
rect 25132 116790 25184 116842
rect 25184 116790 25186 116842
rect 25130 116788 25186 116790
rect 25234 116842 25290 116844
rect 25234 116790 25236 116842
rect 25236 116790 25288 116842
rect 25288 116790 25290 116842
rect 25234 116788 25290 116790
rect 25026 115274 25082 115276
rect 25026 115222 25028 115274
rect 25028 115222 25080 115274
rect 25080 115222 25082 115274
rect 25026 115220 25082 115222
rect 25130 115274 25186 115276
rect 25130 115222 25132 115274
rect 25132 115222 25184 115274
rect 25184 115222 25186 115274
rect 25130 115220 25186 115222
rect 25234 115274 25290 115276
rect 25234 115222 25236 115274
rect 25236 115222 25288 115274
rect 25288 115222 25290 115274
rect 25234 115220 25290 115222
rect 24780 114604 24836 114660
rect 28428 117626 28484 117628
rect 28428 117574 28430 117626
rect 28430 117574 28482 117626
rect 28482 117574 28484 117626
rect 28428 117572 28484 117574
rect 28532 117626 28588 117628
rect 28532 117574 28534 117626
rect 28534 117574 28586 117626
rect 28586 117574 28588 117626
rect 28532 117572 28588 117574
rect 28636 117626 28692 117628
rect 28636 117574 28638 117626
rect 28638 117574 28690 117626
rect 28690 117574 28692 117626
rect 28636 117572 28692 117574
rect 28428 116058 28484 116060
rect 28428 116006 28430 116058
rect 28430 116006 28482 116058
rect 28482 116006 28484 116058
rect 28428 116004 28484 116006
rect 28532 116058 28588 116060
rect 28532 116006 28534 116058
rect 28534 116006 28586 116058
rect 28586 116006 28588 116058
rect 28532 116004 28588 116006
rect 28636 116058 28692 116060
rect 28636 116006 28638 116058
rect 28638 116006 28690 116058
rect 28690 116006 28692 116058
rect 28636 116004 28692 116006
rect 28428 114490 28484 114492
rect 28428 114438 28430 114490
rect 28430 114438 28482 114490
rect 28482 114438 28484 114490
rect 28428 114436 28484 114438
rect 28532 114490 28588 114492
rect 28532 114438 28534 114490
rect 28534 114438 28586 114490
rect 28586 114438 28588 114490
rect 28532 114436 28588 114438
rect 28636 114490 28692 114492
rect 28636 114438 28638 114490
rect 28638 114438 28690 114490
rect 28690 114438 28692 114490
rect 28636 114436 28692 114438
rect 25026 113706 25082 113708
rect 25026 113654 25028 113706
rect 25028 113654 25080 113706
rect 25080 113654 25082 113706
rect 25026 113652 25082 113654
rect 25130 113706 25186 113708
rect 25130 113654 25132 113706
rect 25132 113654 25184 113706
rect 25184 113654 25186 113706
rect 25130 113652 25186 113654
rect 25234 113706 25290 113708
rect 25234 113654 25236 113706
rect 25236 113654 25288 113706
rect 25288 113654 25290 113706
rect 25234 113652 25290 113654
rect 25900 113314 25956 113316
rect 25900 113262 25902 113314
rect 25902 113262 25954 113314
rect 25954 113262 25956 113314
rect 25900 113260 25956 113262
rect 25026 112138 25082 112140
rect 25026 112086 25028 112138
rect 25028 112086 25080 112138
rect 25080 112086 25082 112138
rect 25026 112084 25082 112086
rect 25130 112138 25186 112140
rect 25130 112086 25132 112138
rect 25132 112086 25184 112138
rect 25184 112086 25186 112138
rect 25130 112084 25186 112086
rect 25234 112138 25290 112140
rect 25234 112086 25236 112138
rect 25236 112086 25288 112138
rect 25288 112086 25290 112138
rect 25234 112084 25290 112086
rect 28028 111916 28084 111972
rect 26684 111746 26740 111748
rect 26684 111694 26686 111746
rect 26686 111694 26738 111746
rect 26738 111694 26740 111746
rect 26684 111692 26740 111694
rect 25026 110570 25082 110572
rect 25026 110518 25028 110570
rect 25028 110518 25080 110570
rect 25080 110518 25082 110570
rect 25026 110516 25082 110518
rect 25130 110570 25186 110572
rect 25130 110518 25132 110570
rect 25132 110518 25184 110570
rect 25184 110518 25186 110570
rect 25130 110516 25186 110518
rect 25234 110570 25290 110572
rect 25234 110518 25236 110570
rect 25236 110518 25288 110570
rect 25288 110518 25290 110570
rect 25234 110516 25290 110518
rect 24332 107602 24388 107604
rect 24332 107550 24334 107602
rect 24334 107550 24386 107602
rect 24386 107550 24388 107602
rect 24332 107548 24388 107550
rect 24332 106034 24388 106036
rect 24332 105982 24334 106034
rect 24334 105982 24386 106034
rect 24386 105982 24388 106034
rect 24332 105980 24388 105982
rect 25026 109002 25082 109004
rect 25026 108950 25028 109002
rect 25028 108950 25080 109002
rect 25080 108950 25082 109002
rect 25026 108948 25082 108950
rect 25130 109002 25186 109004
rect 25130 108950 25132 109002
rect 25132 108950 25184 109002
rect 25184 108950 25186 109002
rect 25130 108948 25186 108950
rect 25234 109002 25290 109004
rect 25234 108950 25236 109002
rect 25236 108950 25288 109002
rect 25288 108950 25290 109002
rect 25234 108948 25290 108950
rect 24892 108668 24948 108724
rect 25900 108668 25956 108724
rect 25676 108610 25732 108612
rect 25676 108558 25678 108610
rect 25678 108558 25730 108610
rect 25730 108558 25732 108610
rect 25676 108556 25732 108558
rect 24668 108386 24724 108388
rect 24668 108334 24670 108386
rect 24670 108334 24722 108386
rect 24722 108334 24724 108386
rect 24668 108332 24724 108334
rect 24668 107548 24724 107604
rect 24780 107436 24836 107492
rect 25026 107434 25082 107436
rect 25026 107382 25028 107434
rect 25028 107382 25080 107434
rect 25080 107382 25082 107434
rect 25026 107380 25082 107382
rect 25130 107434 25186 107436
rect 25130 107382 25132 107434
rect 25132 107382 25184 107434
rect 25184 107382 25186 107434
rect 25130 107380 25186 107382
rect 25234 107434 25290 107436
rect 25234 107382 25236 107434
rect 25236 107382 25288 107434
rect 25288 107382 25290 107434
rect 25234 107380 25290 107382
rect 24444 105644 24500 105700
rect 24220 103122 24276 103124
rect 24220 103070 24222 103122
rect 24222 103070 24274 103122
rect 24274 103070 24276 103122
rect 24220 103068 24276 103070
rect 23884 102396 23940 102452
rect 25340 106258 25396 106260
rect 25340 106206 25342 106258
rect 25342 106206 25394 106258
rect 25394 106206 25396 106258
rect 25340 106204 25396 106206
rect 26684 108556 26740 108612
rect 27244 108386 27300 108388
rect 27244 108334 27246 108386
rect 27246 108334 27298 108386
rect 27298 108334 27300 108386
rect 27244 108332 27300 108334
rect 24892 105980 24948 106036
rect 25026 105866 25082 105868
rect 25026 105814 25028 105866
rect 25028 105814 25080 105866
rect 25080 105814 25082 105866
rect 25026 105812 25082 105814
rect 25130 105866 25186 105868
rect 25130 105814 25132 105866
rect 25132 105814 25184 105866
rect 25184 105814 25186 105866
rect 25130 105812 25186 105814
rect 25234 105866 25290 105868
rect 25234 105814 25236 105866
rect 25236 105814 25288 105866
rect 25288 105814 25290 105866
rect 25234 105812 25290 105814
rect 26236 105586 26292 105588
rect 26236 105534 26238 105586
rect 26238 105534 26290 105586
rect 26290 105534 26292 105586
rect 26236 105532 26292 105534
rect 28028 105532 28084 105588
rect 24780 105308 24836 105364
rect 24668 105196 24724 105252
rect 24444 104076 24500 104132
rect 25676 105250 25732 105252
rect 25676 105198 25678 105250
rect 25678 105198 25730 105250
rect 25730 105198 25732 105250
rect 25676 105196 25732 105198
rect 26012 105196 26068 105252
rect 25026 104298 25082 104300
rect 25026 104246 25028 104298
rect 25028 104246 25080 104298
rect 25080 104246 25082 104298
rect 25026 104244 25082 104246
rect 25130 104298 25186 104300
rect 25130 104246 25132 104298
rect 25132 104246 25184 104298
rect 25184 104246 25186 104298
rect 25130 104244 25186 104246
rect 25234 104298 25290 104300
rect 25234 104246 25236 104298
rect 25236 104246 25288 104298
rect 25288 104246 25290 104298
rect 25234 104244 25290 104246
rect 26684 105250 26740 105252
rect 26684 105198 26686 105250
rect 26686 105198 26738 105250
rect 26738 105198 26740 105250
rect 26684 105196 26740 105198
rect 26684 104076 26740 104132
rect 27580 104130 27636 104132
rect 27580 104078 27582 104130
rect 27582 104078 27634 104130
rect 27634 104078 27636 104130
rect 27580 104076 27636 104078
rect 24556 102956 24612 103012
rect 25340 103010 25396 103012
rect 25340 102958 25342 103010
rect 25342 102958 25394 103010
rect 25394 102958 25396 103010
rect 25340 102956 25396 102958
rect 25026 102730 25082 102732
rect 25026 102678 25028 102730
rect 25028 102678 25080 102730
rect 25080 102678 25082 102730
rect 25026 102676 25082 102678
rect 25130 102730 25186 102732
rect 25130 102678 25132 102730
rect 25132 102678 25184 102730
rect 25184 102678 25186 102730
rect 25130 102676 25186 102678
rect 25234 102730 25290 102732
rect 25234 102678 25236 102730
rect 25236 102678 25288 102730
rect 25288 102678 25290 102730
rect 25234 102676 25290 102678
rect 24780 102450 24836 102452
rect 24780 102398 24782 102450
rect 24782 102398 24834 102450
rect 24834 102398 24836 102450
rect 24780 102396 24836 102398
rect 23324 100716 23380 100772
rect 23324 99986 23380 99988
rect 23324 99934 23326 99986
rect 23326 99934 23378 99986
rect 23378 99934 23380 99986
rect 23324 99932 23380 99934
rect 23884 101554 23940 101556
rect 23884 101502 23886 101554
rect 23886 101502 23938 101554
rect 23938 101502 23940 101554
rect 23884 101500 23940 101502
rect 24220 100770 24276 100772
rect 24220 100718 24222 100770
rect 24222 100718 24274 100770
rect 24274 100718 24276 100770
rect 24220 100716 24276 100718
rect 25026 101162 25082 101164
rect 25026 101110 25028 101162
rect 25028 101110 25080 101162
rect 25080 101110 25082 101162
rect 25026 101108 25082 101110
rect 25130 101162 25186 101164
rect 25130 101110 25132 101162
rect 25132 101110 25184 101162
rect 25184 101110 25186 101162
rect 25130 101108 25186 101110
rect 25234 101162 25290 101164
rect 25234 101110 25236 101162
rect 25236 101110 25288 101162
rect 25288 101110 25290 101162
rect 25234 101108 25290 101110
rect 24108 99986 24164 99988
rect 24108 99934 24110 99986
rect 24110 99934 24162 99986
rect 24162 99934 24164 99986
rect 24108 99932 24164 99934
rect 23660 99148 23716 99204
rect 23884 99036 23940 99092
rect 23772 98924 23828 98980
rect 23100 97634 23156 97636
rect 23100 97582 23102 97634
rect 23102 97582 23154 97634
rect 23154 97582 23156 97634
rect 23100 97580 23156 97582
rect 23324 97580 23380 97636
rect 23660 97692 23716 97748
rect 23884 98194 23940 98196
rect 23884 98142 23886 98194
rect 23886 98142 23938 98194
rect 23938 98142 23940 98194
rect 23884 98140 23940 98142
rect 23996 97916 24052 97972
rect 23772 97468 23828 97524
rect 24220 97468 24276 97524
rect 23212 95954 23268 95956
rect 23212 95902 23214 95954
rect 23214 95902 23266 95954
rect 23266 95902 23268 95954
rect 23212 95900 23268 95902
rect 23324 95842 23380 95844
rect 23324 95790 23326 95842
rect 23326 95790 23378 95842
rect 23378 95790 23380 95842
rect 23324 95788 23380 95790
rect 23884 96738 23940 96740
rect 23884 96686 23886 96738
rect 23886 96686 23938 96738
rect 23938 96686 23940 96738
rect 23884 96684 23940 96686
rect 24444 98530 24500 98532
rect 24444 98478 24446 98530
rect 24446 98478 24498 98530
rect 24498 98478 24500 98530
rect 24444 98476 24500 98478
rect 24892 100716 24948 100772
rect 25452 100604 25508 100660
rect 26684 100658 26740 100660
rect 26684 100606 26686 100658
rect 26686 100606 26738 100658
rect 26738 100606 26740 100658
rect 26684 100604 26740 100606
rect 24892 99932 24948 99988
rect 25026 99594 25082 99596
rect 25026 99542 25028 99594
rect 25028 99542 25080 99594
rect 25080 99542 25082 99594
rect 25026 99540 25082 99542
rect 25130 99594 25186 99596
rect 25130 99542 25132 99594
rect 25132 99542 25184 99594
rect 25184 99542 25186 99594
rect 25130 99540 25186 99542
rect 25234 99594 25290 99596
rect 25234 99542 25236 99594
rect 25236 99542 25288 99594
rect 25288 99542 25290 99594
rect 25234 99540 25290 99542
rect 24668 99036 24724 99092
rect 23436 95452 23492 95508
rect 24668 97692 24724 97748
rect 25228 98476 25284 98532
rect 25026 98026 25082 98028
rect 25026 97974 25028 98026
rect 25028 97974 25080 98026
rect 25080 97974 25082 98026
rect 25026 97972 25082 97974
rect 25130 98026 25186 98028
rect 25130 97974 25132 98026
rect 25132 97974 25184 98026
rect 25184 97974 25186 98026
rect 25130 97972 25186 97974
rect 25234 98026 25290 98028
rect 25234 97974 25236 98026
rect 25236 97974 25288 98026
rect 25288 97974 25290 98026
rect 25234 97972 25290 97974
rect 25340 97858 25396 97860
rect 25340 97806 25342 97858
rect 25342 97806 25394 97858
rect 25394 97806 25396 97858
rect 25340 97804 25396 97806
rect 27356 99932 27412 99988
rect 28028 99932 28084 99988
rect 25452 97746 25508 97748
rect 25452 97694 25454 97746
rect 25454 97694 25506 97746
rect 25506 97694 25508 97746
rect 25452 97692 25508 97694
rect 25676 98924 25732 98980
rect 25116 97580 25172 97636
rect 24892 97522 24948 97524
rect 24892 97470 24894 97522
rect 24894 97470 24946 97522
rect 24946 97470 24948 97522
rect 24892 97468 24948 97470
rect 25564 97580 25620 97636
rect 25026 96458 25082 96460
rect 25026 96406 25028 96458
rect 25028 96406 25080 96458
rect 25080 96406 25082 96458
rect 25026 96404 25082 96406
rect 25130 96458 25186 96460
rect 25130 96406 25132 96458
rect 25132 96406 25184 96458
rect 25184 96406 25186 96458
rect 25130 96404 25186 96406
rect 25234 96458 25290 96460
rect 25234 96406 25236 96458
rect 25236 96406 25288 96458
rect 25288 96406 25290 96458
rect 25234 96404 25290 96406
rect 24444 96012 24500 96068
rect 24556 95900 24612 95956
rect 24220 95282 24276 95284
rect 24220 95230 24222 95282
rect 24222 95230 24274 95282
rect 24274 95230 24276 95282
rect 24220 95228 24276 95230
rect 25228 96066 25284 96068
rect 25228 96014 25230 96066
rect 25230 96014 25282 96066
rect 25282 96014 25284 96066
rect 25228 96012 25284 96014
rect 25340 95954 25396 95956
rect 25340 95902 25342 95954
rect 25342 95902 25394 95954
rect 25394 95902 25396 95954
rect 25340 95900 25396 95902
rect 25452 95842 25508 95844
rect 25452 95790 25454 95842
rect 25454 95790 25506 95842
rect 25506 95790 25508 95842
rect 25452 95788 25508 95790
rect 25676 98476 25732 98532
rect 27356 98140 27412 98196
rect 26796 97580 26852 97636
rect 26684 97522 26740 97524
rect 26684 97470 26686 97522
rect 26686 97470 26738 97522
rect 26738 97470 26740 97522
rect 26684 97468 26740 97470
rect 27356 97634 27412 97636
rect 27356 97582 27358 97634
rect 27358 97582 27410 97634
rect 27410 97582 27412 97634
rect 27356 97580 27412 97582
rect 26236 96684 26292 96740
rect 25340 95282 25396 95284
rect 25340 95230 25342 95282
rect 25342 95230 25394 95282
rect 25394 95230 25396 95282
rect 25340 95228 25396 95230
rect 25564 95228 25620 95284
rect 25026 94890 25082 94892
rect 25026 94838 25028 94890
rect 25028 94838 25080 94890
rect 25080 94838 25082 94890
rect 25026 94836 25082 94838
rect 25130 94890 25186 94892
rect 25130 94838 25132 94890
rect 25132 94838 25184 94890
rect 25184 94838 25186 94890
rect 25130 94836 25186 94838
rect 25234 94890 25290 94892
rect 25234 94838 25236 94890
rect 25236 94838 25288 94890
rect 25288 94838 25290 94890
rect 25234 94836 25290 94838
rect 23100 93602 23156 93604
rect 23100 93550 23102 93602
rect 23102 93550 23154 93602
rect 23154 93550 23156 93602
rect 23100 93548 23156 93550
rect 25026 93322 25082 93324
rect 25026 93270 25028 93322
rect 25028 93270 25080 93322
rect 25080 93270 25082 93322
rect 25026 93268 25082 93270
rect 25130 93322 25186 93324
rect 25130 93270 25132 93322
rect 25132 93270 25184 93322
rect 25184 93270 25186 93322
rect 25130 93268 25186 93270
rect 25234 93322 25290 93324
rect 25234 93270 25236 93322
rect 25236 93270 25288 93322
rect 25288 93270 25290 93322
rect 25234 93268 25290 93270
rect 25228 92988 25284 93044
rect 23324 92818 23380 92820
rect 23324 92766 23326 92818
rect 23326 92766 23378 92818
rect 23378 92766 23380 92818
rect 23324 92764 23380 92766
rect 23772 92706 23828 92708
rect 23772 92654 23774 92706
rect 23774 92654 23826 92706
rect 23826 92654 23828 92706
rect 23772 92652 23828 92654
rect 23548 92316 23604 92372
rect 23100 92258 23156 92260
rect 23100 92206 23102 92258
rect 23102 92206 23154 92258
rect 23154 92206 23156 92258
rect 23100 92204 23156 92206
rect 24332 92316 24388 92372
rect 22988 91644 23044 91700
rect 22876 91586 22932 91588
rect 22876 91534 22878 91586
rect 22878 91534 22930 91586
rect 22930 91534 22932 91586
rect 22876 91532 22932 91534
rect 22540 91250 22596 91252
rect 22540 91198 22542 91250
rect 22542 91198 22594 91250
rect 22594 91198 22596 91250
rect 22540 91196 22596 91198
rect 22428 91084 22484 91140
rect 22764 91084 22820 91140
rect 22092 90748 22148 90804
rect 22876 90860 22932 90916
rect 20860 90636 20916 90692
rect 20412 90412 20468 90468
rect 20860 90466 20916 90468
rect 20860 90414 20862 90466
rect 20862 90414 20914 90466
rect 20914 90414 20916 90466
rect 20860 90412 20916 90414
rect 21308 90578 21364 90580
rect 21308 90526 21310 90578
rect 21310 90526 21362 90578
rect 21362 90526 21364 90578
rect 21308 90524 21364 90526
rect 21756 89852 21812 89908
rect 23436 91980 23492 92036
rect 23884 91532 23940 91588
rect 23212 90860 23268 90916
rect 23436 91084 23492 91140
rect 23548 91362 23604 91364
rect 23548 91310 23550 91362
rect 23550 91310 23602 91362
rect 23602 91310 23604 91362
rect 23548 91308 23604 91310
rect 23548 90860 23604 90916
rect 23772 91250 23828 91252
rect 23772 91198 23774 91250
rect 23774 91198 23826 91250
rect 23826 91198 23828 91250
rect 23772 91196 23828 91198
rect 23436 90690 23492 90692
rect 23436 90638 23438 90690
rect 23438 90638 23490 90690
rect 23490 90638 23492 90690
rect 23436 90636 23492 90638
rect 22652 90300 22708 90356
rect 21868 89682 21924 89684
rect 21868 89630 21870 89682
rect 21870 89630 21922 89682
rect 21922 89630 21924 89682
rect 21868 89628 21924 89630
rect 21624 89402 21680 89404
rect 21624 89350 21626 89402
rect 21626 89350 21678 89402
rect 21678 89350 21680 89402
rect 21624 89348 21680 89350
rect 21728 89402 21784 89404
rect 21728 89350 21730 89402
rect 21730 89350 21782 89402
rect 21782 89350 21784 89402
rect 21728 89348 21784 89350
rect 21832 89402 21888 89404
rect 21832 89350 21834 89402
rect 21834 89350 21886 89402
rect 21886 89350 21888 89402
rect 21980 89404 22036 89460
rect 21832 89348 21888 89350
rect 21420 89010 21476 89012
rect 21420 88958 21422 89010
rect 21422 88958 21474 89010
rect 21474 88958 21476 89010
rect 21420 88956 21476 88958
rect 22204 89570 22260 89572
rect 22204 89518 22206 89570
rect 22206 89518 22258 89570
rect 22258 89518 22260 89570
rect 22204 89516 22260 89518
rect 25228 92258 25284 92260
rect 25228 92206 25230 92258
rect 25230 92206 25282 92258
rect 25282 92206 25284 92258
rect 25228 92204 25284 92206
rect 24668 92146 24724 92148
rect 24668 92094 24670 92146
rect 24670 92094 24722 92146
rect 24722 92094 24724 92146
rect 24668 92092 24724 92094
rect 24332 91980 24388 92036
rect 25452 92316 25508 92372
rect 25026 91754 25082 91756
rect 25026 91702 25028 91754
rect 25028 91702 25080 91754
rect 25080 91702 25082 91754
rect 25026 91700 25082 91702
rect 25130 91754 25186 91756
rect 25130 91702 25132 91754
rect 25132 91702 25184 91754
rect 25184 91702 25186 91754
rect 25130 91700 25186 91702
rect 25234 91754 25290 91756
rect 25234 91702 25236 91754
rect 25236 91702 25288 91754
rect 25288 91702 25290 91754
rect 25234 91700 25290 91702
rect 25228 91532 25284 91588
rect 24220 90972 24276 91028
rect 24332 91084 24388 91140
rect 23884 90860 23940 90916
rect 23212 90300 23268 90356
rect 22764 89852 22820 89908
rect 22876 89964 22932 90020
rect 22764 89682 22820 89684
rect 22764 89630 22766 89682
rect 22766 89630 22818 89682
rect 22818 89630 22820 89682
rect 22764 89628 22820 89630
rect 23324 89516 23380 89572
rect 22652 88956 22708 89012
rect 20748 88844 20804 88900
rect 20524 88338 20580 88340
rect 20524 88286 20526 88338
rect 20526 88286 20578 88338
rect 20578 88286 20580 88338
rect 20524 88284 20580 88286
rect 21532 88898 21588 88900
rect 21532 88846 21534 88898
rect 21534 88846 21586 88898
rect 21586 88846 21588 88898
rect 21532 88844 21588 88846
rect 22988 89292 23044 89348
rect 20412 87836 20468 87892
rect 21624 87834 21680 87836
rect 21624 87782 21626 87834
rect 21626 87782 21678 87834
rect 21678 87782 21680 87834
rect 21624 87780 21680 87782
rect 21728 87834 21784 87836
rect 21728 87782 21730 87834
rect 21730 87782 21782 87834
rect 21782 87782 21784 87834
rect 21728 87780 21784 87782
rect 21832 87834 21888 87836
rect 21832 87782 21834 87834
rect 21834 87782 21886 87834
rect 21886 87782 21888 87834
rect 21832 87780 21888 87782
rect 20300 87052 20356 87108
rect 19628 85708 19684 85764
rect 19180 85314 19236 85316
rect 19180 85262 19182 85314
rect 19182 85262 19234 85314
rect 19234 85262 19236 85314
rect 19180 85260 19236 85262
rect 19068 83916 19124 83972
rect 19404 84140 19460 84196
rect 18222 82346 18278 82348
rect 18222 82294 18224 82346
rect 18224 82294 18276 82346
rect 18276 82294 18278 82346
rect 18222 82292 18278 82294
rect 18326 82346 18382 82348
rect 18326 82294 18328 82346
rect 18328 82294 18380 82346
rect 18380 82294 18382 82346
rect 18326 82292 18382 82294
rect 18430 82346 18486 82348
rect 18430 82294 18432 82346
rect 18432 82294 18484 82346
rect 18484 82294 18486 82346
rect 18430 82292 18486 82294
rect 18620 82292 18676 82348
rect 18396 82066 18452 82068
rect 18396 82014 18398 82066
rect 18398 82014 18450 82066
rect 18450 82014 18452 82066
rect 18396 82012 18452 82014
rect 17724 81170 17780 81172
rect 17724 81118 17726 81170
rect 17726 81118 17778 81170
rect 17778 81118 17780 81170
rect 17724 81116 17780 81118
rect 17612 80892 17668 80948
rect 17948 80892 18004 80948
rect 17836 80556 17892 80612
rect 17500 80220 17556 80276
rect 17836 79884 17892 79940
rect 17724 79826 17780 79828
rect 17724 79774 17726 79826
rect 17726 79774 17778 79826
rect 17778 79774 17780 79826
rect 17724 79772 17780 79774
rect 17612 79714 17668 79716
rect 17612 79662 17614 79714
rect 17614 79662 17666 79714
rect 17666 79662 17668 79714
rect 17612 79660 17668 79662
rect 17500 78258 17556 78260
rect 17500 78206 17502 78258
rect 17502 78206 17554 78258
rect 17554 78206 17556 78258
rect 17500 78204 17556 78206
rect 18956 83634 19012 83636
rect 18956 83582 18958 83634
rect 18958 83582 19010 83634
rect 19010 83582 19012 83634
rect 18956 83580 19012 83582
rect 18172 80892 18228 80948
rect 18222 80778 18278 80780
rect 18222 80726 18224 80778
rect 18224 80726 18276 80778
rect 18276 80726 18278 80778
rect 18222 80724 18278 80726
rect 18326 80778 18382 80780
rect 18326 80726 18328 80778
rect 18328 80726 18380 80778
rect 18380 80726 18382 80778
rect 18326 80724 18382 80726
rect 18430 80778 18486 80780
rect 18430 80726 18432 80778
rect 18432 80726 18484 80778
rect 18484 80726 18486 80778
rect 18430 80724 18486 80726
rect 19292 83522 19348 83524
rect 19292 83470 19294 83522
rect 19294 83470 19346 83522
rect 19346 83470 19348 83522
rect 19292 83468 19348 83470
rect 18844 83410 18900 83412
rect 18844 83358 18846 83410
rect 18846 83358 18898 83410
rect 18898 83358 18900 83410
rect 18844 83356 18900 83358
rect 19516 84812 19572 84868
rect 20188 86434 20244 86436
rect 20188 86382 20190 86434
rect 20190 86382 20242 86434
rect 20242 86382 20244 86434
rect 20188 86380 20244 86382
rect 19964 86268 20020 86324
rect 19964 85708 20020 85764
rect 21084 86604 21140 86660
rect 20748 86268 20804 86324
rect 20524 84924 20580 84980
rect 20076 84418 20132 84420
rect 20076 84366 20078 84418
rect 20078 84366 20130 84418
rect 20130 84366 20132 84418
rect 20076 84364 20132 84366
rect 20636 84866 20692 84868
rect 20636 84814 20638 84866
rect 20638 84814 20690 84866
rect 20690 84814 20692 84866
rect 20636 84812 20692 84814
rect 19292 82236 19348 82292
rect 19068 81340 19124 81396
rect 19292 81394 19348 81396
rect 19292 81342 19294 81394
rect 19294 81342 19346 81394
rect 19346 81342 19348 81394
rect 19292 81340 19348 81342
rect 19404 81170 19460 81172
rect 19404 81118 19406 81170
rect 19406 81118 19458 81170
rect 19458 81118 19460 81170
rect 19404 81116 19460 81118
rect 19068 81004 19124 81060
rect 18844 80556 18900 80612
rect 20188 83916 20244 83972
rect 19628 83244 19684 83300
rect 18732 80220 18788 80276
rect 17948 79602 18004 79604
rect 17948 79550 17950 79602
rect 17950 79550 18002 79602
rect 18002 79550 18004 79602
rect 17948 79548 18004 79550
rect 18172 79324 18228 79380
rect 18222 79210 18278 79212
rect 18222 79158 18224 79210
rect 18224 79158 18276 79210
rect 18276 79158 18278 79210
rect 18222 79156 18278 79158
rect 18326 79210 18382 79212
rect 18326 79158 18328 79210
rect 18328 79158 18380 79210
rect 18380 79158 18382 79210
rect 18326 79156 18382 79158
rect 18430 79210 18486 79212
rect 18430 79158 18432 79210
rect 18432 79158 18484 79210
rect 18484 79158 18486 79210
rect 18430 79156 18486 79158
rect 19068 79660 19124 79716
rect 19068 79324 19124 79380
rect 17724 78204 17780 78260
rect 18172 78204 18228 78260
rect 17164 77308 17220 77364
rect 17388 77868 17444 77924
rect 17388 77420 17444 77476
rect 17500 77980 17556 78036
rect 17948 78034 18004 78036
rect 17948 77982 17950 78034
rect 17950 77982 18002 78034
rect 18002 77982 18004 78034
rect 17948 77980 18004 77982
rect 17612 77868 17668 77924
rect 17836 77810 17892 77812
rect 17836 77758 17838 77810
rect 17838 77758 17890 77810
rect 17890 77758 17892 77810
rect 17836 77756 17892 77758
rect 17612 77308 17668 77364
rect 18508 78204 18564 78260
rect 18508 77810 18564 77812
rect 18508 77758 18510 77810
rect 18510 77758 18562 77810
rect 18562 77758 18564 77810
rect 18508 77756 18564 77758
rect 18222 77642 18278 77644
rect 18222 77590 18224 77642
rect 18224 77590 18276 77642
rect 18276 77590 18278 77642
rect 18222 77588 18278 77590
rect 18326 77642 18382 77644
rect 18326 77590 18328 77642
rect 18328 77590 18380 77642
rect 18380 77590 18382 77642
rect 18326 77588 18382 77590
rect 18430 77642 18486 77644
rect 18430 77590 18432 77642
rect 18432 77590 18484 77642
rect 18484 77590 18486 77642
rect 18430 77588 18486 77590
rect 18396 77138 18452 77140
rect 18396 77086 18398 77138
rect 18398 77086 18450 77138
rect 18450 77086 18452 77138
rect 18396 77084 18452 77086
rect 17500 75628 17556 75684
rect 17612 76300 17668 76356
rect 17388 75516 17444 75572
rect 17276 75458 17332 75460
rect 17276 75406 17278 75458
rect 17278 75406 17330 75458
rect 17330 75406 17332 75458
rect 17276 75404 17332 75406
rect 17724 75570 17780 75572
rect 17724 75518 17726 75570
rect 17726 75518 17778 75570
rect 17778 75518 17780 75570
rect 17724 75516 17780 75518
rect 17948 75404 18004 75460
rect 17724 75068 17780 75124
rect 17276 74620 17332 74676
rect 17276 72492 17332 72548
rect 17276 71538 17332 71540
rect 17276 71486 17278 71538
rect 17278 71486 17330 71538
rect 17330 71486 17332 71538
rect 17276 71484 17332 71486
rect 17276 71260 17332 71316
rect 18222 76074 18278 76076
rect 18222 76022 18224 76074
rect 18224 76022 18276 76074
rect 18276 76022 18278 76074
rect 18222 76020 18278 76022
rect 18326 76074 18382 76076
rect 18326 76022 18328 76074
rect 18328 76022 18380 76074
rect 18380 76022 18382 76074
rect 18326 76020 18382 76022
rect 18430 76074 18486 76076
rect 18430 76022 18432 76074
rect 18432 76022 18484 76074
rect 18484 76022 18486 76074
rect 18430 76020 18486 76022
rect 18284 75682 18340 75684
rect 18284 75630 18286 75682
rect 18286 75630 18338 75682
rect 18338 75630 18340 75682
rect 18284 75628 18340 75630
rect 18060 75068 18116 75124
rect 19292 78540 19348 78596
rect 19180 78428 19236 78484
rect 18844 78316 18900 78372
rect 18844 77756 18900 77812
rect 18620 75068 18676 75124
rect 18222 74506 18278 74508
rect 18222 74454 18224 74506
rect 18224 74454 18276 74506
rect 18276 74454 18278 74506
rect 18222 74452 18278 74454
rect 18326 74506 18382 74508
rect 18326 74454 18328 74506
rect 18328 74454 18380 74506
rect 18380 74454 18382 74506
rect 18326 74452 18382 74454
rect 18430 74506 18486 74508
rect 18430 74454 18432 74506
rect 18432 74454 18484 74506
rect 18484 74454 18486 74506
rect 18430 74452 18486 74454
rect 18620 74508 18676 74564
rect 18508 74172 18564 74228
rect 17500 73164 17556 73220
rect 17500 71932 17556 71988
rect 17500 70588 17556 70644
rect 18060 73442 18116 73444
rect 18060 73390 18062 73442
rect 18062 73390 18114 73442
rect 18114 73390 18116 73442
rect 18060 73388 18116 73390
rect 17948 73330 18004 73332
rect 17948 73278 17950 73330
rect 17950 73278 18002 73330
rect 18002 73278 18004 73330
rect 17948 73276 18004 73278
rect 17388 69186 17444 69188
rect 17388 69134 17390 69186
rect 17390 69134 17442 69186
rect 17442 69134 17444 69186
rect 17388 69132 17444 69134
rect 17612 68626 17668 68628
rect 17612 68574 17614 68626
rect 17614 68574 17666 68626
rect 17666 68574 17668 68626
rect 17612 68572 17668 68574
rect 17388 68460 17444 68516
rect 17612 67058 17668 67060
rect 17612 67006 17614 67058
rect 17614 67006 17666 67058
rect 17666 67006 17668 67058
rect 17612 67004 17668 67006
rect 17500 65996 17556 66052
rect 17276 65490 17332 65492
rect 17276 65438 17278 65490
rect 17278 65438 17330 65490
rect 17330 65438 17332 65490
rect 17276 65436 17332 65438
rect 16828 63308 16884 63364
rect 16828 62748 16884 62804
rect 16828 62354 16884 62356
rect 16828 62302 16830 62354
rect 16830 62302 16882 62354
rect 16882 62302 16884 62354
rect 16828 62300 16884 62302
rect 16828 61852 16884 61908
rect 16828 61404 16884 61460
rect 18284 73330 18340 73332
rect 18284 73278 18286 73330
rect 18286 73278 18338 73330
rect 18338 73278 18340 73330
rect 18284 73276 18340 73278
rect 18956 76300 19012 76356
rect 18956 76076 19012 76132
rect 18956 74172 19012 74228
rect 19292 77922 19348 77924
rect 19292 77870 19294 77922
rect 19294 77870 19346 77922
rect 19346 77870 19348 77922
rect 19292 77868 19348 77870
rect 19180 77756 19236 77812
rect 19180 74508 19236 74564
rect 19292 74172 19348 74228
rect 18732 73724 18788 73780
rect 18222 72938 18278 72940
rect 18222 72886 18224 72938
rect 18224 72886 18276 72938
rect 18276 72886 18278 72938
rect 18222 72884 18278 72886
rect 18326 72938 18382 72940
rect 18326 72886 18328 72938
rect 18328 72886 18380 72938
rect 18380 72886 18382 72938
rect 18326 72884 18382 72886
rect 18430 72938 18486 72940
rect 18430 72886 18432 72938
rect 18432 72886 18484 72938
rect 18484 72886 18486 72938
rect 18430 72884 18486 72886
rect 17836 72658 17892 72660
rect 17836 72606 17838 72658
rect 17838 72606 17890 72658
rect 17890 72606 17892 72658
rect 17836 72604 17892 72606
rect 18844 73612 18900 73668
rect 19516 80556 19572 80612
rect 19964 83468 20020 83524
rect 19740 81116 19796 81172
rect 20412 84028 20468 84084
rect 20188 81954 20244 81956
rect 20188 81902 20190 81954
rect 20190 81902 20242 81954
rect 20242 81902 20244 81954
rect 20188 81900 20244 81902
rect 20300 83356 20356 83412
rect 20300 81788 20356 81844
rect 19852 80556 19908 80612
rect 19964 81116 20020 81172
rect 19740 78706 19796 78708
rect 19740 78654 19742 78706
rect 19742 78654 19794 78706
rect 19794 78654 19796 78706
rect 19740 78652 19796 78654
rect 19628 78540 19684 78596
rect 19964 79660 20020 79716
rect 20188 78818 20244 78820
rect 20188 78766 20190 78818
rect 20190 78766 20242 78818
rect 20242 78766 20244 78818
rect 20188 78764 20244 78766
rect 19740 78034 19796 78036
rect 19740 77982 19742 78034
rect 19742 77982 19794 78034
rect 19794 77982 19796 78034
rect 19740 77980 19796 77982
rect 19628 75570 19684 75572
rect 19628 75518 19630 75570
rect 19630 75518 19682 75570
rect 19682 75518 19684 75570
rect 19628 75516 19684 75518
rect 19516 74002 19572 74004
rect 19516 73950 19518 74002
rect 19518 73950 19570 74002
rect 19570 73950 19572 74002
rect 19516 73948 19572 73950
rect 18620 71932 18676 71988
rect 18956 72380 19012 72436
rect 18060 71820 18116 71876
rect 17948 71372 18004 71428
rect 17948 71148 18004 71204
rect 17836 69356 17892 69412
rect 17836 68908 17892 68964
rect 18284 71650 18340 71652
rect 18284 71598 18286 71650
rect 18286 71598 18338 71650
rect 18338 71598 18340 71650
rect 18284 71596 18340 71598
rect 18222 71370 18278 71372
rect 18222 71318 18224 71370
rect 18224 71318 18276 71370
rect 18276 71318 18278 71370
rect 18222 71316 18278 71318
rect 18326 71370 18382 71372
rect 18326 71318 18328 71370
rect 18328 71318 18380 71370
rect 18380 71318 18382 71370
rect 18326 71316 18382 71318
rect 18430 71370 18486 71372
rect 18430 71318 18432 71370
rect 18432 71318 18484 71370
rect 18484 71318 18486 71370
rect 18430 71316 18486 71318
rect 18284 70754 18340 70756
rect 18284 70702 18286 70754
rect 18286 70702 18338 70754
rect 18338 70702 18340 70754
rect 18284 70700 18340 70702
rect 18172 70588 18228 70644
rect 19180 72546 19236 72548
rect 19180 72494 19182 72546
rect 19182 72494 19234 72546
rect 19234 72494 19236 72546
rect 19180 72492 19236 72494
rect 19068 71932 19124 71988
rect 18844 71148 18900 71204
rect 19068 70924 19124 70980
rect 19068 70588 19124 70644
rect 18396 70252 18452 70308
rect 18222 69802 18278 69804
rect 18222 69750 18224 69802
rect 18224 69750 18276 69802
rect 18276 69750 18278 69802
rect 18222 69748 18278 69750
rect 18326 69802 18382 69804
rect 18326 69750 18328 69802
rect 18328 69750 18380 69802
rect 18380 69750 18382 69802
rect 18326 69748 18382 69750
rect 18430 69802 18486 69804
rect 18430 69750 18432 69802
rect 18432 69750 18484 69802
rect 18484 69750 18486 69802
rect 18430 69748 18486 69750
rect 18732 69298 18788 69300
rect 18732 69246 18734 69298
rect 18734 69246 18786 69298
rect 18786 69246 18788 69298
rect 18732 69244 18788 69246
rect 18284 69020 18340 69076
rect 17948 68796 18004 68852
rect 17836 68738 17892 68740
rect 17836 68686 17838 68738
rect 17838 68686 17890 68738
rect 17890 68686 17892 68738
rect 17836 68684 17892 68686
rect 18222 68234 18278 68236
rect 18222 68182 18224 68234
rect 18224 68182 18276 68234
rect 18276 68182 18278 68234
rect 18222 68180 18278 68182
rect 18326 68234 18382 68236
rect 18326 68182 18328 68234
rect 18328 68182 18380 68234
rect 18380 68182 18382 68234
rect 18326 68180 18382 68182
rect 18430 68234 18486 68236
rect 18430 68182 18432 68234
rect 18432 68182 18484 68234
rect 18484 68182 18486 68234
rect 18430 68180 18486 68182
rect 18060 67340 18116 67396
rect 17948 67170 18004 67172
rect 17948 67118 17950 67170
rect 17950 67118 18002 67170
rect 18002 67118 18004 67170
rect 17948 67116 18004 67118
rect 18732 67900 18788 67956
rect 18620 67116 18676 67172
rect 18956 69468 19012 69524
rect 19516 72492 19572 72548
rect 19516 72322 19572 72324
rect 19516 72270 19518 72322
rect 19518 72270 19570 72322
rect 19570 72270 19572 72322
rect 19516 72268 19572 72270
rect 19292 71484 19348 71540
rect 19516 70754 19572 70756
rect 19516 70702 19518 70754
rect 19518 70702 19570 70754
rect 19570 70702 19572 70754
rect 19516 70700 19572 70702
rect 20972 84252 21028 84308
rect 21196 86492 21252 86548
rect 22764 86828 22820 86884
rect 22876 89180 22932 89236
rect 23324 89292 23380 89348
rect 23212 89180 23268 89236
rect 23548 89010 23604 89012
rect 23548 88958 23550 89010
rect 23550 88958 23602 89010
rect 23602 88958 23604 89010
rect 23548 88956 23604 88958
rect 24220 89292 24276 89348
rect 24108 89068 24164 89124
rect 23996 88956 24052 89012
rect 24556 91196 24612 91252
rect 26236 95842 26292 95844
rect 26236 95790 26238 95842
rect 26238 95790 26290 95842
rect 26290 95790 26292 95842
rect 26236 95788 26292 95790
rect 27132 95788 27188 95844
rect 26012 95282 26068 95284
rect 26012 95230 26014 95282
rect 26014 95230 26066 95282
rect 26066 95230 26068 95282
rect 26012 95228 26068 95230
rect 25900 94108 25956 94164
rect 26908 94108 26964 94164
rect 25788 92876 25844 92932
rect 26124 92988 26180 93044
rect 26348 92930 26404 92932
rect 26348 92878 26350 92930
rect 26350 92878 26402 92930
rect 26402 92878 26404 92930
rect 26348 92876 26404 92878
rect 25788 92428 25844 92484
rect 25788 92146 25844 92148
rect 25788 92094 25790 92146
rect 25790 92094 25842 92146
rect 25842 92094 25844 92146
rect 25788 92092 25844 92094
rect 25564 91644 25620 91700
rect 25676 91532 25732 91588
rect 25564 91362 25620 91364
rect 25564 91310 25566 91362
rect 25566 91310 25618 91362
rect 25618 91310 25620 91362
rect 25564 91308 25620 91310
rect 25788 91308 25844 91364
rect 26012 92652 26068 92708
rect 26012 91980 26068 92036
rect 26572 92652 26628 92708
rect 28428 112922 28484 112924
rect 28428 112870 28430 112922
rect 28430 112870 28482 112922
rect 28482 112870 28484 112922
rect 28428 112868 28484 112870
rect 28532 112922 28588 112924
rect 28532 112870 28534 112922
rect 28534 112870 28586 112922
rect 28586 112870 28588 112922
rect 28532 112868 28588 112870
rect 28636 112922 28692 112924
rect 28636 112870 28638 112922
rect 28638 112870 28690 112922
rect 28690 112870 28692 112922
rect 28636 112868 28692 112870
rect 28252 111916 28308 111972
rect 28428 111354 28484 111356
rect 28428 111302 28430 111354
rect 28430 111302 28482 111354
rect 28482 111302 28484 111354
rect 28428 111300 28484 111302
rect 28532 111354 28588 111356
rect 28532 111302 28534 111354
rect 28534 111302 28586 111354
rect 28586 111302 28588 111354
rect 28532 111300 28588 111302
rect 28636 111354 28692 111356
rect 28636 111302 28638 111354
rect 28638 111302 28690 111354
rect 28690 111302 28692 111354
rect 28636 111300 28692 111302
rect 28428 109786 28484 109788
rect 28428 109734 28430 109786
rect 28430 109734 28482 109786
rect 28482 109734 28484 109786
rect 28428 109732 28484 109734
rect 28532 109786 28588 109788
rect 28532 109734 28534 109786
rect 28534 109734 28586 109786
rect 28586 109734 28588 109786
rect 28532 109732 28588 109734
rect 28636 109786 28692 109788
rect 28636 109734 28638 109786
rect 28638 109734 28690 109786
rect 28690 109734 28692 109786
rect 28636 109732 28692 109734
rect 28252 108332 28308 108388
rect 28428 108218 28484 108220
rect 28428 108166 28430 108218
rect 28430 108166 28482 108218
rect 28482 108166 28484 108218
rect 28428 108164 28484 108166
rect 28532 108218 28588 108220
rect 28532 108166 28534 108218
rect 28534 108166 28586 108218
rect 28586 108166 28588 108218
rect 28532 108164 28588 108166
rect 28636 108218 28692 108220
rect 28636 108166 28638 108218
rect 28638 108166 28690 108218
rect 28690 108166 28692 108218
rect 28636 108164 28692 108166
rect 28428 106650 28484 106652
rect 28428 106598 28430 106650
rect 28430 106598 28482 106650
rect 28482 106598 28484 106650
rect 28428 106596 28484 106598
rect 28532 106650 28588 106652
rect 28532 106598 28534 106650
rect 28534 106598 28586 106650
rect 28586 106598 28588 106650
rect 28532 106596 28588 106598
rect 28636 106650 28692 106652
rect 28636 106598 28638 106650
rect 28638 106598 28690 106650
rect 28690 106598 28692 106650
rect 28636 106596 28692 106598
rect 28252 105532 28308 105588
rect 28428 105082 28484 105084
rect 28428 105030 28430 105082
rect 28430 105030 28482 105082
rect 28482 105030 28484 105082
rect 28428 105028 28484 105030
rect 28532 105082 28588 105084
rect 28532 105030 28534 105082
rect 28534 105030 28586 105082
rect 28586 105030 28588 105082
rect 28532 105028 28588 105030
rect 28636 105082 28692 105084
rect 28636 105030 28638 105082
rect 28638 105030 28690 105082
rect 28690 105030 28692 105082
rect 28636 105028 28692 105030
rect 28428 103514 28484 103516
rect 28428 103462 28430 103514
rect 28430 103462 28482 103514
rect 28482 103462 28484 103514
rect 28428 103460 28484 103462
rect 28532 103514 28588 103516
rect 28532 103462 28534 103514
rect 28534 103462 28586 103514
rect 28586 103462 28588 103514
rect 28532 103460 28588 103462
rect 28636 103514 28692 103516
rect 28636 103462 28638 103514
rect 28638 103462 28690 103514
rect 28690 103462 28692 103514
rect 28636 103460 28692 103462
rect 28428 101946 28484 101948
rect 28428 101894 28430 101946
rect 28430 101894 28482 101946
rect 28482 101894 28484 101946
rect 28428 101892 28484 101894
rect 28532 101946 28588 101948
rect 28532 101894 28534 101946
rect 28534 101894 28586 101946
rect 28586 101894 28588 101946
rect 28532 101892 28588 101894
rect 28636 101946 28692 101948
rect 28636 101894 28638 101946
rect 28638 101894 28690 101946
rect 28690 101894 28692 101946
rect 28636 101892 28692 101894
rect 28428 100378 28484 100380
rect 28428 100326 28430 100378
rect 28430 100326 28482 100378
rect 28482 100326 28484 100378
rect 28428 100324 28484 100326
rect 28532 100378 28588 100380
rect 28532 100326 28534 100378
rect 28534 100326 28586 100378
rect 28586 100326 28588 100378
rect 28532 100324 28588 100326
rect 28636 100378 28692 100380
rect 28636 100326 28638 100378
rect 28638 100326 28690 100378
rect 28690 100326 28692 100378
rect 28636 100324 28692 100326
rect 28428 98810 28484 98812
rect 28428 98758 28430 98810
rect 28430 98758 28482 98810
rect 28482 98758 28484 98810
rect 28428 98756 28484 98758
rect 28532 98810 28588 98812
rect 28532 98758 28534 98810
rect 28534 98758 28586 98810
rect 28586 98758 28588 98810
rect 28532 98756 28588 98758
rect 28636 98810 28692 98812
rect 28636 98758 28638 98810
rect 28638 98758 28690 98810
rect 28690 98758 28692 98810
rect 28636 98756 28692 98758
rect 28428 97242 28484 97244
rect 28428 97190 28430 97242
rect 28430 97190 28482 97242
rect 28482 97190 28484 97242
rect 28428 97188 28484 97190
rect 28532 97242 28588 97244
rect 28532 97190 28534 97242
rect 28534 97190 28586 97242
rect 28586 97190 28588 97242
rect 28532 97188 28588 97190
rect 28636 97242 28692 97244
rect 28636 97190 28638 97242
rect 28638 97190 28690 97242
rect 28690 97190 28692 97242
rect 28636 97188 28692 97190
rect 28428 95674 28484 95676
rect 28428 95622 28430 95674
rect 28430 95622 28482 95674
rect 28482 95622 28484 95674
rect 28428 95620 28484 95622
rect 28532 95674 28588 95676
rect 28532 95622 28534 95674
rect 28534 95622 28586 95674
rect 28586 95622 28588 95674
rect 28532 95620 28588 95622
rect 28636 95674 28692 95676
rect 28636 95622 28638 95674
rect 28638 95622 28690 95674
rect 28690 95622 28692 95674
rect 28636 95620 28692 95622
rect 28140 95340 28196 95396
rect 28428 94106 28484 94108
rect 28428 94054 28430 94106
rect 28430 94054 28482 94106
rect 28482 94054 28484 94106
rect 28428 94052 28484 94054
rect 28532 94106 28588 94108
rect 28532 94054 28534 94106
rect 28534 94054 28586 94106
rect 28586 94054 28588 94106
rect 28532 94052 28588 94054
rect 28636 94106 28692 94108
rect 28636 94054 28638 94106
rect 28638 94054 28690 94106
rect 28690 94054 28692 94106
rect 28636 94052 28692 94054
rect 27020 92428 27076 92484
rect 26460 91586 26516 91588
rect 26460 91534 26462 91586
rect 26462 91534 26514 91586
rect 26514 91534 26516 91586
rect 26460 91532 26516 91534
rect 26684 91868 26740 91924
rect 26908 91756 26964 91812
rect 26908 91362 26964 91364
rect 26908 91310 26910 91362
rect 26910 91310 26962 91362
rect 26962 91310 26964 91362
rect 26908 91308 26964 91310
rect 26012 91250 26068 91252
rect 26012 91198 26014 91250
rect 26014 91198 26066 91250
rect 26066 91198 26068 91250
rect 26012 91196 26068 91198
rect 25676 91084 25732 91140
rect 25116 90748 25172 90804
rect 25026 90186 25082 90188
rect 25026 90134 25028 90186
rect 25028 90134 25080 90186
rect 25080 90134 25082 90186
rect 25026 90132 25082 90134
rect 25130 90186 25186 90188
rect 25130 90134 25132 90186
rect 25132 90134 25184 90186
rect 25184 90134 25186 90186
rect 25130 90132 25186 90134
rect 25234 90186 25290 90188
rect 25234 90134 25236 90186
rect 25236 90134 25288 90186
rect 25288 90134 25290 90186
rect 25234 90132 25290 90134
rect 24332 88844 24388 88900
rect 24556 89180 24612 89236
rect 24556 88898 24612 88900
rect 24556 88846 24558 88898
rect 24558 88846 24610 88898
rect 24610 88846 24612 88898
rect 24556 88844 24612 88846
rect 24332 88396 24388 88452
rect 24556 88226 24612 88228
rect 24556 88174 24558 88226
rect 24558 88174 24610 88226
rect 24610 88174 24612 88226
rect 24556 88172 24612 88174
rect 24108 88060 24164 88116
rect 26012 90972 26068 91028
rect 25788 90412 25844 90468
rect 25788 89628 25844 89684
rect 25116 89404 25172 89460
rect 25564 89516 25620 89572
rect 25340 89010 25396 89012
rect 25340 88958 25342 89010
rect 25342 88958 25394 89010
rect 25394 88958 25396 89010
rect 25340 88956 25396 88958
rect 26348 90524 26404 90580
rect 26012 89570 26068 89572
rect 26012 89518 26014 89570
rect 26014 89518 26066 89570
rect 26066 89518 26068 89570
rect 26012 89516 26068 89518
rect 25564 88844 25620 88900
rect 25026 88618 25082 88620
rect 25026 88566 25028 88618
rect 25028 88566 25080 88618
rect 25080 88566 25082 88618
rect 25026 88564 25082 88566
rect 25130 88618 25186 88620
rect 25130 88566 25132 88618
rect 25132 88566 25184 88618
rect 25184 88566 25186 88618
rect 25130 88564 25186 88566
rect 25234 88618 25290 88620
rect 25234 88566 25236 88618
rect 25236 88566 25288 88618
rect 25288 88566 25290 88618
rect 25234 88564 25290 88566
rect 24780 88450 24836 88452
rect 24780 88398 24782 88450
rect 24782 88398 24834 88450
rect 24834 88398 24836 88450
rect 24780 88396 24836 88398
rect 25004 88060 25060 88116
rect 27132 91138 27188 91140
rect 27132 91086 27134 91138
rect 27134 91086 27186 91138
rect 27186 91086 27188 91138
rect 27132 91084 27188 91086
rect 27580 90578 27636 90580
rect 27580 90526 27582 90578
rect 27582 90526 27634 90578
rect 27634 90526 27636 90578
rect 27580 90524 27636 90526
rect 28428 92538 28484 92540
rect 28428 92486 28430 92538
rect 28430 92486 28482 92538
rect 28482 92486 28484 92538
rect 28428 92484 28484 92486
rect 28532 92538 28588 92540
rect 28532 92486 28534 92538
rect 28534 92486 28586 92538
rect 28586 92486 28588 92538
rect 28532 92484 28588 92486
rect 28636 92538 28692 92540
rect 28636 92486 28638 92538
rect 28638 92486 28690 92538
rect 28690 92486 28692 92538
rect 28636 92484 28692 92486
rect 28140 91532 28196 91588
rect 28428 90970 28484 90972
rect 28428 90918 28430 90970
rect 28430 90918 28482 90970
rect 28482 90918 28484 90970
rect 28428 90916 28484 90918
rect 28532 90970 28588 90972
rect 28532 90918 28534 90970
rect 28534 90918 28586 90970
rect 28586 90918 28588 90970
rect 28532 90916 28588 90918
rect 28636 90970 28692 90972
rect 28636 90918 28638 90970
rect 28638 90918 28690 90970
rect 28690 90918 28692 90970
rect 28636 90916 28692 90918
rect 28028 90466 28084 90468
rect 28028 90414 28030 90466
rect 28030 90414 28082 90466
rect 28082 90414 28084 90466
rect 28028 90412 28084 90414
rect 27020 89628 27076 89684
rect 23996 86882 24052 86884
rect 23996 86830 23998 86882
rect 23998 86830 24050 86882
rect 24050 86830 24052 86882
rect 23996 86828 24052 86830
rect 21980 86546 22036 86548
rect 21980 86494 21982 86546
rect 21982 86494 22034 86546
rect 22034 86494 22036 86546
rect 21980 86492 22036 86494
rect 22876 86546 22932 86548
rect 22876 86494 22878 86546
rect 22878 86494 22930 86546
rect 22930 86494 22932 86546
rect 22876 86492 22932 86494
rect 21532 86434 21588 86436
rect 21532 86382 21534 86434
rect 21534 86382 21586 86434
rect 21586 86382 21588 86434
rect 21532 86380 21588 86382
rect 21624 86266 21680 86268
rect 21624 86214 21626 86266
rect 21626 86214 21678 86266
rect 21678 86214 21680 86266
rect 21624 86212 21680 86214
rect 21728 86266 21784 86268
rect 21728 86214 21730 86266
rect 21730 86214 21782 86266
rect 21782 86214 21784 86266
rect 21728 86212 21784 86214
rect 21832 86266 21888 86268
rect 21832 86214 21834 86266
rect 21834 86214 21886 86266
rect 21886 86214 21888 86266
rect 21832 86212 21888 86214
rect 24332 86716 24388 86772
rect 24444 87276 24500 87332
rect 23548 86604 23604 86660
rect 20748 84140 20804 84196
rect 21308 84978 21364 84980
rect 21308 84926 21310 84978
rect 21310 84926 21362 84978
rect 21362 84926 21364 84978
rect 21308 84924 21364 84926
rect 21624 84698 21680 84700
rect 21624 84646 21626 84698
rect 21626 84646 21678 84698
rect 21678 84646 21680 84698
rect 21624 84644 21680 84646
rect 21728 84698 21784 84700
rect 21728 84646 21730 84698
rect 21730 84646 21782 84698
rect 21782 84646 21784 84698
rect 21728 84644 21784 84646
rect 21832 84698 21888 84700
rect 21832 84646 21834 84698
rect 21834 84646 21886 84698
rect 21886 84646 21888 84698
rect 21832 84644 21888 84646
rect 21308 84364 21364 84420
rect 21196 84028 21252 84084
rect 21532 84028 21588 84084
rect 20748 83692 20804 83748
rect 21644 83916 21700 83972
rect 21980 83522 22036 83524
rect 21980 83470 21982 83522
rect 21982 83470 22034 83522
rect 22034 83470 22036 83522
rect 21980 83468 22036 83470
rect 20860 83020 20916 83076
rect 20524 81842 20580 81844
rect 20524 81790 20526 81842
rect 20526 81790 20578 81842
rect 20578 81790 20580 81842
rect 20524 81788 20580 81790
rect 20748 81730 20804 81732
rect 20748 81678 20750 81730
rect 20750 81678 20802 81730
rect 20802 81678 20804 81730
rect 20748 81676 20804 81678
rect 20636 81228 20692 81284
rect 20748 81340 20804 81396
rect 20524 80274 20580 80276
rect 20524 80222 20526 80274
rect 20526 80222 20578 80274
rect 20578 80222 20580 80274
rect 20524 80220 20580 80222
rect 21308 83244 21364 83300
rect 21084 82850 21140 82852
rect 21084 82798 21086 82850
rect 21086 82798 21138 82850
rect 21138 82798 21140 82850
rect 21084 82796 21140 82798
rect 21308 81788 21364 81844
rect 21196 80220 21252 80276
rect 20860 79660 20916 79716
rect 21624 83130 21680 83132
rect 21624 83078 21626 83130
rect 21626 83078 21678 83130
rect 21678 83078 21680 83130
rect 21624 83076 21680 83078
rect 21728 83130 21784 83132
rect 21728 83078 21730 83130
rect 21730 83078 21782 83130
rect 21782 83078 21784 83130
rect 21728 83076 21784 83078
rect 21832 83130 21888 83132
rect 21832 83078 21834 83130
rect 21834 83078 21886 83130
rect 21886 83078 21888 83130
rect 21832 83076 21888 83078
rect 22764 83916 22820 83972
rect 22876 84812 22932 84868
rect 22652 83804 22708 83860
rect 22652 83634 22708 83636
rect 22652 83582 22654 83634
rect 22654 83582 22706 83634
rect 22706 83582 22708 83634
rect 22652 83580 22708 83582
rect 22428 83468 22484 83524
rect 22092 82850 22148 82852
rect 22092 82798 22094 82850
rect 22094 82798 22146 82850
rect 22146 82798 22148 82850
rect 22092 82796 22148 82798
rect 21532 81954 21588 81956
rect 21532 81902 21534 81954
rect 21534 81902 21586 81954
rect 21586 81902 21588 81954
rect 21532 81900 21588 81902
rect 21980 81676 22036 81732
rect 21624 81562 21680 81564
rect 21624 81510 21626 81562
rect 21626 81510 21678 81562
rect 21678 81510 21680 81562
rect 21624 81508 21680 81510
rect 21728 81562 21784 81564
rect 21728 81510 21730 81562
rect 21730 81510 21782 81562
rect 21782 81510 21784 81562
rect 21728 81508 21784 81510
rect 21832 81562 21888 81564
rect 21832 81510 21834 81562
rect 21834 81510 21886 81562
rect 21886 81510 21888 81562
rect 21832 81508 21888 81510
rect 21980 81116 22036 81172
rect 22540 81900 22596 81956
rect 22652 81788 22708 81844
rect 22988 82460 23044 82516
rect 22764 81340 22820 81396
rect 22988 81170 23044 81172
rect 22988 81118 22990 81170
rect 22990 81118 23042 81170
rect 23042 81118 23044 81170
rect 22988 81116 23044 81118
rect 22540 80556 22596 80612
rect 22092 80444 22148 80500
rect 21624 79994 21680 79996
rect 21624 79942 21626 79994
rect 21626 79942 21678 79994
rect 21678 79942 21680 79994
rect 21624 79940 21680 79942
rect 21728 79994 21784 79996
rect 21728 79942 21730 79994
rect 21730 79942 21782 79994
rect 21782 79942 21784 79994
rect 21728 79940 21784 79942
rect 21832 79994 21888 79996
rect 21832 79942 21834 79994
rect 21834 79942 21886 79994
rect 21886 79942 21888 79994
rect 22092 79996 22148 80052
rect 21832 79940 21888 79942
rect 21532 79602 21588 79604
rect 21532 79550 21534 79602
rect 21534 79550 21586 79602
rect 21586 79550 21588 79602
rect 21532 79548 21588 79550
rect 20412 77756 20468 77812
rect 21868 78652 21924 78708
rect 21532 78594 21588 78596
rect 21532 78542 21534 78594
rect 21534 78542 21586 78594
rect 21586 78542 21588 78594
rect 21532 78540 21588 78542
rect 22092 78594 22148 78596
rect 22092 78542 22094 78594
rect 22094 78542 22146 78594
rect 22146 78542 22148 78594
rect 22092 78540 22148 78542
rect 21308 78428 21364 78484
rect 21624 78426 21680 78428
rect 21624 78374 21626 78426
rect 21626 78374 21678 78426
rect 21678 78374 21680 78426
rect 21624 78372 21680 78374
rect 21728 78426 21784 78428
rect 21728 78374 21730 78426
rect 21730 78374 21782 78426
rect 21782 78374 21784 78426
rect 21728 78372 21784 78374
rect 21832 78426 21888 78428
rect 21832 78374 21834 78426
rect 21834 78374 21886 78426
rect 21886 78374 21888 78426
rect 21832 78372 21888 78374
rect 20636 77420 20692 77476
rect 20524 77308 20580 77364
rect 21084 77196 21140 77252
rect 21420 77196 21476 77252
rect 20188 77084 20244 77140
rect 19964 77026 20020 77028
rect 19964 76974 19966 77026
rect 19966 76974 20018 77026
rect 20018 76974 20020 77026
rect 19964 76972 20020 76974
rect 22092 77756 22148 77812
rect 21980 77250 22036 77252
rect 21980 77198 21982 77250
rect 21982 77198 22034 77250
rect 22034 77198 22036 77250
rect 21980 77196 22036 77198
rect 21624 76858 21680 76860
rect 21624 76806 21626 76858
rect 21626 76806 21678 76858
rect 21678 76806 21680 76858
rect 21624 76804 21680 76806
rect 21728 76858 21784 76860
rect 21728 76806 21730 76858
rect 21730 76806 21782 76858
rect 21782 76806 21784 76858
rect 21728 76804 21784 76806
rect 21832 76858 21888 76860
rect 21832 76806 21834 76858
rect 21834 76806 21886 76858
rect 21886 76806 21888 76858
rect 21832 76804 21888 76806
rect 20636 76300 20692 76356
rect 21420 76300 21476 76356
rect 20748 75740 20804 75796
rect 20188 75682 20244 75684
rect 20188 75630 20190 75682
rect 20190 75630 20242 75682
rect 20242 75630 20244 75682
rect 20188 75628 20244 75630
rect 20412 75404 20468 75460
rect 19964 74732 20020 74788
rect 19852 74114 19908 74116
rect 19852 74062 19854 74114
rect 19854 74062 19906 74114
rect 19906 74062 19908 74114
rect 19852 74060 19908 74062
rect 20300 74114 20356 74116
rect 20300 74062 20302 74114
rect 20302 74062 20354 74114
rect 20354 74062 20356 74114
rect 20300 74060 20356 74062
rect 20300 73554 20356 73556
rect 20300 73502 20302 73554
rect 20302 73502 20354 73554
rect 20354 73502 20356 73554
rect 20300 73500 20356 73502
rect 19740 70924 19796 70980
rect 19516 70252 19572 70308
rect 19404 69522 19460 69524
rect 19404 69470 19406 69522
rect 19406 69470 19458 69522
rect 19458 69470 19460 69522
rect 19404 69468 19460 69470
rect 19068 68796 19124 68852
rect 19516 69132 19572 69188
rect 19404 68850 19460 68852
rect 19404 68798 19406 68850
rect 19406 68798 19458 68850
rect 19458 68798 19460 68850
rect 19404 68796 19460 68798
rect 18956 67842 19012 67844
rect 18956 67790 18958 67842
rect 18958 67790 19010 67842
rect 19010 67790 19012 67842
rect 18956 67788 19012 67790
rect 19292 68460 19348 68516
rect 19292 67900 19348 67956
rect 19068 67676 19124 67732
rect 18396 67058 18452 67060
rect 18396 67006 18398 67058
rect 18398 67006 18450 67058
rect 18450 67006 18452 67058
rect 18396 67004 18452 67006
rect 19404 67618 19460 67620
rect 19404 67566 19406 67618
rect 19406 67566 19458 67618
rect 19458 67566 19460 67618
rect 19404 67564 19460 67566
rect 17836 66892 17892 66948
rect 18222 66666 18278 66668
rect 18222 66614 18224 66666
rect 18224 66614 18276 66666
rect 18276 66614 18278 66666
rect 18222 66612 18278 66614
rect 18326 66666 18382 66668
rect 18326 66614 18328 66666
rect 18328 66614 18380 66666
rect 18380 66614 18382 66666
rect 18326 66612 18382 66614
rect 18430 66666 18486 66668
rect 18430 66614 18432 66666
rect 18432 66614 18484 66666
rect 18484 66614 18486 66666
rect 18430 66612 18486 66614
rect 18060 65602 18116 65604
rect 18060 65550 18062 65602
rect 18062 65550 18114 65602
rect 18114 65550 18116 65602
rect 18060 65548 18116 65550
rect 21756 76354 21812 76356
rect 21756 76302 21758 76354
rect 21758 76302 21810 76354
rect 21810 76302 21812 76354
rect 21756 76300 21812 76302
rect 21532 76076 21588 76132
rect 22204 77138 22260 77140
rect 22204 77086 22206 77138
rect 22206 77086 22258 77138
rect 22258 77086 22260 77138
rect 22204 77084 22260 77086
rect 20748 73442 20804 73444
rect 20748 73390 20750 73442
rect 20750 73390 20802 73442
rect 20802 73390 20804 73442
rect 20748 73388 20804 73390
rect 20524 72268 20580 72324
rect 20188 70978 20244 70980
rect 20188 70926 20190 70978
rect 20190 70926 20242 70978
rect 20242 70926 20244 70978
rect 20188 70924 20244 70926
rect 20524 70924 20580 70980
rect 20188 70700 20244 70756
rect 19852 68796 19908 68852
rect 20076 69132 20132 69188
rect 19852 67676 19908 67732
rect 19740 67564 19796 67620
rect 18956 66108 19012 66164
rect 18508 65436 18564 65492
rect 18284 65378 18340 65380
rect 18284 65326 18286 65378
rect 18286 65326 18338 65378
rect 18338 65326 18340 65378
rect 18284 65324 18340 65326
rect 17276 64652 17332 64708
rect 16940 61068 16996 61124
rect 17388 64482 17444 64484
rect 17388 64430 17390 64482
rect 17390 64430 17442 64482
rect 17442 64430 17444 64482
rect 17388 64428 17444 64430
rect 17388 63868 17444 63924
rect 17724 63980 17780 64036
rect 17164 63138 17220 63140
rect 17164 63086 17166 63138
rect 17166 63086 17218 63138
rect 17218 63086 17220 63138
rect 17164 63084 17220 63086
rect 17500 62748 17556 62804
rect 17164 62636 17220 62692
rect 17724 62636 17780 62692
rect 17500 62242 17556 62244
rect 17500 62190 17502 62242
rect 17502 62190 17554 62242
rect 17554 62190 17556 62242
rect 17500 62188 17556 62190
rect 17612 62076 17668 62132
rect 17724 61740 17780 61796
rect 17164 60956 17220 61012
rect 17388 60396 17444 60452
rect 17276 60172 17332 60228
rect 16828 59218 16884 59220
rect 16828 59166 16830 59218
rect 16830 59166 16882 59218
rect 16882 59166 16884 59218
rect 16828 59164 16884 59166
rect 16380 58434 16436 58436
rect 16380 58382 16382 58434
rect 16382 58382 16434 58434
rect 16434 58382 16436 58434
rect 16380 58380 16436 58382
rect 16492 57596 16548 57652
rect 16492 57036 16548 57092
rect 16268 53730 16324 53732
rect 16268 53678 16270 53730
rect 16270 53678 16322 53730
rect 16322 53678 16324 53730
rect 16268 53676 16324 53678
rect 16268 53452 16324 53508
rect 16268 52892 16324 52948
rect 16268 51660 16324 51716
rect 16156 51378 16212 51380
rect 16156 51326 16158 51378
rect 16158 51326 16210 51378
rect 16210 51326 16212 51378
rect 16156 51324 16212 51326
rect 16156 50764 16212 50820
rect 16604 56924 16660 56980
rect 16828 57596 16884 57652
rect 16604 56252 16660 56308
rect 16604 55468 16660 55524
rect 16716 53676 16772 53732
rect 16492 53004 16548 53060
rect 17052 58268 17108 58324
rect 17052 56866 17108 56868
rect 17052 56814 17054 56866
rect 17054 56814 17106 56866
rect 17106 56814 17108 56866
rect 17052 56812 17108 56814
rect 16940 56364 16996 56420
rect 16940 55970 16996 55972
rect 16940 55918 16942 55970
rect 16942 55918 16994 55970
rect 16994 55918 16996 55970
rect 16940 55916 16996 55918
rect 17164 55186 17220 55188
rect 17164 55134 17166 55186
rect 17166 55134 17218 55186
rect 17218 55134 17220 55186
rect 17164 55132 17220 55134
rect 17500 59836 17556 59892
rect 17612 60396 17668 60452
rect 17500 57708 17556 57764
rect 17388 56364 17444 56420
rect 17836 61180 17892 61236
rect 17948 60786 18004 60788
rect 17948 60734 17950 60786
rect 17950 60734 18002 60786
rect 18002 60734 18004 60786
rect 17948 60732 18004 60734
rect 17836 60508 17892 60564
rect 17836 57596 17892 57652
rect 18222 65098 18278 65100
rect 18222 65046 18224 65098
rect 18224 65046 18276 65098
rect 18276 65046 18278 65098
rect 18222 65044 18278 65046
rect 18326 65098 18382 65100
rect 18326 65046 18328 65098
rect 18328 65046 18380 65098
rect 18380 65046 18382 65098
rect 18326 65044 18382 65046
rect 18430 65098 18486 65100
rect 18430 65046 18432 65098
rect 18432 65046 18484 65098
rect 18484 65046 18486 65098
rect 18430 65044 18486 65046
rect 18222 63530 18278 63532
rect 18222 63478 18224 63530
rect 18224 63478 18276 63530
rect 18276 63478 18278 63530
rect 18222 63476 18278 63478
rect 18326 63530 18382 63532
rect 18326 63478 18328 63530
rect 18328 63478 18380 63530
rect 18380 63478 18382 63530
rect 18326 63476 18382 63478
rect 18430 63530 18486 63532
rect 18430 63478 18432 63530
rect 18432 63478 18484 63530
rect 18484 63478 18486 63530
rect 18430 63476 18486 63478
rect 18172 63362 18228 63364
rect 18172 63310 18174 63362
rect 18174 63310 18226 63362
rect 18226 63310 18228 63362
rect 18172 63308 18228 63310
rect 18732 65602 18788 65604
rect 18732 65550 18734 65602
rect 18734 65550 18786 65602
rect 18786 65550 18788 65602
rect 18732 65548 18788 65550
rect 19068 65996 19124 66052
rect 19404 66050 19460 66052
rect 19404 65998 19406 66050
rect 19406 65998 19458 66050
rect 19458 65998 19460 66050
rect 19404 65996 19460 65998
rect 20300 70252 20356 70308
rect 20412 69186 20468 69188
rect 20412 69134 20414 69186
rect 20414 69134 20466 69186
rect 20466 69134 20468 69186
rect 20412 69132 20468 69134
rect 20188 68124 20244 68180
rect 20188 67676 20244 67732
rect 20300 67788 20356 67844
rect 20748 71820 20804 71876
rect 21624 75290 21680 75292
rect 21624 75238 21626 75290
rect 21626 75238 21678 75290
rect 21678 75238 21680 75290
rect 21624 75236 21680 75238
rect 21728 75290 21784 75292
rect 21728 75238 21730 75290
rect 21730 75238 21782 75290
rect 21782 75238 21784 75290
rect 21728 75236 21784 75238
rect 21832 75290 21888 75292
rect 21832 75238 21834 75290
rect 21834 75238 21886 75290
rect 21886 75238 21888 75290
rect 21832 75236 21888 75238
rect 21084 72940 21140 72996
rect 23884 86380 23940 86436
rect 25564 87330 25620 87332
rect 25564 87278 25566 87330
rect 25566 87278 25618 87330
rect 25618 87278 25620 87330
rect 25564 87276 25620 87278
rect 24892 87164 24948 87220
rect 24668 85820 24724 85876
rect 24556 85762 24612 85764
rect 24556 85710 24558 85762
rect 24558 85710 24610 85762
rect 24610 85710 24612 85762
rect 24556 85708 24612 85710
rect 23996 85650 24052 85652
rect 23996 85598 23998 85650
rect 23998 85598 24050 85650
rect 24050 85598 24052 85650
rect 23996 85596 24052 85598
rect 25026 87050 25082 87052
rect 25026 86998 25028 87050
rect 25028 86998 25080 87050
rect 25080 86998 25082 87050
rect 25026 86996 25082 86998
rect 25130 87050 25186 87052
rect 25130 86998 25132 87050
rect 25132 86998 25184 87050
rect 25184 86998 25186 87050
rect 25130 86996 25186 86998
rect 25234 87050 25290 87052
rect 25234 86998 25236 87050
rect 25236 86998 25288 87050
rect 25288 86998 25290 87050
rect 25234 86996 25290 86998
rect 25004 86044 25060 86100
rect 25788 87442 25844 87444
rect 25788 87390 25790 87442
rect 25790 87390 25842 87442
rect 25842 87390 25844 87442
rect 25788 87388 25844 87390
rect 26348 87276 26404 87332
rect 26460 87388 26516 87444
rect 26012 87052 26068 87108
rect 26796 88226 26852 88228
rect 26796 88174 26798 88226
rect 26798 88174 26850 88226
rect 26850 88174 26852 88226
rect 26796 88172 26852 88174
rect 25788 86098 25844 86100
rect 25788 86046 25790 86098
rect 25790 86046 25842 86098
rect 25842 86046 25844 86098
rect 25788 86044 25844 86046
rect 25452 85874 25508 85876
rect 25452 85822 25454 85874
rect 25454 85822 25506 85874
rect 25506 85822 25508 85874
rect 25452 85820 25508 85822
rect 26348 85708 26404 85764
rect 26460 85596 26516 85652
rect 25026 85482 25082 85484
rect 25026 85430 25028 85482
rect 25028 85430 25080 85482
rect 25080 85430 25082 85482
rect 25026 85428 25082 85430
rect 25130 85482 25186 85484
rect 25130 85430 25132 85482
rect 25132 85430 25184 85482
rect 25184 85430 25186 85482
rect 25130 85428 25186 85430
rect 25234 85482 25290 85484
rect 25234 85430 25236 85482
rect 25236 85430 25288 85482
rect 25288 85430 25290 85482
rect 25234 85428 25290 85430
rect 25452 85314 25508 85316
rect 25452 85262 25454 85314
rect 25454 85262 25506 85314
rect 25506 85262 25508 85314
rect 25452 85260 25508 85262
rect 24220 85202 24276 85204
rect 24220 85150 24222 85202
rect 24222 85150 24274 85202
rect 24274 85150 24276 85202
rect 24220 85148 24276 85150
rect 25564 85148 25620 85204
rect 23212 83692 23268 83748
rect 24668 84866 24724 84868
rect 24668 84814 24670 84866
rect 24670 84814 24722 84866
rect 24722 84814 24724 84866
rect 24668 84812 24724 84814
rect 23660 84140 23716 84196
rect 23548 83580 23604 83636
rect 23660 83916 23716 83972
rect 24444 84306 24500 84308
rect 24444 84254 24446 84306
rect 24446 84254 24498 84306
rect 24498 84254 24500 84306
rect 24444 84252 24500 84254
rect 25676 85090 25732 85092
rect 25676 85038 25678 85090
rect 25678 85038 25730 85090
rect 25730 85038 25732 85090
rect 25676 85036 25732 85038
rect 26124 85036 26180 85092
rect 26572 85260 26628 85316
rect 24780 84028 24836 84084
rect 25564 84306 25620 84308
rect 25564 84254 25566 84306
rect 25566 84254 25618 84306
rect 25618 84254 25620 84306
rect 25564 84252 25620 84254
rect 25026 83914 25082 83916
rect 23772 83468 23828 83524
rect 24220 83804 24276 83860
rect 25026 83862 25028 83914
rect 25028 83862 25080 83914
rect 25080 83862 25082 83914
rect 25026 83860 25082 83862
rect 25130 83914 25186 83916
rect 25130 83862 25132 83914
rect 25132 83862 25184 83914
rect 25184 83862 25186 83914
rect 25130 83860 25186 83862
rect 25234 83914 25290 83916
rect 25234 83862 25236 83914
rect 25236 83862 25288 83914
rect 25288 83862 25290 83914
rect 25234 83860 25290 83862
rect 24332 83634 24388 83636
rect 24332 83582 24334 83634
rect 24334 83582 24386 83634
rect 24386 83582 24388 83634
rect 24332 83580 24388 83582
rect 24444 83522 24500 83524
rect 24444 83470 24446 83522
rect 24446 83470 24498 83522
rect 24498 83470 24500 83522
rect 24444 83468 24500 83470
rect 24556 82796 24612 82852
rect 23212 81954 23268 81956
rect 23212 81902 23214 81954
rect 23214 81902 23266 81954
rect 23266 81902 23268 81954
rect 23212 81900 23268 81902
rect 22652 80108 22708 80164
rect 22540 78540 22596 78596
rect 22764 78594 22820 78596
rect 22764 78542 22766 78594
rect 22766 78542 22818 78594
rect 22818 78542 22820 78594
rect 22764 78540 22820 78542
rect 22540 76300 22596 76356
rect 21308 73052 21364 73108
rect 22316 75794 22372 75796
rect 22316 75742 22318 75794
rect 22318 75742 22370 75794
rect 22370 75742 22372 75794
rect 22316 75740 22372 75742
rect 21624 73722 21680 73724
rect 21624 73670 21626 73722
rect 21626 73670 21678 73722
rect 21678 73670 21680 73722
rect 21624 73668 21680 73670
rect 21728 73722 21784 73724
rect 21728 73670 21730 73722
rect 21730 73670 21782 73722
rect 21782 73670 21784 73722
rect 21728 73668 21784 73670
rect 21832 73722 21888 73724
rect 21832 73670 21834 73722
rect 21834 73670 21886 73722
rect 21886 73670 21888 73722
rect 21832 73668 21888 73670
rect 24668 82684 24724 82740
rect 23772 82012 23828 82068
rect 25026 82346 25082 82348
rect 25026 82294 25028 82346
rect 25028 82294 25080 82346
rect 25080 82294 25082 82346
rect 25026 82292 25082 82294
rect 25130 82346 25186 82348
rect 25130 82294 25132 82346
rect 25132 82294 25184 82346
rect 25184 82294 25186 82346
rect 25130 82292 25186 82294
rect 25234 82346 25290 82348
rect 25234 82294 25236 82346
rect 25236 82294 25288 82346
rect 25288 82294 25290 82346
rect 25234 82292 25290 82294
rect 25228 82178 25284 82180
rect 25228 82126 25230 82178
rect 25230 82126 25282 82178
rect 25282 82126 25284 82178
rect 25228 82124 25284 82126
rect 24220 81788 24276 81844
rect 23884 81282 23940 81284
rect 23884 81230 23886 81282
rect 23886 81230 23938 81282
rect 23938 81230 23940 81282
rect 23884 81228 23940 81230
rect 24780 82012 24836 82068
rect 26236 84418 26292 84420
rect 26236 84366 26238 84418
rect 26238 84366 26290 84418
rect 26290 84366 26292 84418
rect 26236 84364 26292 84366
rect 26124 84306 26180 84308
rect 26124 84254 26126 84306
rect 26126 84254 26178 84306
rect 26178 84254 26180 84306
rect 26124 84252 26180 84254
rect 24556 81788 24612 81844
rect 24668 81340 24724 81396
rect 24108 81004 24164 81060
rect 24556 80946 24612 80948
rect 24556 80894 24558 80946
rect 24558 80894 24610 80946
rect 24610 80894 24612 80946
rect 24556 80892 24612 80894
rect 24556 80610 24612 80612
rect 24556 80558 24558 80610
rect 24558 80558 24610 80610
rect 24610 80558 24612 80610
rect 24556 80556 24612 80558
rect 23436 80498 23492 80500
rect 23436 80446 23438 80498
rect 23438 80446 23490 80498
rect 23490 80446 23492 80498
rect 23436 80444 23492 80446
rect 24444 80444 24500 80500
rect 23324 80162 23380 80164
rect 23324 80110 23326 80162
rect 23326 80110 23378 80162
rect 23378 80110 23380 80162
rect 23324 80108 23380 80110
rect 23996 79772 24052 79828
rect 24556 79772 24612 79828
rect 23772 79602 23828 79604
rect 23772 79550 23774 79602
rect 23774 79550 23826 79602
rect 23826 79550 23828 79602
rect 23772 79548 23828 79550
rect 24220 79602 24276 79604
rect 24220 79550 24222 79602
rect 24222 79550 24274 79602
rect 24274 79550 24276 79602
rect 24220 79548 24276 79550
rect 23772 78818 23828 78820
rect 23772 78766 23774 78818
rect 23774 78766 23826 78818
rect 23826 78766 23828 78818
rect 23772 78764 23828 78766
rect 23324 78706 23380 78708
rect 23324 78654 23326 78706
rect 23326 78654 23378 78706
rect 23378 78654 23380 78706
rect 23324 78652 23380 78654
rect 23212 78540 23268 78596
rect 23212 77756 23268 77812
rect 24220 78540 24276 78596
rect 23660 77138 23716 77140
rect 23660 77086 23662 77138
rect 23662 77086 23714 77138
rect 23714 77086 23716 77138
rect 23660 77084 23716 77086
rect 22876 76636 22932 76692
rect 22652 76076 22708 76132
rect 22540 75740 22596 75796
rect 23772 76636 23828 76692
rect 23100 75628 23156 75684
rect 22540 74786 22596 74788
rect 22540 74734 22542 74786
rect 22542 74734 22594 74786
rect 22594 74734 22596 74786
rect 22540 74732 22596 74734
rect 22540 74172 22596 74228
rect 21868 73164 21924 73220
rect 21644 73106 21700 73108
rect 21644 73054 21646 73106
rect 21646 73054 21698 73106
rect 21698 73054 21700 73106
rect 21644 73052 21700 73054
rect 21868 72940 21924 72996
rect 22316 73052 22372 73108
rect 22428 73164 22484 73220
rect 22204 72940 22260 72996
rect 21196 72492 21252 72548
rect 21084 72268 21140 72324
rect 20860 70588 20916 70644
rect 20748 70082 20804 70084
rect 20748 70030 20750 70082
rect 20750 70030 20802 70082
rect 20802 70030 20804 70082
rect 20748 70028 20804 70030
rect 20748 69020 20804 69076
rect 20748 68850 20804 68852
rect 20748 68798 20750 68850
rect 20750 68798 20802 68850
rect 20802 68798 20804 68850
rect 20748 68796 20804 68798
rect 19516 65548 19572 65604
rect 18732 63532 18788 63588
rect 19180 64316 19236 64372
rect 19404 64204 19460 64260
rect 19628 64652 19684 64708
rect 19292 63532 19348 63588
rect 18956 63308 19012 63364
rect 18620 63026 18676 63028
rect 18620 62974 18622 63026
rect 18622 62974 18674 63026
rect 18674 62974 18676 63026
rect 18620 62972 18676 62974
rect 18396 62412 18452 62468
rect 18620 62300 18676 62356
rect 18222 61962 18278 61964
rect 18222 61910 18224 61962
rect 18224 61910 18276 61962
rect 18276 61910 18278 61962
rect 18222 61908 18278 61910
rect 18326 61962 18382 61964
rect 18326 61910 18328 61962
rect 18328 61910 18380 61962
rect 18380 61910 18382 61962
rect 18326 61908 18382 61910
rect 18430 61962 18486 61964
rect 18430 61910 18432 61962
rect 18432 61910 18484 61962
rect 18484 61910 18486 61962
rect 18430 61908 18486 61910
rect 18172 61068 18228 61124
rect 18732 60732 18788 60788
rect 18620 60508 18676 60564
rect 18222 60394 18278 60396
rect 18222 60342 18224 60394
rect 18224 60342 18276 60394
rect 18276 60342 18278 60394
rect 18222 60340 18278 60342
rect 18326 60394 18382 60396
rect 18326 60342 18328 60394
rect 18328 60342 18380 60394
rect 18380 60342 18382 60394
rect 18326 60340 18382 60342
rect 18430 60394 18486 60396
rect 18430 60342 18432 60394
rect 18432 60342 18484 60394
rect 18484 60342 18486 60394
rect 18430 60340 18486 60342
rect 18172 59948 18228 60004
rect 18508 59778 18564 59780
rect 18508 59726 18510 59778
rect 18510 59726 18562 59778
rect 18562 59726 18564 59778
rect 18508 59724 18564 59726
rect 18172 59164 18228 59220
rect 18222 58826 18278 58828
rect 18222 58774 18224 58826
rect 18224 58774 18276 58826
rect 18276 58774 18278 58826
rect 18222 58772 18278 58774
rect 18326 58826 18382 58828
rect 18326 58774 18328 58826
rect 18328 58774 18380 58826
rect 18380 58774 18382 58826
rect 18326 58772 18382 58774
rect 18430 58826 18486 58828
rect 18430 58774 18432 58826
rect 18432 58774 18484 58826
rect 18484 58774 18486 58826
rect 18430 58772 18486 58774
rect 18396 58268 18452 58324
rect 18222 57258 18278 57260
rect 18222 57206 18224 57258
rect 18224 57206 18276 57258
rect 18276 57206 18278 57258
rect 18222 57204 18278 57206
rect 18326 57258 18382 57260
rect 18326 57206 18328 57258
rect 18328 57206 18380 57258
rect 18380 57206 18382 57258
rect 18326 57204 18382 57206
rect 18430 57258 18486 57260
rect 18430 57206 18432 57258
rect 18432 57206 18484 57258
rect 18484 57206 18486 57258
rect 18430 57204 18486 57206
rect 17612 55970 17668 55972
rect 17612 55918 17614 55970
rect 17614 55918 17666 55970
rect 17666 55918 17668 55970
rect 17612 55916 17668 55918
rect 16828 52892 16884 52948
rect 17388 55468 17444 55524
rect 16716 52668 16772 52724
rect 17052 52668 17108 52724
rect 16716 51548 16772 51604
rect 16828 51660 16884 51716
rect 16492 50482 16548 50484
rect 16492 50430 16494 50482
rect 16494 50430 16546 50482
rect 16546 50430 16548 50482
rect 16492 50428 16548 50430
rect 16268 49084 16324 49140
rect 16380 49532 16436 49588
rect 15932 46620 15988 46676
rect 16268 48300 16324 48356
rect 16828 49922 16884 49924
rect 16828 49870 16830 49922
rect 16830 49870 16882 49922
rect 16882 49870 16884 49922
rect 16828 49868 16884 49870
rect 17052 48914 17108 48916
rect 17052 48862 17054 48914
rect 17054 48862 17106 48914
rect 17106 48862 17108 48914
rect 17052 48860 17108 48862
rect 16716 48636 16772 48692
rect 15708 45276 15764 45332
rect 15820 45890 15876 45892
rect 15820 45838 15822 45890
rect 15822 45838 15874 45890
rect 15874 45838 15876 45890
rect 15820 45836 15876 45838
rect 15372 44828 15428 44884
rect 14252 43932 14308 43988
rect 14820 43930 14876 43932
rect 14364 43820 14420 43876
rect 14364 43260 14420 43316
rect 14588 43820 14644 43876
rect 14820 43878 14822 43930
rect 14822 43878 14874 43930
rect 14874 43878 14876 43930
rect 14820 43876 14876 43878
rect 14924 43930 14980 43932
rect 14924 43878 14926 43930
rect 14926 43878 14978 43930
rect 14978 43878 14980 43930
rect 14924 43876 14980 43878
rect 15028 43930 15084 43932
rect 15028 43878 15030 43930
rect 15030 43878 15082 43930
rect 15082 43878 15084 43930
rect 15028 43876 15084 43878
rect 15260 43820 15316 43876
rect 14140 42530 14196 42532
rect 14140 42478 14142 42530
rect 14142 42478 14194 42530
rect 14194 42478 14196 42530
rect 14140 42476 14196 42478
rect 13804 41074 13860 41076
rect 13804 41022 13806 41074
rect 13806 41022 13858 41074
rect 13858 41022 13860 41074
rect 13804 41020 13860 41022
rect 14364 42530 14420 42532
rect 14364 42478 14366 42530
rect 14366 42478 14418 42530
rect 14418 42478 14420 42530
rect 14364 42476 14420 42478
rect 14588 41580 14644 41636
rect 14700 43484 14756 43540
rect 15036 43538 15092 43540
rect 15036 43486 15038 43538
rect 15038 43486 15090 43538
rect 15090 43486 15092 43538
rect 15036 43484 15092 43486
rect 14820 42362 14876 42364
rect 14820 42310 14822 42362
rect 14822 42310 14874 42362
rect 14874 42310 14876 42362
rect 14820 42308 14876 42310
rect 14924 42362 14980 42364
rect 14924 42310 14926 42362
rect 14926 42310 14978 42362
rect 14978 42310 14980 42362
rect 14924 42308 14980 42310
rect 15028 42362 15084 42364
rect 15028 42310 15030 42362
rect 15030 42310 15082 42362
rect 15082 42310 15084 42362
rect 15028 42308 15084 42310
rect 15260 42476 15316 42532
rect 14812 41916 14868 41972
rect 15372 41804 15428 41860
rect 14924 41580 14980 41636
rect 13580 40236 13636 40292
rect 13580 39116 13636 39172
rect 13580 38220 13636 38276
rect 13580 37490 13636 37492
rect 13580 37438 13582 37490
rect 13582 37438 13634 37490
rect 13634 37438 13636 37490
rect 13580 37436 13636 37438
rect 13580 36988 13636 37044
rect 14028 40626 14084 40628
rect 14028 40574 14030 40626
rect 14030 40574 14082 40626
rect 14082 40574 14084 40626
rect 14028 40572 14084 40574
rect 14028 39788 14084 39844
rect 14140 39618 14196 39620
rect 14140 39566 14142 39618
rect 14142 39566 14194 39618
rect 14194 39566 14196 39618
rect 14140 39564 14196 39566
rect 13916 37490 13972 37492
rect 13916 37438 13918 37490
rect 13918 37438 13970 37490
rect 13970 37438 13972 37490
rect 13916 37436 13972 37438
rect 13692 36876 13748 36932
rect 16156 45276 16212 45332
rect 16156 44044 16212 44100
rect 16156 43538 16212 43540
rect 16156 43486 16158 43538
rect 16158 43486 16210 43538
rect 16210 43486 16212 43538
rect 16156 43484 16212 43486
rect 16044 43260 16100 43316
rect 15708 42082 15764 42084
rect 15708 42030 15710 42082
rect 15710 42030 15762 42082
rect 15762 42030 15764 42082
rect 15708 42028 15764 42030
rect 15596 41468 15652 41524
rect 15372 41244 15428 41300
rect 15932 41692 15988 41748
rect 15148 40908 15204 40964
rect 14820 40794 14876 40796
rect 14820 40742 14822 40794
rect 14822 40742 14874 40794
rect 14874 40742 14876 40794
rect 14820 40740 14876 40742
rect 14924 40794 14980 40796
rect 14924 40742 14926 40794
rect 14926 40742 14978 40794
rect 14978 40742 14980 40794
rect 14924 40740 14980 40742
rect 15028 40794 15084 40796
rect 15028 40742 15030 40794
rect 15030 40742 15082 40794
rect 15082 40742 15084 40794
rect 15028 40740 15084 40742
rect 14700 39788 14756 39844
rect 16604 43708 16660 43764
rect 16380 43596 16436 43652
rect 16492 42812 16548 42868
rect 16044 41132 16100 41188
rect 16156 40236 16212 40292
rect 16828 47964 16884 48020
rect 16828 47740 16884 47796
rect 17164 47964 17220 48020
rect 17612 55244 17668 55300
rect 17388 52946 17444 52948
rect 17388 52894 17390 52946
rect 17390 52894 17442 52946
rect 17442 52894 17444 52946
rect 17388 52892 17444 52894
rect 17612 52668 17668 52724
rect 17724 54460 17780 54516
rect 17724 52444 17780 52500
rect 17612 52220 17668 52276
rect 17500 51660 17556 51716
rect 17388 49868 17444 49924
rect 17724 50428 17780 50484
rect 17388 48860 17444 48916
rect 17612 50316 17668 50372
rect 17500 48524 17556 48580
rect 17724 49868 17780 49924
rect 17724 48748 17780 48804
rect 17500 48354 17556 48356
rect 17500 48302 17502 48354
rect 17502 48302 17554 48354
rect 17554 48302 17556 48354
rect 17500 48300 17556 48302
rect 17276 47740 17332 47796
rect 17612 47964 17668 48020
rect 17052 45948 17108 46004
rect 17276 47012 17332 47068
rect 16940 44380 16996 44436
rect 16828 42252 16884 42308
rect 16716 41020 16772 41076
rect 16828 42028 16884 42084
rect 16716 40684 16772 40740
rect 16380 40124 16436 40180
rect 16380 39788 16436 39844
rect 15148 39618 15204 39620
rect 15148 39566 15150 39618
rect 15150 39566 15202 39618
rect 15202 39566 15204 39618
rect 15148 39564 15204 39566
rect 14924 39506 14980 39508
rect 14924 39454 14926 39506
rect 14926 39454 14978 39506
rect 14978 39454 14980 39506
rect 14924 39452 14980 39454
rect 15484 39506 15540 39508
rect 15484 39454 15486 39506
rect 15486 39454 15538 39506
rect 15538 39454 15540 39506
rect 15484 39452 15540 39454
rect 14820 39226 14876 39228
rect 14820 39174 14822 39226
rect 14822 39174 14874 39226
rect 14874 39174 14876 39226
rect 14820 39172 14876 39174
rect 14924 39226 14980 39228
rect 14924 39174 14926 39226
rect 14926 39174 14978 39226
rect 14978 39174 14980 39226
rect 14924 39172 14980 39174
rect 15028 39226 15084 39228
rect 15028 39174 15030 39226
rect 15030 39174 15082 39226
rect 15082 39174 15084 39226
rect 15028 39172 15084 39174
rect 16044 39228 16100 39284
rect 15372 39004 15428 39060
rect 14820 37658 14876 37660
rect 14820 37606 14822 37658
rect 14822 37606 14874 37658
rect 14874 37606 14876 37658
rect 14820 37604 14876 37606
rect 14924 37658 14980 37660
rect 14924 37606 14926 37658
rect 14926 37606 14978 37658
rect 14978 37606 14980 37658
rect 14924 37604 14980 37606
rect 15028 37658 15084 37660
rect 15028 37606 15030 37658
rect 15030 37606 15082 37658
rect 15082 37606 15084 37658
rect 15028 37604 15084 37606
rect 14364 37436 14420 37492
rect 14028 36652 14084 36708
rect 13692 36482 13748 36484
rect 13692 36430 13694 36482
rect 13694 36430 13746 36482
rect 13746 36430 13748 36482
rect 13692 36428 13748 36430
rect 13468 36370 13524 36372
rect 13468 36318 13470 36370
rect 13470 36318 13522 36370
rect 13522 36318 13524 36370
rect 13468 36316 13524 36318
rect 13356 35756 13412 35812
rect 13916 36482 13972 36484
rect 13916 36430 13918 36482
rect 13918 36430 13970 36482
rect 13970 36430 13972 36482
rect 13916 36428 13972 36430
rect 15260 37490 15316 37492
rect 15260 37438 15262 37490
rect 15262 37438 15314 37490
rect 15314 37438 15316 37490
rect 15260 37436 15316 37438
rect 14364 36706 14420 36708
rect 14364 36654 14366 36706
rect 14366 36654 14418 36706
rect 14418 36654 14420 36706
rect 14364 36652 14420 36654
rect 14588 37266 14644 37268
rect 14588 37214 14590 37266
rect 14590 37214 14642 37266
rect 14642 37214 14644 37266
rect 14588 37212 14644 37214
rect 15036 37266 15092 37268
rect 15036 37214 15038 37266
rect 15038 37214 15090 37266
rect 15090 37214 15092 37266
rect 15036 37212 15092 37214
rect 15148 36764 15204 36820
rect 13804 36316 13860 36372
rect 13132 27356 13188 27412
rect 13244 33516 13300 33572
rect 12460 26348 12516 26404
rect 12348 24780 12404 24836
rect 12460 25228 12516 25284
rect 13132 26124 13188 26180
rect 12796 25564 12852 25620
rect 12908 26012 12964 26068
rect 13468 32956 13524 33012
rect 14140 35586 14196 35588
rect 14140 35534 14142 35586
rect 14142 35534 14194 35586
rect 14194 35534 14196 35586
rect 14140 35532 14196 35534
rect 13916 34860 13972 34916
rect 14140 33964 14196 34020
rect 13468 31948 13524 32004
rect 13468 31612 13524 31668
rect 14700 36482 14756 36484
rect 14700 36430 14702 36482
rect 14702 36430 14754 36482
rect 14754 36430 14756 36482
rect 14700 36428 14756 36430
rect 15932 38050 15988 38052
rect 15932 37998 15934 38050
rect 15934 37998 15986 38050
rect 15986 37998 15988 38050
rect 15932 37996 15988 37998
rect 15932 37548 15988 37604
rect 17164 45276 17220 45332
rect 16492 38162 16548 38164
rect 16492 38110 16494 38162
rect 16494 38110 16546 38162
rect 16546 38110 16548 38162
rect 16492 38108 16548 38110
rect 16044 37884 16100 37940
rect 15596 37154 15652 37156
rect 15596 37102 15598 37154
rect 15598 37102 15650 37154
rect 15650 37102 15652 37154
rect 15596 37100 15652 37102
rect 15484 36988 15540 37044
rect 15372 36258 15428 36260
rect 15372 36206 15374 36258
rect 15374 36206 15426 36258
rect 15426 36206 15428 36258
rect 15372 36204 15428 36206
rect 14820 36090 14876 36092
rect 14820 36038 14822 36090
rect 14822 36038 14874 36090
rect 14874 36038 14876 36090
rect 14820 36036 14876 36038
rect 14924 36090 14980 36092
rect 14924 36038 14926 36090
rect 14926 36038 14978 36090
rect 14978 36038 14980 36090
rect 14924 36036 14980 36038
rect 15028 36090 15084 36092
rect 15028 36038 15030 36090
rect 15030 36038 15082 36090
rect 15082 36038 15084 36090
rect 15028 36036 15084 36038
rect 15260 35868 15316 35924
rect 14364 35308 14420 35364
rect 14812 35532 14868 35588
rect 14588 35252 14644 35308
rect 14924 34972 14980 35028
rect 14364 33180 14420 33236
rect 14700 34914 14756 34916
rect 14700 34862 14702 34914
rect 14702 34862 14754 34914
rect 14754 34862 14756 34914
rect 14700 34860 14756 34862
rect 13356 29036 13412 29092
rect 13356 28700 13412 28756
rect 13356 28364 13412 28420
rect 14140 30940 14196 30996
rect 14252 30828 14308 30884
rect 14252 30268 14308 30324
rect 13916 28700 13972 28756
rect 14028 29036 14084 29092
rect 14140 28812 14196 28868
rect 14252 28924 14308 28980
rect 14140 28642 14196 28644
rect 14140 28590 14142 28642
rect 14142 28590 14194 28642
rect 14194 28590 14196 28642
rect 14140 28588 14196 28590
rect 13692 28530 13748 28532
rect 13692 28478 13694 28530
rect 13694 28478 13746 28530
rect 13746 28478 13748 28530
rect 13692 28476 13748 28478
rect 13356 27468 13412 27524
rect 13692 27468 13748 27524
rect 13580 27074 13636 27076
rect 13580 27022 13582 27074
rect 13582 27022 13634 27074
rect 13634 27022 13636 27074
rect 13580 27020 13636 27022
rect 13692 26796 13748 26852
rect 13356 26012 13412 26068
rect 12796 24220 12852 24276
rect 12236 22988 12292 23044
rect 12460 22876 12516 22932
rect 12348 21756 12404 21812
rect 12460 21474 12516 21476
rect 12460 21422 12462 21474
rect 12462 21422 12514 21474
rect 12514 21422 12516 21474
rect 12460 21420 12516 21422
rect 12460 20636 12516 20692
rect 12460 19964 12516 20020
rect 12460 19740 12516 19796
rect 12460 19180 12516 19236
rect 12348 18396 12404 18452
rect 12012 17388 12068 17444
rect 12796 23772 12852 23828
rect 12684 23548 12740 23604
rect 12908 23548 12964 23604
rect 13020 23660 13076 23716
rect 13020 23324 13076 23380
rect 12684 22316 12740 22372
rect 12908 21810 12964 21812
rect 12908 21758 12910 21810
rect 12910 21758 12962 21810
rect 12962 21758 12964 21810
rect 12908 21756 12964 21758
rect 13356 25564 13412 25620
rect 13244 23660 13300 23716
rect 13468 24220 13524 24276
rect 13356 22988 13412 23044
rect 14028 27804 14084 27860
rect 14252 28140 14308 28196
rect 14364 27468 14420 27524
rect 14140 26796 14196 26852
rect 14364 26460 14420 26516
rect 13804 25618 13860 25620
rect 13804 25566 13806 25618
rect 13806 25566 13858 25618
rect 13858 25566 13860 25618
rect 13804 25564 13860 25566
rect 14820 34522 14876 34524
rect 14820 34470 14822 34522
rect 14822 34470 14874 34522
rect 14874 34470 14876 34522
rect 14820 34468 14876 34470
rect 14924 34522 14980 34524
rect 14924 34470 14926 34522
rect 14926 34470 14978 34522
rect 14978 34470 14980 34522
rect 14924 34468 14980 34470
rect 15028 34522 15084 34524
rect 15028 34470 15030 34522
rect 15030 34470 15082 34522
rect 15082 34470 15084 34522
rect 15028 34468 15084 34470
rect 14588 33292 14644 33348
rect 14588 31164 14644 31220
rect 14588 30994 14644 30996
rect 14588 30942 14590 30994
rect 14590 30942 14642 30994
rect 14642 30942 14644 30994
rect 14588 30940 14644 30942
rect 15484 35756 15540 35812
rect 16044 36764 16100 36820
rect 15708 36652 15764 36708
rect 16156 36428 16212 36484
rect 15708 36204 15764 36260
rect 14812 33234 14868 33236
rect 14812 33182 14814 33234
rect 14814 33182 14866 33234
rect 14866 33182 14868 33234
rect 14812 33180 14868 33182
rect 14820 32954 14876 32956
rect 14820 32902 14822 32954
rect 14822 32902 14874 32954
rect 14874 32902 14876 32954
rect 14820 32900 14876 32902
rect 14924 32954 14980 32956
rect 14924 32902 14926 32954
rect 14926 32902 14978 32954
rect 14978 32902 14980 32954
rect 14924 32900 14980 32902
rect 15028 32954 15084 32956
rect 15028 32902 15030 32954
rect 15030 32902 15082 32954
rect 15082 32902 15084 32954
rect 15028 32900 15084 32902
rect 15148 32396 15204 32452
rect 15708 35420 15764 35476
rect 16044 35868 16100 35924
rect 16044 35644 16100 35700
rect 14820 31386 14876 31388
rect 14820 31334 14822 31386
rect 14822 31334 14874 31386
rect 14874 31334 14876 31386
rect 14820 31332 14876 31334
rect 14924 31386 14980 31388
rect 14924 31334 14926 31386
rect 14926 31334 14978 31386
rect 14978 31334 14980 31386
rect 14924 31332 14980 31334
rect 15028 31386 15084 31388
rect 15028 31334 15030 31386
rect 15030 31334 15082 31386
rect 15082 31334 15084 31386
rect 15028 31332 15084 31334
rect 14812 31164 14868 31220
rect 15596 34860 15652 34916
rect 15372 34018 15428 34020
rect 15372 33966 15374 34018
rect 15374 33966 15426 34018
rect 15426 33966 15428 34018
rect 15372 33964 15428 33966
rect 15932 33292 15988 33348
rect 15596 33234 15652 33236
rect 15596 33182 15598 33234
rect 15598 33182 15650 33234
rect 15650 33182 15652 33234
rect 15596 33180 15652 33182
rect 15820 32450 15876 32452
rect 15820 32398 15822 32450
rect 15822 32398 15874 32450
rect 15874 32398 15876 32450
rect 15820 32396 15876 32398
rect 16492 36482 16548 36484
rect 16492 36430 16494 36482
rect 16494 36430 16546 36482
rect 16546 36430 16548 36482
rect 16492 36428 16548 36430
rect 16604 36370 16660 36372
rect 16604 36318 16606 36370
rect 16606 36318 16658 36370
rect 16658 36318 16660 36370
rect 16604 36316 16660 36318
rect 16268 36258 16324 36260
rect 16268 36206 16270 36258
rect 16270 36206 16322 36258
rect 16322 36206 16324 36258
rect 16268 36204 16324 36206
rect 16940 39004 16996 39060
rect 16828 38722 16884 38724
rect 16828 38670 16830 38722
rect 16830 38670 16882 38722
rect 16882 38670 16884 38722
rect 16828 38668 16884 38670
rect 16380 35420 16436 35476
rect 16828 38108 16884 38164
rect 16380 35138 16436 35140
rect 16380 35086 16382 35138
rect 16382 35086 16434 35138
rect 16434 35086 16436 35138
rect 16380 35084 16436 35086
rect 17388 45836 17444 45892
rect 17500 45724 17556 45780
rect 17948 56082 18004 56084
rect 17948 56030 17950 56082
rect 17950 56030 18002 56082
rect 18002 56030 18004 56082
rect 17948 56028 18004 56030
rect 17948 53058 18004 53060
rect 17948 53006 17950 53058
rect 17950 53006 18002 53058
rect 18002 53006 18004 53058
rect 17948 53004 18004 53006
rect 17948 52556 18004 52612
rect 17948 49756 18004 49812
rect 18284 56082 18340 56084
rect 18284 56030 18286 56082
rect 18286 56030 18338 56082
rect 18338 56030 18340 56082
rect 18284 56028 18340 56030
rect 18172 55916 18228 55972
rect 18222 55690 18278 55692
rect 18222 55638 18224 55690
rect 18224 55638 18276 55690
rect 18276 55638 18278 55690
rect 18222 55636 18278 55638
rect 18326 55690 18382 55692
rect 18326 55638 18328 55690
rect 18328 55638 18380 55690
rect 18380 55638 18382 55690
rect 18326 55636 18382 55638
rect 18430 55690 18486 55692
rect 18430 55638 18432 55690
rect 18432 55638 18484 55690
rect 18484 55638 18486 55690
rect 18430 55636 18486 55638
rect 18222 54122 18278 54124
rect 18222 54070 18224 54122
rect 18224 54070 18276 54122
rect 18276 54070 18278 54122
rect 18222 54068 18278 54070
rect 18326 54122 18382 54124
rect 18326 54070 18328 54122
rect 18328 54070 18380 54122
rect 18380 54070 18382 54122
rect 18326 54068 18382 54070
rect 18430 54122 18486 54124
rect 18430 54070 18432 54122
rect 18432 54070 18484 54122
rect 18484 54070 18486 54122
rect 18430 54068 18486 54070
rect 18396 53730 18452 53732
rect 18396 53678 18398 53730
rect 18398 53678 18450 53730
rect 18450 53678 18452 53730
rect 18396 53676 18452 53678
rect 18508 53618 18564 53620
rect 18508 53566 18510 53618
rect 18510 53566 18562 53618
rect 18562 53566 18564 53618
rect 18508 53564 18564 53566
rect 18396 53228 18452 53284
rect 18620 52892 18676 52948
rect 18620 52668 18676 52724
rect 18222 52554 18278 52556
rect 18222 52502 18224 52554
rect 18224 52502 18276 52554
rect 18276 52502 18278 52554
rect 18222 52500 18278 52502
rect 18326 52554 18382 52556
rect 18326 52502 18328 52554
rect 18328 52502 18380 52554
rect 18380 52502 18382 52554
rect 18326 52500 18382 52502
rect 18430 52554 18486 52556
rect 18430 52502 18432 52554
rect 18432 52502 18484 52554
rect 18484 52502 18486 52554
rect 18430 52500 18486 52502
rect 18172 52050 18228 52052
rect 18172 51998 18174 52050
rect 18174 51998 18226 52050
rect 18226 51998 18228 52050
rect 18172 51996 18228 51998
rect 18396 51884 18452 51940
rect 18732 51884 18788 51940
rect 18732 51490 18788 51492
rect 18732 51438 18734 51490
rect 18734 51438 18786 51490
rect 18786 51438 18788 51490
rect 18732 51436 18788 51438
rect 18172 51100 18228 51156
rect 18222 50986 18278 50988
rect 18222 50934 18224 50986
rect 18224 50934 18276 50986
rect 18276 50934 18278 50986
rect 18222 50932 18278 50934
rect 18326 50986 18382 50988
rect 18326 50934 18328 50986
rect 18328 50934 18380 50986
rect 18380 50934 18382 50986
rect 18326 50932 18382 50934
rect 18430 50986 18486 50988
rect 18430 50934 18432 50986
rect 18432 50934 18484 50986
rect 18484 50934 18486 50986
rect 18430 50932 18486 50934
rect 18508 50764 18564 50820
rect 19180 63138 19236 63140
rect 19180 63086 19182 63138
rect 19182 63086 19234 63138
rect 19234 63086 19236 63138
rect 19180 63084 19236 63086
rect 19292 62578 19348 62580
rect 19292 62526 19294 62578
rect 19294 62526 19346 62578
rect 19346 62526 19348 62578
rect 19292 62524 19348 62526
rect 19180 62412 19236 62468
rect 19628 63138 19684 63140
rect 19628 63086 19630 63138
rect 19630 63086 19682 63138
rect 19682 63086 19684 63138
rect 19628 63084 19684 63086
rect 19964 65548 20020 65604
rect 19964 64594 20020 64596
rect 19964 64542 19966 64594
rect 19966 64542 20018 64594
rect 20018 64542 20020 64594
rect 19964 64540 20020 64542
rect 20300 64876 20356 64932
rect 19180 59890 19236 59892
rect 19180 59838 19182 59890
rect 19182 59838 19234 59890
rect 19234 59838 19236 59890
rect 19180 59836 19236 59838
rect 18956 59276 19012 59332
rect 19180 59612 19236 59668
rect 19180 57148 19236 57204
rect 19516 61964 19572 62020
rect 19516 61404 19572 61460
rect 19404 60898 19460 60900
rect 19404 60846 19406 60898
rect 19406 60846 19458 60898
rect 19458 60846 19460 60898
rect 19404 60844 19460 60846
rect 19628 60732 19684 60788
rect 19740 62636 19796 62692
rect 20524 65996 20580 66052
rect 20524 64706 20580 64708
rect 20524 64654 20526 64706
rect 20526 64654 20578 64706
rect 20578 64654 20580 64706
rect 20524 64652 20580 64654
rect 20524 63756 20580 63812
rect 20748 66556 20804 66612
rect 20748 66050 20804 66052
rect 20748 65998 20750 66050
rect 20750 65998 20802 66050
rect 20802 65998 20804 66050
rect 20748 65996 20804 65998
rect 21868 72434 21924 72436
rect 21868 72382 21870 72434
rect 21870 72382 21922 72434
rect 21922 72382 21924 72434
rect 21868 72380 21924 72382
rect 22092 72268 22148 72324
rect 21624 72154 21680 72156
rect 21624 72102 21626 72154
rect 21626 72102 21678 72154
rect 21678 72102 21680 72154
rect 21624 72100 21680 72102
rect 21728 72154 21784 72156
rect 21728 72102 21730 72154
rect 21730 72102 21782 72154
rect 21782 72102 21784 72154
rect 21728 72100 21784 72102
rect 21832 72154 21888 72156
rect 21832 72102 21834 72154
rect 21834 72102 21886 72154
rect 21886 72102 21888 72154
rect 21832 72100 21888 72102
rect 21980 72156 22036 72212
rect 21532 71932 21588 71988
rect 21420 71484 21476 71540
rect 21308 70418 21364 70420
rect 21308 70366 21310 70418
rect 21310 70366 21362 70418
rect 21362 70366 21364 70418
rect 21308 70364 21364 70366
rect 21084 66892 21140 66948
rect 21532 70978 21588 70980
rect 21532 70926 21534 70978
rect 21534 70926 21586 70978
rect 21586 70926 21588 70978
rect 21532 70924 21588 70926
rect 22540 72492 22596 72548
rect 22316 72044 22372 72100
rect 22764 73724 22820 73780
rect 23548 76354 23604 76356
rect 23548 76302 23550 76354
rect 23550 76302 23602 76354
rect 23602 76302 23604 76354
rect 23548 76300 23604 76302
rect 23548 74396 23604 74452
rect 23660 75516 23716 75572
rect 23884 75852 23940 75908
rect 24108 74956 24164 75012
rect 24444 77868 24500 77924
rect 24332 77138 24388 77140
rect 24332 77086 24334 77138
rect 24334 77086 24386 77138
rect 24386 77086 24388 77138
rect 24332 77084 24388 77086
rect 25228 81058 25284 81060
rect 25228 81006 25230 81058
rect 25230 81006 25282 81058
rect 25282 81006 25284 81058
rect 25228 81004 25284 81006
rect 25452 80946 25508 80948
rect 25452 80894 25454 80946
rect 25454 80894 25506 80946
rect 25506 80894 25508 80946
rect 25452 80892 25508 80894
rect 25026 80778 25082 80780
rect 25026 80726 25028 80778
rect 25028 80726 25080 80778
rect 25080 80726 25082 80778
rect 25026 80724 25082 80726
rect 25130 80778 25186 80780
rect 25130 80726 25132 80778
rect 25132 80726 25184 80778
rect 25184 80726 25186 80778
rect 25130 80724 25186 80726
rect 25234 80778 25290 80780
rect 25234 80726 25236 80778
rect 25236 80726 25288 80778
rect 25288 80726 25290 80778
rect 25234 80724 25290 80726
rect 24780 80332 24836 80388
rect 25788 82124 25844 82180
rect 25788 81004 25844 81060
rect 26348 84252 26404 84308
rect 26572 84924 26628 84980
rect 27132 88060 27188 88116
rect 26908 87218 26964 87220
rect 26908 87166 26910 87218
rect 26910 87166 26962 87218
rect 26962 87166 26964 87218
rect 26908 87164 26964 87166
rect 26796 87052 26852 87108
rect 28428 89402 28484 89404
rect 28428 89350 28430 89402
rect 28430 89350 28482 89402
rect 28482 89350 28484 89402
rect 28428 89348 28484 89350
rect 28532 89402 28588 89404
rect 28532 89350 28534 89402
rect 28534 89350 28586 89402
rect 28586 89350 28588 89402
rect 28532 89348 28588 89350
rect 28636 89402 28692 89404
rect 28636 89350 28638 89402
rect 28638 89350 28690 89402
rect 28690 89350 28692 89402
rect 28636 89348 28692 89350
rect 27580 88172 27636 88228
rect 28428 87834 28484 87836
rect 28428 87782 28430 87834
rect 28430 87782 28482 87834
rect 28482 87782 28484 87834
rect 28428 87780 28484 87782
rect 28532 87834 28588 87836
rect 28532 87782 28534 87834
rect 28534 87782 28586 87834
rect 28586 87782 28588 87834
rect 28532 87780 28588 87782
rect 28636 87834 28692 87836
rect 28636 87782 28638 87834
rect 28638 87782 28690 87834
rect 28690 87782 28692 87834
rect 28636 87780 28692 87782
rect 27244 86658 27300 86660
rect 27244 86606 27246 86658
rect 27246 86606 27298 86658
rect 27298 86606 27300 86658
rect 27244 86604 27300 86606
rect 26796 85484 26852 85540
rect 27468 87330 27524 87332
rect 27468 87278 27470 87330
rect 27470 87278 27522 87330
rect 27522 87278 27524 87330
rect 27468 87276 27524 87278
rect 27692 86716 27748 86772
rect 27468 85650 27524 85652
rect 27468 85598 27470 85650
rect 27470 85598 27522 85650
rect 27522 85598 27524 85650
rect 27468 85596 27524 85598
rect 27356 85484 27412 85540
rect 26908 84588 26964 84644
rect 27692 85484 27748 85540
rect 27692 84866 27748 84868
rect 27692 84814 27694 84866
rect 27694 84814 27746 84866
rect 27746 84814 27748 84866
rect 27692 84812 27748 84814
rect 27132 84364 27188 84420
rect 26460 84028 26516 84084
rect 26236 82850 26292 82852
rect 26236 82798 26238 82850
rect 26238 82798 26290 82850
rect 26290 82798 26292 82850
rect 26236 82796 26292 82798
rect 26124 82738 26180 82740
rect 26124 82686 26126 82738
rect 26126 82686 26178 82738
rect 26178 82686 26180 82738
rect 26124 82684 26180 82686
rect 26236 82124 26292 82180
rect 26348 81900 26404 81956
rect 27580 84306 27636 84308
rect 27580 84254 27582 84306
rect 27582 84254 27634 84306
rect 27634 84254 27636 84306
rect 27580 84252 27636 84254
rect 26684 83916 26740 83972
rect 26572 81900 26628 81956
rect 26460 81116 26516 81172
rect 26348 81004 26404 81060
rect 25228 80556 25284 80612
rect 26236 80892 26292 80948
rect 25564 80386 25620 80388
rect 25564 80334 25566 80386
rect 25566 80334 25618 80386
rect 25618 80334 25620 80386
rect 25564 80332 25620 80334
rect 26572 80892 26628 80948
rect 26460 80556 26516 80612
rect 26572 80668 26628 80724
rect 26684 80108 26740 80164
rect 26908 82236 26964 82292
rect 27244 82738 27300 82740
rect 27244 82686 27246 82738
rect 27246 82686 27298 82738
rect 27298 82686 27300 82738
rect 27244 82684 27300 82686
rect 27244 82124 27300 82180
rect 27020 81228 27076 81284
rect 27132 81170 27188 81172
rect 27132 81118 27134 81170
rect 27134 81118 27186 81170
rect 27186 81118 27188 81170
rect 27132 81116 27188 81118
rect 26908 80668 26964 80724
rect 27468 82236 27524 82292
rect 28428 86266 28484 86268
rect 28428 86214 28430 86266
rect 28430 86214 28482 86266
rect 28482 86214 28484 86266
rect 28428 86212 28484 86214
rect 28532 86266 28588 86268
rect 28532 86214 28534 86266
rect 28534 86214 28586 86266
rect 28586 86214 28588 86266
rect 28532 86212 28588 86214
rect 28636 86266 28692 86268
rect 28636 86214 28638 86266
rect 28638 86214 28690 86266
rect 28690 86214 28692 86266
rect 28636 86212 28692 86214
rect 28140 85148 28196 85204
rect 27916 84978 27972 84980
rect 27916 84926 27918 84978
rect 27918 84926 27970 84978
rect 27970 84926 27972 84978
rect 27916 84924 27972 84926
rect 28428 84698 28484 84700
rect 28140 84588 28196 84644
rect 28428 84646 28430 84698
rect 28430 84646 28482 84698
rect 28482 84646 28484 84698
rect 28428 84644 28484 84646
rect 28532 84698 28588 84700
rect 28532 84646 28534 84698
rect 28534 84646 28586 84698
rect 28586 84646 28588 84698
rect 28532 84644 28588 84646
rect 28636 84698 28692 84700
rect 28636 84646 28638 84698
rect 28638 84646 28690 84698
rect 28690 84646 28692 84698
rect 28636 84644 28692 84646
rect 28028 82796 28084 82852
rect 27468 81954 27524 81956
rect 27468 81902 27470 81954
rect 27470 81902 27522 81954
rect 27522 81902 27524 81954
rect 27468 81900 27524 81902
rect 27356 81116 27412 81172
rect 27468 80780 27524 80836
rect 27020 80498 27076 80500
rect 27020 80446 27022 80498
rect 27022 80446 27074 80498
rect 27074 80446 27076 80498
rect 27020 80444 27076 80446
rect 26236 79826 26292 79828
rect 26236 79774 26238 79826
rect 26238 79774 26290 79826
rect 26290 79774 26292 79826
rect 26236 79772 26292 79774
rect 27132 79996 27188 80052
rect 25004 79548 25060 79604
rect 25026 79210 25082 79212
rect 25026 79158 25028 79210
rect 25028 79158 25080 79210
rect 25080 79158 25082 79210
rect 25026 79156 25082 79158
rect 25130 79210 25186 79212
rect 25130 79158 25132 79210
rect 25132 79158 25184 79210
rect 25184 79158 25186 79210
rect 25130 79156 25186 79158
rect 25234 79210 25290 79212
rect 25234 79158 25236 79210
rect 25236 79158 25288 79210
rect 25288 79158 25290 79210
rect 25234 79156 25290 79158
rect 24668 77756 24724 77812
rect 25116 78594 25172 78596
rect 25116 78542 25118 78594
rect 25118 78542 25170 78594
rect 25170 78542 25172 78594
rect 25116 78540 25172 78542
rect 25026 77642 25082 77644
rect 25026 77590 25028 77642
rect 25028 77590 25080 77642
rect 25080 77590 25082 77642
rect 25026 77588 25082 77590
rect 25130 77642 25186 77644
rect 25130 77590 25132 77642
rect 25132 77590 25184 77642
rect 25184 77590 25186 77642
rect 25130 77588 25186 77590
rect 25234 77642 25290 77644
rect 25234 77590 25236 77642
rect 25236 77590 25288 77642
rect 25288 77590 25290 77642
rect 25234 77588 25290 77590
rect 25788 79602 25844 79604
rect 25788 79550 25790 79602
rect 25790 79550 25842 79602
rect 25842 79550 25844 79602
rect 25788 79548 25844 79550
rect 25564 78876 25620 78932
rect 28028 80780 28084 80836
rect 28428 83130 28484 83132
rect 28428 83078 28430 83130
rect 28430 83078 28482 83130
rect 28482 83078 28484 83130
rect 28428 83076 28484 83078
rect 28532 83130 28588 83132
rect 28532 83078 28534 83130
rect 28534 83078 28586 83130
rect 28586 83078 28588 83130
rect 28532 83076 28588 83078
rect 28636 83130 28692 83132
rect 28636 83078 28638 83130
rect 28638 83078 28690 83130
rect 28690 83078 28692 83130
rect 28636 83076 28692 83078
rect 28428 81562 28484 81564
rect 28428 81510 28430 81562
rect 28430 81510 28482 81562
rect 28482 81510 28484 81562
rect 28428 81508 28484 81510
rect 28532 81562 28588 81564
rect 28532 81510 28534 81562
rect 28534 81510 28586 81562
rect 28586 81510 28588 81562
rect 28532 81508 28588 81510
rect 28636 81562 28692 81564
rect 28636 81510 28638 81562
rect 28638 81510 28690 81562
rect 28690 81510 28692 81562
rect 28636 81508 28692 81510
rect 27916 79772 27972 79828
rect 28428 79994 28484 79996
rect 28428 79942 28430 79994
rect 28430 79942 28482 79994
rect 28482 79942 28484 79994
rect 28428 79940 28484 79942
rect 28532 79994 28588 79996
rect 28532 79942 28534 79994
rect 28534 79942 28586 79994
rect 28586 79942 28588 79994
rect 28532 79940 28588 79942
rect 28636 79994 28692 79996
rect 28636 79942 28638 79994
rect 28638 79942 28690 79994
rect 28690 79942 28692 79994
rect 28636 79940 28692 79942
rect 24780 77196 24836 77252
rect 24668 76972 24724 77028
rect 24892 76636 24948 76692
rect 25340 76748 25396 76804
rect 25026 76074 25082 76076
rect 25026 76022 25028 76074
rect 25028 76022 25080 76074
rect 25080 76022 25082 76074
rect 25026 76020 25082 76022
rect 25130 76074 25186 76076
rect 25130 76022 25132 76074
rect 25132 76022 25184 76074
rect 25184 76022 25186 76074
rect 25130 76020 25186 76022
rect 25234 76074 25290 76076
rect 25234 76022 25236 76074
rect 25236 76022 25288 76074
rect 25288 76022 25290 76074
rect 25234 76020 25290 76022
rect 24556 75852 24612 75908
rect 24780 75740 24836 75796
rect 24220 74226 24276 74228
rect 24220 74174 24222 74226
rect 24222 74174 24274 74226
rect 24274 74174 24276 74226
rect 24220 74172 24276 74174
rect 23212 73836 23268 73892
rect 22988 73388 23044 73444
rect 22988 73218 23044 73220
rect 22988 73166 22990 73218
rect 22990 73166 23042 73218
rect 23042 73166 23044 73218
rect 22988 73164 23044 73166
rect 22764 72940 22820 72996
rect 23212 73052 23268 73108
rect 22988 72546 23044 72548
rect 22988 72494 22990 72546
rect 22990 72494 23042 72546
rect 23042 72494 23044 72546
rect 22988 72492 23044 72494
rect 23212 72546 23268 72548
rect 23212 72494 23214 72546
rect 23214 72494 23266 72546
rect 23266 72494 23268 72546
rect 23212 72492 23268 72494
rect 23660 73836 23716 73892
rect 23884 73836 23940 73892
rect 23548 73612 23604 73668
rect 23660 73500 23716 73556
rect 23436 72716 23492 72772
rect 23548 73276 23604 73332
rect 22540 71484 22596 71540
rect 21624 70586 21680 70588
rect 21624 70534 21626 70586
rect 21626 70534 21678 70586
rect 21678 70534 21680 70586
rect 21624 70532 21680 70534
rect 21728 70586 21784 70588
rect 21728 70534 21730 70586
rect 21730 70534 21782 70586
rect 21782 70534 21784 70586
rect 21728 70532 21784 70534
rect 21832 70586 21888 70588
rect 21832 70534 21834 70586
rect 21834 70534 21886 70586
rect 21886 70534 21888 70586
rect 21980 70588 22036 70644
rect 21832 70532 21888 70534
rect 21644 70364 21700 70420
rect 21756 70082 21812 70084
rect 21756 70030 21758 70082
rect 21758 70030 21810 70082
rect 21810 70030 21812 70082
rect 21756 70028 21812 70030
rect 21624 69018 21680 69020
rect 21624 68966 21626 69018
rect 21626 68966 21678 69018
rect 21678 68966 21680 69018
rect 21624 68964 21680 68966
rect 21728 69018 21784 69020
rect 21728 68966 21730 69018
rect 21730 68966 21782 69018
rect 21782 68966 21784 69018
rect 21728 68964 21784 68966
rect 21832 69018 21888 69020
rect 21832 68966 21834 69018
rect 21834 68966 21886 69018
rect 21886 68966 21888 69018
rect 21832 68964 21888 68966
rect 21756 68514 21812 68516
rect 21756 68462 21758 68514
rect 21758 68462 21810 68514
rect 21810 68462 21812 68514
rect 21756 68460 21812 68462
rect 21420 68124 21476 68180
rect 21868 67842 21924 67844
rect 21868 67790 21870 67842
rect 21870 67790 21922 67842
rect 21922 67790 21924 67842
rect 21868 67788 21924 67790
rect 21532 67730 21588 67732
rect 21532 67678 21534 67730
rect 21534 67678 21586 67730
rect 21586 67678 21588 67730
rect 21532 67676 21588 67678
rect 22204 67676 22260 67732
rect 21624 67450 21680 67452
rect 21624 67398 21626 67450
rect 21626 67398 21678 67450
rect 21678 67398 21680 67450
rect 21624 67396 21680 67398
rect 21728 67450 21784 67452
rect 21728 67398 21730 67450
rect 21730 67398 21782 67450
rect 21782 67398 21784 67450
rect 21728 67396 21784 67398
rect 21832 67450 21888 67452
rect 21832 67398 21834 67450
rect 21834 67398 21886 67450
rect 21886 67398 21888 67450
rect 21832 67396 21888 67398
rect 21196 66556 21252 66612
rect 21084 66220 21140 66276
rect 20748 64540 20804 64596
rect 20748 64204 20804 64260
rect 20748 63644 20804 63700
rect 20076 63138 20132 63140
rect 20076 63086 20078 63138
rect 20078 63086 20130 63138
rect 20130 63086 20132 63138
rect 20076 63084 20132 63086
rect 19628 60562 19684 60564
rect 19628 60510 19630 60562
rect 19630 60510 19682 60562
rect 19682 60510 19684 60562
rect 19628 60508 19684 60510
rect 19516 60284 19572 60340
rect 20636 62578 20692 62580
rect 20636 62526 20638 62578
rect 20638 62526 20690 62578
rect 20690 62526 20692 62578
rect 20636 62524 20692 62526
rect 20972 64428 21028 64484
rect 21308 65660 21364 65716
rect 21532 65996 21588 66052
rect 21624 65882 21680 65884
rect 21624 65830 21626 65882
rect 21626 65830 21678 65882
rect 21678 65830 21680 65882
rect 21624 65828 21680 65830
rect 21728 65882 21784 65884
rect 21728 65830 21730 65882
rect 21730 65830 21782 65882
rect 21782 65830 21784 65882
rect 21728 65828 21784 65830
rect 21832 65882 21888 65884
rect 21832 65830 21834 65882
rect 21834 65830 21886 65882
rect 21886 65830 21888 65882
rect 21832 65828 21888 65830
rect 20972 63644 21028 63700
rect 20412 61180 20468 61236
rect 20188 60844 20244 60900
rect 19964 60732 20020 60788
rect 19516 58828 19572 58884
rect 19404 57708 19460 57764
rect 19068 56642 19124 56644
rect 19068 56590 19070 56642
rect 19070 56590 19122 56642
rect 19122 56590 19124 56642
rect 19068 56588 19124 56590
rect 18956 56028 19012 56084
rect 19068 56364 19124 56420
rect 19292 56028 19348 56084
rect 19180 54796 19236 54852
rect 18956 53506 19012 53508
rect 18956 53454 18958 53506
rect 18958 53454 19010 53506
rect 19010 53454 19012 53506
rect 18956 53452 19012 53454
rect 19180 53452 19236 53508
rect 19180 51996 19236 52052
rect 19068 51772 19124 51828
rect 19516 56754 19572 56756
rect 19516 56702 19518 56754
rect 19518 56702 19570 56754
rect 19570 56702 19572 56754
rect 19516 56700 19572 56702
rect 20300 60562 20356 60564
rect 20300 60510 20302 60562
rect 20302 60510 20354 60562
rect 20354 60510 20356 60562
rect 20300 60508 20356 60510
rect 20412 60396 20468 60452
rect 20076 60284 20132 60340
rect 20076 60002 20132 60004
rect 20076 59950 20078 60002
rect 20078 59950 20130 60002
rect 20130 59950 20132 60002
rect 20076 59948 20132 59950
rect 20300 59330 20356 59332
rect 20300 59278 20302 59330
rect 20302 59278 20354 59330
rect 20354 59278 20356 59330
rect 20300 59276 20356 59278
rect 20188 58156 20244 58212
rect 19964 57762 20020 57764
rect 19964 57710 19966 57762
rect 19966 57710 20018 57762
rect 20018 57710 20020 57762
rect 19964 57708 20020 57710
rect 20188 57708 20244 57764
rect 19852 57484 19908 57540
rect 19628 55916 19684 55972
rect 19852 57148 19908 57204
rect 19516 55692 19572 55748
rect 20188 55970 20244 55972
rect 20188 55918 20190 55970
rect 20190 55918 20242 55970
rect 20242 55918 20244 55970
rect 20188 55916 20244 55918
rect 19964 55468 20020 55524
rect 20188 55692 20244 55748
rect 19628 54796 19684 54852
rect 19740 54684 19796 54740
rect 19404 53506 19460 53508
rect 19404 53454 19406 53506
rect 19406 53454 19458 53506
rect 19458 53454 19460 53506
rect 19404 53452 19460 53454
rect 20076 54124 20132 54180
rect 21308 64876 21364 64932
rect 21980 65660 22036 65716
rect 22092 66162 22148 66164
rect 22092 66110 22094 66162
rect 22094 66110 22146 66162
rect 22146 66110 22148 66162
rect 22092 66108 22148 66110
rect 21868 65100 21924 65156
rect 21532 64876 21588 64932
rect 22092 64594 22148 64596
rect 22092 64542 22094 64594
rect 22094 64542 22146 64594
rect 22146 64542 22148 64594
rect 22092 64540 22148 64542
rect 22540 66162 22596 66164
rect 22540 66110 22542 66162
rect 22542 66110 22594 66162
rect 22594 66110 22596 66162
rect 22540 66108 22596 66110
rect 22428 65772 22484 65828
rect 22316 65548 22372 65604
rect 22316 64764 22372 64820
rect 22428 65436 22484 65492
rect 21624 64314 21680 64316
rect 21624 64262 21626 64314
rect 21626 64262 21678 64314
rect 21678 64262 21680 64314
rect 21624 64260 21680 64262
rect 21728 64314 21784 64316
rect 21728 64262 21730 64314
rect 21730 64262 21782 64314
rect 21782 64262 21784 64314
rect 21728 64260 21784 64262
rect 21832 64314 21888 64316
rect 21832 64262 21834 64314
rect 21834 64262 21886 64314
rect 21886 64262 21888 64314
rect 21832 64260 21888 64262
rect 21868 64146 21924 64148
rect 21868 64094 21870 64146
rect 21870 64094 21922 64146
rect 21922 64094 21924 64146
rect 21868 64092 21924 64094
rect 21308 63980 21364 64036
rect 21756 63756 21812 63812
rect 21644 63698 21700 63700
rect 21644 63646 21646 63698
rect 21646 63646 21698 63698
rect 21698 63646 21700 63698
rect 21644 63644 21700 63646
rect 22092 63644 22148 63700
rect 22316 64204 22372 64260
rect 21624 62746 21680 62748
rect 21624 62694 21626 62746
rect 21626 62694 21678 62746
rect 21678 62694 21680 62746
rect 21624 62692 21680 62694
rect 21728 62746 21784 62748
rect 21728 62694 21730 62746
rect 21730 62694 21782 62746
rect 21782 62694 21784 62746
rect 21728 62692 21784 62694
rect 21832 62746 21888 62748
rect 21832 62694 21834 62746
rect 21834 62694 21886 62746
rect 21886 62694 21888 62746
rect 21832 62692 21888 62694
rect 22092 62242 22148 62244
rect 22092 62190 22094 62242
rect 22094 62190 22146 62242
rect 22146 62190 22148 62242
rect 22092 62188 22148 62190
rect 20636 60562 20692 60564
rect 20636 60510 20638 60562
rect 20638 60510 20690 60562
rect 20690 60510 20692 60562
rect 20636 60508 20692 60510
rect 20636 59836 20692 59892
rect 20636 58604 20692 58660
rect 20748 57708 20804 57764
rect 20972 60844 21028 60900
rect 20636 56252 20692 56308
rect 20076 53564 20132 53620
rect 19740 52780 19796 52836
rect 20076 52332 20132 52388
rect 19964 52220 20020 52276
rect 19180 51548 19236 51604
rect 19404 51772 19460 51828
rect 19740 51602 19796 51604
rect 19740 51550 19742 51602
rect 19742 51550 19794 51602
rect 19794 51550 19796 51602
rect 19740 51548 19796 51550
rect 19180 50652 19236 50708
rect 19628 51324 19684 51380
rect 20524 54572 20580 54628
rect 20524 54236 20580 54292
rect 20300 54012 20356 54068
rect 20748 55356 20804 55412
rect 21624 61178 21680 61180
rect 21624 61126 21626 61178
rect 21626 61126 21678 61178
rect 21678 61126 21680 61178
rect 21624 61124 21680 61126
rect 21728 61178 21784 61180
rect 21728 61126 21730 61178
rect 21730 61126 21782 61178
rect 21782 61126 21784 61178
rect 21728 61124 21784 61126
rect 21832 61178 21888 61180
rect 21832 61126 21834 61178
rect 21834 61126 21886 61178
rect 21886 61126 21888 61178
rect 21832 61124 21888 61126
rect 21308 60732 21364 60788
rect 21084 58156 21140 58212
rect 21196 60620 21252 60676
rect 21196 56140 21252 56196
rect 21420 60508 21476 60564
rect 21868 60508 21924 60564
rect 22092 60620 22148 60676
rect 21644 60114 21700 60116
rect 21644 60062 21646 60114
rect 21646 60062 21698 60114
rect 21698 60062 21700 60114
rect 21644 60060 21700 60062
rect 21624 59610 21680 59612
rect 21624 59558 21626 59610
rect 21626 59558 21678 59610
rect 21678 59558 21680 59610
rect 21624 59556 21680 59558
rect 21728 59610 21784 59612
rect 21728 59558 21730 59610
rect 21730 59558 21782 59610
rect 21782 59558 21784 59610
rect 21728 59556 21784 59558
rect 21832 59610 21888 59612
rect 21832 59558 21834 59610
rect 21834 59558 21886 59610
rect 21886 59558 21888 59610
rect 21832 59556 21888 59558
rect 21532 58828 21588 58884
rect 21624 58042 21680 58044
rect 21624 57990 21626 58042
rect 21626 57990 21678 58042
rect 21678 57990 21680 58042
rect 21624 57988 21680 57990
rect 21728 58042 21784 58044
rect 21728 57990 21730 58042
rect 21730 57990 21782 58042
rect 21782 57990 21784 58042
rect 21728 57988 21784 57990
rect 21832 58042 21888 58044
rect 21832 57990 21834 58042
rect 21834 57990 21886 58042
rect 21886 57990 21888 58042
rect 21832 57988 21888 57990
rect 21644 57762 21700 57764
rect 21644 57710 21646 57762
rect 21646 57710 21698 57762
rect 21698 57710 21700 57762
rect 21644 57708 21700 57710
rect 21980 57148 22036 57204
rect 21980 56866 22036 56868
rect 21980 56814 21982 56866
rect 21982 56814 22034 56866
rect 22034 56814 22036 56866
rect 21980 56812 22036 56814
rect 21420 56754 21476 56756
rect 21420 56702 21422 56754
rect 21422 56702 21474 56754
rect 21474 56702 21476 56754
rect 21420 56700 21476 56702
rect 21624 56474 21680 56476
rect 21624 56422 21626 56474
rect 21626 56422 21678 56474
rect 21678 56422 21680 56474
rect 21624 56420 21680 56422
rect 21728 56474 21784 56476
rect 21728 56422 21730 56474
rect 21730 56422 21782 56474
rect 21782 56422 21784 56474
rect 21728 56420 21784 56422
rect 21832 56474 21888 56476
rect 21832 56422 21834 56474
rect 21834 56422 21886 56474
rect 21886 56422 21888 56474
rect 21832 56420 21888 56422
rect 21532 56252 21588 56308
rect 20972 55244 21028 55300
rect 21420 55916 21476 55972
rect 20860 55020 20916 55076
rect 21308 55468 21364 55524
rect 21868 55692 21924 55748
rect 22428 64034 22484 64036
rect 22428 63982 22430 64034
rect 22430 63982 22482 64034
rect 22482 63982 22484 64034
rect 22428 63980 22484 63982
rect 22316 63532 22372 63588
rect 22428 62188 22484 62244
rect 22316 61180 22372 61236
rect 22428 60674 22484 60676
rect 22428 60622 22430 60674
rect 22430 60622 22482 60674
rect 22482 60622 22484 60674
rect 22428 60620 22484 60622
rect 23772 72268 23828 72324
rect 23660 71650 23716 71652
rect 23660 71598 23662 71650
rect 23662 71598 23714 71650
rect 23714 71598 23716 71650
rect 23660 71596 23716 71598
rect 23436 71484 23492 71540
rect 23436 71260 23492 71316
rect 23324 70924 23380 70980
rect 23100 70812 23156 70868
rect 22876 68012 22932 68068
rect 22988 68460 23044 68516
rect 22876 67842 22932 67844
rect 22876 67790 22878 67842
rect 22878 67790 22930 67842
rect 22930 67790 22932 67842
rect 22876 67788 22932 67790
rect 23324 70028 23380 70084
rect 23996 73442 24052 73444
rect 23996 73390 23998 73442
rect 23998 73390 24050 73442
rect 24050 73390 24052 73442
rect 23996 73388 24052 73390
rect 24108 72322 24164 72324
rect 24108 72270 24110 72322
rect 24110 72270 24162 72322
rect 24162 72270 24164 72322
rect 24108 72268 24164 72270
rect 25228 75628 25284 75684
rect 25228 75404 25284 75460
rect 24892 74620 24948 74676
rect 25026 74506 25082 74508
rect 25026 74454 25028 74506
rect 25028 74454 25080 74506
rect 25080 74454 25082 74506
rect 25026 74452 25082 74454
rect 25130 74506 25186 74508
rect 25130 74454 25132 74506
rect 25132 74454 25184 74506
rect 25184 74454 25186 74506
rect 25130 74452 25186 74454
rect 25234 74506 25290 74508
rect 25234 74454 25236 74506
rect 25236 74454 25288 74506
rect 25288 74454 25290 74506
rect 25234 74452 25290 74454
rect 24556 73890 24612 73892
rect 24556 73838 24558 73890
rect 24558 73838 24610 73890
rect 24610 73838 24612 73890
rect 24556 73836 24612 73838
rect 24332 73724 24388 73780
rect 24332 73388 24388 73444
rect 25004 74172 25060 74228
rect 24892 73836 24948 73892
rect 24668 72940 24724 72996
rect 24556 72322 24612 72324
rect 24556 72270 24558 72322
rect 24558 72270 24610 72322
rect 24610 72270 24612 72322
rect 24556 72268 24612 72270
rect 24556 72044 24612 72100
rect 24668 71708 24724 71764
rect 23548 68796 23604 68852
rect 23436 68460 23492 68516
rect 23212 67730 23268 67732
rect 23212 67678 23214 67730
rect 23214 67678 23266 67730
rect 23266 67678 23268 67730
rect 23212 67676 23268 67678
rect 23100 67618 23156 67620
rect 23100 67566 23102 67618
rect 23102 67566 23154 67618
rect 23154 67566 23156 67618
rect 23100 67564 23156 67566
rect 23324 67618 23380 67620
rect 23324 67566 23326 67618
rect 23326 67566 23378 67618
rect 23378 67566 23380 67618
rect 23324 67564 23380 67566
rect 22876 66274 22932 66276
rect 22876 66222 22878 66274
rect 22878 66222 22930 66274
rect 22930 66222 22932 66274
rect 22876 66220 22932 66222
rect 23324 66780 23380 66836
rect 23436 66220 23492 66276
rect 23100 65602 23156 65604
rect 23100 65550 23102 65602
rect 23102 65550 23154 65602
rect 23154 65550 23156 65602
rect 23100 65548 23156 65550
rect 22764 64652 22820 64708
rect 23212 65212 23268 65268
rect 22876 64764 22932 64820
rect 23548 65212 23604 65268
rect 23436 64204 23492 64260
rect 22876 64092 22932 64148
rect 23100 63922 23156 63924
rect 23100 63870 23102 63922
rect 23102 63870 23154 63922
rect 23154 63870 23156 63922
rect 23100 63868 23156 63870
rect 22876 63644 22932 63700
rect 23436 63756 23492 63812
rect 23100 63420 23156 63476
rect 22876 62972 22932 63028
rect 22652 61570 22708 61572
rect 22652 61518 22654 61570
rect 22654 61518 22706 61570
rect 22706 61518 22708 61570
rect 22652 61516 22708 61518
rect 23100 62524 23156 62580
rect 23436 62860 23492 62916
rect 23100 60620 23156 60676
rect 23212 62188 23268 62244
rect 23100 60396 23156 60452
rect 22764 60284 22820 60340
rect 22428 59724 22484 59780
rect 22764 59836 22820 59892
rect 22316 58492 22372 58548
rect 22652 59388 22708 59444
rect 22316 58210 22372 58212
rect 22316 58158 22318 58210
rect 22318 58158 22370 58210
rect 22370 58158 22372 58210
rect 22316 58156 22372 58158
rect 22316 56812 22372 56868
rect 22204 56252 22260 56308
rect 22988 59218 23044 59220
rect 22988 59166 22990 59218
rect 22990 59166 23042 59218
rect 23042 59166 23044 59218
rect 22988 59164 23044 59166
rect 22540 57538 22596 57540
rect 22540 57486 22542 57538
rect 22542 57486 22594 57538
rect 22594 57486 22596 57538
rect 22540 57484 22596 57486
rect 22876 58492 22932 58548
rect 22540 56252 22596 56308
rect 22652 56140 22708 56196
rect 22092 55580 22148 55636
rect 22316 55468 22372 55524
rect 21644 55186 21700 55188
rect 21644 55134 21646 55186
rect 21646 55134 21698 55186
rect 21698 55134 21700 55186
rect 21644 55132 21700 55134
rect 21084 54572 21140 54628
rect 20860 54348 20916 54404
rect 21196 54514 21252 54516
rect 21196 54462 21198 54514
rect 21198 54462 21250 54514
rect 21250 54462 21252 54514
rect 21196 54460 21252 54462
rect 21084 54348 21140 54404
rect 20748 54236 20804 54292
rect 21196 54236 21252 54292
rect 20300 53730 20356 53732
rect 20300 53678 20302 53730
rect 20302 53678 20354 53730
rect 20354 53678 20356 53730
rect 20300 53676 20356 53678
rect 20636 53730 20692 53732
rect 20636 53678 20638 53730
rect 20638 53678 20690 53730
rect 20690 53678 20692 53730
rect 20636 53676 20692 53678
rect 20300 53452 20356 53508
rect 20300 53116 20356 53172
rect 20524 53058 20580 53060
rect 20524 53006 20526 53058
rect 20526 53006 20578 53058
rect 20578 53006 20580 53058
rect 20524 53004 20580 53006
rect 20636 52892 20692 52948
rect 19628 50764 19684 50820
rect 19964 51100 20020 51156
rect 19180 50316 19236 50372
rect 18508 49922 18564 49924
rect 18508 49870 18510 49922
rect 18510 49870 18562 49922
rect 18562 49870 18564 49922
rect 18508 49868 18564 49870
rect 18222 49418 18278 49420
rect 18222 49366 18224 49418
rect 18224 49366 18276 49418
rect 18276 49366 18278 49418
rect 18222 49364 18278 49366
rect 18326 49418 18382 49420
rect 18326 49366 18328 49418
rect 18328 49366 18380 49418
rect 18380 49366 18382 49418
rect 18326 49364 18382 49366
rect 18430 49418 18486 49420
rect 18430 49366 18432 49418
rect 18432 49366 18484 49418
rect 18484 49366 18486 49418
rect 18430 49364 18486 49366
rect 18956 49810 19012 49812
rect 18956 49758 18958 49810
rect 18958 49758 19010 49810
rect 19010 49758 19012 49810
rect 18956 49756 19012 49758
rect 18956 49026 19012 49028
rect 18956 48974 18958 49026
rect 18958 48974 19010 49026
rect 19010 48974 19012 49026
rect 18956 48972 19012 48974
rect 19068 49644 19124 49700
rect 18222 47850 18278 47852
rect 18222 47798 18224 47850
rect 18224 47798 18276 47850
rect 18276 47798 18278 47850
rect 18222 47796 18278 47798
rect 18326 47850 18382 47852
rect 18326 47798 18328 47850
rect 18328 47798 18380 47850
rect 18380 47798 18382 47850
rect 18326 47796 18382 47798
rect 18430 47850 18486 47852
rect 18430 47798 18432 47850
rect 18432 47798 18484 47850
rect 18484 47798 18486 47850
rect 18430 47796 18486 47798
rect 18396 47628 18452 47684
rect 17612 45276 17668 45332
rect 17948 47180 18004 47236
rect 17500 44492 17556 44548
rect 17500 44044 17556 44100
rect 17612 42252 17668 42308
rect 17836 46956 17892 47012
rect 18620 47404 18676 47460
rect 17836 45724 17892 45780
rect 17836 44492 17892 44548
rect 17948 44604 18004 44660
rect 17948 43596 18004 43652
rect 17612 41970 17668 41972
rect 17612 41918 17614 41970
rect 17614 41918 17666 41970
rect 17666 41918 17668 41970
rect 17612 41916 17668 41918
rect 17724 41468 17780 41524
rect 17500 39564 17556 39620
rect 17388 39452 17444 39508
rect 17724 39340 17780 39396
rect 17836 38892 17892 38948
rect 18222 46282 18278 46284
rect 18222 46230 18224 46282
rect 18224 46230 18276 46282
rect 18276 46230 18278 46282
rect 18222 46228 18278 46230
rect 18326 46282 18382 46284
rect 18326 46230 18328 46282
rect 18328 46230 18380 46282
rect 18380 46230 18382 46282
rect 18326 46228 18382 46230
rect 18430 46282 18486 46284
rect 18430 46230 18432 46282
rect 18432 46230 18484 46282
rect 18484 46230 18486 46282
rect 18430 46228 18486 46230
rect 18956 48748 19012 48804
rect 18396 45164 18452 45220
rect 18222 44714 18278 44716
rect 18222 44662 18224 44714
rect 18224 44662 18276 44714
rect 18276 44662 18278 44714
rect 18222 44660 18278 44662
rect 18326 44714 18382 44716
rect 18326 44662 18328 44714
rect 18328 44662 18380 44714
rect 18380 44662 18382 44714
rect 18326 44660 18382 44662
rect 18430 44714 18486 44716
rect 18430 44662 18432 44714
rect 18432 44662 18484 44714
rect 18484 44662 18486 44714
rect 18430 44660 18486 44662
rect 18172 43426 18228 43428
rect 18172 43374 18174 43426
rect 18174 43374 18226 43426
rect 18226 43374 18228 43426
rect 18172 43372 18228 43374
rect 18508 43372 18564 43428
rect 18222 43146 18278 43148
rect 18222 43094 18224 43146
rect 18224 43094 18276 43146
rect 18276 43094 18278 43146
rect 18222 43092 18278 43094
rect 18326 43146 18382 43148
rect 18326 43094 18328 43146
rect 18328 43094 18380 43146
rect 18380 43094 18382 43146
rect 18326 43092 18382 43094
rect 18430 43146 18486 43148
rect 18430 43094 18432 43146
rect 18432 43094 18484 43146
rect 18484 43094 18486 43146
rect 18430 43092 18486 43094
rect 18844 45164 18900 45220
rect 18284 42476 18340 42532
rect 18732 42252 18788 42308
rect 18508 42028 18564 42084
rect 18396 41970 18452 41972
rect 18396 41918 18398 41970
rect 18398 41918 18450 41970
rect 18450 41918 18452 41970
rect 18396 41916 18452 41918
rect 18844 41916 18900 41972
rect 18222 41578 18278 41580
rect 18222 41526 18224 41578
rect 18224 41526 18276 41578
rect 18276 41526 18278 41578
rect 18222 41524 18278 41526
rect 18326 41578 18382 41580
rect 18326 41526 18328 41578
rect 18328 41526 18380 41578
rect 18380 41526 18382 41578
rect 18326 41524 18382 41526
rect 18430 41578 18486 41580
rect 18430 41526 18432 41578
rect 18432 41526 18484 41578
rect 18484 41526 18486 41578
rect 18430 41524 18486 41526
rect 18284 41356 18340 41412
rect 18844 41244 18900 41300
rect 18284 40348 18340 40404
rect 18222 40010 18278 40012
rect 18222 39958 18224 40010
rect 18224 39958 18276 40010
rect 18276 39958 18278 40010
rect 18222 39956 18278 39958
rect 18326 40010 18382 40012
rect 18326 39958 18328 40010
rect 18328 39958 18380 40010
rect 18380 39958 18382 40010
rect 18326 39956 18382 39958
rect 18430 40010 18486 40012
rect 18430 39958 18432 40010
rect 18432 39958 18484 40010
rect 18484 39958 18486 40010
rect 18430 39956 18486 39958
rect 18844 40236 18900 40292
rect 18620 39564 18676 39620
rect 18172 39394 18228 39396
rect 18172 39342 18174 39394
rect 18174 39342 18226 39394
rect 18226 39342 18228 39394
rect 18172 39340 18228 39342
rect 17500 38108 17556 38164
rect 17612 38668 17668 38724
rect 18508 38834 18564 38836
rect 18508 38782 18510 38834
rect 18510 38782 18562 38834
rect 18562 38782 18564 38834
rect 18508 38780 18564 38782
rect 17948 38556 18004 38612
rect 17388 37100 17444 37156
rect 17948 36988 18004 37044
rect 18222 38442 18278 38444
rect 18222 38390 18224 38442
rect 18224 38390 18276 38442
rect 18276 38390 18278 38442
rect 18222 38388 18278 38390
rect 18326 38442 18382 38444
rect 18326 38390 18328 38442
rect 18328 38390 18380 38442
rect 18380 38390 18382 38442
rect 18326 38388 18382 38390
rect 18430 38442 18486 38444
rect 18430 38390 18432 38442
rect 18432 38390 18484 38442
rect 18484 38390 18486 38442
rect 18430 38388 18486 38390
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 18396 37100 18452 37156
rect 18222 36874 18278 36876
rect 18222 36822 18224 36874
rect 18224 36822 18276 36874
rect 18276 36822 18278 36874
rect 18222 36820 18278 36822
rect 18326 36874 18382 36876
rect 18326 36822 18328 36874
rect 18328 36822 18380 36874
rect 18380 36822 18382 36874
rect 18326 36820 18382 36822
rect 18430 36874 18486 36876
rect 18430 36822 18432 36874
rect 18432 36822 18484 36874
rect 18484 36822 18486 36874
rect 18430 36820 18486 36822
rect 16604 35756 16660 35812
rect 16604 33516 16660 33572
rect 16716 35644 16772 35700
rect 17164 36258 17220 36260
rect 17164 36206 17166 36258
rect 17166 36206 17218 36258
rect 17218 36206 17220 36258
rect 17164 36204 17220 36206
rect 17612 36370 17668 36372
rect 17612 36318 17614 36370
rect 17614 36318 17666 36370
rect 17666 36318 17668 36370
rect 17612 36316 17668 36318
rect 17500 36092 17556 36148
rect 16604 32732 16660 32788
rect 17052 33628 17108 33684
rect 16940 33516 16996 33572
rect 16828 32450 16884 32452
rect 16828 32398 16830 32450
rect 16830 32398 16882 32450
rect 16882 32398 16884 32450
rect 16828 32396 16884 32398
rect 15372 31052 15428 31108
rect 15484 31164 15540 31220
rect 14588 29596 14644 29652
rect 14588 28140 14644 28196
rect 14924 29986 14980 29988
rect 14924 29934 14926 29986
rect 14926 29934 14978 29986
rect 14978 29934 14980 29986
rect 14924 29932 14980 29934
rect 14820 29818 14876 29820
rect 14820 29766 14822 29818
rect 14822 29766 14874 29818
rect 14874 29766 14876 29818
rect 14820 29764 14876 29766
rect 14924 29818 14980 29820
rect 14924 29766 14926 29818
rect 14926 29766 14978 29818
rect 14978 29766 14980 29818
rect 14924 29764 14980 29766
rect 15028 29818 15084 29820
rect 15028 29766 15030 29818
rect 15030 29766 15082 29818
rect 15082 29766 15084 29818
rect 15028 29764 15084 29766
rect 14812 29596 14868 29652
rect 14812 29260 14868 29316
rect 15372 30044 15428 30100
rect 15148 29148 15204 29204
rect 15036 28812 15092 28868
rect 14812 28754 14868 28756
rect 14812 28702 14814 28754
rect 14814 28702 14866 28754
rect 14866 28702 14868 28754
rect 14812 28700 14868 28702
rect 14924 28642 14980 28644
rect 14924 28590 14926 28642
rect 14926 28590 14978 28642
rect 14978 28590 14980 28642
rect 14924 28588 14980 28590
rect 15260 29932 15316 29988
rect 15260 28700 15316 28756
rect 14820 28250 14876 28252
rect 14820 28198 14822 28250
rect 14822 28198 14874 28250
rect 14874 28198 14876 28250
rect 14820 28196 14876 28198
rect 14924 28250 14980 28252
rect 14924 28198 14926 28250
rect 14926 28198 14978 28250
rect 14978 28198 14980 28250
rect 14924 28196 14980 28198
rect 15028 28250 15084 28252
rect 15028 28198 15030 28250
rect 15030 28198 15082 28250
rect 15082 28198 15084 28250
rect 15028 28196 15084 28198
rect 14924 27858 14980 27860
rect 14924 27806 14926 27858
rect 14926 27806 14978 27858
rect 14978 27806 14980 27858
rect 14924 27804 14980 27806
rect 15036 27692 15092 27748
rect 15260 28028 15316 28084
rect 15260 27746 15316 27748
rect 15260 27694 15262 27746
rect 15262 27694 15314 27746
rect 15314 27694 15316 27746
rect 15260 27692 15316 27694
rect 15260 27020 15316 27076
rect 14820 26682 14876 26684
rect 14820 26630 14822 26682
rect 14822 26630 14874 26682
rect 14874 26630 14876 26682
rect 14820 26628 14876 26630
rect 14924 26682 14980 26684
rect 14924 26630 14926 26682
rect 14926 26630 14978 26682
rect 14978 26630 14980 26682
rect 14924 26628 14980 26630
rect 15028 26682 15084 26684
rect 15028 26630 15030 26682
rect 15030 26630 15082 26682
rect 15082 26630 15084 26682
rect 15028 26628 15084 26630
rect 15372 26236 15428 26292
rect 15148 26066 15204 26068
rect 15148 26014 15150 26066
rect 15150 26014 15202 26066
rect 15202 26014 15204 26066
rect 15148 26012 15204 26014
rect 14364 25282 14420 25284
rect 14364 25230 14366 25282
rect 14366 25230 14418 25282
rect 14418 25230 14420 25282
rect 14364 25228 14420 25230
rect 14820 25114 14876 25116
rect 14820 25062 14822 25114
rect 14822 25062 14874 25114
rect 14874 25062 14876 25114
rect 14820 25060 14876 25062
rect 14924 25114 14980 25116
rect 14924 25062 14926 25114
rect 14926 25062 14978 25114
rect 14978 25062 14980 25114
rect 14924 25060 14980 25062
rect 15028 25114 15084 25116
rect 15028 25062 15030 25114
rect 15030 25062 15082 25114
rect 15082 25062 15084 25114
rect 15028 25060 15084 25062
rect 13916 24108 13972 24164
rect 13692 23772 13748 23828
rect 13580 22428 13636 22484
rect 12908 20914 12964 20916
rect 12908 20862 12910 20914
rect 12910 20862 12962 20914
rect 12962 20862 12964 20914
rect 12908 20860 12964 20862
rect 13692 22988 13748 23044
rect 13580 21756 13636 21812
rect 13132 20748 13188 20804
rect 13692 20690 13748 20692
rect 13692 20638 13694 20690
rect 13694 20638 13746 20690
rect 13746 20638 13748 20690
rect 13692 20636 13748 20638
rect 13468 20524 13524 20580
rect 12908 20076 12964 20132
rect 14476 24108 14532 24164
rect 14028 24050 14084 24052
rect 14028 23998 14030 24050
rect 14030 23998 14082 24050
rect 14082 23998 14084 24050
rect 14028 23996 14084 23998
rect 15148 24556 15204 24612
rect 15372 25676 15428 25732
rect 15372 24108 15428 24164
rect 14812 23772 14868 23828
rect 14820 23546 14876 23548
rect 14820 23494 14822 23546
rect 14822 23494 14874 23546
rect 14874 23494 14876 23546
rect 14820 23492 14876 23494
rect 14924 23546 14980 23548
rect 14924 23494 14926 23546
rect 14926 23494 14978 23546
rect 14978 23494 14980 23546
rect 14924 23492 14980 23494
rect 15028 23546 15084 23548
rect 15028 23494 15030 23546
rect 15030 23494 15082 23546
rect 15082 23494 15084 23546
rect 15028 23492 15084 23494
rect 15148 23324 15204 23380
rect 14476 23100 14532 23156
rect 14476 21698 14532 21700
rect 14476 21646 14478 21698
rect 14478 21646 14530 21698
rect 14530 21646 14532 21698
rect 14476 21644 14532 21646
rect 14252 21474 14308 21476
rect 14252 21422 14254 21474
rect 14254 21422 14306 21474
rect 14306 21422 14308 21474
rect 14252 21420 14308 21422
rect 14252 20860 14308 20916
rect 14700 22428 14756 22484
rect 15708 30268 15764 30324
rect 15596 30210 15652 30212
rect 15596 30158 15598 30210
rect 15598 30158 15650 30210
rect 15650 30158 15652 30210
rect 15596 30156 15652 30158
rect 16044 31500 16100 31556
rect 16268 31388 16324 31444
rect 16492 31218 16548 31220
rect 16492 31166 16494 31218
rect 16494 31166 16546 31218
rect 16546 31166 16548 31218
rect 16492 31164 16548 31166
rect 16380 30156 16436 30212
rect 16940 30940 16996 30996
rect 16828 30828 16884 30884
rect 16716 30044 16772 30100
rect 15596 29148 15652 29204
rect 15708 28754 15764 28756
rect 15708 28702 15710 28754
rect 15710 28702 15762 28754
rect 15762 28702 15764 28754
rect 15708 28700 15764 28702
rect 15708 28476 15764 28532
rect 15596 27356 15652 27412
rect 15708 26348 15764 26404
rect 16044 28642 16100 28644
rect 16044 28590 16046 28642
rect 16046 28590 16098 28642
rect 16098 28590 16100 28642
rect 16044 28588 16100 28590
rect 16380 27804 16436 27860
rect 16156 27746 16212 27748
rect 16156 27694 16158 27746
rect 16158 27694 16210 27746
rect 16210 27694 16212 27746
rect 16156 27692 16212 27694
rect 16940 27916 16996 27972
rect 17052 28028 17108 28084
rect 16716 27132 16772 27188
rect 17388 35698 17444 35700
rect 17388 35646 17390 35698
rect 17390 35646 17442 35698
rect 17442 35646 17444 35698
rect 17388 35644 17444 35646
rect 17612 34802 17668 34804
rect 17612 34750 17614 34802
rect 17614 34750 17666 34802
rect 17666 34750 17668 34802
rect 17612 34748 17668 34750
rect 17612 33628 17668 33684
rect 17500 32732 17556 32788
rect 18396 36594 18452 36596
rect 18396 36542 18398 36594
rect 18398 36542 18450 36594
rect 18450 36542 18452 36594
rect 18396 36540 18452 36542
rect 19292 48860 19348 48916
rect 19292 48076 19348 48132
rect 19180 47628 19236 47684
rect 19180 46562 19236 46564
rect 19180 46510 19182 46562
rect 19182 46510 19234 46562
rect 19234 46510 19236 46562
rect 19180 46508 19236 46510
rect 19180 44156 19236 44212
rect 19516 49980 19572 50036
rect 20412 52780 20468 52836
rect 20076 50370 20132 50372
rect 20076 50318 20078 50370
rect 20078 50318 20130 50370
rect 20130 50318 20132 50370
rect 20076 50316 20132 50318
rect 19516 49810 19572 49812
rect 19516 49758 19518 49810
rect 19518 49758 19570 49810
rect 19570 49758 19572 49810
rect 19516 49756 19572 49758
rect 19740 48636 19796 48692
rect 19516 47404 19572 47460
rect 19740 47852 19796 47908
rect 19740 47068 19796 47124
rect 19516 46508 19572 46564
rect 19628 45612 19684 45668
rect 19740 45388 19796 45444
rect 19404 43650 19460 43652
rect 19404 43598 19406 43650
rect 19406 43598 19458 43650
rect 19458 43598 19460 43650
rect 19404 43596 19460 43598
rect 19292 43538 19348 43540
rect 19292 43486 19294 43538
rect 19294 43486 19346 43538
rect 19346 43486 19348 43538
rect 19292 43484 19348 43486
rect 19180 42476 19236 42532
rect 19404 42082 19460 42084
rect 19404 42030 19406 42082
rect 19406 42030 19458 42082
rect 19458 42030 19460 42082
rect 19404 42028 19460 42030
rect 19068 41970 19124 41972
rect 19068 41918 19070 41970
rect 19070 41918 19122 41970
rect 19122 41918 19124 41970
rect 19068 41916 19124 41918
rect 18844 37660 18900 37716
rect 18732 36428 18788 36484
rect 18844 37100 18900 37156
rect 18956 36988 19012 37044
rect 19180 36764 19236 36820
rect 17836 35420 17892 35476
rect 18222 35306 18278 35308
rect 18222 35254 18224 35306
rect 18224 35254 18276 35306
rect 18276 35254 18278 35306
rect 18222 35252 18278 35254
rect 18326 35306 18382 35308
rect 18326 35254 18328 35306
rect 18328 35254 18380 35306
rect 18380 35254 18382 35306
rect 18326 35252 18382 35254
rect 18430 35306 18486 35308
rect 18430 35254 18432 35306
rect 18432 35254 18484 35306
rect 18484 35254 18486 35306
rect 18430 35252 18486 35254
rect 18732 35252 18788 35308
rect 17948 34914 18004 34916
rect 17948 34862 17950 34914
rect 17950 34862 18002 34914
rect 18002 34862 18004 34914
rect 17948 34860 18004 34862
rect 18172 34748 18228 34804
rect 17724 32732 17780 32788
rect 17388 32674 17444 32676
rect 17388 32622 17390 32674
rect 17390 32622 17442 32674
rect 17442 32622 17444 32674
rect 17388 32620 17444 32622
rect 17724 32396 17780 32452
rect 17500 31388 17556 31444
rect 17276 31164 17332 31220
rect 18620 34636 18676 34692
rect 18060 34018 18116 34020
rect 18060 33966 18062 34018
rect 18062 33966 18114 34018
rect 18114 33966 18116 34018
rect 18060 33964 18116 33966
rect 18222 33738 18278 33740
rect 18222 33686 18224 33738
rect 18224 33686 18276 33738
rect 18276 33686 18278 33738
rect 18222 33684 18278 33686
rect 18326 33738 18382 33740
rect 18326 33686 18328 33738
rect 18328 33686 18380 33738
rect 18380 33686 18382 33738
rect 18326 33684 18382 33686
rect 18430 33738 18486 33740
rect 18430 33686 18432 33738
rect 18432 33686 18484 33738
rect 18484 33686 18486 33738
rect 18430 33684 18486 33686
rect 18060 33516 18116 33572
rect 18508 32732 18564 32788
rect 18956 35308 19012 35364
rect 19180 35532 19236 35588
rect 19180 35138 19236 35140
rect 19180 35086 19182 35138
rect 19182 35086 19234 35138
rect 19234 35086 19236 35138
rect 19180 35084 19236 35086
rect 18844 32732 18900 32788
rect 18956 34860 19012 34916
rect 18060 32508 18116 32564
rect 18396 32396 18452 32452
rect 18222 32170 18278 32172
rect 18222 32118 18224 32170
rect 18224 32118 18276 32170
rect 18276 32118 18278 32170
rect 18222 32116 18278 32118
rect 18326 32170 18382 32172
rect 18326 32118 18328 32170
rect 18328 32118 18380 32170
rect 18380 32118 18382 32170
rect 18326 32116 18382 32118
rect 18430 32170 18486 32172
rect 18430 32118 18432 32170
rect 18432 32118 18484 32170
rect 18484 32118 18486 32170
rect 18430 32116 18486 32118
rect 17388 31052 17444 31108
rect 17388 29932 17444 29988
rect 18172 31106 18228 31108
rect 18172 31054 18174 31106
rect 18174 31054 18226 31106
rect 18226 31054 18228 31106
rect 18172 31052 18228 31054
rect 17836 30994 17892 30996
rect 17836 30942 17838 30994
rect 17838 30942 17890 30994
rect 17890 30942 17892 30994
rect 17836 30940 17892 30942
rect 17612 30268 17668 30324
rect 17836 29260 17892 29316
rect 17836 28364 17892 28420
rect 17836 28028 17892 28084
rect 18844 32562 18900 32564
rect 18844 32510 18846 32562
rect 18846 32510 18898 32562
rect 18898 32510 18900 32562
rect 18844 32508 18900 32510
rect 18620 30940 18676 30996
rect 18732 31948 18788 32004
rect 18222 30602 18278 30604
rect 18222 30550 18224 30602
rect 18224 30550 18276 30602
rect 18276 30550 18278 30602
rect 18222 30548 18278 30550
rect 18326 30602 18382 30604
rect 18326 30550 18328 30602
rect 18328 30550 18380 30602
rect 18380 30550 18382 30602
rect 18326 30548 18382 30550
rect 18430 30602 18486 30604
rect 18430 30550 18432 30602
rect 18432 30550 18484 30602
rect 18484 30550 18486 30602
rect 18430 30548 18486 30550
rect 18396 30322 18452 30324
rect 18396 30270 18398 30322
rect 18398 30270 18450 30322
rect 18450 30270 18452 30322
rect 18396 30268 18452 30270
rect 19068 34354 19124 34356
rect 19068 34302 19070 34354
rect 19070 34302 19122 34354
rect 19122 34302 19124 34354
rect 19068 34300 19124 34302
rect 19068 33234 19124 33236
rect 19068 33182 19070 33234
rect 19070 33182 19122 33234
rect 19122 33182 19124 33234
rect 19068 33180 19124 33182
rect 19068 32172 19124 32228
rect 19068 31724 19124 31780
rect 19404 41356 19460 41412
rect 19516 41298 19572 41300
rect 19516 41246 19518 41298
rect 19518 41246 19570 41298
rect 19570 41246 19572 41298
rect 19516 41244 19572 41246
rect 19404 40796 19460 40852
rect 19740 40908 19796 40964
rect 20076 48972 20132 49028
rect 20188 48860 20244 48916
rect 20188 47180 20244 47236
rect 20300 47068 20356 47124
rect 20860 53900 20916 53956
rect 20860 53004 20916 53060
rect 20524 52162 20580 52164
rect 20524 52110 20526 52162
rect 20526 52110 20578 52162
rect 20578 52110 20580 52162
rect 20524 52108 20580 52110
rect 20748 51996 20804 52052
rect 20524 49868 20580 49924
rect 20636 49084 20692 49140
rect 20524 47740 20580 47796
rect 20524 47516 20580 47572
rect 20524 47234 20580 47236
rect 20524 47182 20526 47234
rect 20526 47182 20578 47234
rect 20578 47182 20580 47234
rect 20524 47180 20580 47182
rect 22204 55074 22260 55076
rect 22204 55022 22206 55074
rect 22206 55022 22258 55074
rect 22258 55022 22260 55074
rect 22204 55020 22260 55022
rect 21624 54906 21680 54908
rect 21624 54854 21626 54906
rect 21626 54854 21678 54906
rect 21678 54854 21680 54906
rect 21624 54852 21680 54854
rect 21728 54906 21784 54908
rect 21728 54854 21730 54906
rect 21730 54854 21782 54906
rect 21782 54854 21784 54906
rect 21728 54852 21784 54854
rect 21832 54906 21888 54908
rect 21832 54854 21834 54906
rect 21834 54854 21886 54906
rect 21886 54854 21888 54906
rect 21832 54852 21888 54854
rect 21644 54572 21700 54628
rect 22428 54402 22484 54404
rect 22428 54350 22430 54402
rect 22430 54350 22482 54402
rect 22482 54350 22484 54402
rect 22428 54348 22484 54350
rect 21980 54124 22036 54180
rect 22764 55356 22820 55412
rect 22876 55132 22932 55188
rect 22652 54796 22708 54852
rect 21644 53564 21700 53620
rect 22204 53618 22260 53620
rect 22204 53566 22206 53618
rect 22206 53566 22258 53618
rect 22258 53566 22260 53618
rect 22204 53564 22260 53566
rect 21980 53506 22036 53508
rect 21980 53454 21982 53506
rect 21982 53454 22034 53506
rect 22034 53454 22036 53506
rect 21980 53452 22036 53454
rect 21624 53338 21680 53340
rect 21624 53286 21626 53338
rect 21626 53286 21678 53338
rect 21678 53286 21680 53338
rect 21624 53284 21680 53286
rect 21728 53338 21784 53340
rect 21728 53286 21730 53338
rect 21730 53286 21782 53338
rect 21782 53286 21784 53338
rect 21728 53284 21784 53286
rect 21832 53338 21888 53340
rect 21832 53286 21834 53338
rect 21834 53286 21886 53338
rect 21886 53286 21888 53338
rect 21832 53284 21888 53286
rect 21308 52780 21364 52836
rect 21644 53004 21700 53060
rect 23324 61570 23380 61572
rect 23324 61518 23326 61570
rect 23326 61518 23378 61570
rect 23378 61518 23380 61570
rect 23324 61516 23380 61518
rect 23772 63922 23828 63924
rect 23772 63870 23774 63922
rect 23774 63870 23826 63922
rect 23826 63870 23828 63922
rect 23772 63868 23828 63870
rect 23660 62972 23716 63028
rect 23548 62188 23604 62244
rect 23772 60172 23828 60228
rect 23436 59388 23492 59444
rect 23660 60060 23716 60116
rect 23772 59890 23828 59892
rect 23772 59838 23774 59890
rect 23774 59838 23826 59890
rect 23826 59838 23828 59890
rect 23772 59836 23828 59838
rect 23548 59218 23604 59220
rect 23548 59166 23550 59218
rect 23550 59166 23602 59218
rect 23602 59166 23604 59218
rect 23548 59164 23604 59166
rect 23436 59052 23492 59108
rect 23772 58546 23828 58548
rect 23772 58494 23774 58546
rect 23774 58494 23826 58546
rect 23826 58494 23828 58546
rect 23772 58492 23828 58494
rect 24220 68684 24276 68740
rect 23996 65772 24052 65828
rect 23996 65490 24052 65492
rect 23996 65438 23998 65490
rect 23998 65438 24050 65490
rect 24050 65438 24052 65490
rect 23996 65436 24052 65438
rect 24780 70754 24836 70756
rect 24780 70702 24782 70754
rect 24782 70702 24834 70754
rect 24834 70702 24836 70754
rect 24780 70700 24836 70702
rect 24444 68460 24500 68516
rect 24444 67676 24500 67732
rect 24556 68348 24612 68404
rect 24668 67170 24724 67172
rect 24668 67118 24670 67170
rect 24670 67118 24722 67170
rect 24722 67118 24724 67170
rect 24668 67116 24724 67118
rect 24444 65490 24500 65492
rect 24444 65438 24446 65490
rect 24446 65438 24498 65490
rect 24498 65438 24500 65490
rect 24444 65436 24500 65438
rect 24444 65212 24500 65268
rect 24220 64818 24276 64820
rect 24220 64766 24222 64818
rect 24222 64766 24274 64818
rect 24274 64766 24276 64818
rect 24220 64764 24276 64766
rect 24220 63922 24276 63924
rect 24220 63870 24222 63922
rect 24222 63870 24274 63922
rect 24274 63870 24276 63922
rect 24220 63868 24276 63870
rect 24108 63756 24164 63812
rect 24332 62972 24388 63028
rect 24220 62242 24276 62244
rect 24220 62190 24222 62242
rect 24222 62190 24274 62242
rect 24274 62190 24276 62242
rect 24220 62188 24276 62190
rect 24108 61628 24164 61684
rect 23996 61404 24052 61460
rect 23436 57932 23492 57988
rect 23212 57484 23268 57540
rect 23212 57148 23268 57204
rect 23436 57650 23492 57652
rect 23436 57598 23438 57650
rect 23438 57598 23490 57650
rect 23490 57598 23492 57650
rect 23436 57596 23492 57598
rect 23436 56028 23492 56084
rect 23212 55410 23268 55412
rect 23212 55358 23214 55410
rect 23214 55358 23266 55410
rect 23266 55358 23268 55410
rect 23212 55356 23268 55358
rect 23100 54796 23156 54852
rect 23436 54684 23492 54740
rect 21644 51996 21700 52052
rect 21868 51996 21924 52052
rect 21624 51770 21680 51772
rect 21624 51718 21626 51770
rect 21626 51718 21678 51770
rect 21678 51718 21680 51770
rect 21624 51716 21680 51718
rect 21728 51770 21784 51772
rect 21728 51718 21730 51770
rect 21730 51718 21782 51770
rect 21782 51718 21784 51770
rect 21728 51716 21784 51718
rect 21832 51770 21888 51772
rect 21832 51718 21834 51770
rect 21834 51718 21886 51770
rect 21886 51718 21888 51770
rect 21832 51716 21888 51718
rect 21980 51660 22036 51716
rect 21308 50876 21364 50932
rect 20972 49980 21028 50036
rect 20860 47852 20916 47908
rect 20860 47682 20916 47684
rect 20860 47630 20862 47682
rect 20862 47630 20914 47682
rect 20914 47630 20916 47682
rect 20860 47628 20916 47630
rect 20748 47068 20804 47124
rect 20300 46674 20356 46676
rect 20300 46622 20302 46674
rect 20302 46622 20354 46674
rect 20354 46622 20356 46674
rect 20300 46620 20356 46622
rect 20412 45666 20468 45668
rect 20412 45614 20414 45666
rect 20414 45614 20466 45666
rect 20466 45614 20468 45666
rect 20412 45612 20468 45614
rect 20188 44098 20244 44100
rect 20188 44046 20190 44098
rect 20190 44046 20242 44098
rect 20242 44046 20244 44098
rect 20188 44044 20244 44046
rect 20188 43762 20244 43764
rect 20188 43710 20190 43762
rect 20190 43710 20242 43762
rect 20242 43710 20244 43762
rect 20188 43708 20244 43710
rect 20524 45164 20580 45220
rect 20524 44044 20580 44100
rect 20300 43260 20356 43316
rect 20860 46844 20916 46900
rect 21624 50202 21680 50204
rect 21624 50150 21626 50202
rect 21626 50150 21678 50202
rect 21678 50150 21680 50202
rect 21624 50148 21680 50150
rect 21728 50202 21784 50204
rect 21728 50150 21730 50202
rect 21730 50150 21782 50202
rect 21782 50150 21784 50202
rect 21728 50148 21784 50150
rect 21832 50202 21888 50204
rect 21832 50150 21834 50202
rect 21834 50150 21886 50202
rect 21886 50150 21888 50202
rect 21832 50148 21888 50150
rect 21420 49138 21476 49140
rect 21420 49086 21422 49138
rect 21422 49086 21474 49138
rect 21474 49086 21476 49138
rect 21420 49084 21476 49086
rect 21868 48860 21924 48916
rect 21624 48634 21680 48636
rect 21624 48582 21626 48634
rect 21626 48582 21678 48634
rect 21678 48582 21680 48634
rect 21624 48580 21680 48582
rect 21728 48634 21784 48636
rect 21728 48582 21730 48634
rect 21730 48582 21782 48634
rect 21782 48582 21784 48634
rect 21728 48580 21784 48582
rect 21832 48634 21888 48636
rect 21832 48582 21834 48634
rect 21834 48582 21886 48634
rect 21886 48582 21888 48634
rect 21832 48580 21888 48582
rect 21644 48242 21700 48244
rect 21644 48190 21646 48242
rect 21646 48190 21698 48242
rect 21698 48190 21700 48242
rect 21644 48188 21700 48190
rect 21532 47628 21588 47684
rect 21420 47404 21476 47460
rect 22540 53228 22596 53284
rect 22428 52162 22484 52164
rect 22428 52110 22430 52162
rect 22430 52110 22482 52162
rect 22482 52110 22484 52162
rect 22428 52108 22484 52110
rect 22204 49196 22260 49252
rect 22316 50540 22372 50596
rect 22428 50428 22484 50484
rect 23100 54124 23156 54180
rect 22988 53506 23044 53508
rect 22988 53454 22990 53506
rect 22990 53454 23042 53506
rect 23042 53454 23044 53506
rect 22988 53452 23044 53454
rect 22652 53116 22708 53172
rect 23212 53676 23268 53732
rect 23324 53788 23380 53844
rect 23100 53116 23156 53172
rect 22652 52556 22708 52612
rect 22652 50764 22708 50820
rect 22540 49698 22596 49700
rect 22540 49646 22542 49698
rect 22542 49646 22594 49698
rect 22594 49646 22596 49698
rect 22540 49644 22596 49646
rect 22204 48748 22260 48804
rect 22092 48412 22148 48468
rect 21980 47404 22036 47460
rect 22428 48636 22484 48692
rect 22316 47346 22372 47348
rect 22316 47294 22318 47346
rect 22318 47294 22370 47346
rect 22370 47294 22372 47346
rect 22316 47292 22372 47294
rect 21624 47066 21680 47068
rect 21624 47014 21626 47066
rect 21626 47014 21678 47066
rect 21678 47014 21680 47066
rect 21624 47012 21680 47014
rect 21728 47066 21784 47068
rect 21728 47014 21730 47066
rect 21730 47014 21782 47066
rect 21782 47014 21784 47066
rect 21728 47012 21784 47014
rect 21832 47066 21888 47068
rect 21832 47014 21834 47066
rect 21834 47014 21886 47066
rect 21886 47014 21888 47066
rect 21832 47012 21888 47014
rect 21420 46674 21476 46676
rect 21420 46622 21422 46674
rect 21422 46622 21474 46674
rect 21474 46622 21476 46674
rect 21420 46620 21476 46622
rect 21644 46898 21700 46900
rect 21644 46846 21646 46898
rect 21646 46846 21698 46898
rect 21698 46846 21700 46898
rect 21644 46844 21700 46846
rect 22092 46786 22148 46788
rect 22092 46734 22094 46786
rect 22094 46734 22146 46786
rect 22146 46734 22148 46786
rect 22092 46732 22148 46734
rect 20860 45388 20916 45444
rect 21196 45106 21252 45108
rect 21196 45054 21198 45106
rect 21198 45054 21250 45106
rect 21250 45054 21252 45106
rect 21196 45052 21252 45054
rect 20076 42754 20132 42756
rect 20076 42702 20078 42754
rect 20078 42702 20130 42754
rect 20130 42702 20132 42754
rect 20076 42700 20132 42702
rect 19964 41916 20020 41972
rect 20300 42140 20356 42196
rect 20860 43484 20916 43540
rect 20748 42754 20804 42756
rect 20748 42702 20750 42754
rect 20750 42702 20802 42754
rect 20802 42702 20804 42754
rect 20748 42700 20804 42702
rect 19964 40908 20020 40964
rect 19628 40236 19684 40292
rect 20076 40796 20132 40852
rect 19964 40460 20020 40516
rect 19404 38668 19460 38724
rect 19852 39394 19908 39396
rect 19852 39342 19854 39394
rect 19854 39342 19906 39394
rect 19906 39342 19908 39394
rect 19852 39340 19908 39342
rect 19852 38946 19908 38948
rect 19852 38894 19854 38946
rect 19854 38894 19906 38946
rect 19906 38894 19908 38946
rect 19852 38892 19908 38894
rect 19740 38834 19796 38836
rect 19740 38782 19742 38834
rect 19742 38782 19794 38834
rect 19794 38782 19796 38834
rect 19740 38780 19796 38782
rect 19516 37100 19572 37156
rect 19404 36876 19460 36932
rect 19516 35532 19572 35588
rect 19852 37884 19908 37940
rect 19740 34972 19796 35028
rect 20076 38780 20132 38836
rect 20300 41970 20356 41972
rect 20300 41918 20302 41970
rect 20302 41918 20354 41970
rect 20354 41918 20356 41970
rect 20300 41916 20356 41918
rect 20412 41692 20468 41748
rect 20188 38444 20244 38500
rect 20300 40572 20356 40628
rect 20076 38108 20132 38164
rect 20412 40460 20468 40516
rect 20636 41804 20692 41860
rect 20972 42028 21028 42084
rect 21084 41970 21140 41972
rect 21084 41918 21086 41970
rect 21086 41918 21138 41970
rect 21138 41918 21140 41970
rect 21084 41916 21140 41918
rect 20972 41580 21028 41636
rect 20748 40348 20804 40404
rect 20636 40290 20692 40292
rect 20636 40238 20638 40290
rect 20638 40238 20690 40290
rect 20690 40238 20692 40290
rect 20636 40236 20692 40238
rect 20412 39730 20468 39732
rect 20412 39678 20414 39730
rect 20414 39678 20466 39730
rect 20466 39678 20468 39730
rect 20412 39676 20468 39678
rect 20748 39116 20804 39172
rect 20636 38668 20692 38724
rect 20748 38444 20804 38500
rect 21624 45498 21680 45500
rect 21624 45446 21626 45498
rect 21626 45446 21678 45498
rect 21678 45446 21680 45498
rect 21624 45444 21680 45446
rect 21728 45498 21784 45500
rect 21728 45446 21730 45498
rect 21730 45446 21782 45498
rect 21782 45446 21784 45498
rect 21728 45444 21784 45446
rect 21832 45498 21888 45500
rect 21832 45446 21834 45498
rect 21834 45446 21886 45498
rect 21886 45446 21888 45498
rect 21832 45444 21888 45446
rect 22092 45388 22148 45444
rect 21756 44994 21812 44996
rect 21756 44942 21758 44994
rect 21758 44942 21810 44994
rect 21810 44942 21812 44994
rect 21756 44940 21812 44942
rect 21420 44322 21476 44324
rect 21420 44270 21422 44322
rect 21422 44270 21474 44322
rect 21474 44270 21476 44322
rect 21420 44268 21476 44270
rect 21868 44156 21924 44212
rect 21980 44940 22036 44996
rect 21624 43930 21680 43932
rect 21624 43878 21626 43930
rect 21626 43878 21678 43930
rect 21678 43878 21680 43930
rect 21624 43876 21680 43878
rect 21728 43930 21784 43932
rect 21728 43878 21730 43930
rect 21730 43878 21782 43930
rect 21782 43878 21784 43930
rect 21728 43876 21784 43878
rect 21832 43930 21888 43932
rect 21832 43878 21834 43930
rect 21834 43878 21886 43930
rect 21886 43878 21888 43930
rect 21832 43876 21888 43878
rect 21308 43650 21364 43652
rect 21308 43598 21310 43650
rect 21310 43598 21362 43650
rect 21362 43598 21364 43650
rect 21308 43596 21364 43598
rect 21308 42476 21364 42532
rect 22316 44828 22372 44884
rect 22092 44044 22148 44100
rect 22092 43596 22148 43652
rect 21644 43148 21700 43204
rect 22204 42476 22260 42532
rect 21624 42362 21680 42364
rect 21624 42310 21626 42362
rect 21626 42310 21678 42362
rect 21678 42310 21680 42362
rect 21624 42308 21680 42310
rect 21728 42362 21784 42364
rect 21728 42310 21730 42362
rect 21730 42310 21782 42362
rect 21782 42310 21784 42362
rect 21728 42308 21784 42310
rect 21832 42362 21888 42364
rect 21832 42310 21834 42362
rect 21834 42310 21886 42362
rect 21886 42310 21888 42362
rect 21832 42308 21888 42310
rect 21868 42194 21924 42196
rect 21868 42142 21870 42194
rect 21870 42142 21922 42194
rect 21922 42142 21924 42194
rect 21868 42140 21924 42142
rect 22092 42028 22148 42084
rect 21420 41916 21476 41972
rect 21644 41746 21700 41748
rect 21644 41694 21646 41746
rect 21646 41694 21698 41746
rect 21698 41694 21700 41746
rect 21644 41692 21700 41694
rect 21420 41356 21476 41412
rect 21868 41132 21924 41188
rect 21420 40796 21476 40852
rect 22204 41746 22260 41748
rect 22204 41694 22206 41746
rect 22206 41694 22258 41746
rect 22258 41694 22260 41746
rect 22204 41692 22260 41694
rect 22316 41580 22372 41636
rect 23996 57820 24052 57876
rect 24332 61346 24388 61348
rect 24332 61294 24334 61346
rect 24334 61294 24386 61346
rect 24386 61294 24388 61346
rect 24332 61292 24388 61294
rect 24108 58156 24164 58212
rect 23884 57762 23940 57764
rect 23884 57710 23886 57762
rect 23886 57710 23938 57762
rect 23938 57710 23940 57762
rect 23884 57708 23940 57710
rect 23772 57372 23828 57428
rect 24108 57260 24164 57316
rect 24668 65772 24724 65828
rect 24668 64146 24724 64148
rect 24668 64094 24670 64146
rect 24670 64094 24722 64146
rect 24722 64094 24724 64146
rect 24668 64092 24724 64094
rect 24780 65436 24836 65492
rect 24780 63532 24836 63588
rect 24668 62188 24724 62244
rect 24556 60002 24612 60004
rect 24556 59950 24558 60002
rect 24558 59950 24610 60002
rect 24610 59950 24612 60002
rect 24556 59948 24612 59950
rect 24556 59388 24612 59444
rect 24444 59106 24500 59108
rect 24444 59054 24446 59106
rect 24446 59054 24498 59106
rect 24498 59054 24500 59106
rect 24444 59052 24500 59054
rect 24444 58268 24500 58324
rect 24444 57820 24500 57876
rect 24444 57372 24500 57428
rect 24668 57148 24724 57204
rect 24780 60172 24836 60228
rect 25340 73836 25396 73892
rect 25564 76972 25620 77028
rect 26012 77922 26068 77924
rect 26012 77870 26014 77922
rect 26014 77870 26066 77922
rect 26066 77870 26068 77922
rect 26012 77868 26068 77870
rect 25900 77084 25956 77140
rect 25676 75794 25732 75796
rect 25676 75742 25678 75794
rect 25678 75742 25730 75794
rect 25730 75742 25732 75794
rect 25676 75740 25732 75742
rect 26236 77084 26292 77140
rect 26684 76860 26740 76916
rect 26460 76748 26516 76804
rect 26348 76466 26404 76468
rect 26348 76414 26350 76466
rect 26350 76414 26402 76466
rect 26402 76414 26404 76466
rect 26348 76412 26404 76414
rect 26572 75628 26628 75684
rect 25676 74172 25732 74228
rect 25676 74002 25732 74004
rect 25676 73950 25678 74002
rect 25678 73950 25730 74002
rect 25730 73950 25732 74002
rect 25676 73948 25732 73950
rect 25452 73500 25508 73556
rect 25026 72938 25082 72940
rect 25026 72886 25028 72938
rect 25028 72886 25080 72938
rect 25080 72886 25082 72938
rect 25026 72884 25082 72886
rect 25130 72938 25186 72940
rect 25130 72886 25132 72938
rect 25132 72886 25184 72938
rect 25184 72886 25186 72938
rect 25130 72884 25186 72886
rect 25234 72938 25290 72940
rect 25234 72886 25236 72938
rect 25236 72886 25288 72938
rect 25288 72886 25290 72938
rect 25234 72884 25290 72886
rect 25004 72156 25060 72212
rect 25340 71484 25396 71540
rect 25026 71370 25082 71372
rect 25026 71318 25028 71370
rect 25028 71318 25080 71370
rect 25080 71318 25082 71370
rect 25026 71316 25082 71318
rect 25130 71370 25186 71372
rect 25130 71318 25132 71370
rect 25132 71318 25184 71370
rect 25184 71318 25186 71370
rect 25130 71316 25186 71318
rect 25234 71370 25290 71372
rect 25234 71318 25236 71370
rect 25236 71318 25288 71370
rect 25288 71318 25290 71370
rect 25234 71316 25290 71318
rect 26124 74786 26180 74788
rect 26124 74734 26126 74786
rect 26126 74734 26178 74786
rect 26178 74734 26180 74786
rect 26124 74732 26180 74734
rect 25788 72828 25844 72884
rect 25564 71820 25620 71876
rect 25676 72044 25732 72100
rect 25026 69802 25082 69804
rect 25026 69750 25028 69802
rect 25028 69750 25080 69802
rect 25080 69750 25082 69802
rect 25026 69748 25082 69750
rect 25130 69802 25186 69804
rect 25130 69750 25132 69802
rect 25132 69750 25184 69802
rect 25184 69750 25186 69802
rect 25130 69748 25186 69750
rect 25234 69802 25290 69804
rect 25234 69750 25236 69802
rect 25236 69750 25288 69802
rect 25288 69750 25290 69802
rect 25234 69748 25290 69750
rect 26348 74844 26404 74900
rect 26012 71036 26068 71092
rect 25788 70028 25844 70084
rect 25340 68684 25396 68740
rect 25788 69244 25844 69300
rect 25228 68514 25284 68516
rect 25228 68462 25230 68514
rect 25230 68462 25282 68514
rect 25282 68462 25284 68514
rect 25228 68460 25284 68462
rect 25026 68234 25082 68236
rect 25026 68182 25028 68234
rect 25028 68182 25080 68234
rect 25080 68182 25082 68234
rect 25026 68180 25082 68182
rect 25130 68234 25186 68236
rect 25130 68182 25132 68234
rect 25132 68182 25184 68234
rect 25184 68182 25186 68234
rect 25130 68180 25186 68182
rect 25234 68234 25290 68236
rect 25234 68182 25236 68234
rect 25236 68182 25288 68234
rect 25288 68182 25290 68234
rect 25234 68180 25290 68182
rect 25340 67116 25396 67172
rect 25228 66780 25284 66836
rect 25026 66666 25082 66668
rect 25026 66614 25028 66666
rect 25028 66614 25080 66666
rect 25080 66614 25082 66666
rect 25026 66612 25082 66614
rect 25130 66666 25186 66668
rect 25130 66614 25132 66666
rect 25132 66614 25184 66666
rect 25184 66614 25186 66666
rect 25130 66612 25186 66614
rect 25234 66666 25290 66668
rect 25234 66614 25236 66666
rect 25236 66614 25288 66666
rect 25288 66614 25290 66666
rect 25234 66612 25290 66614
rect 25452 65548 25508 65604
rect 25026 65098 25082 65100
rect 25026 65046 25028 65098
rect 25028 65046 25080 65098
rect 25080 65046 25082 65098
rect 25026 65044 25082 65046
rect 25130 65098 25186 65100
rect 25130 65046 25132 65098
rect 25132 65046 25184 65098
rect 25184 65046 25186 65098
rect 25130 65044 25186 65046
rect 25234 65098 25290 65100
rect 25234 65046 25236 65098
rect 25236 65046 25288 65098
rect 25288 65046 25290 65098
rect 25234 65044 25290 65046
rect 25564 65324 25620 65380
rect 26012 68684 26068 68740
rect 26012 67842 26068 67844
rect 26012 67790 26014 67842
rect 26014 67790 26066 67842
rect 26066 67790 26068 67842
rect 26012 67788 26068 67790
rect 25788 65490 25844 65492
rect 25788 65438 25790 65490
rect 25790 65438 25842 65490
rect 25842 65438 25844 65490
rect 25788 65436 25844 65438
rect 25564 64428 25620 64484
rect 25116 64092 25172 64148
rect 25676 64146 25732 64148
rect 25676 64094 25678 64146
rect 25678 64094 25730 64146
rect 25730 64094 25732 64146
rect 25676 64092 25732 64094
rect 26124 65324 26180 65380
rect 25788 63922 25844 63924
rect 25788 63870 25790 63922
rect 25790 63870 25842 63922
rect 25842 63870 25844 63922
rect 25788 63868 25844 63870
rect 25900 64428 25956 64484
rect 25676 63756 25732 63812
rect 25026 63530 25082 63532
rect 25026 63478 25028 63530
rect 25028 63478 25080 63530
rect 25080 63478 25082 63530
rect 25026 63476 25082 63478
rect 25130 63530 25186 63532
rect 25130 63478 25132 63530
rect 25132 63478 25184 63530
rect 25184 63478 25186 63530
rect 25130 63476 25186 63478
rect 25234 63530 25290 63532
rect 25234 63478 25236 63530
rect 25236 63478 25288 63530
rect 25288 63478 25290 63530
rect 25234 63476 25290 63478
rect 25228 62242 25284 62244
rect 25228 62190 25230 62242
rect 25230 62190 25282 62242
rect 25282 62190 25284 62242
rect 25228 62188 25284 62190
rect 25026 61962 25082 61964
rect 25026 61910 25028 61962
rect 25028 61910 25080 61962
rect 25080 61910 25082 61962
rect 25026 61908 25082 61910
rect 25130 61962 25186 61964
rect 25130 61910 25132 61962
rect 25132 61910 25184 61962
rect 25184 61910 25186 61962
rect 25130 61908 25186 61910
rect 25234 61962 25290 61964
rect 25234 61910 25236 61962
rect 25236 61910 25288 61962
rect 25288 61910 25290 61962
rect 25234 61908 25290 61910
rect 25340 61740 25396 61796
rect 25116 61180 25172 61236
rect 26012 64092 26068 64148
rect 25676 60844 25732 60900
rect 25026 60394 25082 60396
rect 25026 60342 25028 60394
rect 25028 60342 25080 60394
rect 25080 60342 25082 60394
rect 25026 60340 25082 60342
rect 25130 60394 25186 60396
rect 25130 60342 25132 60394
rect 25132 60342 25184 60394
rect 25184 60342 25186 60394
rect 25130 60340 25186 60342
rect 25234 60394 25290 60396
rect 25234 60342 25236 60394
rect 25236 60342 25288 60394
rect 25288 60342 25290 60394
rect 25234 60340 25290 60342
rect 25340 60002 25396 60004
rect 25340 59950 25342 60002
rect 25342 59950 25394 60002
rect 25394 59950 25396 60002
rect 25340 59948 25396 59950
rect 25026 58826 25082 58828
rect 25026 58774 25028 58826
rect 25028 58774 25080 58826
rect 25080 58774 25082 58826
rect 25026 58772 25082 58774
rect 25130 58826 25186 58828
rect 25130 58774 25132 58826
rect 25132 58774 25184 58826
rect 25184 58774 25186 58826
rect 25130 58772 25186 58774
rect 25234 58826 25290 58828
rect 25234 58774 25236 58826
rect 25236 58774 25288 58826
rect 25288 58774 25290 58826
rect 25234 58772 25290 58774
rect 25452 58828 25508 58884
rect 24892 58492 24948 58548
rect 24892 58210 24948 58212
rect 24892 58158 24894 58210
rect 24894 58158 24946 58210
rect 24946 58158 24948 58210
rect 24892 58156 24948 58158
rect 25340 57372 25396 57428
rect 25026 57258 25082 57260
rect 25026 57206 25028 57258
rect 25028 57206 25080 57258
rect 25080 57206 25082 57258
rect 25026 57204 25082 57206
rect 25130 57258 25186 57260
rect 25130 57206 25132 57258
rect 25132 57206 25184 57258
rect 25184 57206 25186 57258
rect 25130 57204 25186 57206
rect 25234 57258 25290 57260
rect 25234 57206 25236 57258
rect 25236 57206 25288 57258
rect 25288 57206 25290 57258
rect 25234 57204 25290 57206
rect 23996 56924 24052 56980
rect 24556 56924 24612 56980
rect 24332 56588 24388 56644
rect 23772 54572 23828 54628
rect 23884 54796 23940 54852
rect 23660 54460 23716 54516
rect 23772 54012 23828 54068
rect 24108 54684 24164 54740
rect 24220 55692 24276 55748
rect 24556 55132 24612 55188
rect 24668 54908 24724 54964
rect 24108 53842 24164 53844
rect 24108 53790 24110 53842
rect 24110 53790 24162 53842
rect 24162 53790 24164 53842
rect 24108 53788 24164 53790
rect 23996 53618 24052 53620
rect 23996 53566 23998 53618
rect 23998 53566 24050 53618
rect 24050 53566 24052 53618
rect 23996 53564 24052 53566
rect 23884 53452 23940 53508
rect 24220 53506 24276 53508
rect 24220 53454 24222 53506
rect 24222 53454 24274 53506
rect 24274 53454 24276 53506
rect 24220 53452 24276 53454
rect 24556 53340 24612 53396
rect 25564 57708 25620 57764
rect 25564 56978 25620 56980
rect 25564 56926 25566 56978
rect 25566 56926 25618 56978
rect 25618 56926 25620 56978
rect 25564 56924 25620 56926
rect 25676 58604 25732 58660
rect 25676 56140 25732 56196
rect 25900 63196 25956 63252
rect 25900 59052 25956 59108
rect 25900 58492 25956 58548
rect 25900 56700 25956 56756
rect 26012 56642 26068 56644
rect 26012 56590 26014 56642
rect 26014 56590 26066 56642
rect 26066 56590 26068 56642
rect 26012 56588 26068 56590
rect 25788 56028 25844 56084
rect 25676 55916 25732 55972
rect 25026 55690 25082 55692
rect 25026 55638 25028 55690
rect 25028 55638 25080 55690
rect 25080 55638 25082 55690
rect 25026 55636 25082 55638
rect 25130 55690 25186 55692
rect 25130 55638 25132 55690
rect 25132 55638 25184 55690
rect 25184 55638 25186 55690
rect 25130 55636 25186 55638
rect 25234 55690 25290 55692
rect 25234 55638 25236 55690
rect 25236 55638 25288 55690
rect 25288 55638 25290 55690
rect 25234 55636 25290 55638
rect 25116 55132 25172 55188
rect 25340 55244 25396 55300
rect 26012 55970 26068 55972
rect 26012 55918 26014 55970
rect 26014 55918 26066 55970
rect 26066 55918 26068 55970
rect 26012 55916 26068 55918
rect 27356 77138 27412 77140
rect 27356 77086 27358 77138
rect 27358 77086 27410 77138
rect 27410 77086 27412 77138
rect 27356 77084 27412 77086
rect 27020 76860 27076 76916
rect 27132 76972 27188 77028
rect 26796 76412 26852 76468
rect 26796 74396 26852 74452
rect 27020 76690 27076 76692
rect 27020 76638 27022 76690
rect 27022 76638 27074 76690
rect 27074 76638 27076 76690
rect 27020 76636 27076 76638
rect 27020 75682 27076 75684
rect 27020 75630 27022 75682
rect 27022 75630 27074 75682
rect 27074 75630 27076 75682
rect 27020 75628 27076 75630
rect 27132 75516 27188 75572
rect 28140 78930 28196 78932
rect 28140 78878 28142 78930
rect 28142 78878 28194 78930
rect 28194 78878 28196 78930
rect 28140 78876 28196 78878
rect 28428 78426 28484 78428
rect 28428 78374 28430 78426
rect 28430 78374 28482 78426
rect 28482 78374 28484 78426
rect 28428 78372 28484 78374
rect 28532 78426 28588 78428
rect 28532 78374 28534 78426
rect 28534 78374 28586 78426
rect 28586 78374 28588 78426
rect 28532 78372 28588 78374
rect 28636 78426 28692 78428
rect 28636 78374 28638 78426
rect 28638 78374 28690 78426
rect 28690 78374 28692 78426
rect 28636 78372 28692 78374
rect 28140 76972 28196 77028
rect 28428 76858 28484 76860
rect 28428 76806 28430 76858
rect 28430 76806 28482 76858
rect 28482 76806 28484 76858
rect 28428 76804 28484 76806
rect 28532 76858 28588 76860
rect 28532 76806 28534 76858
rect 28534 76806 28586 76858
rect 28586 76806 28588 76858
rect 28532 76804 28588 76806
rect 28636 76858 28692 76860
rect 28636 76806 28638 76858
rect 28638 76806 28690 76858
rect 28690 76806 28692 76858
rect 28636 76804 28692 76806
rect 27580 76412 27636 76468
rect 27356 75628 27412 75684
rect 26908 75404 26964 75460
rect 26572 74114 26628 74116
rect 26572 74062 26574 74114
rect 26574 74062 26626 74114
rect 26626 74062 26628 74114
rect 26572 74060 26628 74062
rect 27020 74114 27076 74116
rect 27020 74062 27022 74114
rect 27022 74062 27074 74114
rect 27074 74062 27076 74114
rect 27020 74060 27076 74062
rect 27804 75458 27860 75460
rect 27804 75406 27806 75458
rect 27806 75406 27858 75458
rect 27858 75406 27860 75458
rect 27804 75404 27860 75406
rect 28428 75290 28484 75292
rect 28428 75238 28430 75290
rect 28430 75238 28482 75290
rect 28482 75238 28484 75290
rect 28428 75236 28484 75238
rect 28532 75290 28588 75292
rect 28532 75238 28534 75290
rect 28534 75238 28586 75290
rect 28586 75238 28588 75290
rect 28532 75236 28588 75238
rect 28636 75290 28692 75292
rect 28636 75238 28638 75290
rect 28638 75238 28690 75290
rect 28690 75238 28692 75290
rect 28636 75236 28692 75238
rect 27132 74002 27188 74004
rect 27132 73950 27134 74002
rect 27134 73950 27186 74002
rect 27186 73950 27188 74002
rect 27132 73948 27188 73950
rect 26460 73500 26516 73556
rect 26460 72828 26516 72884
rect 26684 73612 26740 73668
rect 27580 74284 27636 74340
rect 28028 74172 28084 74228
rect 27244 73612 27300 73668
rect 26684 72044 26740 72100
rect 26348 69298 26404 69300
rect 26348 69246 26350 69298
rect 26350 69246 26402 69298
rect 26402 69246 26404 69298
rect 26348 69244 26404 69246
rect 26684 71036 26740 71092
rect 27020 71036 27076 71092
rect 27468 71986 27524 71988
rect 27468 71934 27470 71986
rect 27470 71934 27522 71986
rect 27522 71934 27524 71986
rect 27468 71932 27524 71934
rect 27132 70364 27188 70420
rect 26572 67340 26628 67396
rect 26348 64652 26404 64708
rect 26572 64092 26628 64148
rect 26460 63644 26516 63700
rect 26348 63196 26404 63252
rect 26572 62860 26628 62916
rect 26236 61740 26292 61796
rect 26796 70028 26852 70084
rect 27468 70082 27524 70084
rect 27468 70030 27470 70082
rect 27470 70030 27522 70082
rect 27522 70030 27524 70082
rect 27468 70028 27524 70030
rect 26908 69970 26964 69972
rect 26908 69918 26910 69970
rect 26910 69918 26962 69970
rect 26962 69918 26964 69970
rect 26908 69916 26964 69918
rect 28140 73948 28196 74004
rect 28252 73836 28308 73892
rect 27244 68348 27300 68404
rect 27356 67788 27412 67844
rect 26796 67116 26852 67172
rect 27356 67340 27412 67396
rect 27132 66780 27188 66836
rect 26908 65490 26964 65492
rect 26908 65438 26910 65490
rect 26910 65438 26962 65490
rect 26962 65438 26964 65490
rect 26908 65436 26964 65438
rect 27356 65378 27412 65380
rect 27356 65326 27358 65378
rect 27358 65326 27410 65378
rect 27410 65326 27412 65378
rect 27356 65324 27412 65326
rect 27020 64876 27076 64932
rect 27132 63810 27188 63812
rect 27132 63758 27134 63810
rect 27134 63758 27186 63810
rect 27186 63758 27188 63810
rect 27132 63756 27188 63758
rect 27244 63644 27300 63700
rect 26796 63532 26852 63588
rect 27020 63250 27076 63252
rect 27020 63198 27022 63250
rect 27022 63198 27074 63250
rect 27074 63198 27076 63250
rect 27020 63196 27076 63198
rect 26796 63084 26852 63140
rect 27468 64034 27524 64036
rect 27468 63982 27470 64034
rect 27470 63982 27522 64034
rect 27522 63982 27524 64034
rect 27468 63980 27524 63982
rect 27244 62972 27300 63028
rect 27356 62860 27412 62916
rect 28428 73722 28484 73724
rect 28428 73670 28430 73722
rect 28430 73670 28482 73722
rect 28482 73670 28484 73722
rect 28428 73668 28484 73670
rect 28532 73722 28588 73724
rect 28532 73670 28534 73722
rect 28534 73670 28586 73722
rect 28586 73670 28588 73722
rect 28532 73668 28588 73670
rect 28636 73722 28692 73724
rect 28636 73670 28638 73722
rect 28638 73670 28690 73722
rect 28690 73670 28692 73722
rect 28636 73668 28692 73670
rect 28428 72154 28484 72156
rect 28428 72102 28430 72154
rect 28430 72102 28482 72154
rect 28482 72102 28484 72154
rect 28428 72100 28484 72102
rect 28532 72154 28588 72156
rect 28532 72102 28534 72154
rect 28534 72102 28586 72154
rect 28586 72102 28588 72154
rect 28532 72100 28588 72102
rect 28636 72154 28692 72156
rect 28636 72102 28638 72154
rect 28638 72102 28690 72154
rect 28690 72102 28692 72154
rect 28636 72100 28692 72102
rect 28140 71090 28196 71092
rect 28140 71038 28142 71090
rect 28142 71038 28194 71090
rect 28194 71038 28196 71090
rect 28140 71036 28196 71038
rect 27916 70418 27972 70420
rect 27916 70366 27918 70418
rect 27918 70366 27970 70418
rect 27970 70366 27972 70418
rect 27916 70364 27972 70366
rect 27804 69298 27860 69300
rect 27804 69246 27806 69298
rect 27806 69246 27858 69298
rect 27858 69246 27860 69298
rect 27804 69244 27860 69246
rect 28428 70586 28484 70588
rect 28428 70534 28430 70586
rect 28430 70534 28482 70586
rect 28482 70534 28484 70586
rect 28428 70532 28484 70534
rect 28532 70586 28588 70588
rect 28532 70534 28534 70586
rect 28534 70534 28586 70586
rect 28586 70534 28588 70586
rect 28532 70532 28588 70534
rect 28636 70586 28692 70588
rect 28636 70534 28638 70586
rect 28638 70534 28690 70586
rect 28690 70534 28692 70586
rect 28636 70532 28692 70534
rect 28428 69018 28484 69020
rect 28428 68966 28430 69018
rect 28430 68966 28482 69018
rect 28482 68966 28484 69018
rect 28428 68964 28484 68966
rect 28532 69018 28588 69020
rect 28532 68966 28534 69018
rect 28534 68966 28586 69018
rect 28586 68966 28588 69018
rect 28532 68964 28588 68966
rect 28636 69018 28692 69020
rect 28636 68966 28638 69018
rect 28638 68966 28690 69018
rect 28690 68966 28692 69018
rect 28636 68964 28692 68966
rect 28428 67450 28484 67452
rect 28428 67398 28430 67450
rect 28430 67398 28482 67450
rect 28482 67398 28484 67450
rect 28428 67396 28484 67398
rect 28532 67450 28588 67452
rect 28532 67398 28534 67450
rect 28534 67398 28586 67450
rect 28586 67398 28588 67450
rect 28532 67396 28588 67398
rect 28636 67450 28692 67452
rect 28636 67398 28638 67450
rect 28638 67398 28690 67450
rect 28690 67398 28692 67450
rect 28636 67396 28692 67398
rect 28428 65882 28484 65884
rect 28428 65830 28430 65882
rect 28430 65830 28482 65882
rect 28482 65830 28484 65882
rect 28428 65828 28484 65830
rect 28532 65882 28588 65884
rect 28532 65830 28534 65882
rect 28534 65830 28586 65882
rect 28586 65830 28588 65882
rect 28532 65828 28588 65830
rect 28636 65882 28692 65884
rect 28636 65830 28638 65882
rect 28638 65830 28690 65882
rect 28690 65830 28692 65882
rect 28636 65828 28692 65830
rect 27916 65548 27972 65604
rect 27804 65490 27860 65492
rect 27804 65438 27806 65490
rect 27806 65438 27858 65490
rect 27858 65438 27860 65490
rect 27804 65436 27860 65438
rect 28028 64034 28084 64036
rect 28028 63982 28030 64034
rect 28030 63982 28082 64034
rect 28082 63982 28084 64034
rect 28028 63980 28084 63982
rect 28428 64314 28484 64316
rect 28428 64262 28430 64314
rect 28430 64262 28482 64314
rect 28482 64262 28484 64314
rect 28428 64260 28484 64262
rect 28532 64314 28588 64316
rect 28532 64262 28534 64314
rect 28534 64262 28586 64314
rect 28586 64262 28588 64314
rect 28532 64260 28588 64262
rect 28636 64314 28692 64316
rect 28636 64262 28638 64314
rect 28638 64262 28690 64314
rect 28690 64262 28692 64314
rect 28636 64260 28692 64262
rect 28140 63644 28196 63700
rect 28428 62746 28484 62748
rect 28428 62694 28430 62746
rect 28430 62694 28482 62746
rect 28482 62694 28484 62746
rect 28428 62692 28484 62694
rect 28532 62746 28588 62748
rect 28532 62694 28534 62746
rect 28534 62694 28586 62746
rect 28586 62694 28588 62746
rect 28532 62692 28588 62694
rect 28636 62746 28692 62748
rect 28636 62694 28638 62746
rect 28638 62694 28690 62746
rect 28690 62694 28692 62746
rect 28636 62692 28692 62694
rect 26908 61740 26964 61796
rect 26684 60844 26740 60900
rect 26236 59388 26292 59444
rect 26348 60060 26404 60116
rect 26236 59218 26292 59220
rect 26236 59166 26238 59218
rect 26238 59166 26290 59218
rect 26290 59166 26292 59218
rect 26236 59164 26292 59166
rect 26236 57762 26292 57764
rect 26236 57710 26238 57762
rect 26238 57710 26290 57762
rect 26290 57710 26292 57762
rect 26236 57708 26292 57710
rect 26684 60172 26740 60228
rect 26572 59164 26628 59220
rect 26460 57650 26516 57652
rect 26460 57598 26462 57650
rect 26462 57598 26514 57650
rect 26514 57598 26516 57650
rect 26460 57596 26516 57598
rect 26460 57372 26516 57428
rect 25564 55298 25620 55300
rect 25564 55246 25566 55298
rect 25566 55246 25618 55298
rect 25618 55246 25620 55298
rect 25564 55244 25620 55246
rect 25788 55186 25844 55188
rect 25788 55134 25790 55186
rect 25790 55134 25842 55186
rect 25842 55134 25844 55186
rect 25788 55132 25844 55134
rect 25340 54684 25396 54740
rect 25788 54796 25844 54852
rect 25676 54572 25732 54628
rect 25340 54402 25396 54404
rect 25340 54350 25342 54402
rect 25342 54350 25394 54402
rect 25394 54350 25396 54402
rect 25340 54348 25396 54350
rect 25026 54122 25082 54124
rect 25026 54070 25028 54122
rect 25028 54070 25080 54122
rect 25080 54070 25082 54122
rect 25026 54068 25082 54070
rect 25130 54122 25186 54124
rect 25130 54070 25132 54122
rect 25132 54070 25184 54122
rect 25184 54070 25186 54122
rect 25130 54068 25186 54070
rect 25234 54122 25290 54124
rect 25234 54070 25236 54122
rect 25236 54070 25288 54122
rect 25288 54070 25290 54122
rect 25234 54068 25290 54070
rect 25116 53116 25172 53172
rect 23660 52892 23716 52948
rect 24556 52946 24612 52948
rect 24556 52894 24558 52946
rect 24558 52894 24610 52946
rect 24610 52894 24612 52946
rect 24556 52892 24612 52894
rect 24332 52332 24388 52388
rect 23436 51938 23492 51940
rect 23436 51886 23438 51938
rect 23438 51886 23490 51938
rect 23490 51886 23492 51938
rect 23436 51884 23492 51886
rect 22988 51324 23044 51380
rect 23212 51212 23268 51268
rect 22764 47516 22820 47572
rect 22876 50764 22932 50820
rect 22652 46172 22708 46228
rect 22988 49196 23044 49252
rect 23548 51378 23604 51380
rect 23548 51326 23550 51378
rect 23550 51326 23602 51378
rect 23602 51326 23604 51378
rect 23548 51324 23604 51326
rect 23436 50876 23492 50932
rect 23436 49644 23492 49700
rect 23660 49026 23716 49028
rect 23660 48974 23662 49026
rect 23662 48974 23714 49026
rect 23714 48974 23716 49026
rect 23660 48972 23716 48974
rect 23212 47068 23268 47124
rect 23436 47516 23492 47572
rect 23548 47458 23604 47460
rect 23548 47406 23550 47458
rect 23550 47406 23602 47458
rect 23602 47406 23604 47458
rect 23548 47404 23604 47406
rect 23324 47292 23380 47348
rect 23100 46844 23156 46900
rect 22988 46732 23044 46788
rect 23100 46674 23156 46676
rect 23100 46622 23102 46674
rect 23102 46622 23154 46674
rect 23154 46622 23156 46674
rect 23100 46620 23156 46622
rect 22764 46060 22820 46116
rect 23324 46508 23380 46564
rect 23100 45612 23156 45668
rect 22988 44268 23044 44324
rect 22764 44156 22820 44212
rect 22540 43260 22596 43316
rect 22540 42700 22596 42756
rect 22316 40962 22372 40964
rect 22316 40910 22318 40962
rect 22318 40910 22370 40962
rect 22370 40910 22372 40962
rect 22316 40908 22372 40910
rect 21624 40794 21680 40796
rect 21624 40742 21626 40794
rect 21626 40742 21678 40794
rect 21678 40742 21680 40794
rect 21624 40740 21680 40742
rect 21728 40794 21784 40796
rect 21728 40742 21730 40794
rect 21730 40742 21782 40794
rect 21782 40742 21784 40794
rect 21728 40740 21784 40742
rect 21832 40794 21888 40796
rect 21832 40742 21834 40794
rect 21834 40742 21886 40794
rect 21886 40742 21888 40794
rect 21832 40740 21888 40742
rect 21980 40514 22036 40516
rect 21980 40462 21982 40514
rect 21982 40462 22034 40514
rect 22034 40462 22036 40514
rect 21980 40460 22036 40462
rect 21308 39340 21364 39396
rect 21868 39394 21924 39396
rect 21868 39342 21870 39394
rect 21870 39342 21922 39394
rect 21922 39342 21924 39394
rect 21868 39340 21924 39342
rect 21420 39228 21476 39284
rect 21624 39226 21680 39228
rect 21624 39174 21626 39226
rect 21626 39174 21678 39226
rect 21678 39174 21680 39226
rect 21624 39172 21680 39174
rect 21728 39226 21784 39228
rect 21728 39174 21730 39226
rect 21730 39174 21782 39226
rect 21782 39174 21784 39226
rect 21728 39172 21784 39174
rect 21832 39226 21888 39228
rect 21832 39174 21834 39226
rect 21834 39174 21886 39226
rect 21886 39174 21888 39226
rect 21832 39172 21888 39174
rect 21756 38780 21812 38836
rect 21196 38444 21252 38500
rect 20300 37548 20356 37604
rect 20076 37324 20132 37380
rect 19964 36876 20020 36932
rect 19852 36204 19908 36260
rect 20524 37548 20580 37604
rect 20412 37378 20468 37380
rect 20412 37326 20414 37378
rect 20414 37326 20466 37378
rect 20466 37326 20468 37378
rect 20412 37324 20468 37326
rect 20300 35586 20356 35588
rect 20300 35534 20302 35586
rect 20302 35534 20354 35586
rect 20354 35534 20356 35586
rect 20300 35532 20356 35534
rect 20188 34914 20244 34916
rect 20188 34862 20190 34914
rect 20190 34862 20242 34914
rect 20242 34862 20244 34914
rect 20188 34860 20244 34862
rect 19852 34636 19908 34692
rect 19740 34524 19796 34580
rect 20076 34300 20132 34356
rect 20188 34636 20244 34692
rect 19852 34130 19908 34132
rect 19852 34078 19854 34130
rect 19854 34078 19906 34130
rect 19906 34078 19908 34130
rect 19852 34076 19908 34078
rect 19964 33628 20020 33684
rect 20188 33516 20244 33572
rect 20188 33346 20244 33348
rect 20188 33294 20190 33346
rect 20190 33294 20242 33346
rect 20242 33294 20244 33346
rect 20188 33292 20244 33294
rect 19964 32956 20020 33012
rect 20188 33068 20244 33124
rect 19516 32562 19572 32564
rect 19516 32510 19518 32562
rect 19518 32510 19570 32562
rect 19570 32510 19572 32562
rect 19516 32508 19572 32510
rect 19964 32396 20020 32452
rect 19404 31778 19460 31780
rect 19404 31726 19406 31778
rect 19406 31726 19458 31778
rect 19458 31726 19460 31778
rect 19404 31724 19460 31726
rect 19516 31666 19572 31668
rect 19516 31614 19518 31666
rect 19518 31614 19570 31666
rect 19570 31614 19572 31666
rect 19516 31612 19572 31614
rect 19180 31276 19236 31332
rect 19516 31218 19572 31220
rect 19516 31166 19518 31218
rect 19518 31166 19570 31218
rect 19570 31166 19572 31218
rect 19516 31164 19572 31166
rect 18956 31052 19012 31108
rect 19852 31276 19908 31332
rect 19068 30940 19124 30996
rect 18508 29202 18564 29204
rect 18508 29150 18510 29202
rect 18510 29150 18562 29202
rect 18562 29150 18564 29202
rect 18508 29148 18564 29150
rect 18222 29034 18278 29036
rect 18222 28982 18224 29034
rect 18224 28982 18276 29034
rect 18276 28982 18278 29034
rect 18222 28980 18278 28982
rect 18326 29034 18382 29036
rect 18326 28982 18328 29034
rect 18328 28982 18380 29034
rect 18380 28982 18382 29034
rect 18326 28980 18382 28982
rect 18430 29034 18486 29036
rect 18430 28982 18432 29034
rect 18432 28982 18484 29034
rect 18484 28982 18486 29034
rect 18430 28980 18486 28982
rect 18396 28700 18452 28756
rect 17388 27580 17444 27636
rect 16380 26796 16436 26852
rect 17724 27468 17780 27524
rect 17388 27020 17444 27076
rect 16716 26124 16772 26180
rect 17388 26402 17444 26404
rect 17388 26350 17390 26402
rect 17390 26350 17442 26402
rect 17442 26350 17444 26402
rect 17388 26348 17444 26350
rect 16044 25228 16100 25284
rect 15708 24946 15764 24948
rect 15708 24894 15710 24946
rect 15710 24894 15762 24946
rect 15762 24894 15764 24946
rect 15708 24892 15764 24894
rect 15484 22876 15540 22932
rect 15708 23826 15764 23828
rect 15708 23774 15710 23826
rect 15710 23774 15762 23826
rect 15762 23774 15764 23826
rect 15708 23772 15764 23774
rect 15260 22764 15316 22820
rect 15596 22764 15652 22820
rect 15708 22652 15764 22708
rect 15820 23100 15876 23156
rect 16268 24892 16324 24948
rect 16156 24108 16212 24164
rect 16268 24556 16324 24612
rect 16716 23938 16772 23940
rect 16716 23886 16718 23938
rect 16718 23886 16770 23938
rect 16770 23886 16772 23938
rect 16716 23884 16772 23886
rect 16604 23772 16660 23828
rect 16380 23100 16436 23156
rect 15148 22092 15204 22148
rect 15596 22146 15652 22148
rect 15596 22094 15598 22146
rect 15598 22094 15650 22146
rect 15650 22094 15652 22146
rect 15596 22092 15652 22094
rect 14820 21978 14876 21980
rect 14820 21926 14822 21978
rect 14822 21926 14874 21978
rect 14874 21926 14876 21978
rect 14820 21924 14876 21926
rect 14924 21978 14980 21980
rect 14924 21926 14926 21978
rect 14926 21926 14978 21978
rect 14978 21926 14980 21978
rect 14924 21924 14980 21926
rect 15028 21978 15084 21980
rect 15028 21926 15030 21978
rect 15030 21926 15082 21978
rect 15082 21926 15084 21978
rect 15028 21924 15084 21926
rect 15148 21644 15204 21700
rect 15036 21474 15092 21476
rect 15036 21422 15038 21474
rect 15038 21422 15090 21474
rect 15090 21422 15092 21474
rect 15036 21420 15092 21422
rect 14820 20410 14876 20412
rect 14820 20358 14822 20410
rect 14822 20358 14874 20410
rect 14874 20358 14876 20410
rect 14820 20356 14876 20358
rect 14924 20410 14980 20412
rect 14924 20358 14926 20410
rect 14926 20358 14978 20410
rect 14978 20358 14980 20410
rect 14924 20356 14980 20358
rect 15028 20410 15084 20412
rect 15028 20358 15030 20410
rect 15030 20358 15082 20410
rect 15082 20358 15084 20410
rect 15028 20356 15084 20358
rect 13916 20076 13972 20132
rect 13804 19234 13860 19236
rect 13804 19182 13806 19234
rect 13806 19182 13858 19234
rect 13858 19182 13860 19234
rect 13804 19180 13860 19182
rect 12796 18956 12852 19012
rect 12572 17612 12628 17668
rect 12124 16268 12180 16324
rect 12348 17500 12404 17556
rect 12460 17442 12516 17444
rect 12460 17390 12462 17442
rect 12462 17390 12514 17442
rect 12514 17390 12516 17442
rect 12460 17388 12516 17390
rect 12460 15874 12516 15876
rect 12460 15822 12462 15874
rect 12462 15822 12514 15874
rect 12514 15822 12516 15874
rect 12460 15820 12516 15822
rect 12348 15708 12404 15764
rect 13580 19010 13636 19012
rect 13580 18958 13582 19010
rect 13582 18958 13634 19010
rect 13634 18958 13636 19010
rect 13580 18956 13636 18958
rect 13580 18396 13636 18452
rect 12908 17276 12964 17332
rect 12796 16044 12852 16100
rect 12796 15820 12852 15876
rect 13692 17948 13748 18004
rect 14028 19068 14084 19124
rect 14028 17666 14084 17668
rect 14028 17614 14030 17666
rect 14030 17614 14082 17666
rect 14082 17614 14084 17666
rect 14028 17612 14084 17614
rect 14252 17276 14308 17332
rect 14252 16828 14308 16884
rect 13804 16156 13860 16212
rect 13020 15708 13076 15764
rect 13356 15538 13412 15540
rect 13356 15486 13358 15538
rect 13358 15486 13410 15538
rect 13410 15486 13412 15538
rect 13356 15484 13412 15486
rect 11452 12796 11508 12852
rect 11788 12738 11844 12740
rect 11788 12686 11790 12738
rect 11790 12686 11842 12738
rect 11842 12686 11844 12738
rect 11788 12684 11844 12686
rect 11004 12290 11060 12292
rect 11004 12238 11006 12290
rect 11006 12238 11058 12290
rect 11058 12238 11060 12290
rect 11004 12236 11060 12238
rect 11418 11786 11474 11788
rect 11418 11734 11420 11786
rect 11420 11734 11472 11786
rect 11472 11734 11474 11786
rect 11418 11732 11474 11734
rect 11522 11786 11578 11788
rect 11522 11734 11524 11786
rect 11524 11734 11576 11786
rect 11576 11734 11578 11786
rect 11522 11732 11578 11734
rect 11626 11786 11682 11788
rect 11626 11734 11628 11786
rect 11628 11734 11680 11786
rect 11680 11734 11682 11786
rect 11626 11732 11682 11734
rect 11228 11282 11284 11284
rect 11228 11230 11230 11282
rect 11230 11230 11282 11282
rect 11282 11230 11284 11282
rect 11228 11228 11284 11230
rect 10780 10780 10836 10836
rect 11676 11116 11732 11172
rect 12012 14252 12068 14308
rect 12684 13356 12740 13412
rect 12236 13132 12292 13188
rect 12124 13020 12180 13076
rect 11900 11564 11956 11620
rect 11788 10892 11844 10948
rect 11900 11340 11956 11396
rect 12124 10834 12180 10836
rect 12124 10782 12126 10834
rect 12126 10782 12178 10834
rect 12178 10782 12180 10834
rect 12124 10780 12180 10782
rect 11116 10610 11172 10612
rect 11116 10558 11118 10610
rect 11118 10558 11170 10610
rect 11170 10558 11172 10610
rect 11116 10556 11172 10558
rect 11788 10610 11844 10612
rect 11788 10558 11790 10610
rect 11790 10558 11842 10610
rect 11842 10558 11844 10610
rect 11788 10556 11844 10558
rect 11418 10218 11474 10220
rect 11418 10166 11420 10218
rect 11420 10166 11472 10218
rect 11472 10166 11474 10218
rect 11418 10164 11474 10166
rect 11522 10218 11578 10220
rect 11522 10166 11524 10218
rect 11524 10166 11576 10218
rect 11576 10166 11578 10218
rect 11522 10164 11578 10166
rect 11626 10218 11682 10220
rect 11626 10166 11628 10218
rect 11628 10166 11680 10218
rect 11680 10166 11682 10218
rect 11626 10164 11682 10166
rect 9772 9826 9828 9828
rect 9772 9774 9774 9826
rect 9774 9774 9826 9826
rect 9826 9774 9828 9826
rect 9772 9772 9828 9774
rect 6300 8428 6356 8484
rect 6188 7644 6244 7700
rect 6636 8092 6692 8148
rect 7420 7868 7476 7924
rect 8092 8146 8148 8148
rect 8092 8094 8094 8146
rect 8094 8094 8146 8146
rect 8146 8094 8148 8146
rect 8092 8092 8148 8094
rect 5404 6636 5460 6692
rect 4060 6524 4116 6580
rect 3836 6076 3892 6132
rect 2380 1762 2436 1764
rect 2380 1710 2382 1762
rect 2382 1710 2434 1762
rect 2434 1710 2436 1762
rect 2380 1708 2436 1710
rect 3276 1874 3332 1876
rect 3276 1822 3278 1874
rect 3278 1822 3330 1874
rect 3330 1822 3332 1874
rect 3276 1820 3332 1822
rect 4396 6578 4452 6580
rect 4396 6526 4398 6578
rect 4398 6526 4450 6578
rect 4450 6526 4452 6578
rect 4396 6524 4452 6526
rect 8016 7866 8072 7868
rect 8016 7814 8018 7866
rect 8018 7814 8070 7866
rect 8070 7814 8072 7866
rect 8016 7812 8072 7814
rect 8120 7866 8176 7868
rect 8120 7814 8122 7866
rect 8122 7814 8174 7866
rect 8174 7814 8176 7866
rect 8120 7812 8176 7814
rect 8224 7866 8280 7868
rect 8224 7814 8226 7866
rect 8226 7814 8278 7866
rect 8278 7814 8280 7866
rect 8224 7812 8280 7814
rect 12572 11340 12628 11396
rect 12460 11170 12516 11172
rect 12460 11118 12462 11170
rect 12462 11118 12514 11170
rect 12514 11118 12516 11170
rect 12460 11116 12516 11118
rect 13692 15874 13748 15876
rect 13692 15822 13694 15874
rect 13694 15822 13746 15874
rect 13746 15822 13748 15874
rect 13692 15820 13748 15822
rect 14140 14252 14196 14308
rect 15484 20076 15540 20132
rect 15708 20860 15764 20916
rect 16044 22316 16100 22372
rect 17500 26178 17556 26180
rect 17500 26126 17502 26178
rect 17502 26126 17554 26178
rect 17554 26126 17556 26178
rect 17500 26124 17556 26126
rect 16940 25116 16996 25172
rect 17052 24556 17108 24612
rect 16940 24162 16996 24164
rect 16940 24110 16942 24162
rect 16942 24110 16994 24162
rect 16994 24110 16996 24162
rect 16940 24108 16996 24110
rect 16828 23042 16884 23044
rect 16828 22990 16830 23042
rect 16830 22990 16882 23042
rect 16882 22990 16884 23042
rect 16828 22988 16884 22990
rect 16604 22482 16660 22484
rect 16604 22430 16606 22482
rect 16606 22430 16658 22482
rect 16658 22430 16660 22482
rect 16604 22428 16660 22430
rect 16492 21644 16548 21700
rect 16604 20860 16660 20916
rect 15372 19852 15428 19908
rect 15372 19346 15428 19348
rect 15372 19294 15374 19346
rect 15374 19294 15426 19346
rect 15426 19294 15428 19346
rect 15372 19292 15428 19294
rect 15596 19122 15652 19124
rect 15596 19070 15598 19122
rect 15598 19070 15650 19122
rect 15650 19070 15652 19122
rect 15596 19068 15652 19070
rect 14588 17948 14644 18004
rect 16044 20130 16100 20132
rect 16044 20078 16046 20130
rect 16046 20078 16098 20130
rect 16098 20078 16100 20130
rect 16044 20076 16100 20078
rect 16268 20018 16324 20020
rect 16268 19966 16270 20018
rect 16270 19966 16322 20018
rect 16322 19966 16324 20018
rect 16268 19964 16324 19966
rect 16604 19404 16660 19460
rect 16044 19068 16100 19124
rect 16492 19068 16548 19124
rect 15820 18956 15876 19012
rect 14820 18842 14876 18844
rect 14820 18790 14822 18842
rect 14822 18790 14874 18842
rect 14874 18790 14876 18842
rect 14820 18788 14876 18790
rect 14924 18842 14980 18844
rect 14924 18790 14926 18842
rect 14926 18790 14978 18842
rect 14978 18790 14980 18842
rect 14924 18788 14980 18790
rect 15028 18842 15084 18844
rect 15028 18790 15030 18842
rect 15030 18790 15082 18842
rect 15082 18790 15084 18842
rect 15028 18788 15084 18790
rect 16268 18284 16324 18340
rect 15820 18172 15876 18228
rect 14588 17612 14644 17668
rect 15260 17778 15316 17780
rect 15260 17726 15262 17778
rect 15262 17726 15314 17778
rect 15314 17726 15316 17778
rect 15260 17724 15316 17726
rect 14924 17666 14980 17668
rect 14924 17614 14926 17666
rect 14926 17614 14978 17666
rect 14978 17614 14980 17666
rect 14924 17612 14980 17614
rect 14700 17554 14756 17556
rect 14700 17502 14702 17554
rect 14702 17502 14754 17554
rect 14754 17502 14756 17554
rect 14700 17500 14756 17502
rect 14820 17274 14876 17276
rect 14820 17222 14822 17274
rect 14822 17222 14874 17274
rect 14874 17222 14876 17274
rect 14820 17220 14876 17222
rect 14924 17274 14980 17276
rect 14924 17222 14926 17274
rect 14926 17222 14978 17274
rect 14978 17222 14980 17274
rect 14924 17220 14980 17222
rect 15028 17274 15084 17276
rect 15028 17222 15030 17274
rect 15030 17222 15082 17274
rect 15082 17222 15084 17274
rect 15028 17220 15084 17222
rect 15708 17612 15764 17668
rect 15372 17164 15428 17220
rect 15484 17500 15540 17556
rect 15932 17836 15988 17892
rect 16828 18284 16884 18340
rect 17612 23884 17668 23940
rect 17388 23772 17444 23828
rect 17052 23714 17108 23716
rect 17052 23662 17054 23714
rect 17054 23662 17106 23714
rect 17106 23662 17108 23714
rect 17052 23660 17108 23662
rect 17052 22370 17108 22372
rect 17052 22318 17054 22370
rect 17054 22318 17106 22370
rect 17106 22318 17108 22370
rect 17052 22316 17108 22318
rect 17052 20076 17108 20132
rect 16940 17948 16996 18004
rect 17612 22988 17668 23044
rect 17388 22764 17444 22820
rect 17500 22146 17556 22148
rect 17500 22094 17502 22146
rect 17502 22094 17554 22146
rect 17554 22094 17556 22146
rect 17500 22092 17556 22094
rect 19292 29986 19348 29988
rect 19292 29934 19294 29986
rect 19294 29934 19346 29986
rect 19346 29934 19348 29986
rect 19292 29932 19348 29934
rect 19292 29708 19348 29764
rect 19292 29314 19348 29316
rect 19292 29262 19294 29314
rect 19294 29262 19346 29314
rect 19346 29262 19348 29314
rect 19292 29260 19348 29262
rect 18844 28700 18900 28756
rect 19292 29036 19348 29092
rect 18844 27580 18900 27636
rect 18222 27466 18278 27468
rect 18222 27414 18224 27466
rect 18224 27414 18276 27466
rect 18276 27414 18278 27466
rect 18222 27412 18278 27414
rect 18326 27466 18382 27468
rect 18326 27414 18328 27466
rect 18328 27414 18380 27466
rect 18380 27414 18382 27466
rect 18326 27412 18382 27414
rect 18430 27466 18486 27468
rect 18430 27414 18432 27466
rect 18432 27414 18484 27466
rect 18484 27414 18486 27466
rect 18430 27412 18486 27414
rect 18172 27132 18228 27188
rect 18284 26962 18340 26964
rect 18284 26910 18286 26962
rect 18286 26910 18338 26962
rect 18338 26910 18340 26962
rect 18284 26908 18340 26910
rect 18172 26796 18228 26852
rect 17836 26066 17892 26068
rect 17836 26014 17838 26066
rect 17838 26014 17890 26066
rect 17890 26014 17892 26066
rect 17836 26012 17892 26014
rect 18620 27074 18676 27076
rect 18620 27022 18622 27074
rect 18622 27022 18674 27074
rect 18674 27022 18676 27074
rect 18620 27020 18676 27022
rect 18508 26066 18564 26068
rect 18508 26014 18510 26066
rect 18510 26014 18562 26066
rect 18562 26014 18564 26066
rect 18508 26012 18564 26014
rect 18222 25898 18278 25900
rect 18222 25846 18224 25898
rect 18224 25846 18276 25898
rect 18276 25846 18278 25898
rect 18222 25844 18278 25846
rect 18326 25898 18382 25900
rect 18326 25846 18328 25898
rect 18328 25846 18380 25898
rect 18380 25846 18382 25898
rect 18326 25844 18382 25846
rect 18430 25898 18486 25900
rect 18430 25846 18432 25898
rect 18432 25846 18484 25898
rect 18484 25846 18486 25898
rect 18430 25844 18486 25846
rect 18732 25900 18788 25956
rect 18844 25788 18900 25844
rect 18620 25340 18676 25396
rect 18396 24610 18452 24612
rect 18396 24558 18398 24610
rect 18398 24558 18450 24610
rect 18450 24558 18452 24610
rect 18396 24556 18452 24558
rect 17948 24444 18004 24500
rect 18222 24330 18278 24332
rect 18222 24278 18224 24330
rect 18224 24278 18276 24330
rect 18276 24278 18278 24330
rect 18222 24276 18278 24278
rect 18326 24330 18382 24332
rect 18326 24278 18328 24330
rect 18328 24278 18380 24330
rect 18380 24278 18382 24330
rect 18326 24276 18382 24278
rect 18430 24330 18486 24332
rect 18430 24278 18432 24330
rect 18432 24278 18484 24330
rect 18484 24278 18486 24330
rect 18430 24276 18486 24278
rect 18060 23772 18116 23828
rect 18508 24162 18564 24164
rect 18508 24110 18510 24162
rect 18510 24110 18562 24162
rect 18562 24110 18564 24162
rect 18508 24108 18564 24110
rect 17948 23042 18004 23044
rect 17948 22990 17950 23042
rect 17950 22990 18002 23042
rect 18002 22990 18004 23042
rect 17948 22988 18004 22990
rect 18732 24946 18788 24948
rect 18732 24894 18734 24946
rect 18734 24894 18786 24946
rect 18786 24894 18788 24946
rect 18732 24892 18788 24894
rect 19068 28588 19124 28644
rect 19068 27186 19124 27188
rect 19068 27134 19070 27186
rect 19070 27134 19122 27186
rect 19122 27134 19124 27186
rect 19068 27132 19124 27134
rect 19292 27746 19348 27748
rect 19292 27694 19294 27746
rect 19294 27694 19346 27746
rect 19346 27694 19348 27746
rect 19292 27692 19348 27694
rect 19292 27020 19348 27076
rect 19628 30716 19684 30772
rect 19852 30210 19908 30212
rect 19852 30158 19854 30210
rect 19854 30158 19906 30210
rect 19906 30158 19908 30210
rect 19852 30156 19908 30158
rect 19628 29708 19684 29764
rect 19852 29426 19908 29428
rect 19852 29374 19854 29426
rect 19854 29374 19906 29426
rect 19906 29374 19908 29426
rect 19852 29372 19908 29374
rect 19516 27020 19572 27076
rect 19628 27916 19684 27972
rect 19180 26684 19236 26740
rect 19180 26236 19236 26292
rect 20300 32562 20356 32564
rect 20300 32510 20302 32562
rect 20302 32510 20354 32562
rect 20354 32510 20356 32562
rect 20300 32508 20356 32510
rect 20860 37884 20916 37940
rect 21084 37660 21140 37716
rect 21980 38668 22036 38724
rect 21756 38050 21812 38052
rect 21756 37998 21758 38050
rect 21758 37998 21810 38050
rect 21810 37998 21812 38050
rect 21756 37996 21812 37998
rect 21420 37938 21476 37940
rect 21420 37886 21422 37938
rect 21422 37886 21474 37938
rect 21474 37886 21476 37938
rect 21420 37884 21476 37886
rect 21980 37772 22036 37828
rect 20636 35196 20692 35252
rect 20636 34802 20692 34804
rect 20636 34750 20638 34802
rect 20638 34750 20690 34802
rect 20690 34750 20692 34802
rect 20636 34748 20692 34750
rect 20748 34636 20804 34692
rect 20524 33740 20580 33796
rect 20860 35308 20916 35364
rect 20636 33628 20692 33684
rect 20748 34354 20804 34356
rect 20748 34302 20750 34354
rect 20750 34302 20802 34354
rect 20802 34302 20804 34354
rect 20748 34300 20804 34302
rect 20524 32060 20580 32116
rect 20412 31948 20468 32004
rect 20748 32956 20804 33012
rect 20636 31948 20692 32004
rect 20188 31388 20244 31444
rect 20188 30156 20244 30212
rect 20188 29986 20244 29988
rect 20188 29934 20190 29986
rect 20190 29934 20242 29986
rect 20242 29934 20244 29986
rect 20188 29932 20244 29934
rect 20636 31500 20692 31556
rect 20748 30210 20804 30212
rect 20748 30158 20750 30210
rect 20750 30158 20802 30210
rect 20802 30158 20804 30210
rect 20748 30156 20804 30158
rect 20300 29372 20356 29428
rect 20524 28418 20580 28420
rect 20524 28366 20526 28418
rect 20526 28366 20578 28418
rect 20578 28366 20580 28418
rect 20524 28364 20580 28366
rect 20076 27356 20132 27412
rect 20076 27020 20132 27076
rect 19740 26402 19796 26404
rect 19740 26350 19742 26402
rect 19742 26350 19794 26402
rect 19794 26350 19796 26402
rect 19740 26348 19796 26350
rect 19628 26236 19684 26292
rect 19180 26012 19236 26068
rect 18222 22762 18278 22764
rect 18222 22710 18224 22762
rect 18224 22710 18276 22762
rect 18276 22710 18278 22762
rect 18222 22708 18278 22710
rect 18326 22762 18382 22764
rect 18326 22710 18328 22762
rect 18328 22710 18380 22762
rect 18380 22710 18382 22762
rect 18326 22708 18382 22710
rect 18430 22762 18486 22764
rect 18430 22710 18432 22762
rect 18432 22710 18484 22762
rect 18484 22710 18486 22762
rect 18430 22708 18486 22710
rect 17836 22428 17892 22484
rect 17724 22092 17780 22148
rect 18620 22482 18676 22484
rect 18620 22430 18622 22482
rect 18622 22430 18674 22482
rect 18674 22430 18676 22482
rect 18620 22428 18676 22430
rect 18172 22146 18228 22148
rect 18172 22094 18174 22146
rect 18174 22094 18226 22146
rect 18226 22094 18228 22146
rect 18172 22092 18228 22094
rect 17612 21586 17668 21588
rect 17612 21534 17614 21586
rect 17614 21534 17666 21586
rect 17666 21534 17668 21586
rect 17612 21532 17668 21534
rect 17612 18396 17668 18452
rect 17500 18172 17556 18228
rect 16268 17554 16324 17556
rect 16268 17502 16270 17554
rect 16270 17502 16322 17554
rect 16322 17502 16324 17554
rect 16268 17500 16324 17502
rect 16940 17500 16996 17556
rect 15932 17276 15988 17332
rect 14588 16210 14644 16212
rect 14588 16158 14590 16210
rect 14590 16158 14642 16210
rect 14642 16158 14644 16210
rect 14588 16156 14644 16158
rect 15148 16156 15204 16212
rect 14820 15706 14876 15708
rect 14820 15654 14822 15706
rect 14822 15654 14874 15706
rect 14874 15654 14876 15706
rect 14820 15652 14876 15654
rect 14924 15706 14980 15708
rect 14924 15654 14926 15706
rect 14926 15654 14978 15706
rect 14978 15654 14980 15706
rect 14924 15652 14980 15654
rect 15028 15706 15084 15708
rect 15028 15654 15030 15706
rect 15030 15654 15082 15706
rect 15082 15654 15084 15706
rect 15028 15652 15084 15654
rect 15148 15372 15204 15428
rect 14812 15314 14868 15316
rect 14812 15262 14814 15314
rect 14814 15262 14866 15314
rect 14866 15262 14868 15314
rect 14812 15260 14868 15262
rect 14588 14588 14644 14644
rect 14252 13916 14308 13972
rect 13804 13692 13860 13748
rect 13804 13356 13860 13412
rect 13692 13132 13748 13188
rect 13580 12684 13636 12740
rect 12908 11282 12964 11284
rect 12908 11230 12910 11282
rect 12910 11230 12962 11282
rect 12962 11230 12964 11282
rect 12908 11228 12964 11230
rect 12796 10834 12852 10836
rect 12796 10782 12798 10834
rect 12798 10782 12850 10834
rect 12850 10782 12852 10834
rect 12796 10780 12852 10782
rect 13356 12348 13412 12404
rect 14140 13020 14196 13076
rect 14820 14138 14876 14140
rect 14820 14086 14822 14138
rect 14822 14086 14874 14138
rect 14874 14086 14876 14138
rect 14820 14084 14876 14086
rect 14924 14138 14980 14140
rect 14924 14086 14926 14138
rect 14926 14086 14978 14138
rect 14978 14086 14980 14138
rect 14924 14084 14980 14086
rect 15028 14138 15084 14140
rect 15028 14086 15030 14138
rect 15030 14086 15082 14138
rect 15082 14086 15084 14138
rect 15028 14084 15084 14086
rect 15036 13916 15092 13972
rect 14924 13804 14980 13860
rect 14812 13692 14868 13748
rect 14924 13074 14980 13076
rect 14924 13022 14926 13074
rect 14926 13022 14978 13074
rect 14978 13022 14980 13074
rect 14924 13020 14980 13022
rect 14820 12570 14876 12572
rect 14820 12518 14822 12570
rect 14822 12518 14874 12570
rect 14874 12518 14876 12570
rect 14820 12516 14876 12518
rect 14924 12570 14980 12572
rect 14924 12518 14926 12570
rect 14926 12518 14978 12570
rect 14978 12518 14980 12570
rect 14924 12516 14980 12518
rect 15028 12570 15084 12572
rect 15028 12518 15030 12570
rect 15030 12518 15082 12570
rect 15082 12518 15084 12570
rect 15028 12516 15084 12518
rect 13468 11116 13524 11172
rect 13580 11676 13636 11732
rect 14364 11676 14420 11732
rect 14700 12348 14756 12404
rect 14476 11394 14532 11396
rect 14476 11342 14478 11394
rect 14478 11342 14530 11394
rect 14530 11342 14532 11394
rect 14476 11340 14532 11342
rect 13916 11282 13972 11284
rect 13916 11230 13918 11282
rect 13918 11230 13970 11282
rect 13970 11230 13972 11282
rect 13916 11228 13972 11230
rect 13580 11004 13636 11060
rect 14588 11228 14644 11284
rect 15260 15314 15316 15316
rect 15260 15262 15262 15314
rect 15262 15262 15314 15314
rect 15314 15262 15316 15314
rect 15260 15260 15316 15262
rect 15260 13970 15316 13972
rect 15260 13918 15262 13970
rect 15262 13918 15314 13970
rect 15314 13918 15316 13970
rect 15260 13916 15316 13918
rect 15596 16716 15652 16772
rect 16716 17276 16772 17332
rect 16268 16994 16324 16996
rect 16268 16942 16270 16994
rect 16270 16942 16322 16994
rect 16322 16942 16324 16994
rect 16268 16940 16324 16942
rect 15708 14252 15764 14308
rect 15484 12124 15540 12180
rect 15148 11676 15204 11732
rect 13356 10498 13412 10500
rect 13356 10446 13358 10498
rect 13358 10446 13410 10498
rect 13410 10446 13412 10498
rect 13356 10444 13412 10446
rect 13580 10220 13636 10276
rect 12796 9772 12852 9828
rect 13132 9154 13188 9156
rect 13132 9102 13134 9154
rect 13134 9102 13186 9154
rect 13186 9102 13188 9154
rect 13132 9100 13188 9102
rect 13468 9212 13524 9268
rect 11418 8650 11474 8652
rect 11418 8598 11420 8650
rect 11420 8598 11472 8650
rect 11472 8598 11474 8650
rect 11418 8596 11474 8598
rect 11522 8650 11578 8652
rect 11522 8598 11524 8650
rect 11524 8598 11576 8650
rect 11576 8598 11578 8650
rect 11522 8596 11578 8598
rect 11626 8650 11682 8652
rect 11626 8598 11628 8650
rect 11628 8598 11680 8650
rect 11680 8598 11682 8650
rect 11626 8596 11682 8598
rect 13244 8316 13300 8372
rect 14028 10556 14084 10612
rect 13804 10332 13860 10388
rect 14820 11002 14876 11004
rect 14820 10950 14822 11002
rect 14822 10950 14874 11002
rect 14874 10950 14876 11002
rect 14820 10948 14876 10950
rect 14924 11002 14980 11004
rect 14924 10950 14926 11002
rect 14926 10950 14978 11002
rect 14978 10950 14980 11002
rect 14924 10948 14980 10950
rect 15028 11002 15084 11004
rect 15028 10950 15030 11002
rect 15030 10950 15082 11002
rect 15082 10950 15084 11002
rect 15028 10948 15084 10950
rect 14924 10834 14980 10836
rect 14924 10782 14926 10834
rect 14926 10782 14978 10834
rect 14978 10782 14980 10834
rect 14924 10780 14980 10782
rect 14476 10108 14532 10164
rect 14588 10220 14644 10276
rect 14140 9154 14196 9156
rect 14140 9102 14142 9154
rect 14142 9102 14194 9154
rect 14194 9102 14196 9154
rect 14140 9100 14196 9102
rect 14924 10220 14980 10276
rect 15372 10668 15428 10724
rect 14700 9996 14756 10052
rect 15148 9996 15204 10052
rect 15372 10220 15428 10276
rect 14820 9434 14876 9436
rect 14820 9382 14822 9434
rect 14822 9382 14874 9434
rect 14874 9382 14876 9434
rect 14820 9380 14876 9382
rect 14924 9434 14980 9436
rect 14924 9382 14926 9434
rect 14926 9382 14978 9434
rect 14978 9382 14980 9434
rect 14924 9380 14980 9382
rect 15028 9434 15084 9436
rect 15028 9382 15030 9434
rect 15030 9382 15082 9434
rect 15082 9382 15084 9434
rect 15028 9380 15084 9382
rect 14812 9212 14868 9268
rect 14700 9100 14756 9156
rect 14924 8988 14980 9044
rect 14252 8370 14308 8372
rect 14252 8318 14254 8370
rect 14254 8318 14306 8370
rect 14306 8318 14308 8370
rect 14252 8316 14308 8318
rect 9212 7644 9268 7700
rect 16828 16828 16884 16884
rect 16604 15372 16660 15428
rect 17276 17442 17332 17444
rect 17276 17390 17278 17442
rect 17278 17390 17330 17442
rect 17330 17390 17332 17442
rect 17276 17388 17332 17390
rect 17276 17052 17332 17108
rect 17612 16882 17668 16884
rect 17612 16830 17614 16882
rect 17614 16830 17666 16882
rect 17666 16830 17668 16882
rect 17612 16828 17668 16830
rect 16716 15036 16772 15092
rect 17052 16156 17108 16212
rect 16716 13916 16772 13972
rect 16716 12684 16772 12740
rect 16380 12402 16436 12404
rect 16380 12350 16382 12402
rect 16382 12350 16434 12402
rect 16434 12350 16436 12402
rect 16380 12348 16436 12350
rect 16268 12012 16324 12068
rect 16940 14924 16996 14980
rect 16828 12066 16884 12068
rect 16828 12014 16830 12066
rect 16830 12014 16882 12066
rect 16882 12014 16884 12066
rect 16828 12012 16884 12014
rect 15820 11564 15876 11620
rect 15820 11282 15876 11284
rect 15820 11230 15822 11282
rect 15822 11230 15874 11282
rect 15874 11230 15876 11282
rect 15820 11228 15876 11230
rect 15708 11116 15764 11172
rect 15708 10444 15764 10500
rect 15596 9884 15652 9940
rect 16268 10610 16324 10612
rect 16268 10558 16270 10610
rect 16270 10558 16322 10610
rect 16322 10558 16324 10610
rect 16268 10556 16324 10558
rect 16492 10610 16548 10612
rect 16492 10558 16494 10610
rect 16494 10558 16546 10610
rect 16546 10558 16548 10610
rect 16492 10556 16548 10558
rect 16492 10332 16548 10388
rect 15484 9212 15540 9268
rect 16156 8930 16212 8932
rect 16156 8878 16158 8930
rect 16158 8878 16210 8930
rect 16210 8878 16212 8930
rect 16156 8876 16212 8878
rect 15036 8316 15092 8372
rect 17836 20860 17892 20916
rect 17948 21532 18004 21588
rect 18060 21420 18116 21476
rect 18396 21308 18452 21364
rect 18222 21194 18278 21196
rect 18222 21142 18224 21194
rect 18224 21142 18276 21194
rect 18276 21142 18278 21194
rect 18222 21140 18278 21142
rect 18326 21194 18382 21196
rect 18326 21142 18328 21194
rect 18328 21142 18380 21194
rect 18380 21142 18382 21194
rect 18326 21140 18382 21142
rect 18430 21194 18486 21196
rect 18430 21142 18432 21194
rect 18432 21142 18484 21194
rect 18484 21142 18486 21194
rect 18430 21140 18486 21142
rect 18060 20636 18116 20692
rect 18844 24108 18900 24164
rect 18956 24220 19012 24276
rect 18844 23714 18900 23716
rect 18844 23662 18846 23714
rect 18846 23662 18898 23714
rect 18898 23662 18900 23714
rect 18844 23660 18900 23662
rect 18222 19626 18278 19628
rect 18222 19574 18224 19626
rect 18224 19574 18276 19626
rect 18276 19574 18278 19626
rect 18222 19572 18278 19574
rect 18326 19626 18382 19628
rect 18326 19574 18328 19626
rect 18328 19574 18380 19626
rect 18380 19574 18382 19626
rect 18326 19572 18382 19574
rect 18430 19626 18486 19628
rect 18430 19574 18432 19626
rect 18432 19574 18484 19626
rect 18484 19574 18486 19626
rect 18430 19572 18486 19574
rect 18284 19404 18340 19460
rect 18620 18956 18676 19012
rect 17948 18396 18004 18452
rect 18222 18058 18278 18060
rect 18222 18006 18224 18058
rect 18224 18006 18276 18058
rect 18276 18006 18278 18058
rect 18222 18004 18278 18006
rect 18326 18058 18382 18060
rect 18326 18006 18328 18058
rect 18328 18006 18380 18058
rect 18380 18006 18382 18058
rect 18326 18004 18382 18006
rect 18430 18058 18486 18060
rect 18430 18006 18432 18058
rect 18432 18006 18484 18058
rect 18484 18006 18486 18058
rect 18430 18004 18486 18006
rect 19068 23042 19124 23044
rect 19068 22990 19070 23042
rect 19070 22990 19122 23042
rect 19122 22990 19124 23042
rect 19068 22988 19124 22990
rect 19292 25788 19348 25844
rect 19292 25506 19348 25508
rect 19292 25454 19294 25506
rect 19294 25454 19346 25506
rect 19346 25454 19348 25506
rect 19292 25452 19348 25454
rect 19740 25282 19796 25284
rect 19740 25230 19742 25282
rect 19742 25230 19794 25282
rect 19794 25230 19796 25282
rect 19740 25228 19796 25230
rect 20412 27074 20468 27076
rect 20412 27022 20414 27074
rect 20414 27022 20466 27074
rect 20466 27022 20468 27074
rect 20412 27020 20468 27022
rect 19964 26348 20020 26404
rect 19628 24834 19684 24836
rect 19628 24782 19630 24834
rect 19630 24782 19682 24834
rect 19682 24782 19684 24834
rect 19628 24780 19684 24782
rect 19852 24556 19908 24612
rect 19292 23714 19348 23716
rect 19292 23662 19294 23714
rect 19294 23662 19346 23714
rect 19346 23662 19348 23714
rect 19292 23660 19348 23662
rect 19292 22652 19348 22708
rect 19068 22370 19124 22372
rect 19068 22318 19070 22370
rect 19070 22318 19122 22370
rect 19122 22318 19124 22370
rect 19068 22316 19124 22318
rect 19068 21756 19124 21812
rect 18956 21586 19012 21588
rect 18956 21534 18958 21586
rect 18958 21534 19010 21586
rect 19010 21534 19012 21586
rect 18956 21532 19012 21534
rect 19180 21308 19236 21364
rect 18956 20188 19012 20244
rect 18956 19010 19012 19012
rect 18956 18958 18958 19010
rect 18958 18958 19010 19010
rect 19010 18958 19012 19010
rect 18956 18956 19012 18958
rect 18620 17554 18676 17556
rect 18620 17502 18622 17554
rect 18622 17502 18674 17554
rect 18674 17502 18676 17554
rect 18620 17500 18676 17502
rect 18956 17500 19012 17556
rect 18060 17106 18116 17108
rect 18060 17054 18062 17106
rect 18062 17054 18114 17106
rect 18114 17054 18116 17106
rect 18060 17052 18116 17054
rect 18620 16940 18676 16996
rect 18222 16490 18278 16492
rect 18222 16438 18224 16490
rect 18224 16438 18276 16490
rect 18276 16438 18278 16490
rect 18222 16436 18278 16438
rect 18326 16490 18382 16492
rect 18326 16438 18328 16490
rect 18328 16438 18380 16490
rect 18380 16438 18382 16490
rect 18326 16436 18382 16438
rect 18430 16490 18486 16492
rect 18430 16438 18432 16490
rect 18432 16438 18484 16490
rect 18484 16438 18486 16490
rect 18430 16436 18486 16438
rect 18396 16210 18452 16212
rect 18396 16158 18398 16210
rect 18398 16158 18450 16210
rect 18450 16158 18452 16210
rect 18396 16156 18452 16158
rect 18844 17276 18900 17332
rect 19068 17276 19124 17332
rect 19516 23042 19572 23044
rect 19516 22990 19518 23042
rect 19518 22990 19570 23042
rect 19570 22990 19572 23042
rect 19516 22988 19572 22990
rect 19852 24332 19908 24388
rect 19740 22988 19796 23044
rect 19852 23324 19908 23380
rect 19852 22370 19908 22372
rect 19852 22318 19854 22370
rect 19854 22318 19906 22370
rect 19906 22318 19908 22370
rect 19852 22316 19908 22318
rect 19628 21756 19684 21812
rect 19516 21026 19572 21028
rect 19516 20974 19518 21026
rect 19518 20974 19570 21026
rect 19570 20974 19572 21026
rect 19516 20972 19572 20974
rect 19516 20802 19572 20804
rect 19516 20750 19518 20802
rect 19518 20750 19570 20802
rect 19570 20750 19572 20802
rect 19516 20748 19572 20750
rect 20300 25788 20356 25844
rect 20412 26796 20468 26852
rect 20188 24946 20244 24948
rect 20188 24894 20190 24946
rect 20190 24894 20242 24946
rect 20242 24894 20244 24946
rect 20188 24892 20244 24894
rect 20076 24444 20132 24500
rect 20188 24050 20244 24052
rect 20188 23998 20190 24050
rect 20190 23998 20242 24050
rect 20242 23998 20244 24050
rect 20188 23996 20244 23998
rect 20076 23660 20132 23716
rect 20748 29820 20804 29876
rect 20748 27468 20804 27524
rect 20748 27020 20804 27076
rect 20636 26236 20692 26292
rect 20748 25900 20804 25956
rect 20748 25340 20804 25396
rect 20972 32450 21028 32452
rect 20972 32398 20974 32450
rect 20974 32398 21026 32450
rect 21026 32398 21028 32450
rect 20972 32396 21028 32398
rect 21624 37658 21680 37660
rect 21624 37606 21626 37658
rect 21626 37606 21678 37658
rect 21678 37606 21680 37658
rect 21624 37604 21680 37606
rect 21728 37658 21784 37660
rect 21728 37606 21730 37658
rect 21730 37606 21782 37658
rect 21782 37606 21784 37658
rect 21728 37604 21784 37606
rect 21832 37658 21888 37660
rect 21832 37606 21834 37658
rect 21834 37606 21886 37658
rect 21886 37606 21888 37658
rect 21832 37604 21888 37606
rect 22092 37436 22148 37492
rect 22204 37996 22260 38052
rect 21756 37154 21812 37156
rect 21756 37102 21758 37154
rect 21758 37102 21810 37154
rect 21810 37102 21812 37154
rect 21756 37100 21812 37102
rect 23548 45388 23604 45444
rect 23996 52108 24052 52164
rect 23884 51436 23940 51492
rect 24220 51660 24276 51716
rect 24220 51436 24276 51492
rect 24108 51378 24164 51380
rect 24108 51326 24110 51378
rect 24110 51326 24162 51378
rect 24162 51326 24164 51378
rect 24108 51324 24164 51326
rect 24444 51154 24500 51156
rect 24444 51102 24446 51154
rect 24446 51102 24498 51154
rect 24498 51102 24500 51154
rect 24444 51100 24500 51102
rect 24332 50706 24388 50708
rect 24332 50654 24334 50706
rect 24334 50654 24386 50706
rect 24386 50654 24388 50706
rect 24332 50652 24388 50654
rect 24444 50540 24500 50596
rect 24332 50428 24388 50484
rect 24220 49980 24276 50036
rect 24108 49532 24164 49588
rect 23884 49250 23940 49252
rect 23884 49198 23886 49250
rect 23886 49198 23938 49250
rect 23938 49198 23940 49250
rect 23884 49196 23940 49198
rect 23996 48972 24052 49028
rect 23996 46844 24052 46900
rect 23884 45388 23940 45444
rect 23996 45330 24052 45332
rect 23996 45278 23998 45330
rect 23998 45278 24050 45330
rect 24050 45278 24052 45330
rect 23996 45276 24052 45278
rect 23436 43820 23492 43876
rect 23772 44322 23828 44324
rect 23772 44270 23774 44322
rect 23774 44270 23826 44322
rect 23826 44270 23828 44322
rect 23772 44268 23828 44270
rect 24332 48972 24388 49028
rect 24220 48860 24276 48916
rect 24892 52892 24948 52948
rect 24780 52556 24836 52612
rect 25228 52946 25284 52948
rect 25228 52894 25230 52946
rect 25230 52894 25282 52946
rect 25282 52894 25284 52946
rect 25228 52892 25284 52894
rect 25026 52554 25082 52556
rect 25026 52502 25028 52554
rect 25028 52502 25080 52554
rect 25080 52502 25082 52554
rect 25026 52500 25082 52502
rect 25130 52554 25186 52556
rect 25130 52502 25132 52554
rect 25132 52502 25184 52554
rect 25184 52502 25186 52554
rect 25130 52500 25186 52502
rect 25234 52554 25290 52556
rect 25234 52502 25236 52554
rect 25236 52502 25288 52554
rect 25288 52502 25290 52554
rect 25234 52500 25290 52502
rect 25228 52162 25284 52164
rect 25228 52110 25230 52162
rect 25230 52110 25282 52162
rect 25282 52110 25284 52162
rect 25228 52108 25284 52110
rect 25340 51100 25396 51156
rect 25026 50986 25082 50988
rect 25026 50934 25028 50986
rect 25028 50934 25080 50986
rect 25080 50934 25082 50986
rect 25026 50932 25082 50934
rect 25130 50986 25186 50988
rect 25130 50934 25132 50986
rect 25132 50934 25184 50986
rect 25184 50934 25186 50986
rect 25130 50932 25186 50934
rect 25234 50986 25290 50988
rect 25234 50934 25236 50986
rect 25236 50934 25288 50986
rect 25288 50934 25290 50986
rect 25234 50932 25290 50934
rect 25676 52108 25732 52164
rect 25788 53116 25844 53172
rect 25788 51490 25844 51492
rect 25788 51438 25790 51490
rect 25790 51438 25842 51490
rect 25842 51438 25844 51490
rect 25788 51436 25844 51438
rect 24668 49026 24724 49028
rect 24668 48974 24670 49026
rect 24670 48974 24722 49026
rect 24722 48974 24724 49026
rect 24668 48972 24724 48974
rect 24332 48802 24388 48804
rect 24332 48750 24334 48802
rect 24334 48750 24386 48802
rect 24386 48750 24388 48802
rect 24332 48748 24388 48750
rect 24332 46844 24388 46900
rect 24220 46620 24276 46676
rect 24332 45612 24388 45668
rect 24444 46732 24500 46788
rect 24556 46674 24612 46676
rect 24556 46622 24558 46674
rect 24558 46622 24610 46674
rect 24610 46622 24612 46674
rect 24556 46620 24612 46622
rect 24668 45666 24724 45668
rect 24668 45614 24670 45666
rect 24670 45614 24722 45666
rect 24722 45614 24724 45666
rect 24668 45612 24724 45614
rect 24444 44994 24500 44996
rect 24444 44942 24446 44994
rect 24446 44942 24498 44994
rect 24498 44942 24500 44994
rect 24444 44940 24500 44942
rect 23660 42476 23716 42532
rect 23436 42140 23492 42196
rect 22876 41244 22932 41300
rect 22876 40460 22932 40516
rect 23212 41132 23268 41188
rect 23548 41132 23604 41188
rect 23548 40962 23604 40964
rect 23548 40910 23550 40962
rect 23550 40910 23602 40962
rect 23602 40910 23604 40962
rect 23548 40908 23604 40910
rect 23324 40626 23380 40628
rect 23324 40574 23326 40626
rect 23326 40574 23378 40626
rect 23378 40574 23380 40626
rect 23324 40572 23380 40574
rect 23660 40460 23716 40516
rect 23212 40124 23268 40180
rect 22764 38780 22820 38836
rect 22988 39788 23044 39844
rect 22652 38556 22708 38612
rect 21980 37154 22036 37156
rect 21980 37102 21982 37154
rect 21982 37102 22034 37154
rect 22034 37102 22036 37154
rect 21980 37100 22036 37102
rect 22764 38050 22820 38052
rect 22764 37998 22766 38050
rect 22766 37998 22818 38050
rect 22818 37998 22820 38050
rect 22764 37996 22820 37998
rect 23212 39004 23268 39060
rect 22652 37100 22708 37156
rect 22764 37324 22820 37380
rect 21532 36428 21588 36484
rect 21644 36204 21700 36260
rect 21308 35868 21364 35924
rect 21420 36092 21476 36148
rect 21624 36090 21680 36092
rect 21624 36038 21626 36090
rect 21626 36038 21678 36090
rect 21678 36038 21680 36090
rect 21624 36036 21680 36038
rect 21728 36090 21784 36092
rect 21728 36038 21730 36090
rect 21730 36038 21782 36090
rect 21782 36038 21784 36090
rect 21728 36036 21784 36038
rect 21832 36090 21888 36092
rect 21832 36038 21834 36090
rect 21834 36038 21886 36090
rect 21886 36038 21888 36090
rect 21832 36036 21888 36038
rect 22988 37490 23044 37492
rect 22988 37438 22990 37490
rect 22990 37438 23042 37490
rect 23042 37438 23044 37490
rect 22988 37436 23044 37438
rect 22876 37212 22932 37268
rect 23548 40236 23604 40292
rect 23660 38834 23716 38836
rect 23660 38782 23662 38834
rect 23662 38782 23714 38834
rect 23714 38782 23716 38834
rect 23660 38780 23716 38782
rect 23884 42588 23940 42644
rect 23996 42140 24052 42196
rect 24108 42028 24164 42084
rect 24444 42476 24500 42532
rect 23884 41916 23940 41972
rect 23996 41580 24052 41636
rect 24668 42140 24724 42196
rect 24668 41970 24724 41972
rect 24668 41918 24670 41970
rect 24670 41918 24722 41970
rect 24722 41918 24724 41970
rect 24668 41916 24724 41918
rect 24556 41804 24612 41860
rect 24220 40908 24276 40964
rect 24108 40514 24164 40516
rect 24108 40462 24110 40514
rect 24110 40462 24162 40514
rect 24162 40462 24164 40514
rect 24108 40460 24164 40462
rect 24108 39452 24164 39508
rect 24108 39004 24164 39060
rect 24444 39788 24500 39844
rect 24668 41580 24724 41636
rect 23996 38780 24052 38836
rect 23436 37996 23492 38052
rect 23660 38050 23716 38052
rect 23660 37998 23662 38050
rect 23662 37998 23714 38050
rect 23714 37998 23716 38050
rect 23660 37996 23716 37998
rect 23212 37436 23268 37492
rect 23436 37660 23492 37716
rect 22092 35196 22148 35252
rect 21868 34748 21924 34804
rect 21624 34522 21680 34524
rect 21624 34470 21626 34522
rect 21626 34470 21678 34522
rect 21678 34470 21680 34522
rect 21624 34468 21680 34470
rect 21728 34522 21784 34524
rect 21728 34470 21730 34522
rect 21730 34470 21782 34522
rect 21782 34470 21784 34522
rect 21728 34468 21784 34470
rect 21832 34522 21888 34524
rect 21832 34470 21834 34522
rect 21834 34470 21886 34522
rect 21886 34470 21888 34522
rect 21832 34468 21888 34470
rect 22092 34690 22148 34692
rect 22092 34638 22094 34690
rect 22094 34638 22146 34690
rect 22146 34638 22148 34690
rect 22092 34636 22148 34638
rect 22204 34524 22260 34580
rect 22316 35868 22372 35924
rect 21980 34412 22036 34468
rect 21196 34354 21252 34356
rect 21196 34302 21198 34354
rect 21198 34302 21250 34354
rect 21250 34302 21252 34354
rect 21196 34300 21252 34302
rect 21756 34354 21812 34356
rect 21756 34302 21758 34354
rect 21758 34302 21810 34354
rect 21810 34302 21812 34354
rect 21756 34300 21812 34302
rect 21980 34188 22036 34244
rect 21308 33346 21364 33348
rect 21308 33294 21310 33346
rect 21310 33294 21362 33346
rect 21362 33294 21364 33346
rect 21308 33292 21364 33294
rect 21420 33122 21476 33124
rect 21420 33070 21422 33122
rect 21422 33070 21474 33122
rect 21474 33070 21476 33122
rect 21420 33068 21476 33070
rect 21624 32954 21680 32956
rect 21624 32902 21626 32954
rect 21626 32902 21678 32954
rect 21678 32902 21680 32954
rect 21624 32900 21680 32902
rect 21728 32954 21784 32956
rect 21728 32902 21730 32954
rect 21730 32902 21782 32954
rect 21782 32902 21784 32954
rect 21728 32900 21784 32902
rect 21832 32954 21888 32956
rect 21832 32902 21834 32954
rect 21834 32902 21886 32954
rect 21886 32902 21888 32954
rect 21832 32900 21888 32902
rect 23212 36764 23268 36820
rect 22764 35196 22820 35252
rect 22764 34860 22820 34916
rect 22540 34300 22596 34356
rect 22988 36428 23044 36484
rect 21420 32450 21476 32452
rect 21420 32398 21422 32450
rect 21422 32398 21474 32450
rect 21474 32398 21476 32450
rect 21420 32396 21476 32398
rect 21084 31836 21140 31892
rect 21308 31778 21364 31780
rect 21308 31726 21310 31778
rect 21310 31726 21362 31778
rect 21362 31726 21364 31778
rect 21308 31724 21364 31726
rect 21196 31052 21252 31108
rect 21084 30940 21140 30996
rect 21532 31500 21588 31556
rect 21624 31386 21680 31388
rect 21624 31334 21626 31386
rect 21626 31334 21678 31386
rect 21678 31334 21680 31386
rect 21624 31332 21680 31334
rect 21728 31386 21784 31388
rect 21728 31334 21730 31386
rect 21730 31334 21782 31386
rect 21782 31334 21784 31386
rect 21728 31332 21784 31334
rect 21832 31386 21888 31388
rect 21832 31334 21834 31386
rect 21834 31334 21886 31386
rect 21886 31334 21888 31386
rect 21832 31332 21888 31334
rect 21644 31218 21700 31220
rect 21644 31166 21646 31218
rect 21646 31166 21698 31218
rect 21698 31166 21700 31218
rect 21644 31164 21700 31166
rect 21980 30994 22036 30996
rect 21980 30942 21982 30994
rect 21982 30942 22034 30994
rect 22034 30942 22036 30994
rect 21980 30940 22036 30942
rect 21420 30380 21476 30436
rect 21868 29986 21924 29988
rect 21868 29934 21870 29986
rect 21870 29934 21922 29986
rect 21922 29934 21924 29986
rect 21868 29932 21924 29934
rect 21420 29820 21476 29876
rect 21624 29818 21680 29820
rect 21624 29766 21626 29818
rect 21626 29766 21678 29818
rect 21678 29766 21680 29818
rect 21624 29764 21680 29766
rect 21728 29818 21784 29820
rect 21728 29766 21730 29818
rect 21730 29766 21782 29818
rect 21782 29766 21784 29818
rect 21728 29764 21784 29766
rect 21832 29818 21888 29820
rect 21832 29766 21834 29818
rect 21834 29766 21886 29818
rect 21886 29766 21888 29818
rect 21832 29764 21888 29766
rect 21308 29372 21364 29428
rect 21868 29596 21924 29652
rect 21980 28364 22036 28420
rect 21624 28250 21680 28252
rect 21624 28198 21626 28250
rect 21626 28198 21678 28250
rect 21678 28198 21680 28250
rect 21624 28196 21680 28198
rect 21728 28250 21784 28252
rect 21728 28198 21730 28250
rect 21730 28198 21782 28250
rect 21782 28198 21784 28250
rect 21728 28196 21784 28198
rect 21832 28250 21888 28252
rect 21832 28198 21834 28250
rect 21834 28198 21886 28250
rect 21886 28198 21888 28250
rect 21832 28196 21888 28198
rect 21308 27356 21364 27412
rect 20972 27244 21028 27300
rect 21308 27020 21364 27076
rect 21308 26514 21364 26516
rect 21308 26462 21310 26514
rect 21310 26462 21362 26514
rect 21362 26462 21364 26514
rect 21308 26460 21364 26462
rect 21624 26682 21680 26684
rect 21624 26630 21626 26682
rect 21626 26630 21678 26682
rect 21678 26630 21680 26682
rect 21624 26628 21680 26630
rect 21728 26682 21784 26684
rect 21728 26630 21730 26682
rect 21730 26630 21782 26682
rect 21782 26630 21784 26682
rect 21728 26628 21784 26630
rect 21832 26682 21888 26684
rect 21832 26630 21834 26682
rect 21834 26630 21886 26682
rect 21886 26630 21888 26682
rect 21832 26628 21888 26630
rect 21644 26236 21700 26292
rect 20972 25900 21028 25956
rect 20412 23884 20468 23940
rect 20972 25564 21028 25620
rect 21980 26012 22036 26068
rect 21420 25340 21476 25396
rect 21084 25116 21140 25172
rect 20636 24050 20692 24052
rect 20636 23998 20638 24050
rect 20638 23998 20690 24050
rect 20690 23998 20692 24050
rect 20636 23996 20692 23998
rect 20300 23324 20356 23380
rect 20636 23100 20692 23156
rect 20860 23996 20916 24052
rect 20972 24668 21028 24724
rect 20412 22930 20468 22932
rect 20412 22878 20414 22930
rect 20414 22878 20466 22930
rect 20466 22878 20468 22930
rect 20412 22876 20468 22878
rect 20300 22428 20356 22484
rect 20076 21026 20132 21028
rect 20076 20974 20078 21026
rect 20078 20974 20130 21026
rect 20130 20974 20132 21026
rect 20076 20972 20132 20974
rect 19516 19404 19572 19460
rect 19404 18956 19460 19012
rect 19180 16994 19236 16996
rect 19180 16942 19182 16994
rect 19182 16942 19234 16994
rect 19234 16942 19236 16994
rect 19180 16940 19236 16942
rect 19740 18396 19796 18452
rect 19740 17276 19796 17332
rect 18732 16156 18788 16212
rect 18060 16044 18116 16100
rect 18956 15538 19012 15540
rect 18956 15486 18958 15538
rect 18958 15486 19010 15538
rect 19010 15486 19012 15538
rect 18956 15484 19012 15486
rect 18732 15314 18788 15316
rect 18732 15262 18734 15314
rect 18734 15262 18786 15314
rect 18786 15262 18788 15314
rect 18732 15260 18788 15262
rect 18222 14922 18278 14924
rect 18222 14870 18224 14922
rect 18224 14870 18276 14922
rect 18276 14870 18278 14922
rect 18222 14868 18278 14870
rect 18326 14922 18382 14924
rect 18326 14870 18328 14922
rect 18328 14870 18380 14922
rect 18380 14870 18382 14922
rect 18326 14868 18382 14870
rect 18430 14922 18486 14924
rect 18430 14870 18432 14922
rect 18432 14870 18484 14922
rect 18484 14870 18486 14922
rect 18430 14868 18486 14870
rect 17948 13804 18004 13860
rect 20972 21644 21028 21700
rect 20748 21420 20804 21476
rect 20412 20690 20468 20692
rect 20412 20638 20414 20690
rect 20414 20638 20466 20690
rect 20466 20638 20468 20690
rect 20412 20636 20468 20638
rect 20076 19852 20132 19908
rect 20300 19404 20356 19460
rect 20076 18956 20132 19012
rect 20524 19346 20580 19348
rect 20524 19294 20526 19346
rect 20526 19294 20578 19346
rect 20578 19294 20580 19346
rect 20524 19292 20580 19294
rect 20636 18956 20692 19012
rect 19292 15820 19348 15876
rect 20300 16940 20356 16996
rect 20748 18396 20804 18452
rect 20524 17052 20580 17108
rect 20188 16828 20244 16884
rect 19964 15484 20020 15540
rect 19292 15372 19348 15428
rect 19740 15426 19796 15428
rect 19740 15374 19742 15426
rect 19742 15374 19794 15426
rect 19794 15374 19796 15426
rect 19740 15372 19796 15374
rect 19180 14700 19236 14756
rect 20076 16156 20132 16212
rect 20300 16098 20356 16100
rect 20300 16046 20302 16098
rect 20302 16046 20354 16098
rect 20354 16046 20356 16098
rect 20300 16044 20356 16046
rect 20188 15314 20244 15316
rect 20188 15262 20190 15314
rect 20190 15262 20242 15314
rect 20242 15262 20244 15314
rect 20188 15260 20244 15262
rect 20972 17052 21028 17108
rect 20636 15538 20692 15540
rect 20636 15486 20638 15538
rect 20638 15486 20690 15538
rect 20690 15486 20692 15538
rect 20636 15484 20692 15486
rect 19068 14364 19124 14420
rect 19068 13858 19124 13860
rect 19068 13806 19070 13858
rect 19070 13806 19122 13858
rect 19122 13806 19124 13858
rect 19068 13804 19124 13806
rect 17052 13580 17108 13636
rect 17724 13634 17780 13636
rect 17724 13582 17726 13634
rect 17726 13582 17778 13634
rect 17778 13582 17780 13634
rect 17724 13580 17780 13582
rect 18396 13580 18452 13636
rect 18222 13354 18278 13356
rect 18222 13302 18224 13354
rect 18224 13302 18276 13354
rect 18276 13302 18278 13354
rect 18222 13300 18278 13302
rect 18326 13354 18382 13356
rect 18326 13302 18328 13354
rect 18328 13302 18380 13354
rect 18380 13302 18382 13354
rect 18326 13300 18382 13302
rect 18430 13354 18486 13356
rect 18430 13302 18432 13354
rect 18432 13302 18484 13354
rect 18484 13302 18486 13354
rect 18430 13300 18486 13302
rect 17948 12850 18004 12852
rect 17948 12798 17950 12850
rect 17950 12798 18002 12850
rect 18002 12798 18004 12850
rect 17948 12796 18004 12798
rect 17388 12684 17444 12740
rect 18172 12684 18228 12740
rect 17724 12402 17780 12404
rect 17724 12350 17726 12402
rect 17726 12350 17778 12402
rect 17778 12350 17780 12402
rect 17724 12348 17780 12350
rect 18396 12850 18452 12852
rect 18396 12798 18398 12850
rect 18398 12798 18450 12850
rect 18450 12798 18452 12850
rect 18396 12796 18452 12798
rect 18284 12572 18340 12628
rect 17724 12124 17780 12180
rect 17388 11788 17444 11844
rect 16940 11116 16996 11172
rect 16716 10668 16772 10724
rect 16716 10220 16772 10276
rect 16604 9996 16660 10052
rect 16828 9436 16884 9492
rect 16940 10556 16996 10612
rect 16828 9154 16884 9156
rect 16828 9102 16830 9154
rect 16830 9102 16882 9154
rect 16882 9102 16884 9154
rect 16828 9100 16884 9102
rect 16716 8876 16772 8932
rect 17052 9884 17108 9940
rect 8988 7532 9044 7588
rect 14820 7866 14876 7868
rect 14820 7814 14822 7866
rect 14822 7814 14874 7866
rect 14874 7814 14876 7866
rect 14820 7812 14876 7814
rect 14924 7866 14980 7868
rect 14924 7814 14926 7866
rect 14926 7814 14978 7866
rect 14978 7814 14980 7866
rect 14924 7812 14980 7814
rect 15028 7866 15084 7868
rect 15028 7814 15030 7866
rect 15030 7814 15082 7866
rect 15082 7814 15084 7866
rect 15028 7812 15084 7814
rect 16156 7308 16212 7364
rect 11418 7082 11474 7084
rect 11418 7030 11420 7082
rect 11420 7030 11472 7082
rect 11472 7030 11474 7082
rect 11418 7028 11474 7030
rect 11522 7082 11578 7084
rect 11522 7030 11524 7082
rect 11524 7030 11576 7082
rect 11576 7030 11578 7082
rect 11522 7028 11578 7030
rect 11626 7082 11682 7084
rect 11626 7030 11628 7082
rect 11628 7030 11680 7082
rect 11680 7030 11682 7082
rect 11626 7028 11682 7030
rect 17612 10556 17668 10612
rect 17388 10444 17444 10500
rect 17388 9714 17444 9716
rect 17388 9662 17390 9714
rect 17390 9662 17442 9714
rect 17442 9662 17444 9714
rect 17388 9660 17444 9662
rect 17388 9436 17444 9492
rect 17612 9436 17668 9492
rect 17388 8204 17444 8260
rect 17276 7980 17332 8036
rect 18956 12402 19012 12404
rect 18956 12350 18958 12402
rect 18958 12350 19010 12402
rect 19010 12350 19012 12402
rect 18956 12348 19012 12350
rect 18508 12012 18564 12068
rect 18620 12236 18676 12292
rect 18620 11900 18676 11956
rect 18222 11786 18278 11788
rect 18222 11734 18224 11786
rect 18224 11734 18276 11786
rect 18276 11734 18278 11786
rect 18222 11732 18278 11734
rect 18326 11786 18382 11788
rect 18326 11734 18328 11786
rect 18328 11734 18380 11786
rect 18380 11734 18382 11786
rect 18326 11732 18382 11734
rect 18430 11786 18486 11788
rect 18430 11734 18432 11786
rect 18432 11734 18484 11786
rect 18484 11734 18486 11786
rect 18430 11732 18486 11734
rect 18620 11676 18676 11732
rect 17948 10834 18004 10836
rect 17948 10782 17950 10834
rect 17950 10782 18002 10834
rect 18002 10782 18004 10834
rect 17948 10780 18004 10782
rect 18508 10332 18564 10388
rect 18222 10218 18278 10220
rect 18222 10166 18224 10218
rect 18224 10166 18276 10218
rect 18276 10166 18278 10218
rect 18222 10164 18278 10166
rect 18326 10218 18382 10220
rect 18326 10166 18328 10218
rect 18328 10166 18380 10218
rect 18380 10166 18382 10218
rect 18326 10164 18382 10166
rect 18430 10218 18486 10220
rect 18430 10166 18432 10218
rect 18432 10166 18484 10218
rect 18484 10166 18486 10218
rect 18430 10164 18486 10166
rect 17836 9996 17892 10052
rect 18620 9938 18676 9940
rect 18620 9886 18622 9938
rect 18622 9886 18674 9938
rect 18674 9886 18676 9938
rect 18620 9884 18676 9886
rect 18060 9660 18116 9716
rect 20188 12908 20244 12964
rect 19292 12236 19348 12292
rect 19628 12684 19684 12740
rect 19292 12012 19348 12068
rect 20188 12572 20244 12628
rect 19740 11788 19796 11844
rect 20188 11788 20244 11844
rect 19068 10668 19124 10724
rect 19964 11452 20020 11508
rect 20748 14642 20804 14644
rect 20748 14590 20750 14642
rect 20750 14590 20802 14642
rect 20802 14590 20804 14642
rect 20748 14588 20804 14590
rect 20524 12908 20580 12964
rect 19516 10108 19572 10164
rect 19068 9436 19124 9492
rect 17948 9154 18004 9156
rect 17948 9102 17950 9154
rect 17950 9102 18002 9154
rect 18002 9102 18004 9154
rect 17948 9100 18004 9102
rect 18844 9100 18900 9156
rect 17836 8876 17892 8932
rect 18222 8650 18278 8652
rect 18222 8598 18224 8650
rect 18224 8598 18276 8650
rect 18276 8598 18278 8650
rect 18222 8596 18278 8598
rect 18326 8650 18382 8652
rect 18326 8598 18328 8650
rect 18328 8598 18380 8650
rect 18380 8598 18382 8650
rect 18326 8596 18382 8598
rect 18430 8650 18486 8652
rect 18430 8598 18432 8650
rect 18432 8598 18484 8650
rect 18484 8598 18486 8650
rect 18430 8596 18486 8598
rect 18172 8370 18228 8372
rect 18172 8318 18174 8370
rect 18174 8318 18226 8370
rect 18226 8318 18228 8370
rect 18172 8316 18228 8318
rect 18620 8204 18676 8260
rect 17724 7532 17780 7588
rect 18222 7082 18278 7084
rect 18222 7030 18224 7082
rect 18224 7030 18276 7082
rect 18276 7030 18278 7082
rect 18222 7028 18278 7030
rect 18326 7082 18382 7084
rect 18326 7030 18328 7082
rect 18328 7030 18380 7082
rect 18380 7030 18382 7082
rect 18326 7028 18382 7030
rect 18430 7082 18486 7084
rect 18430 7030 18432 7082
rect 18432 7030 18484 7082
rect 18484 7030 18486 7082
rect 18430 7028 18486 7030
rect 20076 11394 20132 11396
rect 20076 11342 20078 11394
rect 20078 11342 20130 11394
rect 20130 11342 20132 11394
rect 20076 11340 20132 11342
rect 20300 10834 20356 10836
rect 20300 10782 20302 10834
rect 20302 10782 20354 10834
rect 20354 10782 20356 10834
rect 20300 10780 20356 10782
rect 20188 10556 20244 10612
rect 20300 10444 20356 10500
rect 19852 9884 19908 9940
rect 19628 9436 19684 9492
rect 19292 8258 19348 8260
rect 19292 8206 19294 8258
rect 19294 8206 19346 8258
rect 19346 8206 19348 8258
rect 19292 8204 19348 8206
rect 19740 8146 19796 8148
rect 19740 8094 19742 8146
rect 19742 8094 19794 8146
rect 19794 8094 19796 8146
rect 19740 8092 19796 8094
rect 20300 7644 20356 7700
rect 19068 7362 19124 7364
rect 19068 7310 19070 7362
rect 19070 7310 19122 7362
rect 19122 7310 19124 7362
rect 19068 7308 19124 7310
rect 19516 6636 19572 6692
rect 7644 6300 7700 6356
rect 8016 6298 8072 6300
rect 8016 6246 8018 6298
rect 8018 6246 8070 6298
rect 8070 6246 8072 6298
rect 8016 6244 8072 6246
rect 8120 6298 8176 6300
rect 8120 6246 8122 6298
rect 8122 6246 8174 6298
rect 8174 6246 8176 6298
rect 8120 6244 8176 6246
rect 8224 6298 8280 6300
rect 8224 6246 8226 6298
rect 8226 6246 8278 6298
rect 8278 6246 8280 6298
rect 8224 6244 8280 6246
rect 14820 6298 14876 6300
rect 14820 6246 14822 6298
rect 14822 6246 14874 6298
rect 14874 6246 14876 6298
rect 14820 6244 14876 6246
rect 14924 6298 14980 6300
rect 14924 6246 14926 6298
rect 14926 6246 14978 6298
rect 14978 6246 14980 6298
rect 14924 6244 14980 6246
rect 15028 6298 15084 6300
rect 15028 6246 15030 6298
rect 15030 6246 15082 6298
rect 15082 6246 15084 6298
rect 15028 6244 15084 6246
rect 18732 6130 18788 6132
rect 18732 6078 18734 6130
rect 18734 6078 18786 6130
rect 18786 6078 18788 6130
rect 18732 6076 18788 6078
rect 19852 5740 19908 5796
rect 4614 5514 4670 5516
rect 4614 5462 4616 5514
rect 4616 5462 4668 5514
rect 4668 5462 4670 5514
rect 4614 5460 4670 5462
rect 4718 5514 4774 5516
rect 4718 5462 4720 5514
rect 4720 5462 4772 5514
rect 4772 5462 4774 5514
rect 4718 5460 4774 5462
rect 4822 5514 4878 5516
rect 4822 5462 4824 5514
rect 4824 5462 4876 5514
rect 4876 5462 4878 5514
rect 4822 5460 4878 5462
rect 11418 5514 11474 5516
rect 11418 5462 11420 5514
rect 11420 5462 11472 5514
rect 11472 5462 11474 5514
rect 11418 5460 11474 5462
rect 11522 5514 11578 5516
rect 11522 5462 11524 5514
rect 11524 5462 11576 5514
rect 11576 5462 11578 5514
rect 11522 5460 11578 5462
rect 11626 5514 11682 5516
rect 11626 5462 11628 5514
rect 11628 5462 11680 5514
rect 11680 5462 11682 5514
rect 11626 5460 11682 5462
rect 18222 5514 18278 5516
rect 18222 5462 18224 5514
rect 18224 5462 18276 5514
rect 18276 5462 18278 5514
rect 18222 5460 18278 5462
rect 18326 5514 18382 5516
rect 18326 5462 18328 5514
rect 18328 5462 18380 5514
rect 18380 5462 18382 5514
rect 18326 5460 18382 5462
rect 18430 5514 18486 5516
rect 18430 5462 18432 5514
rect 18432 5462 18484 5514
rect 18484 5462 18486 5514
rect 18430 5460 18486 5462
rect 18732 5122 18788 5124
rect 18732 5070 18734 5122
rect 18734 5070 18786 5122
rect 18786 5070 18788 5122
rect 18732 5068 18788 5070
rect 8016 4730 8072 4732
rect 8016 4678 8018 4730
rect 8018 4678 8070 4730
rect 8070 4678 8072 4730
rect 8016 4676 8072 4678
rect 8120 4730 8176 4732
rect 8120 4678 8122 4730
rect 8122 4678 8174 4730
rect 8174 4678 8176 4730
rect 8120 4676 8176 4678
rect 8224 4730 8280 4732
rect 8224 4678 8226 4730
rect 8226 4678 8278 4730
rect 8278 4678 8280 4730
rect 8224 4676 8280 4678
rect 14820 4730 14876 4732
rect 14820 4678 14822 4730
rect 14822 4678 14874 4730
rect 14874 4678 14876 4730
rect 14820 4676 14876 4678
rect 14924 4730 14980 4732
rect 14924 4678 14926 4730
rect 14926 4678 14978 4730
rect 14978 4678 14980 4730
rect 14924 4676 14980 4678
rect 15028 4730 15084 4732
rect 15028 4678 15030 4730
rect 15030 4678 15082 4730
rect 15082 4678 15084 4730
rect 15028 4676 15084 4678
rect 4614 3946 4670 3948
rect 4614 3894 4616 3946
rect 4616 3894 4668 3946
rect 4668 3894 4670 3946
rect 4614 3892 4670 3894
rect 4718 3946 4774 3948
rect 4718 3894 4720 3946
rect 4720 3894 4772 3946
rect 4772 3894 4774 3946
rect 4718 3892 4774 3894
rect 4822 3946 4878 3948
rect 4822 3894 4824 3946
rect 4824 3894 4876 3946
rect 4876 3894 4878 3946
rect 4822 3892 4878 3894
rect 4956 3388 5012 3444
rect 4284 2716 4340 2772
rect 3612 2156 3668 2212
rect 3948 1820 4004 1876
rect 4614 2378 4670 2380
rect 4614 2326 4616 2378
rect 4616 2326 4668 2378
rect 4668 2326 4670 2378
rect 4614 2324 4670 2326
rect 4718 2378 4774 2380
rect 4718 2326 4720 2378
rect 4720 2326 4772 2378
rect 4772 2326 4774 2378
rect 4718 2324 4774 2326
rect 4822 2378 4878 2380
rect 4822 2326 4824 2378
rect 4824 2326 4876 2378
rect 4876 2326 4878 2378
rect 4822 2324 4878 2326
rect 4732 1820 4788 1876
rect 5404 1820 5460 1876
rect 5740 3442 5796 3444
rect 5740 3390 5742 3442
rect 5742 3390 5794 3442
rect 5794 3390 5796 3442
rect 5740 3388 5796 3390
rect 6412 3388 6468 3444
rect 6188 2770 6244 2772
rect 6188 2718 6190 2770
rect 6190 2718 6242 2770
rect 6242 2718 6244 2770
rect 6188 2716 6244 2718
rect 6300 2156 6356 2212
rect 8764 3500 8820 3556
rect 8016 3162 8072 3164
rect 8016 3110 8018 3162
rect 8018 3110 8070 3162
rect 8070 3110 8072 3162
rect 8016 3108 8072 3110
rect 8120 3162 8176 3164
rect 8120 3110 8122 3162
rect 8122 3110 8174 3162
rect 8174 3110 8176 3162
rect 8120 3108 8176 3110
rect 8224 3162 8280 3164
rect 8224 3110 8226 3162
rect 8226 3110 8278 3162
rect 8278 3110 8280 3162
rect 8224 3108 8280 3110
rect 8092 2940 8148 2996
rect 8016 1594 8072 1596
rect 8016 1542 8018 1594
rect 8018 1542 8070 1594
rect 8070 1542 8072 1594
rect 8016 1540 8072 1542
rect 8120 1594 8176 1596
rect 8120 1542 8122 1594
rect 8122 1542 8174 1594
rect 8174 1542 8176 1594
rect 8120 1540 8176 1542
rect 8224 1594 8280 1596
rect 8224 1542 8226 1594
rect 8226 1542 8278 1594
rect 8278 1542 8280 1594
rect 8224 1540 8280 1542
rect 9660 3554 9716 3556
rect 9660 3502 9662 3554
rect 9662 3502 9714 3554
rect 9714 3502 9716 3554
rect 9660 3500 9716 3502
rect 11676 4226 11732 4228
rect 11676 4174 11678 4226
rect 11678 4174 11730 4226
rect 11730 4174 11732 4226
rect 11676 4172 11732 4174
rect 11564 4060 11620 4116
rect 11418 3946 11474 3948
rect 11418 3894 11420 3946
rect 11420 3894 11472 3946
rect 11472 3894 11474 3946
rect 11418 3892 11474 3894
rect 11522 3946 11578 3948
rect 11522 3894 11524 3946
rect 11524 3894 11576 3946
rect 11576 3894 11578 3946
rect 11522 3892 11578 3894
rect 11626 3946 11682 3948
rect 11626 3894 11628 3946
rect 11628 3894 11680 3946
rect 11680 3894 11682 3946
rect 11626 3892 11682 3894
rect 11004 3500 11060 3556
rect 11788 3554 11844 3556
rect 11788 3502 11790 3554
rect 11790 3502 11842 3554
rect 11842 3502 11844 3554
rect 11788 3500 11844 3502
rect 10220 3164 10276 3220
rect 12124 3948 12180 4004
rect 12124 3442 12180 3444
rect 12124 3390 12126 3442
rect 12126 3390 12178 3442
rect 12178 3390 12180 3442
rect 12124 3388 12180 3390
rect 13020 3724 13076 3780
rect 9996 2716 10052 2772
rect 10556 2770 10612 2772
rect 10556 2718 10558 2770
rect 10558 2718 10610 2770
rect 10610 2718 10612 2770
rect 10556 2716 10612 2718
rect 11676 2940 11732 2996
rect 12572 2994 12628 2996
rect 12572 2942 12574 2994
rect 12574 2942 12626 2994
rect 12626 2942 12628 2994
rect 12572 2940 12628 2942
rect 10780 2156 10836 2212
rect 11228 2380 11284 2436
rect 11418 2378 11474 2380
rect 11418 2326 11420 2378
rect 11420 2326 11472 2378
rect 11472 2326 11474 2378
rect 11418 2324 11474 2326
rect 11522 2378 11578 2380
rect 11522 2326 11524 2378
rect 11524 2326 11576 2378
rect 11576 2326 11578 2378
rect 11522 2324 11578 2326
rect 11626 2378 11682 2380
rect 11626 2326 11628 2378
rect 11628 2326 11680 2378
rect 11680 2326 11682 2378
rect 11626 2324 11682 2326
rect 10892 1762 10948 1764
rect 10892 1710 10894 1762
rect 10894 1710 10946 1762
rect 10946 1710 10948 1762
rect 10892 1708 10948 1710
rect 14820 3162 14876 3164
rect 14820 3110 14822 3162
rect 14822 3110 14874 3162
rect 14874 3110 14876 3162
rect 14820 3108 14876 3110
rect 14924 3162 14980 3164
rect 14924 3110 14926 3162
rect 14926 3110 14978 3162
rect 14978 3110 14980 3162
rect 14924 3108 14980 3110
rect 15028 3162 15084 3164
rect 15028 3110 15030 3162
rect 15030 3110 15082 3162
rect 15082 3110 15084 3162
rect 15028 3108 15084 3110
rect 13580 2604 13636 2660
rect 12348 2156 12404 2212
rect 12908 2546 12964 2548
rect 12908 2494 12910 2546
rect 12910 2494 12962 2546
rect 12962 2494 12964 2546
rect 12908 2492 12964 2494
rect 12796 2156 12852 2212
rect 13468 1986 13524 1988
rect 13468 1934 13470 1986
rect 13470 1934 13522 1986
rect 13522 1934 13524 1986
rect 13468 1932 13524 1934
rect 14140 2156 14196 2212
rect 14364 2492 14420 2548
rect 14140 1932 14196 1988
rect 14700 1986 14756 1988
rect 14700 1934 14702 1986
rect 14702 1934 14754 1986
rect 14754 1934 14756 1986
rect 14700 1932 14756 1934
rect 14820 1594 14876 1596
rect 14820 1542 14822 1594
rect 14822 1542 14874 1594
rect 14874 1542 14876 1594
rect 14820 1540 14876 1542
rect 14924 1594 14980 1596
rect 14924 1542 14926 1594
rect 14926 1542 14978 1594
rect 14978 1542 14980 1594
rect 14924 1540 14980 1542
rect 15028 1594 15084 1596
rect 15028 1542 15030 1594
rect 15030 1542 15082 1594
rect 15082 1542 15084 1594
rect 15028 1540 15084 1542
rect 16268 2658 16324 2660
rect 16268 2606 16270 2658
rect 16270 2606 16322 2658
rect 16322 2606 16324 2658
rect 16268 2604 16324 2606
rect 16156 1820 16212 1876
rect 17052 2604 17108 2660
rect 16940 1874 16996 1876
rect 16940 1822 16942 1874
rect 16942 1822 16994 1874
rect 16994 1822 16996 1874
rect 16940 1820 16996 1822
rect 17500 3164 17556 3220
rect 17724 3052 17780 3108
rect 17388 2770 17444 2772
rect 17388 2718 17390 2770
rect 17390 2718 17442 2770
rect 17442 2718 17444 2770
rect 17388 2716 17444 2718
rect 17612 2604 17668 2660
rect 17948 3052 18004 3108
rect 18284 4060 18340 4116
rect 18222 3946 18278 3948
rect 18222 3894 18224 3946
rect 18224 3894 18276 3946
rect 18276 3894 18278 3946
rect 18222 3892 18278 3894
rect 18326 3946 18382 3948
rect 18326 3894 18328 3946
rect 18328 3894 18380 3946
rect 18380 3894 18382 3946
rect 18326 3892 18382 3894
rect 18430 3946 18486 3948
rect 18430 3894 18432 3946
rect 18432 3894 18484 3946
rect 18484 3894 18486 3946
rect 18430 3892 18486 3894
rect 18396 2828 18452 2884
rect 18222 2378 18278 2380
rect 18222 2326 18224 2378
rect 18224 2326 18276 2378
rect 18276 2326 18278 2378
rect 18222 2324 18278 2326
rect 18326 2378 18382 2380
rect 18326 2326 18328 2378
rect 18328 2326 18380 2378
rect 18380 2326 18382 2378
rect 18326 2324 18382 2326
rect 18430 2378 18486 2380
rect 18430 2326 18432 2378
rect 18432 2326 18484 2378
rect 18484 2326 18486 2378
rect 18430 2324 18486 2326
rect 18172 2156 18228 2212
rect 18508 1874 18564 1876
rect 18508 1822 18510 1874
rect 18510 1822 18562 1874
rect 18562 1822 18564 1874
rect 18508 1820 18564 1822
rect 19852 4898 19908 4900
rect 19852 4846 19854 4898
rect 19854 4846 19906 4898
rect 19906 4846 19908 4898
rect 19852 4844 19908 4846
rect 19628 4732 19684 4788
rect 19292 4060 19348 4116
rect 19740 3612 19796 3668
rect 21196 24946 21252 24948
rect 21196 24894 21198 24946
rect 21198 24894 21250 24946
rect 21250 24894 21252 24946
rect 21196 24892 21252 24894
rect 21624 25114 21680 25116
rect 21624 25062 21626 25114
rect 21626 25062 21678 25114
rect 21678 25062 21680 25114
rect 21624 25060 21680 25062
rect 21728 25114 21784 25116
rect 21728 25062 21730 25114
rect 21730 25062 21782 25114
rect 21782 25062 21784 25114
rect 21728 25060 21784 25062
rect 21832 25114 21888 25116
rect 21832 25062 21834 25114
rect 21834 25062 21886 25114
rect 21886 25062 21888 25114
rect 21832 25060 21888 25062
rect 22428 33852 22484 33908
rect 22988 35532 23044 35588
rect 22316 33404 22372 33460
rect 22428 33346 22484 33348
rect 22428 33294 22430 33346
rect 22430 33294 22482 33346
rect 22482 33294 22484 33346
rect 22428 33292 22484 33294
rect 22316 33180 22372 33236
rect 22652 33180 22708 33236
rect 22540 33122 22596 33124
rect 22540 33070 22542 33122
rect 22542 33070 22594 33122
rect 22594 33070 22596 33122
rect 22540 33068 22596 33070
rect 22876 33068 22932 33124
rect 23660 35420 23716 35476
rect 23100 32844 23156 32900
rect 23212 35308 23268 35364
rect 22316 31948 22372 32004
rect 22540 29820 22596 29876
rect 22540 29596 22596 29652
rect 22316 29484 22372 29540
rect 22540 28364 22596 28420
rect 22204 25564 22260 25620
rect 22316 26178 22372 26180
rect 22316 26126 22318 26178
rect 22318 26126 22370 26178
rect 22370 26126 22372 26178
rect 22316 26124 22372 26126
rect 22316 25228 22372 25284
rect 21196 23660 21252 23716
rect 21196 22876 21252 22932
rect 21420 24332 21476 24388
rect 21624 23546 21680 23548
rect 21624 23494 21626 23546
rect 21626 23494 21678 23546
rect 21678 23494 21680 23546
rect 21624 23492 21680 23494
rect 21728 23546 21784 23548
rect 21728 23494 21730 23546
rect 21730 23494 21782 23546
rect 21782 23494 21784 23546
rect 21728 23492 21784 23494
rect 21832 23546 21888 23548
rect 21832 23494 21834 23546
rect 21834 23494 21886 23546
rect 21886 23494 21888 23546
rect 21832 23492 21888 23494
rect 21420 23324 21476 23380
rect 21980 23212 22036 23268
rect 21624 21978 21680 21980
rect 21624 21926 21626 21978
rect 21626 21926 21678 21978
rect 21678 21926 21680 21978
rect 21624 21924 21680 21926
rect 21728 21978 21784 21980
rect 21728 21926 21730 21978
rect 21730 21926 21782 21978
rect 21782 21926 21784 21978
rect 21728 21924 21784 21926
rect 21832 21978 21888 21980
rect 21832 21926 21834 21978
rect 21834 21926 21886 21978
rect 21886 21926 21888 21978
rect 21832 21924 21888 21926
rect 21420 21756 21476 21812
rect 21868 21474 21924 21476
rect 21868 21422 21870 21474
rect 21870 21422 21922 21474
rect 21922 21422 21924 21474
rect 21868 21420 21924 21422
rect 21420 20578 21476 20580
rect 21420 20526 21422 20578
rect 21422 20526 21474 20578
rect 21474 20526 21476 20578
rect 21420 20524 21476 20526
rect 21624 20410 21680 20412
rect 21624 20358 21626 20410
rect 21626 20358 21678 20410
rect 21678 20358 21680 20410
rect 21624 20356 21680 20358
rect 21728 20410 21784 20412
rect 21728 20358 21730 20410
rect 21730 20358 21782 20410
rect 21782 20358 21784 20410
rect 21728 20356 21784 20358
rect 21832 20410 21888 20412
rect 21832 20358 21834 20410
rect 21834 20358 21886 20410
rect 21886 20358 21888 20410
rect 21832 20356 21888 20358
rect 21308 19852 21364 19908
rect 21644 19404 21700 19460
rect 21532 19068 21588 19124
rect 21308 17500 21364 17556
rect 21196 17276 21252 17332
rect 21756 19122 21812 19124
rect 21756 19070 21758 19122
rect 21758 19070 21810 19122
rect 21810 19070 21812 19122
rect 21756 19068 21812 19070
rect 21624 18842 21680 18844
rect 21624 18790 21626 18842
rect 21626 18790 21678 18842
rect 21678 18790 21680 18842
rect 21624 18788 21680 18790
rect 21728 18842 21784 18844
rect 21728 18790 21730 18842
rect 21730 18790 21782 18842
rect 21782 18790 21784 18842
rect 21728 18788 21784 18790
rect 21832 18842 21888 18844
rect 21832 18790 21834 18842
rect 21834 18790 21886 18842
rect 21886 18790 21888 18842
rect 21832 18788 21888 18790
rect 21624 17274 21680 17276
rect 21624 17222 21626 17274
rect 21626 17222 21678 17274
rect 21678 17222 21680 17274
rect 21624 17220 21680 17222
rect 21728 17274 21784 17276
rect 21728 17222 21730 17274
rect 21730 17222 21782 17274
rect 21782 17222 21784 17274
rect 21728 17220 21784 17222
rect 21832 17274 21888 17276
rect 21832 17222 21834 17274
rect 21834 17222 21886 17274
rect 21886 17222 21888 17274
rect 21832 17220 21888 17222
rect 22204 23324 22260 23380
rect 22316 23548 22372 23604
rect 22988 32060 23044 32116
rect 22652 26796 22708 26852
rect 22876 31948 22932 32004
rect 22988 29820 23044 29876
rect 23548 35308 23604 35364
rect 23324 34412 23380 34468
rect 23436 34076 23492 34132
rect 23324 33628 23380 33684
rect 23772 35084 23828 35140
rect 23996 38108 24052 38164
rect 24332 37548 24388 37604
rect 24220 36428 24276 36484
rect 24332 37100 24388 37156
rect 24108 35420 24164 35476
rect 24220 35308 24276 35364
rect 24332 35420 24388 35476
rect 23996 35196 24052 35252
rect 23660 34018 23716 34020
rect 23660 33966 23662 34018
rect 23662 33966 23714 34018
rect 23714 33966 23716 34018
rect 23660 33964 23716 33966
rect 23996 34972 24052 35028
rect 23660 33628 23716 33684
rect 23324 33404 23380 33460
rect 23324 31836 23380 31892
rect 23436 32844 23492 32900
rect 23324 31666 23380 31668
rect 23324 31614 23326 31666
rect 23326 31614 23378 31666
rect 23378 31614 23380 31666
rect 23324 31612 23380 31614
rect 23660 33122 23716 33124
rect 23660 33070 23662 33122
rect 23662 33070 23714 33122
rect 23714 33070 23716 33122
rect 23660 33068 23716 33070
rect 23660 32396 23716 32452
rect 23212 29596 23268 29652
rect 22988 28588 23044 28644
rect 22988 28028 23044 28084
rect 23100 27244 23156 27300
rect 23660 30156 23716 30212
rect 23660 29932 23716 29988
rect 23548 28476 23604 28532
rect 23212 27020 23268 27076
rect 22876 26460 22932 26516
rect 23100 26684 23156 26740
rect 22652 26290 22708 26292
rect 22652 26238 22654 26290
rect 22654 26238 22706 26290
rect 22706 26238 22708 26290
rect 22652 26236 22708 26238
rect 22428 23324 22484 23380
rect 22092 22428 22148 22484
rect 22204 22930 22260 22932
rect 22204 22878 22206 22930
rect 22206 22878 22258 22930
rect 22258 22878 22260 22930
rect 22204 22876 22260 22878
rect 22316 22482 22372 22484
rect 22316 22430 22318 22482
rect 22318 22430 22370 22482
rect 22370 22430 22372 22482
rect 22316 22428 22372 22430
rect 22092 20188 22148 20244
rect 22204 20524 22260 20580
rect 22428 20524 22484 20580
rect 22316 20076 22372 20132
rect 23548 27858 23604 27860
rect 23548 27806 23550 27858
rect 23550 27806 23602 27858
rect 23602 27806 23604 27858
rect 23548 27804 23604 27806
rect 23212 26124 23268 26180
rect 24108 34748 24164 34804
rect 24220 34188 24276 34244
rect 23884 32620 23940 32676
rect 23884 32060 23940 32116
rect 24668 39116 24724 39172
rect 24668 38220 24724 38276
rect 25452 50540 25508 50596
rect 25026 49418 25082 49420
rect 25026 49366 25028 49418
rect 25028 49366 25080 49418
rect 25080 49366 25082 49418
rect 25026 49364 25082 49366
rect 25130 49418 25186 49420
rect 25130 49366 25132 49418
rect 25132 49366 25184 49418
rect 25184 49366 25186 49418
rect 25130 49364 25186 49366
rect 25234 49418 25290 49420
rect 25234 49366 25236 49418
rect 25236 49366 25288 49418
rect 25288 49366 25290 49418
rect 25234 49364 25290 49366
rect 25788 50540 25844 50596
rect 25564 49644 25620 49700
rect 25564 49420 25620 49476
rect 25452 49308 25508 49364
rect 25228 49250 25284 49252
rect 25228 49198 25230 49250
rect 25230 49198 25282 49250
rect 25282 49198 25284 49250
rect 25228 49196 25284 49198
rect 24892 48914 24948 48916
rect 24892 48862 24894 48914
rect 24894 48862 24946 48914
rect 24946 48862 24948 48914
rect 24892 48860 24948 48862
rect 24892 48636 24948 48692
rect 24556 37266 24612 37268
rect 24556 37214 24558 37266
rect 24558 37214 24610 37266
rect 24610 37214 24612 37266
rect 24556 37212 24612 37214
rect 24780 37826 24836 37828
rect 24780 37774 24782 37826
rect 24782 37774 24834 37826
rect 24834 37774 24836 37826
rect 24780 37772 24836 37774
rect 24444 33404 24500 33460
rect 24780 37548 24836 37604
rect 24444 33122 24500 33124
rect 24444 33070 24446 33122
rect 24446 33070 24498 33122
rect 24498 33070 24500 33122
rect 24444 33068 24500 33070
rect 24220 31890 24276 31892
rect 24220 31838 24222 31890
rect 24222 31838 24274 31890
rect 24274 31838 24276 31890
rect 24220 31836 24276 31838
rect 24108 31218 24164 31220
rect 24108 31166 24110 31218
rect 24110 31166 24162 31218
rect 24162 31166 24164 31218
rect 24108 31164 24164 31166
rect 24332 31106 24388 31108
rect 24332 31054 24334 31106
rect 24334 31054 24386 31106
rect 24386 31054 24388 31106
rect 24332 31052 24388 31054
rect 23996 30828 24052 30884
rect 23996 30044 24052 30100
rect 23884 29314 23940 29316
rect 23884 29262 23886 29314
rect 23886 29262 23938 29314
rect 23938 29262 23940 29314
rect 23884 29260 23940 29262
rect 23772 28140 23828 28196
rect 24668 35586 24724 35588
rect 24668 35534 24670 35586
rect 24670 35534 24722 35586
rect 24722 35534 24724 35586
rect 24668 35532 24724 35534
rect 24668 35196 24724 35252
rect 25228 49026 25284 49028
rect 25228 48974 25230 49026
rect 25230 48974 25282 49026
rect 25282 48974 25284 49026
rect 25228 48972 25284 48974
rect 25026 47850 25082 47852
rect 25026 47798 25028 47850
rect 25028 47798 25080 47850
rect 25080 47798 25082 47850
rect 25026 47796 25082 47798
rect 25130 47850 25186 47852
rect 25130 47798 25132 47850
rect 25132 47798 25184 47850
rect 25184 47798 25186 47850
rect 25130 47796 25186 47798
rect 25234 47850 25290 47852
rect 25234 47798 25236 47850
rect 25236 47798 25288 47850
rect 25288 47798 25290 47850
rect 25234 47796 25290 47798
rect 25564 47404 25620 47460
rect 25452 47180 25508 47236
rect 25340 46674 25396 46676
rect 25340 46622 25342 46674
rect 25342 46622 25394 46674
rect 25394 46622 25396 46674
rect 25340 46620 25396 46622
rect 25228 46508 25284 46564
rect 25026 46282 25082 46284
rect 25026 46230 25028 46282
rect 25028 46230 25080 46282
rect 25080 46230 25082 46282
rect 25026 46228 25082 46230
rect 25130 46282 25186 46284
rect 25130 46230 25132 46282
rect 25132 46230 25184 46282
rect 25184 46230 25186 46282
rect 25130 46228 25186 46230
rect 25234 46282 25290 46284
rect 25234 46230 25236 46282
rect 25236 46230 25288 46282
rect 25288 46230 25290 46282
rect 25234 46228 25290 46230
rect 25116 46002 25172 46004
rect 25116 45950 25118 46002
rect 25118 45950 25170 46002
rect 25170 45950 25172 46002
rect 25116 45948 25172 45950
rect 25676 47068 25732 47124
rect 26348 57036 26404 57092
rect 26012 55356 26068 55412
rect 26012 55020 26068 55076
rect 26012 54348 26068 54404
rect 26796 60060 26852 60116
rect 26908 59388 26964 59444
rect 26684 58828 26740 58884
rect 28428 61178 28484 61180
rect 28428 61126 28430 61178
rect 28430 61126 28482 61178
rect 28482 61126 28484 61178
rect 28428 61124 28484 61126
rect 28532 61178 28588 61180
rect 28532 61126 28534 61178
rect 28534 61126 28586 61178
rect 28586 61126 28588 61178
rect 28532 61124 28588 61126
rect 28636 61178 28692 61180
rect 28636 61126 28638 61178
rect 28638 61126 28690 61178
rect 28690 61126 28692 61178
rect 28636 61124 28692 61126
rect 28028 60172 28084 60228
rect 28140 60114 28196 60116
rect 28140 60062 28142 60114
rect 28142 60062 28194 60114
rect 28194 60062 28196 60114
rect 28140 60060 28196 60062
rect 28428 59610 28484 59612
rect 28428 59558 28430 59610
rect 28430 59558 28482 59610
rect 28482 59558 28484 59610
rect 28428 59556 28484 59558
rect 28532 59610 28588 59612
rect 28532 59558 28534 59610
rect 28534 59558 28586 59610
rect 28586 59558 28588 59610
rect 28532 59556 28588 59558
rect 28636 59610 28692 59612
rect 28636 59558 28638 59610
rect 28638 59558 28690 59610
rect 28690 59558 28692 59610
rect 28636 59556 28692 59558
rect 27356 59330 27412 59332
rect 27356 59278 27358 59330
rect 27358 59278 27410 59330
rect 27410 59278 27412 59330
rect 27356 59276 27412 59278
rect 27244 58268 27300 58324
rect 26908 57650 26964 57652
rect 26908 57598 26910 57650
rect 26910 57598 26962 57650
rect 26962 57598 26964 57650
rect 26908 57596 26964 57598
rect 26796 57372 26852 57428
rect 26796 57036 26852 57092
rect 27020 57036 27076 57092
rect 26684 56924 26740 56980
rect 27692 56978 27748 56980
rect 27692 56926 27694 56978
rect 27694 56926 27746 56978
rect 27746 56926 27748 56978
rect 27692 56924 27748 56926
rect 26460 55356 26516 55412
rect 26236 54572 26292 54628
rect 26348 54684 26404 54740
rect 26124 53618 26180 53620
rect 26124 53566 26126 53618
rect 26126 53566 26178 53618
rect 26178 53566 26180 53618
rect 26124 53564 26180 53566
rect 26572 55074 26628 55076
rect 26572 55022 26574 55074
rect 26574 55022 26626 55074
rect 26626 55022 26628 55074
rect 26572 55020 26628 55022
rect 26908 56754 26964 56756
rect 26908 56702 26910 56754
rect 26910 56702 26962 56754
rect 26962 56702 26964 56754
rect 26908 56700 26964 56702
rect 27020 55356 27076 55412
rect 27468 56588 27524 56644
rect 26796 55298 26852 55300
rect 26796 55246 26798 55298
rect 26798 55246 26850 55298
rect 26850 55246 26852 55298
rect 26796 55244 26852 55246
rect 27356 55298 27412 55300
rect 27356 55246 27358 55298
rect 27358 55246 27410 55298
rect 27410 55246 27412 55298
rect 27356 55244 27412 55246
rect 27244 55186 27300 55188
rect 27244 55134 27246 55186
rect 27246 55134 27298 55186
rect 27298 55134 27300 55186
rect 27244 55132 27300 55134
rect 26460 53900 26516 53956
rect 26348 53730 26404 53732
rect 26348 53678 26350 53730
rect 26350 53678 26402 53730
rect 26402 53678 26404 53730
rect 26348 53676 26404 53678
rect 26796 53730 26852 53732
rect 26796 53678 26798 53730
rect 26798 53678 26850 53730
rect 26850 53678 26852 53730
rect 26796 53676 26852 53678
rect 26684 53618 26740 53620
rect 26684 53566 26686 53618
rect 26686 53566 26738 53618
rect 26738 53566 26740 53618
rect 26684 53564 26740 53566
rect 26236 52274 26292 52276
rect 26236 52222 26238 52274
rect 26238 52222 26290 52274
rect 26290 52222 26292 52274
rect 26236 52220 26292 52222
rect 26236 52050 26292 52052
rect 26236 51998 26238 52050
rect 26238 51998 26290 52050
rect 26290 51998 26292 52050
rect 26236 51996 26292 51998
rect 26012 51884 26068 51940
rect 26684 53340 26740 53396
rect 26572 53228 26628 53284
rect 26572 52050 26628 52052
rect 26572 51998 26574 52050
rect 26574 51998 26626 52050
rect 26626 51998 26628 52050
rect 26572 51996 26628 51998
rect 26348 51884 26404 51940
rect 26236 51490 26292 51492
rect 26236 51438 26238 51490
rect 26238 51438 26290 51490
rect 26290 51438 26292 51490
rect 26236 51436 26292 51438
rect 26460 51378 26516 51380
rect 26460 51326 26462 51378
rect 26462 51326 26514 51378
rect 26514 51326 26516 51378
rect 26460 51324 26516 51326
rect 26236 50988 26292 51044
rect 27020 53452 27076 53508
rect 26796 52780 26852 52836
rect 27132 54796 27188 54852
rect 27132 53228 27188 53284
rect 27244 53564 27300 53620
rect 27132 52162 27188 52164
rect 27132 52110 27134 52162
rect 27134 52110 27186 52162
rect 27186 52110 27188 52162
rect 27132 52108 27188 52110
rect 28428 58042 28484 58044
rect 28428 57990 28430 58042
rect 28430 57990 28482 58042
rect 28482 57990 28484 58042
rect 28428 57988 28484 57990
rect 28532 58042 28588 58044
rect 28532 57990 28534 58042
rect 28534 57990 28586 58042
rect 28586 57990 28588 58042
rect 28532 57988 28588 57990
rect 28636 58042 28692 58044
rect 28636 57990 28638 58042
rect 28638 57990 28690 58042
rect 28690 57990 28692 58042
rect 28636 57988 28692 57990
rect 27916 57036 27972 57092
rect 28140 56978 28196 56980
rect 28140 56926 28142 56978
rect 28142 56926 28194 56978
rect 28194 56926 28196 56978
rect 28140 56924 28196 56926
rect 28428 56474 28484 56476
rect 28428 56422 28430 56474
rect 28430 56422 28482 56474
rect 28482 56422 28484 56474
rect 28428 56420 28484 56422
rect 28532 56474 28588 56476
rect 28532 56422 28534 56474
rect 28534 56422 28586 56474
rect 28586 56422 28588 56474
rect 28532 56420 28588 56422
rect 28636 56474 28692 56476
rect 28636 56422 28638 56474
rect 28638 56422 28690 56474
rect 28690 56422 28692 56474
rect 28636 56420 28692 56422
rect 27692 54460 27748 54516
rect 27692 53618 27748 53620
rect 27692 53566 27694 53618
rect 27694 53566 27746 53618
rect 27746 53566 27748 53618
rect 27692 53564 27748 53566
rect 27580 53452 27636 53508
rect 27468 52668 27524 52724
rect 27580 52050 27636 52052
rect 27580 51998 27582 52050
rect 27582 51998 27634 52050
rect 27634 51998 27636 52050
rect 27580 51996 27636 51998
rect 26908 51436 26964 51492
rect 25900 49084 25956 49140
rect 26012 49420 26068 49476
rect 26572 49308 26628 49364
rect 26348 49026 26404 49028
rect 26348 48974 26350 49026
rect 26350 48974 26402 49026
rect 26402 48974 26404 49026
rect 26348 48972 26404 48974
rect 26572 48972 26628 49028
rect 25564 45052 25620 45108
rect 25228 44828 25284 44884
rect 25026 44714 25082 44716
rect 25026 44662 25028 44714
rect 25028 44662 25080 44714
rect 25080 44662 25082 44714
rect 25026 44660 25082 44662
rect 25130 44714 25186 44716
rect 25130 44662 25132 44714
rect 25132 44662 25184 44714
rect 25184 44662 25186 44714
rect 25130 44660 25186 44662
rect 25234 44714 25290 44716
rect 25234 44662 25236 44714
rect 25236 44662 25288 44714
rect 25288 44662 25290 44714
rect 25234 44660 25290 44662
rect 25788 46674 25844 46676
rect 25788 46622 25790 46674
rect 25790 46622 25842 46674
rect 25842 46622 25844 46674
rect 25788 46620 25844 46622
rect 25788 45388 25844 45444
rect 25026 43146 25082 43148
rect 25026 43094 25028 43146
rect 25028 43094 25080 43146
rect 25080 43094 25082 43146
rect 25026 43092 25082 43094
rect 25130 43146 25186 43148
rect 25130 43094 25132 43146
rect 25132 43094 25184 43146
rect 25184 43094 25186 43146
rect 25130 43092 25186 43094
rect 25234 43146 25290 43148
rect 25234 43094 25236 43146
rect 25236 43094 25288 43146
rect 25288 43094 25290 43146
rect 25234 43092 25290 43094
rect 25228 41858 25284 41860
rect 25228 41806 25230 41858
rect 25230 41806 25282 41858
rect 25282 41806 25284 41858
rect 25228 41804 25284 41806
rect 25026 41578 25082 41580
rect 25026 41526 25028 41578
rect 25028 41526 25080 41578
rect 25080 41526 25082 41578
rect 25026 41524 25082 41526
rect 25130 41578 25186 41580
rect 25130 41526 25132 41578
rect 25132 41526 25184 41578
rect 25184 41526 25186 41578
rect 25130 41524 25186 41526
rect 25234 41578 25290 41580
rect 25234 41526 25236 41578
rect 25236 41526 25288 41578
rect 25288 41526 25290 41578
rect 25234 41524 25290 41526
rect 25116 41298 25172 41300
rect 25116 41246 25118 41298
rect 25118 41246 25170 41298
rect 25170 41246 25172 41298
rect 25116 41244 25172 41246
rect 25340 40796 25396 40852
rect 25026 40010 25082 40012
rect 25026 39958 25028 40010
rect 25028 39958 25080 40010
rect 25080 39958 25082 40010
rect 25026 39956 25082 39958
rect 25130 40010 25186 40012
rect 25130 39958 25132 40010
rect 25132 39958 25184 40010
rect 25184 39958 25186 40010
rect 25130 39956 25186 39958
rect 25234 40010 25290 40012
rect 25234 39958 25236 40010
rect 25236 39958 25288 40010
rect 25288 39958 25290 40010
rect 25234 39956 25290 39958
rect 25116 39506 25172 39508
rect 25116 39454 25118 39506
rect 25118 39454 25170 39506
rect 25170 39454 25172 39506
rect 25116 39452 25172 39454
rect 25228 38892 25284 38948
rect 25026 38442 25082 38444
rect 25026 38390 25028 38442
rect 25028 38390 25080 38442
rect 25080 38390 25082 38442
rect 25026 38388 25082 38390
rect 25130 38442 25186 38444
rect 25130 38390 25132 38442
rect 25132 38390 25184 38442
rect 25184 38390 25186 38442
rect 25130 38388 25186 38390
rect 25234 38442 25290 38444
rect 25234 38390 25236 38442
rect 25236 38390 25288 38442
rect 25288 38390 25290 38442
rect 25234 38388 25290 38390
rect 25228 38220 25284 38276
rect 25116 37548 25172 37604
rect 25228 37490 25284 37492
rect 25228 37438 25230 37490
rect 25230 37438 25282 37490
rect 25282 37438 25284 37490
rect 25228 37436 25284 37438
rect 25564 43820 25620 43876
rect 25564 43596 25620 43652
rect 25564 42700 25620 42756
rect 25564 41916 25620 41972
rect 25564 41580 25620 41636
rect 25788 43762 25844 43764
rect 25788 43710 25790 43762
rect 25790 43710 25842 43762
rect 25842 43710 25844 43762
rect 25788 43708 25844 43710
rect 26684 48914 26740 48916
rect 26684 48862 26686 48914
rect 26686 48862 26738 48914
rect 26738 48862 26740 48914
rect 26684 48860 26740 48862
rect 26124 48076 26180 48132
rect 26012 47068 26068 47124
rect 26012 43708 26068 43764
rect 25900 43314 25956 43316
rect 25900 43262 25902 43314
rect 25902 43262 25954 43314
rect 25954 43262 25956 43314
rect 25900 43260 25956 43262
rect 26348 47180 26404 47236
rect 26236 45836 26292 45892
rect 26236 45388 26292 45444
rect 27020 50988 27076 51044
rect 27244 50652 27300 50708
rect 26908 48860 26964 48916
rect 27468 49698 27524 49700
rect 27468 49646 27470 49698
rect 27470 49646 27522 49698
rect 27522 49646 27524 49698
rect 27468 49644 27524 49646
rect 27132 49532 27188 49588
rect 26684 46956 26740 47012
rect 27244 46956 27300 47012
rect 27132 46898 27188 46900
rect 27132 46846 27134 46898
rect 27134 46846 27186 46898
rect 27186 46846 27188 46898
rect 27132 46844 27188 46846
rect 26572 46396 26628 46452
rect 26460 44940 26516 44996
rect 27244 45948 27300 46004
rect 27804 51324 27860 51380
rect 28028 55356 28084 55412
rect 28140 55244 28196 55300
rect 28428 54906 28484 54908
rect 28428 54854 28430 54906
rect 28430 54854 28482 54906
rect 28482 54854 28484 54906
rect 28428 54852 28484 54854
rect 28532 54906 28588 54908
rect 28532 54854 28534 54906
rect 28534 54854 28586 54906
rect 28586 54854 28588 54906
rect 28532 54852 28588 54854
rect 28636 54906 28692 54908
rect 28636 54854 28638 54906
rect 28638 54854 28690 54906
rect 28690 54854 28692 54906
rect 28636 54852 28692 54854
rect 28028 53788 28084 53844
rect 28140 53506 28196 53508
rect 28140 53454 28142 53506
rect 28142 53454 28194 53506
rect 28194 53454 28196 53506
rect 28140 53452 28196 53454
rect 28428 53338 28484 53340
rect 28428 53286 28430 53338
rect 28430 53286 28482 53338
rect 28482 53286 28484 53338
rect 28428 53284 28484 53286
rect 28532 53338 28588 53340
rect 28532 53286 28534 53338
rect 28534 53286 28586 53338
rect 28586 53286 28588 53338
rect 28532 53284 28588 53286
rect 28636 53338 28692 53340
rect 28636 53286 28638 53338
rect 28638 53286 28690 53338
rect 28690 53286 28692 53338
rect 28636 53284 28692 53286
rect 28140 52834 28196 52836
rect 28140 52782 28142 52834
rect 28142 52782 28194 52834
rect 28194 52782 28196 52834
rect 28140 52780 28196 52782
rect 28428 51770 28484 51772
rect 28428 51718 28430 51770
rect 28430 51718 28482 51770
rect 28482 51718 28484 51770
rect 28428 51716 28484 51718
rect 28532 51770 28588 51772
rect 28532 51718 28534 51770
rect 28534 51718 28586 51770
rect 28586 51718 28588 51770
rect 28532 51716 28588 51718
rect 28636 51770 28692 51772
rect 28636 51718 28638 51770
rect 28638 51718 28690 51770
rect 28690 51718 28692 51770
rect 28636 51716 28692 51718
rect 27804 46956 27860 47012
rect 28428 50202 28484 50204
rect 28428 50150 28430 50202
rect 28430 50150 28482 50202
rect 28482 50150 28484 50202
rect 28428 50148 28484 50150
rect 28532 50202 28588 50204
rect 28532 50150 28534 50202
rect 28534 50150 28586 50202
rect 28586 50150 28588 50202
rect 28532 50148 28588 50150
rect 28636 50202 28692 50204
rect 28636 50150 28638 50202
rect 28638 50150 28690 50202
rect 28690 50150 28692 50202
rect 28636 50148 28692 50150
rect 28428 48634 28484 48636
rect 28428 48582 28430 48634
rect 28430 48582 28482 48634
rect 28482 48582 28484 48634
rect 28428 48580 28484 48582
rect 28532 48634 28588 48636
rect 28532 48582 28534 48634
rect 28534 48582 28586 48634
rect 28586 48582 28588 48634
rect 28532 48580 28588 48582
rect 28636 48634 28692 48636
rect 28636 48582 28638 48634
rect 28638 48582 28690 48634
rect 28690 48582 28692 48634
rect 28636 48580 28692 48582
rect 28428 47066 28484 47068
rect 28428 47014 28430 47066
rect 28430 47014 28482 47066
rect 28482 47014 28484 47066
rect 28428 47012 28484 47014
rect 28532 47066 28588 47068
rect 28532 47014 28534 47066
rect 28534 47014 28586 47066
rect 28586 47014 28588 47066
rect 28532 47012 28588 47014
rect 28636 47066 28692 47068
rect 28636 47014 28638 47066
rect 28638 47014 28690 47066
rect 28690 47014 28692 47066
rect 28636 47012 28692 47014
rect 27356 45836 27412 45892
rect 26796 45052 26852 45108
rect 27468 45052 27524 45108
rect 27356 44994 27412 44996
rect 27356 44942 27358 44994
rect 27358 44942 27410 44994
rect 27410 44942 27412 44994
rect 27356 44940 27412 44942
rect 27132 44828 27188 44884
rect 26684 43820 26740 43876
rect 26236 43372 26292 43428
rect 26460 43484 26516 43540
rect 26124 42028 26180 42084
rect 26348 43260 26404 43316
rect 26012 41580 26068 41636
rect 25788 40962 25844 40964
rect 25788 40910 25790 40962
rect 25790 40910 25842 40962
rect 25842 40910 25844 40962
rect 25788 40908 25844 40910
rect 25676 38556 25732 38612
rect 25676 37772 25732 37828
rect 25676 37548 25732 37604
rect 25340 37266 25396 37268
rect 25340 37214 25342 37266
rect 25342 37214 25394 37266
rect 25394 37214 25396 37266
rect 25340 37212 25396 37214
rect 25026 36874 25082 36876
rect 25026 36822 25028 36874
rect 25028 36822 25080 36874
rect 25080 36822 25082 36874
rect 25026 36820 25082 36822
rect 25130 36874 25186 36876
rect 25130 36822 25132 36874
rect 25132 36822 25184 36874
rect 25184 36822 25186 36874
rect 25130 36820 25186 36822
rect 25234 36874 25290 36876
rect 25234 36822 25236 36874
rect 25236 36822 25288 36874
rect 25288 36822 25290 36874
rect 25234 36820 25290 36822
rect 25452 36652 25508 36708
rect 25228 36540 25284 36596
rect 25026 35306 25082 35308
rect 25026 35254 25028 35306
rect 25028 35254 25080 35306
rect 25080 35254 25082 35306
rect 25026 35252 25082 35254
rect 25130 35306 25186 35308
rect 25130 35254 25132 35306
rect 25132 35254 25184 35306
rect 25184 35254 25186 35306
rect 25130 35252 25186 35254
rect 25234 35306 25290 35308
rect 25234 35254 25236 35306
rect 25236 35254 25288 35306
rect 25288 35254 25290 35306
rect 25234 35252 25290 35254
rect 25004 35084 25060 35140
rect 24668 34636 24724 34692
rect 24668 32450 24724 32452
rect 24668 32398 24670 32450
rect 24670 32398 24722 32450
rect 24722 32398 24724 32450
rect 24668 32396 24724 32398
rect 24668 31666 24724 31668
rect 24668 31614 24670 31666
rect 24670 31614 24722 31666
rect 24722 31614 24724 31666
rect 24668 31612 24724 31614
rect 24668 30828 24724 30884
rect 24668 30044 24724 30100
rect 25116 34690 25172 34692
rect 25116 34638 25118 34690
rect 25118 34638 25170 34690
rect 25170 34638 25172 34690
rect 25116 34636 25172 34638
rect 25340 34748 25396 34804
rect 25026 33738 25082 33740
rect 25026 33686 25028 33738
rect 25028 33686 25080 33738
rect 25080 33686 25082 33738
rect 25026 33684 25082 33686
rect 25130 33738 25186 33740
rect 25130 33686 25132 33738
rect 25132 33686 25184 33738
rect 25184 33686 25186 33738
rect 25130 33684 25186 33686
rect 25234 33738 25290 33740
rect 25234 33686 25236 33738
rect 25236 33686 25288 33738
rect 25288 33686 25290 33738
rect 25234 33684 25290 33686
rect 25340 33516 25396 33572
rect 25228 33292 25284 33348
rect 25452 32732 25508 32788
rect 25026 32170 25082 32172
rect 25026 32118 25028 32170
rect 25028 32118 25080 32170
rect 25080 32118 25082 32170
rect 25026 32116 25082 32118
rect 25130 32170 25186 32172
rect 25130 32118 25132 32170
rect 25132 32118 25184 32170
rect 25184 32118 25186 32170
rect 25130 32116 25186 32118
rect 25234 32170 25290 32172
rect 25234 32118 25236 32170
rect 25236 32118 25288 32170
rect 25288 32118 25290 32170
rect 25234 32116 25290 32118
rect 25900 40236 25956 40292
rect 25788 37436 25844 37492
rect 25676 35532 25732 35588
rect 25900 35138 25956 35140
rect 25900 35086 25902 35138
rect 25902 35086 25954 35138
rect 25954 35086 25956 35138
rect 25900 35084 25956 35086
rect 25676 34300 25732 34356
rect 25900 34636 25956 34692
rect 25900 34130 25956 34132
rect 25900 34078 25902 34130
rect 25902 34078 25954 34130
rect 25954 34078 25956 34130
rect 25900 34076 25956 34078
rect 26236 41132 26292 41188
rect 26572 43260 26628 43316
rect 26796 43538 26852 43540
rect 26796 43486 26798 43538
rect 26798 43486 26850 43538
rect 26850 43486 26852 43538
rect 26796 43484 26852 43486
rect 26684 42642 26740 42644
rect 26684 42590 26686 42642
rect 26686 42590 26738 42642
rect 26738 42590 26740 42642
rect 26684 42588 26740 42590
rect 26572 41132 26628 41188
rect 26796 41132 26852 41188
rect 27020 41804 27076 41860
rect 26236 40572 26292 40628
rect 26348 40514 26404 40516
rect 26348 40462 26350 40514
rect 26350 40462 26402 40514
rect 26402 40462 26404 40514
rect 26348 40460 26404 40462
rect 26460 40236 26516 40292
rect 26572 40124 26628 40180
rect 26236 38668 26292 38724
rect 26572 39004 26628 39060
rect 26348 38108 26404 38164
rect 26460 37996 26516 38052
rect 26796 40962 26852 40964
rect 26796 40910 26798 40962
rect 26798 40910 26850 40962
rect 26850 40910 26852 40962
rect 26796 40908 26852 40910
rect 27020 40908 27076 40964
rect 26908 40572 26964 40628
rect 27244 43538 27300 43540
rect 27244 43486 27246 43538
rect 27246 43486 27298 43538
rect 27298 43486 27300 43538
rect 27244 43484 27300 43486
rect 27356 43372 27412 43428
rect 27132 40460 27188 40516
rect 26796 40402 26852 40404
rect 26796 40350 26798 40402
rect 26798 40350 26850 40402
rect 26850 40350 26852 40402
rect 26796 40348 26852 40350
rect 26908 40124 26964 40180
rect 26796 39842 26852 39844
rect 26796 39790 26798 39842
rect 26798 39790 26850 39842
rect 26850 39790 26852 39842
rect 26796 39788 26852 39790
rect 27020 39394 27076 39396
rect 27020 39342 27022 39394
rect 27022 39342 27074 39394
rect 27074 39342 27076 39394
rect 27020 39340 27076 39342
rect 26908 38780 26964 38836
rect 26236 36876 26292 36932
rect 26348 37436 26404 37492
rect 26236 36652 26292 36708
rect 26236 35026 26292 35028
rect 26236 34974 26238 35026
rect 26238 34974 26290 35026
rect 26290 34974 26292 35026
rect 26236 34972 26292 34974
rect 26572 36764 26628 36820
rect 26572 35532 26628 35588
rect 26460 34860 26516 34916
rect 27468 41916 27524 41972
rect 27356 41858 27412 41860
rect 27356 41806 27358 41858
rect 27358 41806 27410 41858
rect 27410 41806 27412 41858
rect 27356 41804 27412 41806
rect 27804 45890 27860 45892
rect 27804 45838 27806 45890
rect 27806 45838 27858 45890
rect 27858 45838 27860 45890
rect 27804 45836 27860 45838
rect 27692 43372 27748 43428
rect 27580 41244 27636 41300
rect 27692 42700 27748 42756
rect 27580 41020 27636 41076
rect 27356 39842 27412 39844
rect 27356 39790 27358 39842
rect 27358 39790 27410 39842
rect 27410 39790 27412 39842
rect 27356 39788 27412 39790
rect 27356 39340 27412 39396
rect 27468 38892 27524 38948
rect 26796 37324 26852 37380
rect 26908 36540 26964 36596
rect 27356 37884 27412 37940
rect 28428 45498 28484 45500
rect 28428 45446 28430 45498
rect 28430 45446 28482 45498
rect 28482 45446 28484 45498
rect 28428 45444 28484 45446
rect 28532 45498 28588 45500
rect 28532 45446 28534 45498
rect 28534 45446 28586 45498
rect 28586 45446 28588 45498
rect 28532 45444 28588 45446
rect 28636 45498 28692 45500
rect 28636 45446 28638 45498
rect 28638 45446 28690 45498
rect 28690 45446 28692 45498
rect 28636 45444 28692 45446
rect 28140 45106 28196 45108
rect 28140 45054 28142 45106
rect 28142 45054 28194 45106
rect 28194 45054 28196 45106
rect 28140 45052 28196 45054
rect 28428 43930 28484 43932
rect 28428 43878 28430 43930
rect 28430 43878 28482 43930
rect 28482 43878 28484 43930
rect 28428 43876 28484 43878
rect 28532 43930 28588 43932
rect 28532 43878 28534 43930
rect 28534 43878 28586 43930
rect 28586 43878 28588 43930
rect 28532 43876 28588 43878
rect 28636 43930 28692 43932
rect 28636 43878 28638 43930
rect 28638 43878 28690 43930
rect 28690 43878 28692 43930
rect 28636 43876 28692 43878
rect 28140 43650 28196 43652
rect 28140 43598 28142 43650
rect 28142 43598 28194 43650
rect 28194 43598 28196 43650
rect 28140 43596 28196 43598
rect 27692 39842 27748 39844
rect 27692 39790 27694 39842
rect 27694 39790 27746 39842
rect 27746 39790 27748 39842
rect 27692 39788 27748 39790
rect 27692 37660 27748 37716
rect 28428 42362 28484 42364
rect 28428 42310 28430 42362
rect 28430 42310 28482 42362
rect 28482 42310 28484 42362
rect 28428 42308 28484 42310
rect 28532 42362 28588 42364
rect 28532 42310 28534 42362
rect 28534 42310 28586 42362
rect 28586 42310 28588 42362
rect 28532 42308 28588 42310
rect 28636 42362 28692 42364
rect 28636 42310 28638 42362
rect 28638 42310 28690 42362
rect 28690 42310 28692 42362
rect 28636 42308 28692 42310
rect 28028 41970 28084 41972
rect 28028 41918 28030 41970
rect 28030 41918 28082 41970
rect 28082 41918 28084 41970
rect 28028 41916 28084 41918
rect 28428 40794 28484 40796
rect 28428 40742 28430 40794
rect 28430 40742 28482 40794
rect 28482 40742 28484 40794
rect 28428 40740 28484 40742
rect 28532 40794 28588 40796
rect 28532 40742 28534 40794
rect 28534 40742 28586 40794
rect 28586 40742 28588 40794
rect 28532 40740 28588 40742
rect 28636 40794 28692 40796
rect 28636 40742 28638 40794
rect 28638 40742 28690 40794
rect 28690 40742 28692 40794
rect 28636 40740 28692 40742
rect 28140 40626 28196 40628
rect 28140 40574 28142 40626
rect 28142 40574 28194 40626
rect 28194 40574 28196 40626
rect 28140 40572 28196 40574
rect 28140 39788 28196 39844
rect 28428 39226 28484 39228
rect 28428 39174 28430 39226
rect 28430 39174 28482 39226
rect 28482 39174 28484 39226
rect 28428 39172 28484 39174
rect 28532 39226 28588 39228
rect 28532 39174 28534 39226
rect 28534 39174 28586 39226
rect 28586 39174 28588 39226
rect 28532 39172 28588 39174
rect 28636 39226 28692 39228
rect 28636 39174 28638 39226
rect 28638 39174 28690 39226
rect 28690 39174 28692 39226
rect 28636 39172 28692 39174
rect 27020 36482 27076 36484
rect 27020 36430 27022 36482
rect 27022 36430 27074 36482
rect 27074 36430 27076 36482
rect 27020 36428 27076 36430
rect 26684 34972 26740 35028
rect 26796 36316 26852 36372
rect 26572 34748 26628 34804
rect 26124 34412 26180 34468
rect 26348 34300 26404 34356
rect 25676 33964 25732 34020
rect 26460 33906 26516 33908
rect 26460 33854 26462 33906
rect 26462 33854 26514 33906
rect 26514 33854 26516 33906
rect 26460 33852 26516 33854
rect 26348 32732 26404 32788
rect 25564 32620 25620 32676
rect 26124 32396 26180 32452
rect 26460 32396 26516 32452
rect 24780 29820 24836 29876
rect 24892 31164 24948 31220
rect 24556 29260 24612 29316
rect 24444 28812 24500 28868
rect 23660 27074 23716 27076
rect 23660 27022 23662 27074
rect 23662 27022 23714 27074
rect 23714 27022 23716 27074
rect 23660 27020 23716 27022
rect 23548 26236 23604 26292
rect 23660 26460 23716 26516
rect 23100 25452 23156 25508
rect 22988 25340 23044 25396
rect 23548 25900 23604 25956
rect 22764 23714 22820 23716
rect 22764 23662 22766 23714
rect 22766 23662 22818 23714
rect 22818 23662 22820 23714
rect 22764 23660 22820 23662
rect 22652 23266 22708 23268
rect 22652 23214 22654 23266
rect 22654 23214 22706 23266
rect 22706 23214 22708 23266
rect 22652 23212 22708 23214
rect 23436 23660 23492 23716
rect 23100 23324 23156 23380
rect 22652 22876 22708 22932
rect 22988 22652 23044 22708
rect 22876 22428 22932 22484
rect 22764 21868 22820 21924
rect 22652 21532 22708 21588
rect 22652 20802 22708 20804
rect 22652 20750 22654 20802
rect 22654 20750 22706 20802
rect 22706 20750 22708 20802
rect 22652 20748 22708 20750
rect 22540 19404 22596 19460
rect 22652 19346 22708 19348
rect 22652 19294 22654 19346
rect 22654 19294 22706 19346
rect 22706 19294 22708 19346
rect 22652 19292 22708 19294
rect 22428 19180 22484 19236
rect 22316 18956 22372 19012
rect 23100 21756 23156 21812
rect 22876 20748 22932 20804
rect 22876 20524 22932 20580
rect 22092 18172 22148 18228
rect 21756 17052 21812 17108
rect 22204 16882 22260 16884
rect 22204 16830 22206 16882
rect 22206 16830 22258 16882
rect 22258 16830 22260 16882
rect 22204 16828 22260 16830
rect 21308 16098 21364 16100
rect 21308 16046 21310 16098
rect 21310 16046 21362 16098
rect 21362 16046 21364 16098
rect 21308 16044 21364 16046
rect 21624 15706 21680 15708
rect 21624 15654 21626 15706
rect 21626 15654 21678 15706
rect 21678 15654 21680 15706
rect 21624 15652 21680 15654
rect 21728 15706 21784 15708
rect 21728 15654 21730 15706
rect 21730 15654 21782 15706
rect 21782 15654 21784 15706
rect 21728 15652 21784 15654
rect 21832 15706 21888 15708
rect 21832 15654 21834 15706
rect 21834 15654 21886 15706
rect 21886 15654 21888 15706
rect 21832 15652 21888 15654
rect 21196 15202 21252 15204
rect 21196 15150 21198 15202
rect 21198 15150 21250 15202
rect 21250 15150 21252 15202
rect 21196 15148 21252 15150
rect 21532 14588 21588 14644
rect 21196 14364 21252 14420
rect 22204 15148 22260 15204
rect 21624 14138 21680 14140
rect 21624 14086 21626 14138
rect 21626 14086 21678 14138
rect 21678 14086 21680 14138
rect 21624 14084 21680 14086
rect 21728 14138 21784 14140
rect 21728 14086 21730 14138
rect 21730 14086 21782 14138
rect 21782 14086 21784 14138
rect 21728 14084 21784 14086
rect 21832 14138 21888 14140
rect 21832 14086 21834 14138
rect 21834 14086 21886 14138
rect 21886 14086 21888 14138
rect 21832 14084 21888 14086
rect 21980 13692 22036 13748
rect 20972 12684 21028 12740
rect 20748 11394 20804 11396
rect 20748 11342 20750 11394
rect 20750 11342 20802 11394
rect 20802 11342 20804 11394
rect 20748 11340 20804 11342
rect 21624 12570 21680 12572
rect 21624 12518 21626 12570
rect 21626 12518 21678 12570
rect 21678 12518 21680 12570
rect 21624 12516 21680 12518
rect 21728 12570 21784 12572
rect 21728 12518 21730 12570
rect 21730 12518 21782 12570
rect 21782 12518 21784 12570
rect 21728 12516 21784 12518
rect 21832 12570 21888 12572
rect 21832 12518 21834 12570
rect 21834 12518 21886 12570
rect 21886 12518 21888 12570
rect 21832 12516 21888 12518
rect 21756 12402 21812 12404
rect 21756 12350 21758 12402
rect 21758 12350 21810 12402
rect 21810 12350 21812 12402
rect 21756 12348 21812 12350
rect 22092 14252 22148 14308
rect 22204 12348 22260 12404
rect 21980 12124 22036 12180
rect 21308 11506 21364 11508
rect 21308 11454 21310 11506
rect 21310 11454 21362 11506
rect 21362 11454 21364 11506
rect 21308 11452 21364 11454
rect 22764 17164 22820 17220
rect 22652 16994 22708 16996
rect 22652 16942 22654 16994
rect 22654 16942 22706 16994
rect 22706 16942 22708 16994
rect 22652 16940 22708 16942
rect 22652 15708 22708 15764
rect 23100 20242 23156 20244
rect 23100 20190 23102 20242
rect 23102 20190 23154 20242
rect 23154 20190 23156 20242
rect 23100 20188 23156 20190
rect 23100 18620 23156 18676
rect 22988 17612 23044 17668
rect 23436 22428 23492 22484
rect 23548 21868 23604 21924
rect 23884 26514 23940 26516
rect 23884 26462 23886 26514
rect 23886 26462 23938 26514
rect 23938 26462 23940 26514
rect 23884 26460 23940 26462
rect 23772 25394 23828 25396
rect 23772 25342 23774 25394
rect 23774 25342 23826 25394
rect 23826 25342 23828 25394
rect 23772 25340 23828 25342
rect 23772 25116 23828 25172
rect 24780 28642 24836 28644
rect 24780 28590 24782 28642
rect 24782 28590 24834 28642
rect 24834 28590 24836 28642
rect 24780 28588 24836 28590
rect 25340 30882 25396 30884
rect 25340 30830 25342 30882
rect 25342 30830 25394 30882
rect 25394 30830 25396 30882
rect 25340 30828 25396 30830
rect 25026 30602 25082 30604
rect 25026 30550 25028 30602
rect 25028 30550 25080 30602
rect 25080 30550 25082 30602
rect 25026 30548 25082 30550
rect 25130 30602 25186 30604
rect 25130 30550 25132 30602
rect 25132 30550 25184 30602
rect 25184 30550 25186 30602
rect 25130 30548 25186 30550
rect 25234 30602 25290 30604
rect 25234 30550 25236 30602
rect 25236 30550 25288 30602
rect 25288 30550 25290 30602
rect 25234 30548 25290 30550
rect 25340 29820 25396 29876
rect 25228 29314 25284 29316
rect 25228 29262 25230 29314
rect 25230 29262 25282 29314
rect 25282 29262 25284 29314
rect 25228 29260 25284 29262
rect 25026 29034 25082 29036
rect 25026 28982 25028 29034
rect 25028 28982 25080 29034
rect 25080 28982 25082 29034
rect 25026 28980 25082 28982
rect 25130 29034 25186 29036
rect 25130 28982 25132 29034
rect 25132 28982 25184 29034
rect 25184 28982 25186 29034
rect 25130 28980 25186 28982
rect 25234 29034 25290 29036
rect 25234 28982 25236 29034
rect 25236 28982 25288 29034
rect 25288 28982 25290 29034
rect 25234 28980 25290 28982
rect 25340 28700 25396 28756
rect 25004 28642 25060 28644
rect 25004 28590 25006 28642
rect 25006 28590 25058 28642
rect 25058 28590 25060 28642
rect 25004 28588 25060 28590
rect 24108 25004 24164 25060
rect 24220 27468 24276 27524
rect 23772 23436 23828 23492
rect 24444 27186 24500 27188
rect 24444 27134 24446 27186
rect 24446 27134 24498 27186
rect 24498 27134 24500 27186
rect 24444 27132 24500 27134
rect 23996 23714 24052 23716
rect 23996 23662 23998 23714
rect 23998 23662 24050 23714
rect 24050 23662 24052 23714
rect 23996 23660 24052 23662
rect 23996 23436 24052 23492
rect 23772 23266 23828 23268
rect 23772 23214 23774 23266
rect 23774 23214 23826 23266
rect 23826 23214 23828 23266
rect 23772 23212 23828 23214
rect 23884 22652 23940 22708
rect 23996 22428 24052 22484
rect 23436 21644 23492 21700
rect 23548 20188 23604 20244
rect 22876 15036 22932 15092
rect 23436 18396 23492 18452
rect 22764 12962 22820 12964
rect 22764 12910 22766 12962
rect 22766 12910 22818 12962
rect 22818 12910 22820 12962
rect 22764 12908 22820 12910
rect 22540 12684 22596 12740
rect 22316 11564 22372 11620
rect 22540 11676 22596 11732
rect 22428 11452 22484 11508
rect 22092 11116 22148 11172
rect 22316 11116 22372 11172
rect 21624 11002 21680 11004
rect 21624 10950 21626 11002
rect 21626 10950 21678 11002
rect 21678 10950 21680 11002
rect 21624 10948 21680 10950
rect 21728 11002 21784 11004
rect 21728 10950 21730 11002
rect 21730 10950 21782 11002
rect 21782 10950 21784 11002
rect 21728 10948 21784 10950
rect 21832 11002 21888 11004
rect 21832 10950 21834 11002
rect 21834 10950 21886 11002
rect 21886 10950 21888 11002
rect 21832 10948 21888 10950
rect 20524 9996 20580 10052
rect 21308 10610 21364 10612
rect 21308 10558 21310 10610
rect 21310 10558 21362 10610
rect 21362 10558 21364 10610
rect 21308 10556 21364 10558
rect 21196 10444 21252 10500
rect 22540 10780 22596 10836
rect 21644 10722 21700 10724
rect 21644 10670 21646 10722
rect 21646 10670 21698 10722
rect 21698 10670 21700 10722
rect 21644 10668 21700 10670
rect 22652 10722 22708 10724
rect 22652 10670 22654 10722
rect 22654 10670 22706 10722
rect 22706 10670 22708 10722
rect 22652 10668 22708 10670
rect 21980 10444 22036 10500
rect 21532 9996 21588 10052
rect 21624 9434 21680 9436
rect 21624 9382 21626 9434
rect 21626 9382 21678 9434
rect 21678 9382 21680 9434
rect 21624 9380 21680 9382
rect 21728 9434 21784 9436
rect 21728 9382 21730 9434
rect 21730 9382 21782 9434
rect 21782 9382 21784 9434
rect 21728 9380 21784 9382
rect 21832 9434 21888 9436
rect 21832 9382 21834 9434
rect 21834 9382 21886 9434
rect 21886 9382 21888 9434
rect 21832 9380 21888 9382
rect 20636 8316 20692 8372
rect 20972 8930 21028 8932
rect 20972 8878 20974 8930
rect 20974 8878 21026 8930
rect 21026 8878 21028 8930
rect 20972 8876 21028 8878
rect 20636 7980 20692 8036
rect 20524 7644 20580 7700
rect 20300 7308 20356 7364
rect 20076 6018 20132 6020
rect 20076 5966 20078 6018
rect 20078 5966 20130 6018
rect 20130 5966 20132 6018
rect 20076 5964 20132 5966
rect 21196 8316 21252 8372
rect 21980 9100 22036 9156
rect 22652 8988 22708 9044
rect 20972 6636 21028 6692
rect 20524 6578 20580 6580
rect 20524 6526 20526 6578
rect 20526 6526 20578 6578
rect 20578 6526 20580 6578
rect 20524 6524 20580 6526
rect 20412 5292 20468 5348
rect 20860 5852 20916 5908
rect 21308 6578 21364 6580
rect 21308 6526 21310 6578
rect 21310 6526 21362 6578
rect 21362 6526 21364 6578
rect 21308 6524 21364 6526
rect 21624 7866 21680 7868
rect 21624 7814 21626 7866
rect 21626 7814 21678 7866
rect 21678 7814 21680 7866
rect 21624 7812 21680 7814
rect 21728 7866 21784 7868
rect 21728 7814 21730 7866
rect 21730 7814 21782 7866
rect 21782 7814 21784 7866
rect 21728 7812 21784 7814
rect 21832 7866 21888 7868
rect 21832 7814 21834 7866
rect 21834 7814 21886 7866
rect 21886 7814 21888 7866
rect 21832 7812 21888 7814
rect 22092 7644 22148 7700
rect 21644 6690 21700 6692
rect 21644 6638 21646 6690
rect 21646 6638 21698 6690
rect 21698 6638 21700 6690
rect 21644 6636 21700 6638
rect 21624 6298 21680 6300
rect 21624 6246 21626 6298
rect 21626 6246 21678 6298
rect 21678 6246 21680 6298
rect 21624 6244 21680 6246
rect 21728 6298 21784 6300
rect 21728 6246 21730 6298
rect 21730 6246 21782 6298
rect 21782 6246 21784 6298
rect 21728 6244 21784 6246
rect 21832 6298 21888 6300
rect 21832 6246 21834 6298
rect 21834 6246 21886 6298
rect 21886 6246 21888 6298
rect 21832 6244 21888 6246
rect 20412 5010 20468 5012
rect 20412 4958 20414 5010
rect 20414 4958 20466 5010
rect 20466 4958 20468 5010
rect 20412 4956 20468 4958
rect 20636 4844 20692 4900
rect 20748 5068 20804 5124
rect 20076 4620 20132 4676
rect 20636 4620 20692 4676
rect 19404 3388 19460 3444
rect 19180 3164 19236 3220
rect 19292 3052 19348 3108
rect 18956 2098 19012 2100
rect 18956 2046 18958 2098
rect 18958 2046 19010 2098
rect 19010 2046 19012 2098
rect 18956 2044 19012 2046
rect 18844 1820 18900 1876
rect 19964 3388 20020 3444
rect 20300 3724 20356 3780
rect 19404 1820 19460 1876
rect 19516 1932 19572 1988
rect 20076 2156 20132 2212
rect 19628 1874 19684 1876
rect 19628 1822 19630 1874
rect 19630 1822 19682 1874
rect 19682 1822 19684 1874
rect 19628 1820 19684 1822
rect 20524 3948 20580 4004
rect 20524 1932 20580 1988
rect 20636 3836 20692 3892
rect 20748 3164 20804 3220
rect 21868 5852 21924 5908
rect 21756 5180 21812 5236
rect 23436 17554 23492 17556
rect 23436 17502 23438 17554
rect 23438 17502 23490 17554
rect 23490 17502 23492 17554
rect 23436 17500 23492 17502
rect 23772 22316 23828 22372
rect 23996 20748 24052 20804
rect 23772 20188 23828 20244
rect 24220 24610 24276 24612
rect 24220 24558 24222 24610
rect 24222 24558 24274 24610
rect 24274 24558 24276 24610
rect 24220 24556 24276 24558
rect 24220 24332 24276 24388
rect 24556 26908 24612 26964
rect 24332 23660 24388 23716
rect 24444 25004 24500 25060
rect 25026 27466 25082 27468
rect 25026 27414 25028 27466
rect 25028 27414 25080 27466
rect 25080 27414 25082 27466
rect 25026 27412 25082 27414
rect 25130 27466 25186 27468
rect 25130 27414 25132 27466
rect 25132 27414 25184 27466
rect 25184 27414 25186 27466
rect 25130 27412 25186 27414
rect 25234 27466 25290 27468
rect 25234 27414 25236 27466
rect 25236 27414 25288 27466
rect 25288 27414 25290 27466
rect 25234 27412 25290 27414
rect 25228 27244 25284 27300
rect 25340 27020 25396 27076
rect 24892 26850 24948 26852
rect 24892 26798 24894 26850
rect 24894 26798 24946 26850
rect 24946 26798 24948 26850
rect 24892 26796 24948 26798
rect 26236 31948 26292 32004
rect 26124 31612 26180 31668
rect 26124 31106 26180 31108
rect 26124 31054 26126 31106
rect 26126 31054 26178 31106
rect 26178 31054 26180 31106
rect 26124 31052 26180 31054
rect 25900 30994 25956 30996
rect 25900 30942 25902 30994
rect 25902 30942 25954 30994
rect 25954 30942 25956 30994
rect 25900 30940 25956 30942
rect 26684 33404 26740 33460
rect 26684 32338 26740 32340
rect 26684 32286 26686 32338
rect 26686 32286 26738 32338
rect 26738 32286 26740 32338
rect 26684 32284 26740 32286
rect 27132 34636 27188 34692
rect 27356 34860 27412 34916
rect 27692 34412 27748 34468
rect 27804 34636 27860 34692
rect 27020 33906 27076 33908
rect 27020 33854 27022 33906
rect 27022 33854 27074 33906
rect 27074 33854 27076 33906
rect 27020 33852 27076 33854
rect 27020 33292 27076 33348
rect 27356 33458 27412 33460
rect 27356 33406 27358 33458
rect 27358 33406 27410 33458
rect 27410 33406 27412 33458
rect 27356 33404 27412 33406
rect 26796 32060 26852 32116
rect 26684 31612 26740 31668
rect 26236 30156 26292 30212
rect 25676 28642 25732 28644
rect 25676 28590 25678 28642
rect 25678 28590 25730 28642
rect 25730 28590 25732 28642
rect 25676 28588 25732 28590
rect 26460 28642 26516 28644
rect 26460 28590 26462 28642
rect 26462 28590 26514 28642
rect 26514 28590 26516 28642
rect 26460 28588 26516 28590
rect 25788 28364 25844 28420
rect 24892 26236 24948 26292
rect 25452 26290 25508 26292
rect 25452 26238 25454 26290
rect 25454 26238 25506 26290
rect 25506 26238 25508 26290
rect 25452 26236 25508 26238
rect 25026 25898 25082 25900
rect 25026 25846 25028 25898
rect 25028 25846 25080 25898
rect 25080 25846 25082 25898
rect 25026 25844 25082 25846
rect 25130 25898 25186 25900
rect 25130 25846 25132 25898
rect 25132 25846 25184 25898
rect 25184 25846 25186 25898
rect 25130 25844 25186 25846
rect 25234 25898 25290 25900
rect 25234 25846 25236 25898
rect 25236 25846 25288 25898
rect 25288 25846 25290 25898
rect 25234 25844 25290 25846
rect 24780 24668 24836 24724
rect 25452 24892 25508 24948
rect 24668 24610 24724 24612
rect 24668 24558 24670 24610
rect 24670 24558 24722 24610
rect 24722 24558 24724 24610
rect 24668 24556 24724 24558
rect 24556 24108 24612 24164
rect 25026 24330 25082 24332
rect 25026 24278 25028 24330
rect 25028 24278 25080 24330
rect 25080 24278 25082 24330
rect 25026 24276 25082 24278
rect 25130 24330 25186 24332
rect 25130 24278 25132 24330
rect 25132 24278 25184 24330
rect 25184 24278 25186 24330
rect 25130 24276 25186 24278
rect 25234 24330 25290 24332
rect 25234 24278 25236 24330
rect 25236 24278 25288 24330
rect 25288 24278 25290 24330
rect 25234 24276 25290 24278
rect 25340 24050 25396 24052
rect 25340 23998 25342 24050
rect 25342 23998 25394 24050
rect 25394 23998 25396 24050
rect 25340 23996 25396 23998
rect 24668 23042 24724 23044
rect 24668 22990 24670 23042
rect 24670 22990 24722 23042
rect 24722 22990 24724 23042
rect 24668 22988 24724 22990
rect 25004 23884 25060 23940
rect 24332 21810 24388 21812
rect 24332 21758 24334 21810
rect 24334 21758 24386 21810
rect 24386 21758 24388 21810
rect 24332 21756 24388 21758
rect 24220 21532 24276 21588
rect 23996 17164 24052 17220
rect 24108 17666 24164 17668
rect 24108 17614 24110 17666
rect 24110 17614 24162 17666
rect 24162 17614 24164 17666
rect 24108 17612 24164 17614
rect 24444 20636 24500 20692
rect 24444 19292 24500 19348
rect 24332 18620 24388 18676
rect 24444 18956 24500 19012
rect 23548 15148 23604 15204
rect 23212 14364 23268 14420
rect 23548 13746 23604 13748
rect 23548 13694 23550 13746
rect 23550 13694 23602 13746
rect 23602 13694 23604 13746
rect 23548 13692 23604 13694
rect 22988 12684 23044 12740
rect 24108 15314 24164 15316
rect 24108 15262 24110 15314
rect 24110 15262 24162 15314
rect 24162 15262 24164 15314
rect 24108 15260 24164 15262
rect 24668 20130 24724 20132
rect 24668 20078 24670 20130
rect 24670 20078 24722 20130
rect 24722 20078 24724 20130
rect 24668 20076 24724 20078
rect 24668 19292 24724 19348
rect 24668 18508 24724 18564
rect 24668 17164 24724 17220
rect 24556 15260 24612 15316
rect 24668 15484 24724 15540
rect 24332 14700 24388 14756
rect 24444 14364 24500 14420
rect 24220 13634 24276 13636
rect 24220 13582 24222 13634
rect 24222 13582 24274 13634
rect 24274 13582 24276 13634
rect 24220 13580 24276 13582
rect 23548 12908 23604 12964
rect 24108 13020 24164 13076
rect 23436 12124 23492 12180
rect 24108 10834 24164 10836
rect 24108 10782 24110 10834
rect 24110 10782 24162 10834
rect 24162 10782 24164 10834
rect 24108 10780 24164 10782
rect 23212 10722 23268 10724
rect 23212 10670 23214 10722
rect 23214 10670 23266 10722
rect 23266 10670 23268 10722
rect 23212 10668 23268 10670
rect 23660 10722 23716 10724
rect 23660 10670 23662 10722
rect 23662 10670 23714 10722
rect 23714 10670 23716 10722
rect 23660 10668 23716 10670
rect 24444 13074 24500 13076
rect 24444 13022 24446 13074
rect 24446 13022 24498 13074
rect 24498 13022 24500 13074
rect 24444 13020 24500 13022
rect 24668 12124 24724 12180
rect 23436 9042 23492 9044
rect 23436 8990 23438 9042
rect 23438 8990 23490 9042
rect 23490 8990 23492 9042
rect 23436 8988 23492 8990
rect 23212 7698 23268 7700
rect 23212 7646 23214 7698
rect 23214 7646 23266 7698
rect 23266 7646 23268 7698
rect 23212 7644 23268 7646
rect 22204 5628 22260 5684
rect 23884 7474 23940 7476
rect 23884 7422 23886 7474
rect 23886 7422 23938 7474
rect 23938 7422 23940 7474
rect 23884 7420 23940 7422
rect 23772 6636 23828 6692
rect 26348 28530 26404 28532
rect 26348 28478 26350 28530
rect 26350 28478 26402 28530
rect 26402 28478 26404 28530
rect 26348 28476 26404 28478
rect 26236 28364 26292 28420
rect 26124 28252 26180 28308
rect 25900 27970 25956 27972
rect 25900 27918 25902 27970
rect 25902 27918 25954 27970
rect 25954 27918 25956 27970
rect 25900 27916 25956 27918
rect 26684 28252 26740 28308
rect 26572 28140 26628 28196
rect 26124 27356 26180 27412
rect 26460 27858 26516 27860
rect 26460 27806 26462 27858
rect 26462 27806 26514 27858
rect 26514 27806 26516 27858
rect 26460 27804 26516 27806
rect 26348 27634 26404 27636
rect 26348 27582 26350 27634
rect 26350 27582 26402 27634
rect 26402 27582 26404 27634
rect 26348 27580 26404 27582
rect 26236 27020 26292 27076
rect 26460 27132 26516 27188
rect 25900 26796 25956 26852
rect 25900 26124 25956 26180
rect 25676 25340 25732 25396
rect 25900 24722 25956 24724
rect 25900 24670 25902 24722
rect 25902 24670 25954 24722
rect 25954 24670 25956 24722
rect 25900 24668 25956 24670
rect 25564 24556 25620 24612
rect 26124 24556 26180 24612
rect 25452 23772 25508 23828
rect 25004 23714 25060 23716
rect 25004 23662 25006 23714
rect 25006 23662 25058 23714
rect 25058 23662 25060 23714
rect 25004 23660 25060 23662
rect 26012 23660 26068 23716
rect 25676 23436 25732 23492
rect 25228 23212 25284 23268
rect 25026 22762 25082 22764
rect 25026 22710 25028 22762
rect 25028 22710 25080 22762
rect 25080 22710 25082 22762
rect 25026 22708 25082 22710
rect 25130 22762 25186 22764
rect 25130 22710 25132 22762
rect 25132 22710 25184 22762
rect 25184 22710 25186 22762
rect 25130 22708 25186 22710
rect 25234 22762 25290 22764
rect 25234 22710 25236 22762
rect 25236 22710 25288 22762
rect 25288 22710 25290 22762
rect 25234 22708 25290 22710
rect 25116 22540 25172 22596
rect 25116 22204 25172 22260
rect 25452 21532 25508 21588
rect 25026 21194 25082 21196
rect 25026 21142 25028 21194
rect 25028 21142 25080 21194
rect 25080 21142 25082 21194
rect 25026 21140 25082 21142
rect 25130 21194 25186 21196
rect 25130 21142 25132 21194
rect 25132 21142 25184 21194
rect 25184 21142 25186 21194
rect 25130 21140 25186 21142
rect 25234 21194 25290 21196
rect 25234 21142 25236 21194
rect 25236 21142 25288 21194
rect 25288 21142 25290 21194
rect 25234 21140 25290 21142
rect 25452 20300 25508 20356
rect 25340 20018 25396 20020
rect 25340 19966 25342 20018
rect 25342 19966 25394 20018
rect 25394 19966 25396 20018
rect 25340 19964 25396 19966
rect 25026 19626 25082 19628
rect 25026 19574 25028 19626
rect 25028 19574 25080 19626
rect 25080 19574 25082 19626
rect 25026 19572 25082 19574
rect 25130 19626 25186 19628
rect 25130 19574 25132 19626
rect 25132 19574 25184 19626
rect 25184 19574 25186 19626
rect 25130 19572 25186 19574
rect 25234 19626 25290 19628
rect 25234 19574 25236 19626
rect 25236 19574 25288 19626
rect 25288 19574 25290 19626
rect 25234 19572 25290 19574
rect 25452 19180 25508 19236
rect 25228 18450 25284 18452
rect 25228 18398 25230 18450
rect 25230 18398 25282 18450
rect 25282 18398 25284 18450
rect 25228 18396 25284 18398
rect 25788 21308 25844 21364
rect 25788 20690 25844 20692
rect 25788 20638 25790 20690
rect 25790 20638 25842 20690
rect 25842 20638 25844 20690
rect 25788 20636 25844 20638
rect 26236 24332 26292 24388
rect 26684 27132 26740 27188
rect 26572 24220 26628 24276
rect 27356 31666 27412 31668
rect 27356 31614 27358 31666
rect 27358 31614 27410 31666
rect 27410 31614 27412 31666
rect 27356 31612 27412 31614
rect 27132 30044 27188 30100
rect 27356 28700 27412 28756
rect 27020 27634 27076 27636
rect 27020 27582 27022 27634
rect 27022 27582 27074 27634
rect 27074 27582 27076 27634
rect 27020 27580 27076 27582
rect 28140 37826 28196 37828
rect 28140 37774 28142 37826
rect 28142 37774 28194 37826
rect 28194 37774 28196 37826
rect 28140 37772 28196 37774
rect 27580 30882 27636 30884
rect 27580 30830 27582 30882
rect 27582 30830 27634 30882
rect 27634 30830 27636 30882
rect 27580 30828 27636 30830
rect 28028 34748 28084 34804
rect 27916 32450 27972 32452
rect 27916 32398 27918 32450
rect 27918 32398 27970 32450
rect 27970 32398 27972 32450
rect 27916 32396 27972 32398
rect 28428 37658 28484 37660
rect 28428 37606 28430 37658
rect 28430 37606 28482 37658
rect 28482 37606 28484 37658
rect 28428 37604 28484 37606
rect 28532 37658 28588 37660
rect 28532 37606 28534 37658
rect 28534 37606 28586 37658
rect 28586 37606 28588 37658
rect 28532 37604 28588 37606
rect 28636 37658 28692 37660
rect 28636 37606 28638 37658
rect 28638 37606 28690 37658
rect 28690 37606 28692 37658
rect 28636 37604 28692 37606
rect 28428 36090 28484 36092
rect 28428 36038 28430 36090
rect 28430 36038 28482 36090
rect 28482 36038 28484 36090
rect 28428 36036 28484 36038
rect 28532 36090 28588 36092
rect 28532 36038 28534 36090
rect 28534 36038 28586 36090
rect 28586 36038 28588 36090
rect 28532 36036 28588 36038
rect 28636 36090 28692 36092
rect 28636 36038 28638 36090
rect 28638 36038 28690 36090
rect 28690 36038 28692 36090
rect 28636 36036 28692 36038
rect 28140 34412 28196 34468
rect 28428 34522 28484 34524
rect 28428 34470 28430 34522
rect 28430 34470 28482 34522
rect 28482 34470 28484 34522
rect 28428 34468 28484 34470
rect 28532 34522 28588 34524
rect 28532 34470 28534 34522
rect 28534 34470 28586 34522
rect 28586 34470 28588 34522
rect 28532 34468 28588 34470
rect 28636 34522 28692 34524
rect 28636 34470 28638 34522
rect 28638 34470 28690 34522
rect 28690 34470 28692 34522
rect 28636 34468 28692 34470
rect 28428 32954 28484 32956
rect 28428 32902 28430 32954
rect 28430 32902 28482 32954
rect 28482 32902 28484 32954
rect 28428 32900 28484 32902
rect 28532 32954 28588 32956
rect 28532 32902 28534 32954
rect 28534 32902 28586 32954
rect 28586 32902 28588 32954
rect 28532 32900 28588 32902
rect 28636 32954 28692 32956
rect 28636 32902 28638 32954
rect 28638 32902 28690 32954
rect 28690 32902 28692 32954
rect 28636 32900 28692 32902
rect 28428 31386 28484 31388
rect 28428 31334 28430 31386
rect 28430 31334 28482 31386
rect 28482 31334 28484 31386
rect 28428 31332 28484 31334
rect 28532 31386 28588 31388
rect 28532 31334 28534 31386
rect 28534 31334 28586 31386
rect 28586 31334 28588 31386
rect 28532 31332 28588 31334
rect 28636 31386 28692 31388
rect 28636 31334 28638 31386
rect 28638 31334 28690 31386
rect 28690 31334 28692 31386
rect 28636 31332 28692 31334
rect 27916 30098 27972 30100
rect 27916 30046 27918 30098
rect 27918 30046 27970 30098
rect 27970 30046 27972 30098
rect 27916 30044 27972 30046
rect 28428 29818 28484 29820
rect 28428 29766 28430 29818
rect 28430 29766 28482 29818
rect 28482 29766 28484 29818
rect 28428 29764 28484 29766
rect 28532 29818 28588 29820
rect 28532 29766 28534 29818
rect 28534 29766 28586 29818
rect 28586 29766 28588 29818
rect 28532 29764 28588 29766
rect 28636 29818 28692 29820
rect 28636 29766 28638 29818
rect 28638 29766 28690 29818
rect 28690 29766 28692 29818
rect 28636 29764 28692 29766
rect 27804 28140 27860 28196
rect 27804 27970 27860 27972
rect 27804 27918 27806 27970
rect 27806 27918 27858 27970
rect 27858 27918 27860 27970
rect 27804 27916 27860 27918
rect 27020 27244 27076 27300
rect 27356 27186 27412 27188
rect 27356 27134 27358 27186
rect 27358 27134 27410 27186
rect 27410 27134 27412 27186
rect 27356 27132 27412 27134
rect 27244 27020 27300 27076
rect 27020 25394 27076 25396
rect 27020 25342 27022 25394
rect 27022 25342 27074 25394
rect 27074 25342 27076 25394
rect 27020 25340 27076 25342
rect 26236 23996 26292 24052
rect 26348 23938 26404 23940
rect 26348 23886 26350 23938
rect 26350 23886 26402 23938
rect 26402 23886 26404 23938
rect 26348 23884 26404 23886
rect 26236 21644 26292 21700
rect 26348 21026 26404 21028
rect 26348 20974 26350 21026
rect 26350 20974 26402 21026
rect 26402 20974 26404 21026
rect 26348 20972 26404 20974
rect 26124 20636 26180 20692
rect 25026 18058 25082 18060
rect 25026 18006 25028 18058
rect 25028 18006 25080 18058
rect 25080 18006 25082 18058
rect 25026 18004 25082 18006
rect 25130 18058 25186 18060
rect 25130 18006 25132 18058
rect 25132 18006 25184 18058
rect 25184 18006 25186 18058
rect 25130 18004 25186 18006
rect 25234 18058 25290 18060
rect 25234 18006 25236 18058
rect 25236 18006 25288 18058
rect 25288 18006 25290 18058
rect 25234 18004 25290 18006
rect 25228 17388 25284 17444
rect 25026 16490 25082 16492
rect 25026 16438 25028 16490
rect 25028 16438 25080 16490
rect 25080 16438 25082 16490
rect 25026 16436 25082 16438
rect 25130 16490 25186 16492
rect 25130 16438 25132 16490
rect 25132 16438 25184 16490
rect 25184 16438 25186 16490
rect 25130 16436 25186 16438
rect 25234 16490 25290 16492
rect 25234 16438 25236 16490
rect 25236 16438 25288 16490
rect 25288 16438 25290 16490
rect 25234 16436 25290 16438
rect 25026 14922 25082 14924
rect 25026 14870 25028 14922
rect 25028 14870 25080 14922
rect 25080 14870 25082 14922
rect 25026 14868 25082 14870
rect 25130 14922 25186 14924
rect 25130 14870 25132 14922
rect 25132 14870 25184 14922
rect 25184 14870 25186 14922
rect 25130 14868 25186 14870
rect 25234 14922 25290 14924
rect 25234 14870 25236 14922
rect 25236 14870 25288 14922
rect 25288 14870 25290 14922
rect 25234 14868 25290 14870
rect 25676 18450 25732 18452
rect 25676 18398 25678 18450
rect 25678 18398 25730 18450
rect 25730 18398 25732 18450
rect 25676 18396 25732 18398
rect 25900 17612 25956 17668
rect 26572 23826 26628 23828
rect 26572 23774 26574 23826
rect 26574 23774 26626 23826
rect 26626 23774 26628 23826
rect 26572 23772 26628 23774
rect 26796 23548 26852 23604
rect 26684 23100 26740 23156
rect 26796 23324 26852 23380
rect 26572 20076 26628 20132
rect 26348 18956 26404 19012
rect 26124 18732 26180 18788
rect 26348 18674 26404 18676
rect 26348 18622 26350 18674
rect 26350 18622 26402 18674
rect 26402 18622 26404 18674
rect 26348 18620 26404 18622
rect 26236 18450 26292 18452
rect 26236 18398 26238 18450
rect 26238 18398 26290 18450
rect 26290 18398 26292 18450
rect 26236 18396 26292 18398
rect 26012 17164 26068 17220
rect 26348 16994 26404 16996
rect 26348 16942 26350 16994
rect 26350 16942 26402 16994
rect 26402 16942 26404 16994
rect 26348 16940 26404 16942
rect 26572 16828 26628 16884
rect 26348 15260 26404 15316
rect 25676 14700 25732 14756
rect 25788 13634 25844 13636
rect 25788 13582 25790 13634
rect 25790 13582 25842 13634
rect 25842 13582 25844 13634
rect 25788 13580 25844 13582
rect 25026 13354 25082 13356
rect 25026 13302 25028 13354
rect 25028 13302 25080 13354
rect 25080 13302 25082 13354
rect 25026 13300 25082 13302
rect 25130 13354 25186 13356
rect 25130 13302 25132 13354
rect 25132 13302 25184 13354
rect 25184 13302 25186 13354
rect 25130 13300 25186 13302
rect 25234 13354 25290 13356
rect 25234 13302 25236 13354
rect 25236 13302 25288 13354
rect 25288 13302 25290 13354
rect 25234 13300 25290 13302
rect 26236 13244 26292 13300
rect 27356 26514 27412 26516
rect 27356 26462 27358 26514
rect 27358 26462 27410 26514
rect 27410 26462 27412 26514
rect 27356 26460 27412 26462
rect 28428 28250 28484 28252
rect 28428 28198 28430 28250
rect 28430 28198 28482 28250
rect 28482 28198 28484 28250
rect 28428 28196 28484 28198
rect 28532 28250 28588 28252
rect 28532 28198 28534 28250
rect 28534 28198 28586 28250
rect 28586 28198 28588 28250
rect 28532 28196 28588 28198
rect 28636 28250 28692 28252
rect 28636 28198 28638 28250
rect 28638 28198 28690 28250
rect 28690 28198 28692 28250
rect 28636 28196 28692 28198
rect 28428 26682 28484 26684
rect 28428 26630 28430 26682
rect 28430 26630 28482 26682
rect 28482 26630 28484 26682
rect 28428 26628 28484 26630
rect 28532 26682 28588 26684
rect 28532 26630 28534 26682
rect 28534 26630 28586 26682
rect 28586 26630 28588 26682
rect 28532 26628 28588 26630
rect 28636 26682 28692 26684
rect 28636 26630 28638 26682
rect 28638 26630 28690 26682
rect 28690 26630 28692 26682
rect 28636 26628 28692 26630
rect 28140 26460 28196 26516
rect 27244 24444 27300 24500
rect 27356 24668 27412 24724
rect 27356 23154 27412 23156
rect 27356 23102 27358 23154
rect 27358 23102 27410 23154
rect 27410 23102 27412 23154
rect 27356 23100 27412 23102
rect 27020 22204 27076 22260
rect 26908 21308 26964 21364
rect 27132 21026 27188 21028
rect 27132 20974 27134 21026
rect 27134 20974 27186 21026
rect 27186 20974 27188 21026
rect 27132 20972 27188 20974
rect 27132 20802 27188 20804
rect 27132 20750 27134 20802
rect 27134 20750 27186 20802
rect 27186 20750 27188 20802
rect 27132 20748 27188 20750
rect 27020 20076 27076 20132
rect 27468 20636 27524 20692
rect 26796 15484 26852 15540
rect 27020 18732 27076 18788
rect 28428 25114 28484 25116
rect 28428 25062 28430 25114
rect 28430 25062 28482 25114
rect 28482 25062 28484 25114
rect 28428 25060 28484 25062
rect 28532 25114 28588 25116
rect 28532 25062 28534 25114
rect 28534 25062 28586 25114
rect 28586 25062 28588 25114
rect 28532 25060 28588 25062
rect 28636 25114 28692 25116
rect 28636 25062 28638 25114
rect 28638 25062 28690 25114
rect 28690 25062 28692 25114
rect 28636 25060 28692 25062
rect 27692 23660 27748 23716
rect 28428 23546 28484 23548
rect 28428 23494 28430 23546
rect 28430 23494 28482 23546
rect 28482 23494 28484 23546
rect 28428 23492 28484 23494
rect 28532 23546 28588 23548
rect 28532 23494 28534 23546
rect 28534 23494 28586 23546
rect 28586 23494 28588 23546
rect 28532 23492 28588 23494
rect 28636 23546 28692 23548
rect 28636 23494 28638 23546
rect 28638 23494 28690 23546
rect 28690 23494 28692 23546
rect 28636 23492 28692 23494
rect 28028 22988 28084 23044
rect 27804 18732 27860 18788
rect 27916 20300 27972 20356
rect 27580 18508 27636 18564
rect 28428 21978 28484 21980
rect 28428 21926 28430 21978
rect 28430 21926 28482 21978
rect 28482 21926 28484 21978
rect 28428 21924 28484 21926
rect 28532 21978 28588 21980
rect 28532 21926 28534 21978
rect 28534 21926 28586 21978
rect 28586 21926 28588 21978
rect 28532 21924 28588 21926
rect 28636 21978 28692 21980
rect 28636 21926 28638 21978
rect 28638 21926 28690 21978
rect 28690 21926 28692 21978
rect 28636 21924 28692 21926
rect 28028 19964 28084 20020
rect 28140 20748 28196 20804
rect 28428 20410 28484 20412
rect 28428 20358 28430 20410
rect 28430 20358 28482 20410
rect 28482 20358 28484 20410
rect 28428 20356 28484 20358
rect 28532 20410 28588 20412
rect 28532 20358 28534 20410
rect 28534 20358 28586 20410
rect 28586 20358 28588 20410
rect 28532 20356 28588 20358
rect 28636 20410 28692 20412
rect 28636 20358 28638 20410
rect 28638 20358 28690 20410
rect 28690 20358 28692 20410
rect 28636 20356 28692 20358
rect 27020 17164 27076 17220
rect 27580 16882 27636 16884
rect 27580 16830 27582 16882
rect 27582 16830 27634 16882
rect 27634 16830 27636 16882
rect 27580 16828 27636 16830
rect 26460 13580 26516 13636
rect 26460 13186 26516 13188
rect 26460 13134 26462 13186
rect 26462 13134 26514 13186
rect 26514 13134 26516 13186
rect 26460 13132 26516 13134
rect 26124 12908 26180 12964
rect 25228 12178 25284 12180
rect 25228 12126 25230 12178
rect 25230 12126 25282 12178
rect 25282 12126 25284 12178
rect 25228 12124 25284 12126
rect 28028 17442 28084 17444
rect 28028 17390 28030 17442
rect 28030 17390 28082 17442
rect 28082 17390 28084 17442
rect 28028 17388 28084 17390
rect 28428 18842 28484 18844
rect 28428 18790 28430 18842
rect 28430 18790 28482 18842
rect 28482 18790 28484 18842
rect 28428 18788 28484 18790
rect 28532 18842 28588 18844
rect 28532 18790 28534 18842
rect 28534 18790 28586 18842
rect 28586 18790 28588 18842
rect 28532 18788 28588 18790
rect 28636 18842 28692 18844
rect 28636 18790 28638 18842
rect 28638 18790 28690 18842
rect 28690 18790 28692 18842
rect 28636 18788 28692 18790
rect 28428 17274 28484 17276
rect 28428 17222 28430 17274
rect 28430 17222 28482 17274
rect 28482 17222 28484 17274
rect 28428 17220 28484 17222
rect 28532 17274 28588 17276
rect 28532 17222 28534 17274
rect 28534 17222 28586 17274
rect 28586 17222 28588 17274
rect 28532 17220 28588 17222
rect 28636 17274 28692 17276
rect 28636 17222 28638 17274
rect 28638 17222 28690 17274
rect 28690 17222 28692 17274
rect 28636 17220 28692 17222
rect 28428 15706 28484 15708
rect 28428 15654 28430 15706
rect 28430 15654 28482 15706
rect 28482 15654 28484 15706
rect 28428 15652 28484 15654
rect 28532 15706 28588 15708
rect 28532 15654 28534 15706
rect 28534 15654 28586 15706
rect 28586 15654 28588 15706
rect 28532 15652 28588 15654
rect 28636 15706 28692 15708
rect 28636 15654 28638 15706
rect 28638 15654 28690 15706
rect 28690 15654 28692 15706
rect 28636 15652 28692 15654
rect 28428 14138 28484 14140
rect 28428 14086 28430 14138
rect 28430 14086 28482 14138
rect 28482 14086 28484 14138
rect 28428 14084 28484 14086
rect 28532 14138 28588 14140
rect 28532 14086 28534 14138
rect 28534 14086 28586 14138
rect 28586 14086 28588 14138
rect 28532 14084 28588 14086
rect 28636 14138 28692 14140
rect 28636 14086 28638 14138
rect 28638 14086 28690 14138
rect 28690 14086 28692 14138
rect 28636 14084 28692 14086
rect 27132 13804 27188 13860
rect 26572 12962 26628 12964
rect 26572 12910 26574 12962
rect 26574 12910 26626 12962
rect 26626 12910 26628 12962
rect 26572 12908 26628 12910
rect 26460 12124 26516 12180
rect 28428 12570 28484 12572
rect 28428 12518 28430 12570
rect 28430 12518 28482 12570
rect 28482 12518 28484 12570
rect 28428 12516 28484 12518
rect 28532 12570 28588 12572
rect 28532 12518 28534 12570
rect 28534 12518 28586 12570
rect 28586 12518 28588 12570
rect 28532 12516 28588 12518
rect 28636 12570 28692 12572
rect 28636 12518 28638 12570
rect 28638 12518 28690 12570
rect 28690 12518 28692 12570
rect 28636 12516 28692 12518
rect 25026 11786 25082 11788
rect 25026 11734 25028 11786
rect 25028 11734 25080 11786
rect 25080 11734 25082 11786
rect 25026 11732 25082 11734
rect 25130 11786 25186 11788
rect 25130 11734 25132 11786
rect 25132 11734 25184 11786
rect 25184 11734 25186 11786
rect 25130 11732 25186 11734
rect 25234 11786 25290 11788
rect 25234 11734 25236 11786
rect 25236 11734 25288 11786
rect 25288 11734 25290 11786
rect 25234 11732 25290 11734
rect 28428 11002 28484 11004
rect 28428 10950 28430 11002
rect 28430 10950 28482 11002
rect 28482 10950 28484 11002
rect 28428 10948 28484 10950
rect 28532 11002 28588 11004
rect 28532 10950 28534 11002
rect 28534 10950 28586 11002
rect 28586 10950 28588 11002
rect 28532 10948 28588 10950
rect 28636 11002 28692 11004
rect 28636 10950 28638 11002
rect 28638 10950 28690 11002
rect 28690 10950 28692 11002
rect 28636 10948 28692 10950
rect 25788 10780 25844 10836
rect 25026 10218 25082 10220
rect 25026 10166 25028 10218
rect 25028 10166 25080 10218
rect 25080 10166 25082 10218
rect 25026 10164 25082 10166
rect 25130 10218 25186 10220
rect 25130 10166 25132 10218
rect 25132 10166 25184 10218
rect 25184 10166 25186 10218
rect 25130 10164 25186 10166
rect 25234 10218 25290 10220
rect 25234 10166 25236 10218
rect 25236 10166 25288 10218
rect 25288 10166 25290 10218
rect 25234 10164 25290 10166
rect 24892 9826 24948 9828
rect 24892 9774 24894 9826
rect 24894 9774 24946 9826
rect 24946 9774 24948 9826
rect 24892 9772 24948 9774
rect 24444 6690 24500 6692
rect 24444 6638 24446 6690
rect 24446 6638 24498 6690
rect 24498 6638 24500 6690
rect 24444 6636 24500 6638
rect 22540 6018 22596 6020
rect 22540 5966 22542 6018
rect 22542 5966 22594 6018
rect 22594 5966 22596 6018
rect 22540 5964 22596 5966
rect 22428 5740 22484 5796
rect 21532 5122 21588 5124
rect 21532 5070 21534 5122
rect 21534 5070 21586 5122
rect 21586 5070 21588 5122
rect 21532 5068 21588 5070
rect 21980 4956 22036 5012
rect 20972 3388 21028 3444
rect 20748 2156 20804 2212
rect 21624 4730 21680 4732
rect 21624 4678 21626 4730
rect 21626 4678 21678 4730
rect 21678 4678 21680 4730
rect 21624 4676 21680 4678
rect 21728 4730 21784 4732
rect 21728 4678 21730 4730
rect 21730 4678 21782 4730
rect 21782 4678 21784 4730
rect 21728 4676 21784 4678
rect 21832 4730 21888 4732
rect 21832 4678 21834 4730
rect 21834 4678 21886 4730
rect 21886 4678 21888 4730
rect 21832 4676 21888 4678
rect 21420 3276 21476 3332
rect 22540 5234 22596 5236
rect 22540 5182 22542 5234
rect 22542 5182 22594 5234
rect 22594 5182 22596 5234
rect 22540 5180 22596 5182
rect 23436 5964 23492 6020
rect 23660 5906 23716 5908
rect 23660 5854 23662 5906
rect 23662 5854 23714 5906
rect 23714 5854 23716 5906
rect 23660 5852 23716 5854
rect 23884 5628 23940 5684
rect 24444 6076 24500 6132
rect 24780 7420 24836 7476
rect 24556 5964 24612 6020
rect 24556 5740 24612 5796
rect 26348 10498 26404 10500
rect 26348 10446 26350 10498
rect 26350 10446 26402 10498
rect 26402 10446 26404 10498
rect 26348 10444 26404 10446
rect 25564 9826 25620 9828
rect 25564 9774 25566 9826
rect 25566 9774 25618 9826
rect 25618 9774 25620 9826
rect 25564 9772 25620 9774
rect 26012 9826 26068 9828
rect 26012 9774 26014 9826
rect 26014 9774 26066 9826
rect 26066 9774 26068 9826
rect 26012 9772 26068 9774
rect 28428 9434 28484 9436
rect 28428 9382 28430 9434
rect 28430 9382 28482 9434
rect 28482 9382 28484 9434
rect 28428 9380 28484 9382
rect 28532 9434 28588 9436
rect 28532 9382 28534 9434
rect 28534 9382 28586 9434
rect 28586 9382 28588 9434
rect 28532 9380 28588 9382
rect 28636 9434 28692 9436
rect 28636 9382 28638 9434
rect 28638 9382 28690 9434
rect 28690 9382 28692 9434
rect 28636 9380 28692 9382
rect 25026 8650 25082 8652
rect 25026 8598 25028 8650
rect 25028 8598 25080 8650
rect 25080 8598 25082 8650
rect 25026 8596 25082 8598
rect 25130 8650 25186 8652
rect 25130 8598 25132 8650
rect 25132 8598 25184 8650
rect 25184 8598 25186 8650
rect 25130 8596 25186 8598
rect 25234 8650 25290 8652
rect 25234 8598 25236 8650
rect 25236 8598 25288 8650
rect 25288 8598 25290 8650
rect 25234 8596 25290 8598
rect 28428 7866 28484 7868
rect 28428 7814 28430 7866
rect 28430 7814 28482 7866
rect 28482 7814 28484 7866
rect 28428 7812 28484 7814
rect 28532 7866 28588 7868
rect 28532 7814 28534 7866
rect 28534 7814 28586 7866
rect 28586 7814 28588 7866
rect 28532 7812 28588 7814
rect 28636 7866 28692 7868
rect 28636 7814 28638 7866
rect 28638 7814 28690 7866
rect 28690 7814 28692 7866
rect 28636 7812 28692 7814
rect 25026 7082 25082 7084
rect 25026 7030 25028 7082
rect 25028 7030 25080 7082
rect 25080 7030 25082 7082
rect 25026 7028 25082 7030
rect 25130 7082 25186 7084
rect 25130 7030 25132 7082
rect 25132 7030 25184 7082
rect 25184 7030 25186 7082
rect 25130 7028 25186 7030
rect 25234 7082 25290 7084
rect 25234 7030 25236 7082
rect 25236 7030 25288 7082
rect 25288 7030 25290 7082
rect 25234 7028 25290 7030
rect 28428 6298 28484 6300
rect 28428 6246 28430 6298
rect 28430 6246 28482 6298
rect 28482 6246 28484 6298
rect 28428 6244 28484 6246
rect 28532 6298 28588 6300
rect 28532 6246 28534 6298
rect 28534 6246 28586 6298
rect 28586 6246 28588 6298
rect 28532 6244 28588 6246
rect 28636 6298 28692 6300
rect 28636 6246 28638 6298
rect 28638 6246 28690 6298
rect 28690 6246 28692 6298
rect 28636 6244 28692 6246
rect 24780 5964 24836 6020
rect 23212 4396 23268 4452
rect 23996 4844 24052 4900
rect 23212 4226 23268 4228
rect 23212 4174 23214 4226
rect 23214 4174 23266 4226
rect 23266 4174 23268 4226
rect 23212 4172 23268 4174
rect 22316 3724 22372 3780
rect 21980 3666 22036 3668
rect 21980 3614 21982 3666
rect 21982 3614 22034 3666
rect 22034 3614 22036 3666
rect 21980 3612 22036 3614
rect 22764 3724 22820 3780
rect 21624 3162 21680 3164
rect 21624 3110 21626 3162
rect 21626 3110 21678 3162
rect 21678 3110 21680 3162
rect 21624 3108 21680 3110
rect 21728 3162 21784 3164
rect 21728 3110 21730 3162
rect 21730 3110 21782 3162
rect 21782 3110 21784 3162
rect 21728 3108 21784 3110
rect 21832 3162 21888 3164
rect 21832 3110 21834 3162
rect 21834 3110 21886 3162
rect 21886 3110 21888 3162
rect 21832 3108 21888 3110
rect 22652 2940 22708 2996
rect 21420 2156 21476 2212
rect 22428 2604 22484 2660
rect 21532 1932 21588 1988
rect 22428 1986 22484 1988
rect 22428 1934 22430 1986
rect 22430 1934 22482 1986
rect 22482 1934 22484 1986
rect 22428 1932 22484 1934
rect 21624 1594 21680 1596
rect 21624 1542 21626 1594
rect 21626 1542 21678 1594
rect 21678 1542 21680 1594
rect 21624 1540 21680 1542
rect 21728 1594 21784 1596
rect 21728 1542 21730 1594
rect 21730 1542 21782 1594
rect 21782 1542 21784 1594
rect 21728 1540 21784 1542
rect 21832 1594 21888 1596
rect 21832 1542 21834 1594
rect 21834 1542 21886 1594
rect 21886 1542 21888 1594
rect 21832 1540 21888 1542
rect 23212 3612 23268 3668
rect 22876 2716 22932 2772
rect 23324 3442 23380 3444
rect 23324 3390 23326 3442
rect 23326 3390 23378 3442
rect 23378 3390 23380 3442
rect 23324 3388 23380 3390
rect 23660 4060 23716 4116
rect 23660 3836 23716 3892
rect 24220 4338 24276 4340
rect 24220 4286 24222 4338
rect 24222 4286 24274 4338
rect 24274 4286 24276 4338
rect 24220 4284 24276 4286
rect 23996 3948 24052 4004
rect 23436 2940 23492 2996
rect 23772 3276 23828 3332
rect 23660 2828 23716 2884
rect 22428 476 22484 532
rect 23212 476 23268 532
rect 23548 1932 23604 1988
rect 24108 3554 24164 3556
rect 24108 3502 24110 3554
rect 24110 3502 24162 3554
rect 24162 3502 24164 3554
rect 24108 3500 24164 3502
rect 24108 2770 24164 2772
rect 24108 2718 24110 2770
rect 24110 2718 24162 2770
rect 24162 2718 24164 2770
rect 24108 2716 24164 2718
rect 24668 2828 24724 2884
rect 24220 2044 24276 2100
rect 25452 6130 25508 6132
rect 25452 6078 25454 6130
rect 25454 6078 25506 6130
rect 25506 6078 25508 6130
rect 25452 6076 25508 6078
rect 25026 5514 25082 5516
rect 25026 5462 25028 5514
rect 25028 5462 25080 5514
rect 25080 5462 25082 5514
rect 25026 5460 25082 5462
rect 25130 5514 25186 5516
rect 25130 5462 25132 5514
rect 25132 5462 25184 5514
rect 25184 5462 25186 5514
rect 25130 5460 25186 5462
rect 25234 5514 25290 5516
rect 25234 5462 25236 5514
rect 25236 5462 25288 5514
rect 25288 5462 25290 5514
rect 25234 5460 25290 5462
rect 26012 6018 26068 6020
rect 26012 5966 26014 6018
rect 26014 5966 26066 6018
rect 26066 5966 26068 6018
rect 26012 5964 26068 5966
rect 25900 5906 25956 5908
rect 25900 5854 25902 5906
rect 25902 5854 25954 5906
rect 25954 5854 25956 5906
rect 25900 5852 25956 5854
rect 25564 5794 25620 5796
rect 25564 5742 25566 5794
rect 25566 5742 25618 5794
rect 25618 5742 25620 5794
rect 25564 5740 25620 5742
rect 25228 4450 25284 4452
rect 25228 4398 25230 4450
rect 25230 4398 25282 4450
rect 25282 4398 25284 4450
rect 25228 4396 25284 4398
rect 25340 4338 25396 4340
rect 25340 4286 25342 4338
rect 25342 4286 25394 4338
rect 25394 4286 25396 4338
rect 25340 4284 25396 4286
rect 24892 4172 24948 4228
rect 25026 3946 25082 3948
rect 25026 3894 25028 3946
rect 25028 3894 25080 3946
rect 25080 3894 25082 3946
rect 25026 3892 25082 3894
rect 25130 3946 25186 3948
rect 25130 3894 25132 3946
rect 25132 3894 25184 3946
rect 25184 3894 25186 3946
rect 25130 3892 25186 3894
rect 25234 3946 25290 3948
rect 25234 3894 25236 3946
rect 25236 3894 25288 3946
rect 25288 3894 25290 3946
rect 25234 3892 25290 3894
rect 24892 3724 24948 3780
rect 25676 5292 25732 5348
rect 26012 4898 26068 4900
rect 26012 4846 26014 4898
rect 26014 4846 26066 4898
rect 26066 4846 26068 4898
rect 26012 4844 26068 4846
rect 25340 2994 25396 2996
rect 25340 2942 25342 2994
rect 25342 2942 25394 2994
rect 25394 2942 25396 2994
rect 25340 2940 25396 2942
rect 25676 2940 25732 2996
rect 25452 2882 25508 2884
rect 25452 2830 25454 2882
rect 25454 2830 25506 2882
rect 25506 2830 25508 2882
rect 25452 2828 25508 2830
rect 25788 3500 25844 3556
rect 26908 4226 26964 4228
rect 26908 4174 26910 4226
rect 26910 4174 26962 4226
rect 26962 4174 26964 4226
rect 26908 4172 26964 4174
rect 26460 4060 26516 4116
rect 25900 2716 25956 2772
rect 25026 2378 25082 2380
rect 25026 2326 25028 2378
rect 25028 2326 25080 2378
rect 25080 2326 25082 2378
rect 25026 2324 25082 2326
rect 25130 2378 25186 2380
rect 25130 2326 25132 2378
rect 25132 2326 25184 2378
rect 25184 2326 25186 2378
rect 25130 2324 25186 2326
rect 25234 2378 25290 2380
rect 25234 2326 25236 2378
rect 25236 2326 25288 2378
rect 25288 2326 25290 2378
rect 25234 2324 25290 2326
rect 24332 1820 24388 1876
rect 24892 1708 24948 1764
rect 26124 3388 26180 3444
rect 27132 3442 27188 3444
rect 27132 3390 27134 3442
rect 27134 3390 27186 3442
rect 27186 3390 27188 3442
rect 27132 3388 27188 3390
rect 26236 2940 26292 2996
rect 26684 2716 26740 2772
rect 25676 1932 25732 1988
rect 27580 3500 27636 3556
rect 27356 2882 27412 2884
rect 27356 2830 27358 2882
rect 27358 2830 27410 2882
rect 27410 2830 27412 2882
rect 27356 2828 27412 2830
rect 27356 1874 27412 1876
rect 27356 1822 27358 1874
rect 27358 1822 27410 1874
rect 27410 1822 27412 1874
rect 27356 1820 27412 1822
rect 26908 1708 26964 1764
rect 28428 4730 28484 4732
rect 28428 4678 28430 4730
rect 28430 4678 28482 4730
rect 28482 4678 28484 4730
rect 28428 4676 28484 4678
rect 28532 4730 28588 4732
rect 28532 4678 28534 4730
rect 28534 4678 28586 4730
rect 28586 4678 28588 4730
rect 28532 4676 28588 4678
rect 28636 4730 28692 4732
rect 28636 4678 28638 4730
rect 28638 4678 28690 4730
rect 28690 4678 28692 4730
rect 28636 4676 28692 4678
rect 27916 3666 27972 3668
rect 27916 3614 27918 3666
rect 27918 3614 27970 3666
rect 27970 3614 27972 3666
rect 27916 3612 27972 3614
rect 28428 3162 28484 3164
rect 28428 3110 28430 3162
rect 28430 3110 28482 3162
rect 28482 3110 28484 3162
rect 28428 3108 28484 3110
rect 28532 3162 28588 3164
rect 28532 3110 28534 3162
rect 28534 3110 28586 3162
rect 28586 3110 28588 3162
rect 28532 3108 28588 3110
rect 28636 3162 28692 3164
rect 28636 3110 28638 3162
rect 28638 3110 28690 3162
rect 28690 3110 28692 3162
rect 28636 3108 28692 3110
rect 28140 2658 28196 2660
rect 28140 2606 28142 2658
rect 28142 2606 28194 2658
rect 28194 2606 28196 2658
rect 28140 2604 28196 2606
rect 27580 2044 27636 2100
rect 28428 1594 28484 1596
rect 28428 1542 28430 1594
rect 28430 1542 28482 1594
rect 28482 1542 28484 1594
rect 28428 1540 28484 1542
rect 28532 1594 28588 1596
rect 28532 1542 28534 1594
rect 28534 1542 28586 1594
rect 28586 1542 28588 1594
rect 28532 1540 28588 1542
rect 28636 1594 28692 1596
rect 28636 1542 28638 1594
rect 28638 1542 28690 1594
rect 28690 1542 28692 1594
rect 28636 1540 28692 1542
<< metal3 >>
rect 4604 118356 4614 118412
rect 4670 118356 4718 118412
rect 4774 118356 4822 118412
rect 4878 118356 4888 118412
rect 11408 118356 11418 118412
rect 11474 118356 11522 118412
rect 11578 118356 11626 118412
rect 11682 118356 11692 118412
rect 18212 118356 18222 118412
rect 18278 118356 18326 118412
rect 18382 118356 18430 118412
rect 18486 118356 18496 118412
rect 25016 118356 25026 118412
rect 25082 118356 25130 118412
rect 25186 118356 25234 118412
rect 25290 118356 25300 118412
rect 8006 117572 8016 117628
rect 8072 117572 8120 117628
rect 8176 117572 8224 117628
rect 8280 117572 8290 117628
rect 14810 117572 14820 117628
rect 14876 117572 14924 117628
rect 14980 117572 15028 117628
rect 15084 117572 15094 117628
rect 21614 117572 21624 117628
rect 21680 117572 21728 117628
rect 21784 117572 21832 117628
rect 21888 117572 21898 117628
rect 28418 117572 28428 117628
rect 28484 117572 28532 117628
rect 28588 117572 28636 117628
rect 28692 117572 28702 117628
rect 24658 117180 24668 117236
rect 24724 117180 25340 117236
rect 25396 117180 25406 117236
rect 4604 116788 4614 116844
rect 4670 116788 4718 116844
rect 4774 116788 4822 116844
rect 4878 116788 4888 116844
rect 11408 116788 11418 116844
rect 11474 116788 11522 116844
rect 11578 116788 11626 116844
rect 11682 116788 11692 116844
rect 18212 116788 18222 116844
rect 18278 116788 18326 116844
rect 18382 116788 18430 116844
rect 18486 116788 18496 116844
rect 25016 116788 25026 116844
rect 25082 116788 25130 116844
rect 25186 116788 25234 116844
rect 25290 116788 25300 116844
rect 16818 116508 16828 116564
rect 16884 116508 17780 116564
rect 17724 116452 17780 116508
rect 15138 116396 15148 116452
rect 15204 116396 16268 116452
rect 16324 116396 16334 116452
rect 16706 116396 16716 116452
rect 16772 116396 17388 116452
rect 17444 116396 17454 116452
rect 17714 116396 17724 116452
rect 17780 116396 18396 116452
rect 18452 116396 18462 116452
rect 8006 116004 8016 116060
rect 8072 116004 8120 116060
rect 8176 116004 8224 116060
rect 8280 116004 8290 116060
rect 14810 116004 14820 116060
rect 14876 116004 14924 116060
rect 14980 116004 15028 116060
rect 15084 116004 15094 116060
rect 21614 116004 21624 116060
rect 21680 116004 21728 116060
rect 21784 116004 21832 116060
rect 21888 116004 21898 116060
rect 28418 116004 28428 116060
rect 28484 116004 28532 116060
rect 28588 116004 28636 116060
rect 28692 116004 28702 116060
rect 10770 115612 10780 115668
rect 10836 115612 12236 115668
rect 12292 115612 13356 115668
rect 13412 115612 13916 115668
rect 13972 115612 13982 115668
rect 4604 115220 4614 115276
rect 4670 115220 4718 115276
rect 4774 115220 4822 115276
rect 4878 115220 4888 115276
rect 11408 115220 11418 115276
rect 11474 115220 11522 115276
rect 11578 115220 11626 115276
rect 11682 115220 11692 115276
rect 18212 115220 18222 115276
rect 18278 115220 18326 115276
rect 18382 115220 18430 115276
rect 18486 115220 18496 115276
rect 25016 115220 25026 115276
rect 25082 115220 25130 115276
rect 25186 115220 25234 115276
rect 25290 115220 25300 115276
rect 0 114996 400 115024
rect 0 114940 1708 114996
rect 1764 114940 1774 114996
rect 17266 114940 17276 114996
rect 17332 114940 18620 114996
rect 18676 114940 18686 114996
rect 0 114912 400 114940
rect 17490 114828 17500 114884
rect 17556 114828 18060 114884
rect 18116 114828 20076 114884
rect 20132 114828 20142 114884
rect 22642 114604 22652 114660
rect 22708 114604 24108 114660
rect 24164 114604 24780 114660
rect 24836 114604 24846 114660
rect 8006 114436 8016 114492
rect 8072 114436 8120 114492
rect 8176 114436 8224 114492
rect 8280 114436 8290 114492
rect 14810 114436 14820 114492
rect 14876 114436 14924 114492
rect 14980 114436 15028 114492
rect 15084 114436 15094 114492
rect 21614 114436 21624 114492
rect 21680 114436 21728 114492
rect 21784 114436 21832 114492
rect 21888 114436 21898 114492
rect 28418 114436 28428 114492
rect 28484 114436 28532 114492
rect 28588 114436 28636 114492
rect 28692 114436 28702 114492
rect 22866 114380 22876 114436
rect 22932 114380 24108 114436
rect 24164 114380 24174 114436
rect 20066 114268 20076 114324
rect 20132 114268 21420 114324
rect 21476 114268 21486 114324
rect 10098 114156 10108 114212
rect 10164 114156 11116 114212
rect 11172 114156 11182 114212
rect 10546 114044 10556 114100
rect 10612 114044 12124 114100
rect 12180 114044 12684 114100
rect 12740 114044 12750 114100
rect 4604 113652 4614 113708
rect 4670 113652 4718 113708
rect 4774 113652 4822 113708
rect 4878 113652 4888 113708
rect 11408 113652 11418 113708
rect 11474 113652 11522 113708
rect 11578 113652 11626 113708
rect 11682 113652 11692 113708
rect 18212 113652 18222 113708
rect 18278 113652 18326 113708
rect 18382 113652 18430 113708
rect 18486 113652 18496 113708
rect 25016 113652 25026 113708
rect 25082 113652 25130 113708
rect 25186 113652 25234 113708
rect 25290 113652 25300 113708
rect 18610 113260 18620 113316
rect 18676 113260 19180 113316
rect 19236 113260 20076 113316
rect 20132 113260 20142 113316
rect 24098 113260 24108 113316
rect 24164 113260 25900 113316
rect 25956 113260 25966 113316
rect 7970 113148 7980 113204
rect 8036 113148 9212 113204
rect 9268 113148 10556 113204
rect 10612 113148 10622 113204
rect 12114 113036 12124 113092
rect 12180 113036 12796 113092
rect 12852 113036 13356 113092
rect 13412 113036 13422 113092
rect 8006 112868 8016 112924
rect 8072 112868 8120 112924
rect 8176 112868 8224 112924
rect 8280 112868 8290 112924
rect 14810 112868 14820 112924
rect 14876 112868 14924 112924
rect 14980 112868 15028 112924
rect 15084 112868 15094 112924
rect 21614 112868 21624 112924
rect 21680 112868 21728 112924
rect 21784 112868 21832 112924
rect 21888 112868 21898 112924
rect 28418 112868 28428 112924
rect 28484 112868 28532 112924
rect 28588 112868 28636 112924
rect 28692 112868 28702 112924
rect 8418 112588 8428 112644
rect 8484 112588 8876 112644
rect 8932 112588 10332 112644
rect 10388 112588 11228 112644
rect 11284 112588 11294 112644
rect 11442 112476 11452 112532
rect 11508 112476 13020 112532
rect 13076 112476 13086 112532
rect 14690 112476 14700 112532
rect 14756 112476 15708 112532
rect 15764 112476 16604 112532
rect 16660 112476 17388 112532
rect 17444 112476 17454 112532
rect 19282 112476 19292 112532
rect 19348 112476 19964 112532
rect 20020 112476 20030 112532
rect 0 112308 400 112336
rect 0 112252 3948 112308
rect 4004 112252 4014 112308
rect 0 112224 400 112252
rect 4604 112084 4614 112140
rect 4670 112084 4718 112140
rect 4774 112084 4822 112140
rect 4878 112084 4888 112140
rect 11408 112084 11418 112140
rect 11474 112084 11522 112140
rect 11578 112084 11626 112140
rect 11682 112084 11692 112140
rect 18212 112084 18222 112140
rect 18278 112084 18326 112140
rect 18382 112084 18430 112140
rect 18486 112084 18496 112140
rect 25016 112084 25026 112140
rect 25082 112084 25130 112140
rect 25186 112084 25234 112140
rect 25290 112084 25300 112140
rect 28018 111916 28028 111972
rect 28084 111916 28252 111972
rect 28308 111916 28318 111972
rect 17378 111692 17388 111748
rect 17444 111692 18172 111748
rect 18228 111692 18956 111748
rect 19012 111692 19022 111748
rect 23426 111692 23436 111748
rect 23492 111692 24108 111748
rect 24164 111692 26684 111748
rect 26740 111692 26750 111748
rect 8006 111300 8016 111356
rect 8072 111300 8120 111356
rect 8176 111300 8224 111356
rect 8280 111300 8290 111356
rect 14810 111300 14820 111356
rect 14876 111300 14924 111356
rect 14980 111300 15028 111356
rect 15084 111300 15094 111356
rect 21614 111300 21624 111356
rect 21680 111300 21728 111356
rect 21784 111300 21832 111356
rect 21888 111300 21898 111356
rect 28418 111300 28428 111356
rect 28484 111300 28532 111356
rect 28588 111300 28636 111356
rect 28692 111300 28702 111356
rect 6850 110908 6860 110964
rect 6916 110908 9604 110964
rect 16706 110908 16716 110964
rect 16772 110908 17500 110964
rect 17556 110908 20076 110964
rect 20132 110908 21420 110964
rect 21476 110908 21486 110964
rect 9548 110740 9604 110908
rect 11778 110796 11788 110852
rect 11844 110796 12684 110852
rect 12740 110796 12750 110852
rect 9538 110684 9548 110740
rect 9604 110684 10220 110740
rect 10276 110684 11004 110740
rect 11060 110684 11676 110740
rect 11732 110684 14476 110740
rect 14532 110684 14542 110740
rect 4604 110516 4614 110572
rect 4670 110516 4718 110572
rect 4774 110516 4822 110572
rect 4878 110516 4888 110572
rect 11408 110516 11418 110572
rect 11474 110516 11522 110572
rect 11578 110516 11626 110572
rect 11682 110516 11692 110572
rect 18212 110516 18222 110572
rect 18278 110516 18326 110572
rect 18382 110516 18430 110572
rect 18486 110516 18496 110572
rect 25016 110516 25026 110572
rect 25082 110516 25130 110572
rect 25186 110516 25234 110572
rect 25290 110516 25300 110572
rect 11442 110236 11452 110292
rect 11508 110236 12460 110292
rect 12516 110236 12526 110292
rect 8978 110124 8988 110180
rect 9044 110124 9660 110180
rect 9716 110124 10332 110180
rect 10388 110124 10780 110180
rect 10836 110124 10846 110180
rect 11666 110124 11676 110180
rect 11732 110124 14252 110180
rect 14308 110124 14318 110180
rect 12786 110012 12796 110068
rect 12852 110012 13916 110068
rect 13972 110012 13982 110068
rect 8006 109732 8016 109788
rect 8072 109732 8120 109788
rect 8176 109732 8224 109788
rect 8280 109732 8290 109788
rect 14810 109732 14820 109788
rect 14876 109732 14924 109788
rect 14980 109732 15028 109788
rect 15084 109732 15094 109788
rect 21614 109732 21624 109788
rect 21680 109732 21728 109788
rect 21784 109732 21832 109788
rect 21888 109732 21898 109788
rect 28418 109732 28428 109788
rect 28484 109732 28532 109788
rect 28588 109732 28636 109788
rect 28692 109732 28702 109788
rect 0 109620 400 109648
rect 0 109564 1708 109620
rect 1764 109564 1774 109620
rect 0 109536 400 109564
rect 14018 109340 14028 109396
rect 14084 109340 15372 109396
rect 15428 109340 15820 109396
rect 15876 109340 16716 109396
rect 16772 109340 19516 109396
rect 19572 109340 20188 109396
rect 20132 109284 20188 109340
rect 12450 109228 12460 109284
rect 12516 109228 12908 109284
rect 12964 109228 13468 109284
rect 13524 109228 13534 109284
rect 15026 109228 15036 109284
rect 15092 109228 16156 109284
rect 16212 109228 18732 109284
rect 18788 109228 18798 109284
rect 20132 109228 20412 109284
rect 20468 109228 20478 109284
rect 4604 108948 4614 109004
rect 4670 108948 4718 109004
rect 4774 108948 4822 109004
rect 4878 108948 4888 109004
rect 11408 108948 11418 109004
rect 11474 108948 11522 109004
rect 11578 108948 11626 109004
rect 11682 108948 11692 109004
rect 18212 108948 18222 109004
rect 18278 108948 18326 109004
rect 18382 108948 18430 109004
rect 18486 108948 18496 109004
rect 25016 108948 25026 109004
rect 25082 108948 25130 109004
rect 25186 108948 25234 109004
rect 25290 108948 25300 109004
rect 16930 108780 16940 108836
rect 16996 108780 17948 108836
rect 18004 108780 18014 108836
rect 22306 108668 22316 108724
rect 22372 108668 23212 108724
rect 23268 108668 24892 108724
rect 24948 108668 25900 108724
rect 25956 108668 25966 108724
rect 12562 108556 12572 108612
rect 12628 108556 14924 108612
rect 14980 108556 14990 108612
rect 23090 108556 23100 108612
rect 23156 108556 25676 108612
rect 25732 108556 26684 108612
rect 26740 108556 26750 108612
rect 9202 108444 9212 108500
rect 9268 108444 13692 108500
rect 13748 108444 13758 108500
rect 16034 108444 16044 108500
rect 16100 108444 18172 108500
rect 18228 108444 18238 108500
rect 19170 108444 19180 108500
rect 19236 108444 21420 108500
rect 21476 108444 21486 108500
rect 16930 108332 16940 108388
rect 16996 108332 19068 108388
rect 19124 108332 19134 108388
rect 20178 108332 20188 108388
rect 20244 108332 20524 108388
rect 20580 108332 21868 108388
rect 21924 108332 22204 108388
rect 22260 108332 23996 108388
rect 24052 108332 24668 108388
rect 24724 108332 24734 108388
rect 27234 108332 27244 108388
rect 27300 108332 28252 108388
rect 28308 108332 28318 108388
rect 16594 108220 16604 108276
rect 16660 108220 18508 108276
rect 18564 108220 18574 108276
rect 8006 108164 8016 108220
rect 8072 108164 8120 108220
rect 8176 108164 8224 108220
rect 8280 108164 8290 108220
rect 14810 108164 14820 108220
rect 14876 108164 14924 108220
rect 14980 108164 15028 108220
rect 15084 108164 15094 108220
rect 16604 108052 16660 108220
rect 21614 108164 21624 108220
rect 21680 108164 21728 108220
rect 21784 108164 21832 108220
rect 21888 108164 21898 108220
rect 28418 108164 28428 108220
rect 28484 108164 28532 108220
rect 28588 108164 28636 108220
rect 28692 108164 28702 108220
rect 14914 107996 14924 108052
rect 14980 107996 16660 108052
rect 17388 108108 17500 108164
rect 17556 108108 17566 108164
rect 17388 107940 17444 108108
rect 16268 107884 17444 107940
rect 16268 107828 16324 107884
rect 9762 107772 9772 107828
rect 9828 107772 13580 107828
rect 13636 107772 13646 107828
rect 16258 107772 16268 107828
rect 16324 107772 16334 107828
rect 16818 107772 16828 107828
rect 16884 107772 20748 107828
rect 20804 107772 20814 107828
rect 7522 107660 7532 107716
rect 7588 107660 12236 107716
rect 12292 107660 12302 107716
rect 9874 107548 9884 107604
rect 9940 107548 12124 107604
rect 12180 107548 12190 107604
rect 21634 107548 21644 107604
rect 21700 107548 22428 107604
rect 22484 107548 23492 107604
rect 24322 107548 24332 107604
rect 24388 107548 24668 107604
rect 24724 107548 24734 107604
rect 23436 107492 23492 107548
rect 18946 107436 18956 107492
rect 19012 107436 19852 107492
rect 19908 107436 19918 107492
rect 23436 107436 24780 107492
rect 24836 107436 24846 107492
rect 4604 107380 4614 107436
rect 4670 107380 4718 107436
rect 4774 107380 4822 107436
rect 4878 107380 4888 107436
rect 11408 107380 11418 107436
rect 11474 107380 11522 107436
rect 11578 107380 11626 107436
rect 11682 107380 11692 107436
rect 18212 107380 18222 107436
rect 18278 107380 18326 107436
rect 18382 107380 18430 107436
rect 18486 107380 18496 107436
rect 25016 107380 25026 107436
rect 25082 107380 25130 107436
rect 25186 107380 25234 107436
rect 25290 107380 25300 107436
rect 9986 106988 9996 107044
rect 10052 106988 10780 107044
rect 10836 106988 11452 107044
rect 11508 106988 11518 107044
rect 11778 106988 11788 107044
rect 11844 106988 12460 107044
rect 12516 106988 12526 107044
rect 13570 106988 13580 107044
rect 13636 106988 16156 107044
rect 16212 106988 16222 107044
rect 17714 106988 17724 107044
rect 17780 106988 19964 107044
rect 20020 106988 20030 107044
rect 0 106932 400 106960
rect 0 106876 4284 106932
rect 4340 106876 4350 106932
rect 13458 106876 13468 106932
rect 13524 106876 14588 106932
rect 14644 106876 14654 106932
rect 0 106848 400 106876
rect 9650 106764 9660 106820
rect 9716 106764 10108 106820
rect 10164 106764 10174 106820
rect 17714 106764 17724 106820
rect 17780 106764 19180 106820
rect 19236 106764 19246 106820
rect 8006 106596 8016 106652
rect 8072 106596 8120 106652
rect 8176 106596 8224 106652
rect 8280 106596 8290 106652
rect 14810 106596 14820 106652
rect 14876 106596 14924 106652
rect 14980 106596 15028 106652
rect 15084 106596 15094 106652
rect 21614 106596 21624 106652
rect 21680 106596 21728 106652
rect 21784 106596 21832 106652
rect 21888 106596 21898 106652
rect 28418 106596 28428 106652
rect 28484 106596 28532 106652
rect 28588 106596 28636 106652
rect 28692 106596 28702 106652
rect 3938 106428 3948 106484
rect 4004 106428 5628 106484
rect 5684 106428 5694 106484
rect 21298 106428 21308 106484
rect 21364 106428 22316 106484
rect 22372 106428 22382 106484
rect 9090 106316 9100 106372
rect 9156 106316 12348 106372
rect 12404 106316 12414 106372
rect 8082 106204 8092 106260
rect 8148 106204 9996 106260
rect 10052 106204 10062 106260
rect 18946 106204 18956 106260
rect 19012 106204 22204 106260
rect 22260 106204 25340 106260
rect 25396 106204 25406 106260
rect 3154 106092 3164 106148
rect 3220 106092 3836 106148
rect 3892 106092 4956 106148
rect 5012 106092 5740 106148
rect 5796 106092 5806 106148
rect 7634 106092 7644 106148
rect 7700 106092 8540 106148
rect 8596 106092 8606 106148
rect 22530 106092 22540 106148
rect 22596 106092 23324 106148
rect 23380 106092 23772 106148
rect 23828 106092 23838 106148
rect 4834 105980 4844 106036
rect 4900 105980 5012 106036
rect 16482 105980 16492 106036
rect 16548 105980 17388 106036
rect 17444 105980 17454 106036
rect 24322 105980 24332 106036
rect 24388 105980 24892 106036
rect 24948 105980 24958 106036
rect 4604 105812 4614 105868
rect 4670 105812 4718 105868
rect 4774 105812 4822 105868
rect 4878 105812 4888 105868
rect 4956 105812 5012 105980
rect 12674 105868 12684 105924
rect 12740 105868 13580 105924
rect 13636 105868 13646 105924
rect 14578 105868 14588 105924
rect 14644 105868 15708 105924
rect 15764 105868 15774 105924
rect 11408 105812 11418 105868
rect 11474 105812 11522 105868
rect 11578 105812 11626 105868
rect 11682 105812 11692 105868
rect 18212 105812 18222 105868
rect 18278 105812 18326 105868
rect 18382 105812 18430 105868
rect 18486 105812 18496 105868
rect 25016 105812 25026 105868
rect 25082 105812 25130 105868
rect 25186 105812 25234 105868
rect 25290 105812 25300 105868
rect 4956 105756 7532 105812
rect 7588 105756 7598 105812
rect 4956 105700 5012 105756
rect 4050 105644 4060 105700
rect 4116 105644 5012 105700
rect 12674 105644 12684 105700
rect 12740 105644 20636 105700
rect 20692 105644 20702 105700
rect 24406 105644 24444 105700
rect 24500 105644 24510 105700
rect 6290 105532 6300 105588
rect 6356 105532 7756 105588
rect 7812 105532 7822 105588
rect 12786 105532 12796 105588
rect 12852 105532 17612 105588
rect 17668 105532 17678 105588
rect 20178 105532 20188 105588
rect 20244 105532 22204 105588
rect 22260 105532 26236 105588
rect 26292 105532 26302 105588
rect 26852 105532 28028 105588
rect 28084 105532 28252 105588
rect 28308 105532 28318 105588
rect 4498 105420 4508 105476
rect 4564 105420 5292 105476
rect 5348 105420 5358 105476
rect 8866 105308 8876 105364
rect 8932 105308 10444 105364
rect 10500 105308 10510 105364
rect 20290 105308 20300 105364
rect 20356 105308 21308 105364
rect 21364 105308 21374 105364
rect 23202 105308 23212 105364
rect 23268 105308 23884 105364
rect 23940 105308 24780 105364
rect 24836 105308 26068 105364
rect 26012 105252 26068 105308
rect 26852 105252 26908 105532
rect 4274 105196 4284 105252
rect 4340 105196 5852 105252
rect 5908 105196 5918 105252
rect 24658 105196 24668 105252
rect 24724 105196 25676 105252
rect 25732 105196 25742 105252
rect 26002 105196 26012 105252
rect 26068 105196 26684 105252
rect 26740 105196 26908 105252
rect 7522 105084 7532 105140
rect 7588 105084 7598 105140
rect 7532 104916 7588 105084
rect 8006 105028 8016 105084
rect 8072 105028 8120 105084
rect 8176 105028 8224 105084
rect 8280 105028 8290 105084
rect 14810 105028 14820 105084
rect 14876 105028 14924 105084
rect 14980 105028 15028 105084
rect 15084 105028 15094 105084
rect 21614 105028 21624 105084
rect 21680 105028 21728 105084
rect 21784 105028 21832 105084
rect 21888 105028 21898 105084
rect 28418 105028 28428 105084
rect 28484 105028 28532 105084
rect 28588 105028 28636 105084
rect 28692 105028 28702 105084
rect 1698 104860 1708 104916
rect 1764 104860 3836 104916
rect 3892 104860 3902 104916
rect 6850 104860 6860 104916
rect 6916 104860 8092 104916
rect 8148 104860 8158 104916
rect 8306 104860 8316 104916
rect 8372 104860 12684 104916
rect 12740 104860 18620 104916
rect 18676 104860 18686 104916
rect 4274 104748 4284 104804
rect 4340 104748 12796 104804
rect 12852 104748 12862 104804
rect 19058 104748 19068 104804
rect 19124 104748 20300 104804
rect 20356 104748 20366 104804
rect 3714 104636 3724 104692
rect 3780 104636 5180 104692
rect 5236 104636 6524 104692
rect 6580 104636 7644 104692
rect 7700 104636 7710 104692
rect 8978 104636 8988 104692
rect 9044 104636 11788 104692
rect 11844 104636 11854 104692
rect 14242 104636 14252 104692
rect 14308 104636 18508 104692
rect 18564 104636 18574 104692
rect 3266 104524 3276 104580
rect 3332 104524 4396 104580
rect 4452 104524 4462 104580
rect 7074 104524 7084 104580
rect 7140 104524 15260 104580
rect 15316 104524 15326 104580
rect 7868 104468 7924 104524
rect 5842 104412 5852 104468
rect 5908 104412 7532 104468
rect 7588 104412 7598 104468
rect 7858 104412 7868 104468
rect 7924 104412 7934 104468
rect 11218 104412 11228 104468
rect 11284 104412 12460 104468
rect 12516 104412 12526 104468
rect 13794 104412 13804 104468
rect 13860 104412 13870 104468
rect 8502 104300 8540 104356
rect 8596 104300 8606 104356
rect 0 104244 400 104272
rect 4604 104244 4614 104300
rect 4670 104244 4718 104300
rect 4774 104244 4822 104300
rect 4878 104244 4888 104300
rect 11408 104244 11418 104300
rect 11474 104244 11522 104300
rect 11578 104244 11626 104300
rect 11682 104244 11692 104300
rect 13804 104244 13860 104412
rect 15026 104300 15036 104356
rect 15092 104300 15820 104356
rect 15876 104300 15886 104356
rect 22306 104300 22316 104356
rect 22372 104300 23660 104356
rect 23716 104300 23726 104356
rect 18212 104244 18222 104300
rect 18278 104244 18326 104300
rect 18382 104244 18430 104300
rect 18486 104244 18496 104300
rect 25016 104244 25026 104300
rect 25082 104244 25130 104300
rect 25186 104244 25234 104300
rect 25290 104244 25300 104300
rect 0 104188 1764 104244
rect 8306 104188 8316 104244
rect 8372 104188 8652 104244
rect 8708 104188 8718 104244
rect 13804 104188 16044 104244
rect 16100 104188 16110 104244
rect 23426 104188 23436 104244
rect 23492 104188 23772 104244
rect 23828 104188 23838 104244
rect 0 104160 400 104188
rect 1708 104020 1764 104188
rect 5058 104076 5068 104132
rect 5124 104076 8988 104132
rect 9044 104076 9054 104132
rect 9202 104076 9212 104132
rect 9268 104076 10108 104132
rect 10164 104076 12908 104132
rect 12964 104076 14700 104132
rect 14756 104076 14766 104132
rect 17938 104076 17948 104132
rect 18004 104076 18396 104132
rect 18452 104076 18462 104132
rect 23986 104076 23996 104132
rect 24052 104076 24444 104132
rect 24500 104076 24510 104132
rect 26674 104076 26684 104132
rect 26740 104076 27580 104132
rect 27636 104076 27646 104132
rect 1698 103964 1708 104020
rect 1764 103964 1774 104020
rect 4834 103964 4844 104020
rect 4900 103964 17164 104020
rect 17220 103964 17230 104020
rect 5282 103852 5292 103908
rect 5348 103852 8876 103908
rect 8932 103852 8942 103908
rect 9874 103852 9884 103908
rect 9940 103852 16828 103908
rect 16884 103852 16894 103908
rect 7074 103740 7084 103796
rect 7140 103740 7980 103796
rect 8036 103740 8046 103796
rect 8502 103740 8540 103796
rect 8596 103740 8606 103796
rect 9426 103740 9436 103796
rect 9492 103740 9548 103796
rect 9604 103740 9614 103796
rect 10098 103740 10108 103796
rect 10164 103740 10668 103796
rect 10724 103740 10734 103796
rect 11106 103740 11116 103796
rect 11172 103740 17500 103796
rect 17556 103740 17566 103796
rect 3266 103628 3276 103684
rect 3332 103628 4956 103684
rect 5012 103628 5022 103684
rect 7634 103628 7644 103684
rect 7700 103628 14812 103684
rect 14868 103628 14878 103684
rect 8866 103516 8876 103572
rect 8932 103516 14252 103572
rect 14308 103516 14318 103572
rect 8006 103460 8016 103516
rect 8072 103460 8120 103516
rect 8176 103460 8224 103516
rect 8280 103460 8290 103516
rect 14810 103460 14820 103516
rect 14876 103460 14924 103516
rect 14980 103460 15028 103516
rect 15084 103460 15094 103516
rect 21614 103460 21624 103516
rect 21680 103460 21728 103516
rect 21784 103460 21832 103516
rect 21888 103460 21898 103516
rect 28418 103460 28428 103516
rect 28484 103460 28532 103516
rect 28588 103460 28636 103516
rect 28692 103460 28702 103516
rect 9548 103404 11788 103460
rect 11844 103404 11854 103460
rect 9548 103348 9604 103404
rect 1698 103292 1708 103348
rect 1764 103292 4284 103348
rect 4340 103292 4350 103348
rect 4946 103292 4956 103348
rect 5012 103292 6972 103348
rect 7028 103292 7038 103348
rect 8194 103292 8204 103348
rect 8260 103292 9548 103348
rect 9604 103292 9614 103348
rect 10210 103292 10220 103348
rect 10276 103292 23324 103348
rect 23380 103292 23390 103348
rect 3490 103180 3500 103236
rect 3556 103180 4060 103236
rect 4116 103180 4126 103236
rect 6402 103180 6412 103236
rect 6468 103180 7756 103236
rect 7812 103180 8316 103236
rect 8372 103180 8382 103236
rect 9436 103180 12572 103236
rect 12628 103180 12638 103236
rect 13010 103180 13020 103236
rect 13076 103180 16492 103236
rect 16548 103180 22428 103236
rect 22484 103180 22494 103236
rect 9436 103124 9492 103180
rect 2594 103068 2604 103124
rect 2660 103068 3948 103124
rect 4004 103068 4844 103124
rect 4900 103068 4910 103124
rect 8978 103068 8988 103124
rect 9044 103068 9492 103124
rect 9650 103068 9660 103124
rect 9716 103068 10668 103124
rect 10724 103068 10734 103124
rect 11106 103068 11116 103124
rect 11172 103068 14924 103124
rect 14980 103068 14990 103124
rect 22530 103068 22540 103124
rect 22596 103068 24220 103124
rect 24276 103068 24286 103124
rect 3602 102956 3612 103012
rect 3668 102956 10780 103012
rect 10836 102956 10846 103012
rect 11218 102956 11228 103012
rect 11284 102956 13804 103012
rect 13860 102956 13870 103012
rect 20626 102956 20636 103012
rect 20692 102956 22988 103012
rect 23044 102956 23660 103012
rect 23716 102956 24556 103012
rect 24612 102956 25340 103012
rect 25396 102956 25406 103012
rect 6850 102844 6860 102900
rect 6916 102844 9212 102900
rect 9268 102844 9278 102900
rect 9874 102844 9884 102900
rect 9940 102844 10668 102900
rect 10724 102844 11116 102900
rect 11172 102844 11182 102900
rect 8306 102732 8316 102788
rect 8372 102732 8382 102788
rect 8978 102732 8988 102788
rect 9044 102732 9436 102788
rect 9492 102732 9502 102788
rect 9650 102732 9660 102788
rect 9716 102732 9754 102788
rect 10322 102732 10332 102788
rect 10388 102732 11228 102788
rect 11284 102732 11294 102788
rect 4604 102676 4614 102732
rect 4670 102676 4718 102732
rect 4774 102676 4822 102732
rect 4878 102676 4888 102732
rect 8316 102676 8372 102732
rect 11408 102676 11418 102732
rect 11474 102676 11522 102732
rect 11578 102676 11626 102732
rect 11682 102676 11692 102732
rect 18212 102676 18222 102732
rect 18278 102676 18326 102732
rect 18382 102676 18430 102732
rect 18486 102676 18496 102732
rect 25016 102676 25026 102732
rect 25082 102676 25130 102732
rect 25186 102676 25234 102732
rect 25290 102676 25300 102732
rect 8316 102620 9212 102676
rect 9268 102620 10108 102676
rect 10164 102620 10174 102676
rect 6486 102508 6524 102564
rect 6580 102508 10220 102564
rect 10276 102508 10286 102564
rect 20178 102508 20188 102564
rect 20244 102508 21756 102564
rect 21812 102508 21822 102564
rect 12572 102396 13580 102452
rect 13636 102396 13646 102452
rect 15092 102396 17612 102452
rect 17668 102396 17678 102452
rect 18834 102396 18844 102452
rect 18900 102396 22764 102452
rect 22820 102396 23884 102452
rect 23940 102396 24780 102452
rect 24836 102396 24846 102452
rect 12572 102340 12628 102396
rect 15092 102340 15148 102396
rect 3332 102228 3388 102340
rect 3444 102284 4284 102340
rect 4340 102284 4350 102340
rect 8754 102284 8764 102340
rect 8820 102284 10108 102340
rect 10164 102284 12124 102340
rect 12180 102284 12572 102340
rect 12628 102284 12638 102340
rect 13458 102284 13468 102340
rect 13524 102284 14140 102340
rect 14196 102284 15148 102340
rect 17826 102284 17836 102340
rect 17892 102284 20972 102340
rect 21028 102284 21868 102340
rect 21924 102284 23212 102340
rect 23268 102284 23278 102340
rect 2706 102172 2716 102228
rect 2772 102172 3388 102228
rect 8978 102172 8988 102228
rect 9044 102172 9436 102228
rect 9492 102172 9502 102228
rect 9650 102172 9660 102228
rect 9716 102172 19740 102228
rect 19796 102172 19806 102228
rect 4274 102060 4284 102116
rect 4340 102060 4732 102116
rect 4788 102060 4798 102116
rect 6850 102060 6860 102116
rect 6916 102060 8652 102116
rect 8708 102060 9884 102116
rect 9940 102060 9950 102116
rect 8006 101892 8016 101948
rect 8072 101892 8120 101948
rect 8176 101892 8224 101948
rect 8280 101892 8290 101948
rect 14810 101892 14820 101948
rect 14876 101892 14924 101948
rect 14980 101892 15028 101948
rect 15084 101892 15094 101948
rect 21614 101892 21624 101948
rect 21680 101892 21728 101948
rect 21784 101892 21832 101948
rect 21888 101892 21898 101948
rect 28418 101892 28428 101948
rect 28484 101892 28532 101948
rect 28588 101892 28636 101948
rect 28692 101892 28702 101948
rect 8530 101836 8540 101892
rect 8596 101836 9212 101892
rect 9268 101836 9278 101892
rect 1698 101612 1708 101668
rect 1764 101612 3500 101668
rect 3556 101612 3566 101668
rect 9538 101612 9548 101668
rect 9604 101612 9884 101668
rect 9940 101612 9950 101668
rect 0 101556 400 101584
rect 1708 101556 1764 101612
rect 0 101500 1764 101556
rect 3042 101500 3052 101556
rect 3108 101500 4396 101556
rect 4452 101500 4462 101556
rect 5058 101500 5068 101556
rect 5124 101500 5852 101556
rect 5908 101500 6860 101556
rect 6916 101500 6926 101556
rect 21298 101500 21308 101556
rect 21364 101500 23884 101556
rect 23940 101500 23950 101556
rect 0 101472 400 101500
rect 5170 101388 5180 101444
rect 5236 101388 10220 101444
rect 10276 101388 10286 101444
rect 7746 101276 7756 101332
rect 7812 101276 9772 101332
rect 9828 101276 12012 101332
rect 12068 101276 12796 101332
rect 12852 101276 12862 101332
rect 15092 101276 18844 101332
rect 18900 101276 18910 101332
rect 4604 101108 4614 101164
rect 4670 101108 4718 101164
rect 4774 101108 4822 101164
rect 4878 101108 4888 101164
rect 11408 101108 11418 101164
rect 11474 101108 11522 101164
rect 11578 101108 11626 101164
rect 11682 101108 11692 101164
rect 8866 100940 8876 100996
rect 8932 100940 10780 100996
rect 10836 100940 11116 100996
rect 11172 100940 12236 100996
rect 12292 100940 12908 100996
rect 12964 100940 14028 100996
rect 14084 100940 14094 100996
rect 15092 100884 15148 101276
rect 18212 101108 18222 101164
rect 18278 101108 18326 101164
rect 18382 101108 18430 101164
rect 18486 101108 18496 101164
rect 25016 101108 25026 101164
rect 25082 101108 25130 101164
rect 25186 101108 25234 101164
rect 25290 101108 25300 101164
rect 18274 100940 18284 100996
rect 18340 100940 19404 100996
rect 19460 100940 19470 100996
rect 7410 100828 7420 100884
rect 7476 100828 8764 100884
rect 8820 100828 8830 100884
rect 9314 100828 9324 100884
rect 9380 100828 9772 100884
rect 9828 100828 9838 100884
rect 12562 100828 12572 100884
rect 12628 100828 15148 100884
rect 17938 100828 17948 100884
rect 18004 100828 18732 100884
rect 18788 100828 18798 100884
rect 5618 100716 5628 100772
rect 5684 100716 6524 100772
rect 6580 100716 7700 100772
rect 9202 100716 9212 100772
rect 9268 100716 13468 100772
rect 13524 100716 13534 100772
rect 14578 100716 14588 100772
rect 14644 100716 15540 100772
rect 17490 100716 17500 100772
rect 17556 100716 20076 100772
rect 20132 100716 21868 100772
rect 21924 100716 23324 100772
rect 23380 100716 23390 100772
rect 24210 100716 24220 100772
rect 24276 100716 24892 100772
rect 24948 100716 24958 100772
rect 7644 100660 7700 100716
rect 15484 100660 15540 100716
rect 2594 100604 2604 100660
rect 2660 100604 3388 100660
rect 4834 100604 4844 100660
rect 4900 100604 5740 100660
rect 5796 100604 5964 100660
rect 6020 100604 6030 100660
rect 6402 100604 6412 100660
rect 6468 100604 7420 100660
rect 7476 100604 7486 100660
rect 7644 100604 10444 100660
rect 10500 100604 10510 100660
rect 15474 100604 15484 100660
rect 15540 100604 15550 100660
rect 21410 100604 21420 100660
rect 21476 100604 21486 100660
rect 25442 100604 25452 100660
rect 25508 100604 26684 100660
rect 26740 100604 26750 100660
rect 3332 100548 3388 100604
rect 21420 100548 21476 100604
rect 3332 100492 3948 100548
rect 4004 100492 21476 100548
rect 4946 100380 4956 100436
rect 5012 100380 7308 100436
rect 7364 100380 7374 100436
rect 9538 100380 9548 100436
rect 9604 100380 10108 100436
rect 10164 100380 10668 100436
rect 10724 100380 10734 100436
rect 8006 100324 8016 100380
rect 8072 100324 8120 100380
rect 8176 100324 8224 100380
rect 8280 100324 8290 100380
rect 14810 100324 14820 100380
rect 14876 100324 14924 100380
rect 14980 100324 15028 100380
rect 15084 100324 15094 100380
rect 21614 100324 21624 100380
rect 21680 100324 21728 100380
rect 21784 100324 21832 100380
rect 21888 100324 21898 100380
rect 28418 100324 28428 100380
rect 28484 100324 28532 100380
rect 28588 100324 28636 100380
rect 28692 100324 28702 100380
rect 6178 100268 6188 100324
rect 6244 100268 7756 100324
rect 7812 100268 7822 100324
rect 4274 100156 4284 100212
rect 4340 100156 8988 100212
rect 9044 100156 9884 100212
rect 9940 100156 9950 100212
rect 7522 99932 7532 99988
rect 7588 99932 10108 99988
rect 10164 99932 10174 99988
rect 22306 99932 22316 99988
rect 22372 99932 23324 99988
rect 23380 99932 24108 99988
rect 24164 99932 24174 99988
rect 24882 99932 24892 99988
rect 24948 99932 27356 99988
rect 27412 99932 28028 99988
rect 28084 99932 28094 99988
rect 7074 99820 7084 99876
rect 7140 99820 13580 99876
rect 13636 99820 13646 99876
rect 4604 99540 4614 99596
rect 4670 99540 4718 99596
rect 4774 99540 4822 99596
rect 4878 99540 4888 99596
rect 11408 99540 11418 99596
rect 11474 99540 11522 99596
rect 11578 99540 11626 99596
rect 11682 99540 11692 99596
rect 18212 99540 18222 99596
rect 18278 99540 18326 99596
rect 18382 99540 18430 99596
rect 18486 99540 18496 99596
rect 25016 99540 25026 99596
rect 25082 99540 25130 99596
rect 25186 99540 25234 99596
rect 25290 99540 25300 99596
rect 18834 99484 18844 99540
rect 18900 99484 20636 99540
rect 20692 99484 20702 99540
rect 5170 99372 5180 99428
rect 5236 99372 8540 99428
rect 8596 99372 12572 99428
rect 12628 99372 12638 99428
rect 18162 99372 18172 99428
rect 18228 99372 19964 99428
rect 20020 99372 20030 99428
rect 10994 99260 11004 99316
rect 11060 99260 15484 99316
rect 15540 99260 15550 99316
rect 5730 99148 5740 99204
rect 5796 99148 5806 99204
rect 6626 99148 6636 99204
rect 6692 99148 7644 99204
rect 7700 99148 7710 99204
rect 16706 99148 16716 99204
rect 16772 99148 19180 99204
rect 19236 99148 19246 99204
rect 19730 99148 19740 99204
rect 19796 99148 21084 99204
rect 21140 99148 21756 99204
rect 21812 99148 23660 99204
rect 23716 99148 23726 99204
rect 5740 99092 5796 99148
rect 5740 99036 6860 99092
rect 6916 99036 6926 99092
rect 7410 99036 7420 99092
rect 7476 99036 9884 99092
rect 9940 99036 9950 99092
rect 10546 99036 10556 99092
rect 10612 99036 15148 99092
rect 15204 99036 15214 99092
rect 15474 99036 15484 99092
rect 15540 99036 18060 99092
rect 18116 99036 18126 99092
rect 19282 99036 19292 99092
rect 19348 99036 20748 99092
rect 20804 99036 20814 99092
rect 21970 99036 21980 99092
rect 22036 99036 23884 99092
rect 23940 99036 24668 99092
rect 24724 99036 24734 99092
rect 8754 98924 8764 98980
rect 8820 98924 11900 98980
rect 11956 98924 11966 98980
rect 17378 98924 17388 98980
rect 17444 98924 17836 98980
rect 17892 98924 19516 98980
rect 19572 98924 19582 98980
rect 20066 98924 20076 98980
rect 20132 98924 22764 98980
rect 22820 98924 23772 98980
rect 23828 98924 25676 98980
rect 25732 98924 25742 98980
rect 0 98868 400 98896
rect 0 98812 1708 98868
rect 1764 98812 3276 98868
rect 3332 98812 3342 98868
rect 0 98784 400 98812
rect 8006 98756 8016 98812
rect 8072 98756 8120 98812
rect 8176 98756 8224 98812
rect 8280 98756 8290 98812
rect 14810 98756 14820 98812
rect 14876 98756 14924 98812
rect 14980 98756 15028 98812
rect 15084 98756 15094 98812
rect 21614 98756 21624 98812
rect 21680 98756 21728 98812
rect 21784 98756 21832 98812
rect 21888 98756 21898 98812
rect 28418 98756 28428 98812
rect 28484 98756 28532 98812
rect 28588 98756 28636 98812
rect 28692 98756 28702 98812
rect 2818 98700 2828 98756
rect 2884 98700 3164 98756
rect 3220 98700 4452 98756
rect 17910 98700 17948 98756
rect 18004 98700 18014 98756
rect 4396 98644 4452 98700
rect 4386 98588 4396 98644
rect 4452 98588 6188 98644
rect 6244 98588 6254 98644
rect 19170 98588 19180 98644
rect 19236 98588 21868 98644
rect 21924 98588 21934 98644
rect 4050 98476 4060 98532
rect 4116 98476 5852 98532
rect 5908 98476 5918 98532
rect 9426 98476 9436 98532
rect 9492 98476 11788 98532
rect 11844 98476 11854 98532
rect 17938 98476 17948 98532
rect 18004 98476 18060 98532
rect 18116 98476 18126 98532
rect 21186 98476 21196 98532
rect 21252 98476 22204 98532
rect 22260 98476 24444 98532
rect 24500 98476 25228 98532
rect 25284 98476 25676 98532
rect 25732 98476 25742 98532
rect 2370 98364 2380 98420
rect 2436 98364 2716 98420
rect 2772 98364 3388 98420
rect 3444 98364 3454 98420
rect 5170 98364 5180 98420
rect 5236 98364 8764 98420
rect 8820 98364 9548 98420
rect 9604 98364 9614 98420
rect 18274 98364 18284 98420
rect 18340 98364 20188 98420
rect 20244 98364 20254 98420
rect 4946 98252 4956 98308
rect 5012 98252 5964 98308
rect 6020 98252 12348 98308
rect 12404 98252 12414 98308
rect 7522 98028 7532 98084
rect 7588 98028 10332 98084
rect 10388 98028 10398 98084
rect 4604 97972 4614 98028
rect 4670 97972 4718 98028
rect 4774 97972 4822 98028
rect 4878 97972 4888 98028
rect 10556 97972 10612 98252
rect 15922 98140 15932 98196
rect 15988 98140 18620 98196
rect 18676 98140 21868 98196
rect 21924 98140 21934 98196
rect 23874 98140 23884 98196
rect 23940 98140 27356 98196
rect 27412 98140 27422 98196
rect 11408 97972 11418 98028
rect 11474 97972 11522 98028
rect 11578 97972 11626 98028
rect 11682 97972 11692 98028
rect 18212 97972 18222 98028
rect 18278 97972 18326 98028
rect 18382 97972 18430 98028
rect 18486 97972 18496 98028
rect 25016 97972 25026 98028
rect 25082 97972 25130 98028
rect 25186 97972 25234 98028
rect 25290 97972 25300 98028
rect 10434 97916 10444 97972
rect 10500 97916 10612 97972
rect 23986 97916 23996 97972
rect 24052 97916 24062 97972
rect 23996 97860 24052 97916
rect 4610 97804 4620 97860
rect 4676 97804 7084 97860
rect 7140 97804 7150 97860
rect 19954 97804 19964 97860
rect 20020 97804 21980 97860
rect 22036 97804 22046 97860
rect 23996 97804 25340 97860
rect 25396 97804 25406 97860
rect 2594 97692 2604 97748
rect 2660 97692 3276 97748
rect 3332 97692 4956 97748
rect 5012 97692 5022 97748
rect 6290 97692 6300 97748
rect 6356 97692 6860 97748
rect 6916 97692 6926 97748
rect 15026 97692 15036 97748
rect 15092 97692 15260 97748
rect 15316 97692 17388 97748
rect 17444 97692 17454 97748
rect 19394 97692 19404 97748
rect 19460 97692 22540 97748
rect 22596 97692 22606 97748
rect 23650 97692 23660 97748
rect 23716 97692 24668 97748
rect 24724 97692 25452 97748
rect 25508 97692 25518 97748
rect 3826 97580 3836 97636
rect 3892 97580 5628 97636
rect 5684 97580 5852 97636
rect 5908 97580 5918 97636
rect 6066 97580 6076 97636
rect 6132 97580 6748 97636
rect 6804 97580 6814 97636
rect 9986 97580 9996 97636
rect 10052 97580 14700 97636
rect 14756 97580 14766 97636
rect 15586 97580 15596 97636
rect 15652 97580 15932 97636
rect 15988 97580 15998 97636
rect 18050 97580 18060 97636
rect 18116 97580 18508 97636
rect 18564 97580 18574 97636
rect 20066 97580 20076 97636
rect 20132 97580 20860 97636
rect 20916 97580 20926 97636
rect 22194 97580 22204 97636
rect 22260 97580 23100 97636
rect 23156 97580 23166 97636
rect 23314 97580 23324 97636
rect 23380 97580 25116 97636
rect 25172 97580 25182 97636
rect 25554 97580 25564 97636
rect 25620 97580 26796 97636
rect 26852 97580 27356 97636
rect 27412 97580 27422 97636
rect 24220 97524 24276 97580
rect 5058 97468 5068 97524
rect 5124 97468 6636 97524
rect 6692 97468 6702 97524
rect 14130 97468 14140 97524
rect 14196 97468 14588 97524
rect 14644 97468 14654 97524
rect 18162 97468 18172 97524
rect 18228 97468 18956 97524
rect 19012 97468 19022 97524
rect 19842 97468 19852 97524
rect 19908 97468 21420 97524
rect 21476 97468 21486 97524
rect 22866 97468 22876 97524
rect 22932 97468 23772 97524
rect 23828 97468 23838 97524
rect 24210 97468 24220 97524
rect 24276 97468 24286 97524
rect 24882 97468 24892 97524
rect 24948 97468 26684 97524
rect 26740 97468 26750 97524
rect 7532 97356 24444 97412
rect 24500 97356 24510 97412
rect 7532 97300 7588 97356
rect 7522 97244 7532 97300
rect 7588 97244 7598 97300
rect 8978 97244 8988 97300
rect 9044 97244 10108 97300
rect 10164 97244 10174 97300
rect 14214 97244 14252 97300
rect 14308 97244 14318 97300
rect 16482 97244 16492 97300
rect 16548 97244 18732 97300
rect 18788 97244 18798 97300
rect 8006 97188 8016 97244
rect 8072 97188 8120 97244
rect 8176 97188 8224 97244
rect 8280 97188 8290 97244
rect 14810 97188 14820 97244
rect 14876 97188 14924 97244
rect 14980 97188 15028 97244
rect 15084 97188 15094 97244
rect 21614 97188 21624 97244
rect 21680 97188 21728 97244
rect 21784 97188 21832 97244
rect 21888 97188 21898 97244
rect 28418 97188 28428 97244
rect 28484 97188 28532 97244
rect 28588 97188 28636 97244
rect 28692 97188 28702 97244
rect 9986 97132 9996 97188
rect 10052 97132 10556 97188
rect 10612 97132 12012 97188
rect 12068 97132 12078 97188
rect 14018 97132 14028 97188
rect 14084 97132 14140 97188
rect 14196 97132 14206 97188
rect 14354 97132 14364 97188
rect 14420 97132 14458 97188
rect 16370 97132 16380 97188
rect 16436 97132 17780 97188
rect 17938 97132 17948 97188
rect 18004 97132 19516 97188
rect 19572 97132 19582 97188
rect 17724 97076 17780 97132
rect 8866 97020 8876 97076
rect 8932 97020 9660 97076
rect 9716 97020 9726 97076
rect 12114 97020 12124 97076
rect 12180 97020 12460 97076
rect 12516 97020 12526 97076
rect 13458 97020 13468 97076
rect 13524 97020 16716 97076
rect 16772 97020 16782 97076
rect 16930 97020 16940 97076
rect 16996 97020 17500 97076
rect 17556 97020 17566 97076
rect 17724 97020 18396 97076
rect 18452 97020 18844 97076
rect 18900 97020 18910 97076
rect 10322 96908 10332 96964
rect 10388 96908 13692 96964
rect 13748 96908 13758 96964
rect 13906 96908 13916 96964
rect 13972 96908 14028 96964
rect 14084 96908 14094 96964
rect 14242 96908 14252 96964
rect 14308 96908 20188 96964
rect 20244 96908 20254 96964
rect 8754 96796 8764 96852
rect 8820 96796 8830 96852
rect 12562 96796 12572 96852
rect 12628 96796 16380 96852
rect 16436 96796 16446 96852
rect 17490 96796 17500 96852
rect 17556 96796 17948 96852
rect 18004 96796 18014 96852
rect 21298 96796 21308 96852
rect 21364 96796 22092 96852
rect 22148 96796 22158 96852
rect 8764 96740 8820 96796
rect 3154 96684 3164 96740
rect 3220 96684 3836 96740
rect 3892 96684 3902 96740
rect 4162 96684 4172 96740
rect 4228 96684 5740 96740
rect 5796 96684 5806 96740
rect 8764 96684 17836 96740
rect 17892 96684 17902 96740
rect 18060 96684 19068 96740
rect 19124 96684 19852 96740
rect 19908 96684 19918 96740
rect 23874 96684 23884 96740
rect 23940 96684 26236 96740
rect 26292 96684 26302 96740
rect 4172 96628 4228 96684
rect 3378 96572 3388 96628
rect 3444 96572 4228 96628
rect 10210 96572 10220 96628
rect 10276 96572 13188 96628
rect 13346 96572 13356 96628
rect 13412 96572 15148 96628
rect 15204 96572 16324 96628
rect 13132 96516 13188 96572
rect 16268 96516 16324 96572
rect 18060 96516 18116 96684
rect 20178 96572 20188 96628
rect 20244 96572 20524 96628
rect 20580 96572 20590 96628
rect 13122 96460 13132 96516
rect 13188 96460 15596 96516
rect 15652 96460 15820 96516
rect 15876 96460 15886 96516
rect 16268 96460 18116 96516
rect 4604 96404 4614 96460
rect 4670 96404 4718 96460
rect 4774 96404 4822 96460
rect 4878 96404 4888 96460
rect 11408 96404 11418 96460
rect 11474 96404 11522 96460
rect 11578 96404 11626 96460
rect 11682 96404 11692 96460
rect 18212 96404 18222 96460
rect 18278 96404 18326 96460
rect 18382 96404 18430 96460
rect 18486 96404 18496 96460
rect 25016 96404 25026 96460
rect 25082 96404 25130 96460
rect 25186 96404 25234 96460
rect 25290 96404 25300 96460
rect 5954 96348 5964 96404
rect 6020 96348 10892 96404
rect 10948 96348 10958 96404
rect 12338 96348 12348 96404
rect 12404 96348 14028 96404
rect 14084 96348 14094 96404
rect 14242 96348 14252 96404
rect 14308 96348 15372 96404
rect 15428 96348 15438 96404
rect 12002 96236 12012 96292
rect 12068 96236 13748 96292
rect 13906 96236 13916 96292
rect 13972 96236 15596 96292
rect 15652 96236 15662 96292
rect 16258 96236 16268 96292
rect 16324 96236 19740 96292
rect 19796 96236 19806 96292
rect 0 96180 400 96208
rect 13692 96180 13748 96236
rect 16268 96180 16324 96236
rect 0 96124 1708 96180
rect 1764 96124 2268 96180
rect 2324 96124 2334 96180
rect 5506 96124 5516 96180
rect 5572 96124 6636 96180
rect 6692 96124 6702 96180
rect 10770 96124 10780 96180
rect 10836 96124 12124 96180
rect 12180 96124 12190 96180
rect 13692 96124 14588 96180
rect 14644 96124 14700 96180
rect 14756 96124 14766 96180
rect 15036 96124 16324 96180
rect 16706 96124 16716 96180
rect 16772 96124 20636 96180
rect 20692 96124 20702 96180
rect 0 96096 400 96124
rect 15036 96068 15092 96124
rect 7186 96012 7196 96068
rect 7252 96012 11788 96068
rect 11844 96012 15092 96068
rect 16594 96012 16604 96068
rect 16660 96012 17724 96068
rect 17780 96012 17790 96068
rect 20076 96012 20860 96068
rect 20916 96012 20926 96068
rect 24434 96012 24444 96068
rect 24500 96012 25228 96068
rect 25284 96012 25294 96068
rect 20076 95956 20132 96012
rect 6066 95900 6076 95956
rect 6132 95900 11004 95956
rect 11060 95900 11900 95956
rect 11956 95900 12124 95956
rect 12180 95900 12190 95956
rect 13580 95900 14812 95956
rect 14868 95900 18844 95956
rect 18900 95900 19628 95956
rect 19684 95900 19694 95956
rect 19852 95900 20076 95956
rect 20132 95900 20142 95956
rect 20626 95900 20636 95956
rect 20692 95900 22316 95956
rect 22372 95900 23212 95956
rect 23268 95900 23278 95956
rect 24546 95900 24556 95956
rect 24612 95900 25340 95956
rect 25396 95900 25406 95956
rect 5394 95788 5404 95844
rect 5460 95788 7756 95844
rect 7812 95788 7822 95844
rect 10882 95788 10892 95844
rect 10948 95788 13356 95844
rect 13412 95788 13422 95844
rect 13580 95732 13636 95900
rect 19852 95844 19908 95900
rect 14326 95788 14364 95844
rect 14420 95788 14430 95844
rect 15250 95788 15260 95844
rect 15316 95788 15820 95844
rect 15876 95788 15886 95844
rect 19842 95788 19852 95844
rect 19908 95788 19918 95844
rect 20076 95788 21084 95844
rect 21140 95788 21644 95844
rect 21700 95788 21710 95844
rect 23314 95788 23324 95844
rect 23380 95788 25452 95844
rect 25508 95788 25518 95844
rect 26226 95788 26236 95844
rect 26292 95788 27132 95844
rect 27188 95788 27198 95844
rect 20076 95732 20132 95788
rect 3266 95676 3276 95732
rect 3332 95620 3388 95732
rect 8418 95676 8428 95732
rect 8484 95676 10668 95732
rect 10724 95676 10734 95732
rect 11330 95676 11340 95732
rect 11396 95676 13636 95732
rect 15922 95676 15932 95732
rect 15988 95676 16716 95732
rect 16772 95676 16782 95732
rect 20066 95676 20076 95732
rect 20132 95676 20142 95732
rect 8006 95620 8016 95676
rect 8072 95620 8120 95676
rect 8176 95620 8224 95676
rect 8280 95620 8290 95676
rect 14810 95620 14820 95676
rect 14876 95620 14924 95676
rect 14980 95620 15028 95676
rect 15084 95620 15094 95676
rect 21614 95620 21624 95676
rect 21680 95620 21728 95676
rect 21784 95620 21832 95676
rect 21888 95620 21898 95676
rect 28418 95620 28428 95676
rect 28484 95620 28532 95676
rect 28588 95620 28636 95676
rect 28692 95620 28702 95676
rect 3332 95564 7700 95620
rect 8530 95564 8540 95620
rect 8596 95564 13300 95620
rect 2370 95452 2380 95508
rect 2436 95452 6076 95508
rect 6132 95452 6142 95508
rect 6514 95452 6524 95508
rect 6580 95452 6860 95508
rect 6916 95452 6926 95508
rect 7644 95396 7700 95564
rect 13244 95508 13300 95564
rect 7858 95452 7868 95508
rect 7924 95452 10220 95508
rect 10276 95452 11116 95508
rect 11172 95452 11182 95508
rect 13234 95452 13244 95508
rect 13300 95452 14812 95508
rect 14868 95452 16268 95508
rect 16324 95452 16828 95508
rect 16884 95452 16894 95508
rect 17266 95452 17276 95508
rect 17332 95452 18844 95508
rect 18900 95452 20524 95508
rect 20580 95452 23436 95508
rect 23492 95452 23502 95508
rect 2818 95340 2828 95396
rect 2884 95340 5628 95396
rect 5684 95340 5694 95396
rect 7644 95340 11228 95396
rect 11284 95340 11294 95396
rect 11788 95340 28140 95396
rect 28196 95340 28206 95396
rect 5394 95228 5404 95284
rect 5460 95228 9660 95284
rect 9716 95228 9726 95284
rect 3714 95116 3724 95172
rect 3780 95116 4508 95172
rect 4564 95116 5180 95172
rect 5236 95116 5246 95172
rect 6290 95116 6300 95172
rect 6356 95116 6972 95172
rect 7028 95116 7038 95172
rect 7634 95116 7644 95172
rect 7700 95116 11340 95172
rect 11396 95116 11406 95172
rect 11788 95060 11844 95340
rect 13570 95228 13580 95284
rect 13636 95228 14140 95284
rect 14196 95228 14206 95284
rect 14578 95228 14588 95284
rect 14644 95228 15596 95284
rect 15652 95228 15662 95284
rect 16370 95228 16380 95284
rect 16436 95228 17612 95284
rect 17668 95228 17678 95284
rect 24210 95228 24220 95284
rect 24276 95228 25340 95284
rect 25396 95228 25406 95284
rect 25554 95228 25564 95284
rect 25620 95228 26012 95284
rect 26068 95228 26078 95284
rect 12338 95116 12348 95172
rect 12404 95116 13692 95172
rect 13748 95116 13758 95172
rect 13906 95116 13916 95172
rect 13972 95116 15372 95172
rect 15428 95116 17388 95172
rect 17444 95116 17454 95172
rect 19030 95116 19068 95172
rect 19124 95116 19134 95172
rect 3938 95004 3948 95060
rect 4004 95004 11788 95060
rect 11844 95004 11854 95060
rect 14354 95004 14364 95060
rect 14420 95004 15932 95060
rect 15988 95004 15998 95060
rect 16482 95004 16492 95060
rect 16548 95004 18396 95060
rect 18452 95004 18462 95060
rect 5842 94892 5852 94948
rect 5908 94892 7532 94948
rect 7588 94892 7598 94948
rect 15092 94892 17500 94948
rect 17556 94892 17566 94948
rect 4604 94836 4614 94892
rect 4670 94836 4718 94892
rect 4774 94836 4822 94892
rect 4878 94836 4888 94892
rect 11408 94836 11418 94892
rect 11474 94836 11522 94892
rect 11578 94836 11626 94892
rect 11682 94836 11692 94892
rect 5170 94780 5180 94836
rect 5236 94780 6636 94836
rect 6692 94780 6860 94836
rect 6916 94780 7196 94836
rect 7252 94780 7644 94836
rect 7700 94780 7710 94836
rect 13682 94780 13692 94836
rect 13748 94780 14924 94836
rect 14980 94780 14990 94836
rect 15092 94724 15148 94892
rect 18212 94836 18222 94892
rect 18278 94836 18326 94892
rect 18382 94836 18430 94892
rect 18486 94836 18496 94892
rect 25016 94836 25026 94892
rect 25082 94836 25130 94892
rect 25186 94836 25234 94892
rect 25290 94836 25300 94892
rect 4834 94668 4844 94724
rect 4900 94668 6748 94724
rect 6804 94668 6814 94724
rect 8082 94668 8092 94724
rect 8148 94668 10780 94724
rect 10836 94668 15148 94724
rect 18386 94668 18396 94724
rect 18452 94668 19516 94724
rect 19572 94668 19582 94724
rect 19730 94668 19740 94724
rect 19796 94668 19834 94724
rect 3042 94556 3052 94612
rect 3108 94556 3724 94612
rect 3780 94556 5740 94612
rect 5796 94556 6524 94612
rect 6580 94556 11676 94612
rect 11732 94556 20972 94612
rect 21028 94556 21038 94612
rect 10658 94444 10668 94500
rect 10724 94444 11340 94500
rect 11396 94444 14700 94500
rect 14756 94444 14766 94500
rect 15026 94444 15036 94500
rect 15092 94444 15932 94500
rect 15988 94444 15998 94500
rect 16146 94444 16156 94500
rect 16212 94444 18172 94500
rect 18228 94444 19068 94500
rect 19124 94444 19134 94500
rect 7074 94332 7084 94388
rect 7140 94332 11228 94388
rect 11284 94332 11294 94388
rect 13906 94332 13916 94388
rect 13972 94332 18060 94388
rect 18116 94332 18126 94388
rect 19170 94332 19180 94388
rect 19236 94332 19740 94388
rect 19796 94332 19806 94388
rect 21858 94332 21868 94388
rect 21924 94332 22036 94388
rect 4050 94220 4060 94276
rect 4116 94220 7308 94276
rect 7364 94220 7532 94276
rect 7588 94220 8540 94276
rect 8596 94220 8606 94276
rect 14914 94220 14924 94276
rect 14980 94220 15372 94276
rect 15428 94220 15438 94276
rect 16034 94220 16044 94276
rect 16100 94220 17164 94276
rect 17220 94220 17230 94276
rect 19740 94220 21756 94276
rect 21812 94220 21822 94276
rect 15372 94164 15428 94220
rect 19740 94164 19796 94220
rect 6178 94108 6188 94164
rect 6244 94108 6636 94164
rect 6692 94108 7084 94164
rect 7140 94108 7150 94164
rect 13906 94108 13916 94164
rect 13972 94108 14364 94164
rect 14420 94108 14430 94164
rect 15372 94108 16660 94164
rect 18610 94108 18620 94164
rect 18676 94108 19740 94164
rect 19796 94108 19806 94164
rect 8006 94052 8016 94108
rect 8072 94052 8120 94108
rect 8176 94052 8224 94108
rect 8280 94052 8290 94108
rect 14810 94052 14820 94108
rect 14876 94052 14924 94108
rect 14980 94052 15028 94108
rect 15084 94052 15094 94108
rect 16604 94052 16660 94108
rect 21614 94052 21624 94108
rect 21680 94052 21728 94108
rect 21784 94052 21832 94108
rect 21888 94052 21898 94108
rect 2482 93996 2492 94052
rect 2548 93996 3276 94052
rect 3332 93828 3388 94052
rect 15250 93996 15260 94052
rect 15316 93996 16380 94052
rect 16436 93996 16446 94052
rect 16604 93996 17500 94052
rect 17556 93996 17566 94052
rect 21980 93940 22036 94332
rect 25890 94108 25900 94164
rect 25956 94108 26908 94164
rect 26964 94108 26974 94164
rect 28418 94052 28428 94108
rect 28484 94052 28532 94108
rect 28588 94052 28636 94108
rect 28692 94052 28702 94108
rect 6066 93884 6076 93940
rect 6132 93884 6412 93940
rect 6468 93884 6478 93940
rect 8306 93884 8316 93940
rect 8372 93884 9996 93940
rect 10052 93884 10444 93940
rect 10500 93884 11116 93940
rect 11172 93884 11182 93940
rect 14578 93884 14588 93940
rect 14644 93884 15596 93940
rect 15652 93884 15662 93940
rect 20738 93884 20748 93940
rect 20804 93884 21644 93940
rect 21700 93884 21710 93940
rect 21970 93884 21980 93940
rect 22036 93884 22046 93940
rect 22418 93884 22428 93940
rect 22484 93884 22494 93940
rect 3332 93772 8260 93828
rect 10322 93772 10332 93828
rect 10388 93772 13468 93828
rect 13524 93772 13534 93828
rect 14252 93772 15260 93828
rect 15316 93772 15326 93828
rect 15922 93772 15932 93828
rect 15988 93772 21308 93828
rect 21364 93772 21756 93828
rect 21812 93772 21822 93828
rect 8204 93604 8260 93772
rect 10332 93716 10388 93772
rect 14252 93716 14308 93772
rect 22428 93716 22484 93884
rect 8754 93660 8764 93716
rect 8820 93660 10388 93716
rect 12450 93660 12460 93716
rect 12516 93660 13132 93716
rect 13188 93660 13692 93716
rect 13748 93660 13758 93716
rect 14242 93660 14252 93716
rect 14308 93660 14318 93716
rect 15372 93660 15876 93716
rect 16370 93660 16380 93716
rect 16436 93660 17612 93716
rect 17668 93660 17678 93716
rect 17836 93660 20356 93716
rect 20486 93660 20524 93716
rect 20580 93660 22484 93716
rect 15372 93604 15428 93660
rect 3042 93548 3052 93604
rect 3108 93548 3836 93604
rect 3892 93548 3902 93604
rect 4498 93548 4508 93604
rect 4564 93548 5292 93604
rect 5348 93548 5358 93604
rect 5506 93548 5516 93604
rect 5572 93548 6188 93604
rect 6244 93548 6254 93604
rect 8204 93548 15428 93604
rect 15820 93604 15876 93660
rect 17836 93604 17892 93660
rect 20300 93604 20356 93660
rect 15820 93548 17892 93604
rect 18050 93548 18060 93604
rect 18116 93548 19068 93604
rect 19124 93548 19134 93604
rect 20290 93548 20300 93604
rect 20356 93548 23100 93604
rect 23156 93548 23166 93604
rect 0 93492 400 93520
rect 0 93436 1708 93492
rect 1764 93436 3500 93492
rect 3556 93436 3566 93492
rect 6076 93436 6412 93492
rect 6468 93436 9548 93492
rect 9604 93436 9614 93492
rect 9874 93436 9884 93492
rect 9940 93436 11844 93492
rect 12114 93436 12124 93492
rect 12180 93436 13356 93492
rect 13412 93436 13422 93492
rect 14018 93436 14028 93492
rect 14084 93436 15932 93492
rect 15988 93436 16492 93492
rect 16548 93436 18508 93492
rect 18564 93436 18574 93492
rect 0 93408 400 93436
rect 6076 93380 6132 93436
rect 6066 93324 6076 93380
rect 6132 93324 6142 93380
rect 4604 93268 4614 93324
rect 4670 93268 4718 93324
rect 4774 93268 4822 93324
rect 4878 93268 4888 93324
rect 11408 93268 11418 93324
rect 11474 93268 11522 93324
rect 11578 93268 11626 93324
rect 11682 93268 11692 93324
rect 11788 93156 11844 93436
rect 18212 93268 18222 93324
rect 18278 93268 18326 93324
rect 18382 93268 18430 93324
rect 18486 93268 18496 93324
rect 25016 93268 25026 93324
rect 25082 93268 25130 93324
rect 25186 93268 25234 93324
rect 25290 93268 25300 93324
rect 13794 93212 13804 93268
rect 13860 93212 14476 93268
rect 14532 93212 14542 93268
rect 15558 93212 15596 93268
rect 15652 93212 15662 93268
rect 17602 93212 17612 93268
rect 17668 93212 18060 93268
rect 18116 93212 18126 93268
rect 10994 93100 11004 93156
rect 11060 93100 11564 93156
rect 11620 93100 11630 93156
rect 11788 93100 18452 93156
rect 5170 92988 5180 93044
rect 5236 92988 6524 93044
rect 6580 92988 9884 93044
rect 9940 92988 9950 93044
rect 10322 92988 10332 93044
rect 10388 92988 11340 93044
rect 11396 92988 16156 93044
rect 16212 92988 16222 93044
rect 18396 92932 18452 93100
rect 25218 92988 25228 93044
rect 25284 92988 26124 93044
rect 26180 92988 26190 93044
rect 6962 92876 6972 92932
rect 7028 92876 8316 92932
rect 8372 92876 8382 92932
rect 17266 92876 17276 92932
rect 17332 92876 18340 92932
rect 18396 92876 18956 92932
rect 19012 92876 19180 92932
rect 19236 92876 19852 92932
rect 19908 92876 19918 92932
rect 25778 92876 25788 92932
rect 25844 92876 25854 92932
rect 26338 92876 26348 92932
rect 26404 92876 26414 92932
rect 18284 92820 18340 92876
rect 13346 92764 13356 92820
rect 13412 92764 14364 92820
rect 14420 92764 14430 92820
rect 15922 92764 15932 92820
rect 15988 92764 16380 92820
rect 16436 92764 16446 92820
rect 16930 92764 16940 92820
rect 16996 92764 17948 92820
rect 18004 92764 18014 92820
rect 18284 92764 18620 92820
rect 18676 92764 18686 92820
rect 20850 92764 20860 92820
rect 20916 92764 21532 92820
rect 21588 92764 21598 92820
rect 22530 92764 22540 92820
rect 22596 92764 23324 92820
rect 23380 92764 23390 92820
rect 25788 92708 25844 92876
rect 11890 92652 11900 92708
rect 11956 92652 17164 92708
rect 17220 92652 17230 92708
rect 20150 92652 20188 92708
rect 20244 92652 20254 92708
rect 20626 92652 20636 92708
rect 20692 92652 23772 92708
rect 23828 92652 23838 92708
rect 25788 92652 26012 92708
rect 26068 92652 26078 92708
rect 17164 92596 17220 92652
rect 16818 92540 16828 92596
rect 16884 92540 17220 92596
rect 8006 92484 8016 92540
rect 8072 92484 8120 92540
rect 8176 92484 8224 92540
rect 8280 92484 8290 92540
rect 14810 92484 14820 92540
rect 14876 92484 14924 92540
rect 14980 92484 15028 92540
rect 15084 92484 15094 92540
rect 21614 92484 21624 92540
rect 21680 92484 21728 92540
rect 21784 92484 21832 92540
rect 21888 92484 21898 92540
rect 26348 92484 26404 92876
rect 26562 92652 26572 92708
rect 26628 92652 26638 92708
rect 14018 92428 14028 92484
rect 14084 92428 14094 92484
rect 16146 92428 16156 92484
rect 16212 92428 17164 92484
rect 17220 92428 17230 92484
rect 19394 92428 19404 92484
rect 19460 92428 19740 92484
rect 19796 92428 20748 92484
rect 20804 92428 20814 92484
rect 25778 92428 25788 92484
rect 25844 92428 26404 92484
rect 14028 92372 14084 92428
rect 26572 92372 26628 92652
rect 28418 92484 28428 92540
rect 28484 92484 28532 92540
rect 28588 92484 28636 92540
rect 28692 92484 28702 92540
rect 27010 92428 27020 92484
rect 27076 92428 27086 92484
rect 2930 92316 2940 92372
rect 2996 92316 4284 92372
rect 4340 92316 4350 92372
rect 8978 92316 8988 92372
rect 9044 92316 10220 92372
rect 10276 92316 10286 92372
rect 10882 92316 10892 92372
rect 10948 92316 12348 92372
rect 12404 92316 12414 92372
rect 12786 92316 12796 92372
rect 12852 92316 15148 92372
rect 17798 92316 17836 92372
rect 17892 92316 17902 92372
rect 18498 92316 18508 92372
rect 18564 92316 19628 92372
rect 19684 92316 19694 92372
rect 23538 92316 23548 92372
rect 23604 92316 24332 92372
rect 24388 92316 25452 92372
rect 25508 92316 26628 92372
rect 2482 92204 2492 92260
rect 2548 92204 3276 92260
rect 3332 92204 5404 92260
rect 5460 92204 5852 92260
rect 5908 92204 5918 92260
rect 7522 92204 7532 92260
rect 7588 92204 9772 92260
rect 9828 92204 10444 92260
rect 10500 92204 10510 92260
rect 13570 92204 13580 92260
rect 13636 92204 14588 92260
rect 14644 92204 14654 92260
rect 15092 92148 15148 92316
rect 20290 92204 20300 92260
rect 20356 92204 21196 92260
rect 21252 92204 21262 92260
rect 22082 92204 22092 92260
rect 22148 92204 22316 92260
rect 22372 92204 23100 92260
rect 23156 92204 25228 92260
rect 25284 92204 25294 92260
rect 15092 92092 15596 92148
rect 15652 92092 17500 92148
rect 17556 92092 17566 92148
rect 22418 92092 22428 92148
rect 22484 92092 22876 92148
rect 22932 92092 24388 92148
rect 24658 92092 24668 92148
rect 24724 92092 25788 92148
rect 25844 92092 25854 92148
rect 24332 92036 24388 92092
rect 1810 91980 1820 92036
rect 1876 91980 2828 92036
rect 2884 91980 4620 92036
rect 4676 91980 4686 92036
rect 14354 91980 14364 92036
rect 14420 91980 15484 92036
rect 15540 91980 15932 92036
rect 15988 91980 15998 92036
rect 18834 91980 18844 92036
rect 18900 91980 19292 92036
rect 19348 91980 19358 92036
rect 22642 91980 22652 92036
rect 22708 91980 23436 92036
rect 23492 91980 23502 92036
rect 24322 91980 24332 92036
rect 24388 91980 26012 92036
rect 26068 91980 26908 92036
rect 26852 91924 26908 91980
rect 27020 91924 27076 92428
rect 19170 91868 19180 91924
rect 19236 91868 26684 91924
rect 26740 91868 26750 91924
rect 26852 91868 27076 91924
rect 18946 91756 18956 91812
rect 19012 91756 19022 91812
rect 26460 91756 26908 91812
rect 26964 91756 26974 91812
rect 4604 91700 4614 91756
rect 4670 91700 4718 91756
rect 4774 91700 4822 91756
rect 4878 91700 4888 91756
rect 11408 91700 11418 91756
rect 11474 91700 11522 91756
rect 11578 91700 11626 91756
rect 11682 91700 11692 91756
rect 18212 91700 18222 91756
rect 18278 91700 18326 91756
rect 18382 91700 18430 91756
rect 18486 91700 18496 91756
rect 18956 91588 19012 91756
rect 25016 91700 25026 91756
rect 25082 91700 25130 91756
rect 25186 91700 25234 91756
rect 25290 91700 25300 91756
rect 22950 91644 22988 91700
rect 23044 91644 23054 91700
rect 25526 91644 25564 91700
rect 25620 91644 25630 91700
rect 26460 91588 26516 91756
rect 3378 91532 3388 91588
rect 3444 91532 5740 91588
rect 5796 91532 5806 91588
rect 12674 91532 12684 91588
rect 12740 91532 14252 91588
rect 14308 91532 14318 91588
rect 14578 91532 14588 91588
rect 14644 91532 16268 91588
rect 16324 91532 16334 91588
rect 17826 91532 17836 91588
rect 17892 91532 19012 91588
rect 22838 91532 22876 91588
rect 22932 91532 22942 91588
rect 23874 91532 23884 91588
rect 23940 91532 25228 91588
rect 25284 91532 25294 91588
rect 25666 91532 25676 91588
rect 25732 91532 26460 91588
rect 26516 91532 26526 91588
rect 26852 91532 28140 91588
rect 28196 91532 28206 91588
rect 18956 91476 19012 91532
rect 26852 91476 26908 91532
rect 6066 91420 6076 91476
rect 6132 91420 7308 91476
rect 7364 91420 7374 91476
rect 12898 91420 12908 91476
rect 12964 91420 13580 91476
rect 13636 91420 15372 91476
rect 15428 91420 15438 91476
rect 18956 91420 26908 91476
rect 15474 91308 15484 91364
rect 15540 91308 16828 91364
rect 16884 91308 16894 91364
rect 21970 91308 21980 91364
rect 22036 91308 22316 91364
rect 22372 91308 23548 91364
rect 23604 91308 23614 91364
rect 25554 91308 25564 91364
rect 25620 91308 25788 91364
rect 25844 91308 26908 91364
rect 26964 91308 26974 91364
rect 13682 91196 13692 91252
rect 13748 91196 15708 91252
rect 15764 91196 15774 91252
rect 18946 91196 18956 91252
rect 19012 91196 19628 91252
rect 19684 91196 20300 91252
rect 20356 91196 20366 91252
rect 22530 91196 22540 91252
rect 22596 91196 23772 91252
rect 23828 91196 23838 91252
rect 24546 91196 24556 91252
rect 24612 91196 26012 91252
rect 26068 91196 26078 91252
rect 5058 91084 5068 91140
rect 5124 91084 6748 91140
rect 6804 91084 7420 91140
rect 7476 91084 7486 91140
rect 14690 91084 14700 91140
rect 14756 91084 15540 91140
rect 22418 91084 22428 91140
rect 22484 91084 22764 91140
rect 22820 91084 22830 91140
rect 23426 91084 23436 91140
rect 23492 91084 24332 91140
rect 24388 91084 25676 91140
rect 25732 91084 25742 91140
rect 26852 91084 27132 91140
rect 27188 91084 27198 91140
rect 8006 90916 8016 90972
rect 8072 90916 8120 90972
rect 8176 90916 8224 90972
rect 8280 90916 8290 90972
rect 14810 90916 14820 90972
rect 14876 90916 14924 90972
rect 14980 90916 15028 90972
rect 15084 90916 15094 90972
rect 0 90804 400 90832
rect 15484 90804 15540 91084
rect 26852 91028 26908 91084
rect 24210 90972 24220 91028
rect 24276 90972 26012 91028
rect 26068 90972 26908 91028
rect 21614 90916 21624 90972
rect 21680 90916 21728 90972
rect 21784 90916 21832 90972
rect 21888 90916 21898 90972
rect 28418 90916 28428 90972
rect 28484 90916 28532 90972
rect 28588 90916 28636 90972
rect 28692 90916 28702 90972
rect 22866 90860 22876 90916
rect 22932 90860 23212 90916
rect 23268 90860 23278 90916
rect 23538 90860 23548 90916
rect 23604 90860 23884 90916
rect 23940 90860 23950 90916
rect 0 90748 1764 90804
rect 5282 90748 5292 90804
rect 5348 90748 6524 90804
rect 6580 90748 7196 90804
rect 7252 90748 7812 90804
rect 8418 90748 8428 90804
rect 8484 90748 9660 90804
rect 9716 90748 10108 90804
rect 10164 90748 10556 90804
rect 10612 90748 11452 90804
rect 11508 90748 13468 90804
rect 13524 90748 13534 90804
rect 15474 90748 15484 90804
rect 15540 90748 15550 90804
rect 19394 90748 19404 90804
rect 19460 90748 19964 90804
rect 20020 90748 20030 90804
rect 22082 90748 22092 90804
rect 22148 90748 25116 90804
rect 25172 90748 25182 90804
rect 0 90720 400 90748
rect 1708 90580 1764 90748
rect 5292 90692 5348 90748
rect 7756 90692 7812 90748
rect 4498 90636 4508 90692
rect 4564 90636 5348 90692
rect 5730 90636 5740 90692
rect 5796 90636 7532 90692
rect 7588 90636 7598 90692
rect 7756 90636 8764 90692
rect 8820 90636 8830 90692
rect 8988 90636 10892 90692
rect 10948 90636 10958 90692
rect 12002 90636 12012 90692
rect 12068 90636 14924 90692
rect 14980 90636 14990 90692
rect 17724 90636 20860 90692
rect 20916 90636 20926 90692
rect 23426 90636 23436 90692
rect 23492 90636 23548 90748
rect 8988 90580 9044 90636
rect 17724 90580 17780 90636
rect 1698 90524 1708 90580
rect 1764 90524 1774 90580
rect 8866 90524 8876 90580
rect 8932 90524 9044 90580
rect 9202 90524 9212 90580
rect 9268 90524 9772 90580
rect 9828 90524 9838 90580
rect 10434 90524 10444 90580
rect 10500 90524 11228 90580
rect 11284 90524 11900 90580
rect 11956 90524 11966 90580
rect 12674 90524 12684 90580
rect 12740 90524 13356 90580
rect 13412 90524 13422 90580
rect 15138 90524 15148 90580
rect 15204 90524 17780 90580
rect 18162 90524 18172 90580
rect 18228 90524 18844 90580
rect 18900 90524 19740 90580
rect 19796 90524 21308 90580
rect 21364 90524 21374 90580
rect 26338 90524 26348 90580
rect 26404 90524 27580 90580
rect 27636 90524 27646 90580
rect 8082 90412 8092 90468
rect 8148 90412 9884 90468
rect 9940 90412 12012 90468
rect 12068 90412 12078 90468
rect 15362 90412 15372 90468
rect 15428 90412 16380 90468
rect 16436 90412 16604 90468
rect 16660 90412 17948 90468
rect 18004 90412 18014 90468
rect 20188 90356 20244 90524
rect 20402 90412 20412 90468
rect 20468 90412 20860 90468
rect 20916 90412 20926 90468
rect 25778 90412 25788 90468
rect 25844 90412 28028 90468
rect 28084 90412 28094 90468
rect 20178 90300 20188 90356
rect 20244 90300 20254 90356
rect 22642 90300 22652 90356
rect 22708 90300 23212 90356
rect 23268 90300 23278 90356
rect 4604 90132 4614 90188
rect 4670 90132 4718 90188
rect 4774 90132 4822 90188
rect 4878 90132 4888 90188
rect 11408 90132 11418 90188
rect 11474 90132 11522 90188
rect 11578 90132 11626 90188
rect 11682 90132 11692 90188
rect 18212 90132 18222 90188
rect 18278 90132 18326 90188
rect 18382 90132 18430 90188
rect 18486 90132 18496 90188
rect 25016 90132 25026 90188
rect 25082 90132 25130 90188
rect 25186 90132 25234 90188
rect 25290 90132 25300 90188
rect 12898 89964 12908 90020
rect 12964 89964 13468 90020
rect 13524 89964 15708 90020
rect 15764 89964 16828 90020
rect 16884 89964 16894 90020
rect 17378 89964 17388 90020
rect 17444 89964 18508 90020
rect 18564 89964 18574 90020
rect 22838 89964 22876 90020
rect 22932 89964 22942 90020
rect 9538 89852 9548 89908
rect 9604 89852 10332 89908
rect 10388 89852 10398 89908
rect 13570 89852 13580 89908
rect 13636 89852 14588 89908
rect 14644 89852 14654 89908
rect 15026 89852 15036 89908
rect 15092 89852 17052 89908
rect 17108 89852 17118 89908
rect 21746 89852 21756 89908
rect 21812 89852 22764 89908
rect 22820 89852 22830 89908
rect 11778 89740 11788 89796
rect 11844 89740 12684 89796
rect 12740 89740 13804 89796
rect 13860 89740 13870 89796
rect 17714 89740 17724 89796
rect 17780 89740 26908 89796
rect 26852 89684 26908 89740
rect 14018 89628 14028 89684
rect 14084 89628 15260 89684
rect 15316 89628 15326 89684
rect 16156 89628 17612 89684
rect 17668 89628 17678 89684
rect 17938 89628 17948 89684
rect 18004 89628 18396 89684
rect 18452 89628 18462 89684
rect 19954 89628 19964 89684
rect 20020 89628 21868 89684
rect 21924 89628 21934 89684
rect 22754 89628 22764 89684
rect 22820 89628 25788 89684
rect 25844 89628 25854 89684
rect 26852 89628 27020 89684
rect 27076 89628 27086 89684
rect 16156 89572 16212 89628
rect 13682 89516 13692 89572
rect 13748 89516 14812 89572
rect 14868 89516 16212 89572
rect 16370 89516 16380 89572
rect 16436 89516 18060 89572
rect 18116 89516 18126 89572
rect 22194 89516 22204 89572
rect 22260 89516 23324 89572
rect 23380 89516 23390 89572
rect 25554 89516 25564 89572
rect 25620 89516 26012 89572
rect 26068 89516 26078 89572
rect 21970 89404 21980 89460
rect 22036 89404 25116 89460
rect 25172 89404 25182 89460
rect 8006 89348 8016 89404
rect 8072 89348 8120 89404
rect 8176 89348 8224 89404
rect 8280 89348 8290 89404
rect 14810 89348 14820 89404
rect 14876 89348 14924 89404
rect 14980 89348 15028 89404
rect 15084 89348 15094 89404
rect 21614 89348 21624 89404
rect 21680 89348 21728 89404
rect 21784 89348 21832 89404
rect 21888 89348 21898 89404
rect 28418 89348 28428 89404
rect 28484 89348 28532 89404
rect 28588 89348 28636 89404
rect 28692 89348 28702 89404
rect 16706 89292 16716 89348
rect 16772 89292 17500 89348
rect 17556 89292 19628 89348
rect 19684 89292 19694 89348
rect 22978 89292 22988 89348
rect 23044 89292 23324 89348
rect 23380 89292 24220 89348
rect 24276 89292 24286 89348
rect 6514 89180 6524 89236
rect 6580 89180 6860 89236
rect 6916 89180 7756 89236
rect 7812 89180 7822 89236
rect 15362 89180 15372 89236
rect 15428 89180 15820 89236
rect 15876 89180 15886 89236
rect 18274 89180 18284 89236
rect 18340 89180 18620 89236
rect 18676 89180 18686 89236
rect 22866 89180 22876 89236
rect 22932 89180 22988 89236
rect 23044 89180 23054 89236
rect 23202 89180 23212 89236
rect 23268 89180 24556 89236
rect 24612 89180 24622 89236
rect 15670 89068 15708 89124
rect 15764 89068 15774 89124
rect 17938 89068 17948 89124
rect 18004 89068 24108 89124
rect 24164 89068 24174 89124
rect 6402 88956 6412 89012
rect 6468 88956 7196 89012
rect 7252 88956 7262 89012
rect 7634 88956 7644 89012
rect 7700 88956 10108 89012
rect 10164 88956 10174 89012
rect 14690 88956 14700 89012
rect 14756 88956 16156 89012
rect 16212 88956 16222 89012
rect 16818 88956 16828 89012
rect 16884 88956 19292 89012
rect 19348 88956 19358 89012
rect 21410 88956 21420 89012
rect 21476 88956 22652 89012
rect 22708 88956 22718 89012
rect 23538 88956 23548 89012
rect 23604 88956 23828 89012
rect 23986 88956 23996 89012
rect 24052 88956 25340 89012
rect 25396 88956 25406 89012
rect 16828 88900 16884 88956
rect 23772 88900 23828 88956
rect 2482 88844 2492 88900
rect 2548 88844 3836 88900
rect 3892 88844 3902 88900
rect 6066 88844 6076 88900
rect 6132 88844 8092 88900
rect 8148 88844 8158 88900
rect 11106 88844 11116 88900
rect 11172 88844 13356 88900
rect 13412 88844 13422 88900
rect 13794 88844 13804 88900
rect 13860 88844 15372 88900
rect 15428 88844 16884 88900
rect 18386 88844 18396 88900
rect 18452 88844 19964 88900
rect 20020 88844 20030 88900
rect 20738 88844 20748 88900
rect 20804 88844 21532 88900
rect 21588 88844 21598 88900
rect 23772 88844 24332 88900
rect 24388 88844 24398 88900
rect 24546 88844 24556 88900
rect 24612 88844 25564 88900
rect 25620 88844 25630 88900
rect 9426 88732 9436 88788
rect 9492 88732 15148 88788
rect 15204 88732 15214 88788
rect 18946 88732 18956 88788
rect 19012 88732 19628 88788
rect 19684 88732 19740 88788
rect 19796 88732 19806 88788
rect 4604 88564 4614 88620
rect 4670 88564 4718 88620
rect 4774 88564 4822 88620
rect 4878 88564 4888 88620
rect 11408 88564 11418 88620
rect 11474 88564 11522 88620
rect 11578 88564 11626 88620
rect 11682 88564 11692 88620
rect 18212 88564 18222 88620
rect 18278 88564 18326 88620
rect 18382 88564 18430 88620
rect 18486 88564 18496 88620
rect 25016 88564 25026 88620
rect 25082 88564 25130 88620
rect 25186 88564 25234 88620
rect 25290 88564 25300 88620
rect 9090 88396 9100 88452
rect 9156 88396 14028 88452
rect 14084 88396 14094 88452
rect 24322 88396 24332 88452
rect 24388 88396 24780 88452
rect 24836 88396 24846 88452
rect 5058 88284 5068 88340
rect 5124 88284 5740 88340
rect 5796 88284 5806 88340
rect 20066 88284 20076 88340
rect 20132 88284 20524 88340
rect 20580 88284 20590 88340
rect 12898 88172 12908 88228
rect 12964 88172 13468 88228
rect 13524 88172 13534 88228
rect 16034 88172 16044 88228
rect 16100 88172 16604 88228
rect 16660 88172 16670 88228
rect 19282 88172 19292 88228
rect 19348 88172 24556 88228
rect 24612 88172 24622 88228
rect 26786 88172 26796 88228
rect 26852 88172 27580 88228
rect 27636 88172 27646 88228
rect 0 88116 400 88144
rect 0 88060 1708 88116
rect 1764 88060 1774 88116
rect 7746 88060 7756 88116
rect 7812 88060 9212 88116
rect 9268 88060 12348 88116
rect 12404 88060 13244 88116
rect 13300 88060 13310 88116
rect 15446 88060 15484 88116
rect 15540 88060 15550 88116
rect 16706 88060 16716 88116
rect 16772 88060 17724 88116
rect 17780 88060 17790 88116
rect 18050 88060 18060 88116
rect 18116 88060 18508 88116
rect 18564 88060 19180 88116
rect 19236 88060 19246 88116
rect 24098 88060 24108 88116
rect 24164 88060 25004 88116
rect 25060 88060 27132 88116
rect 27188 88060 27198 88116
rect 0 88032 400 88060
rect 2818 87948 2828 88004
rect 2884 87948 3388 88004
rect 3444 87948 3482 88004
rect 7970 87948 7980 88004
rect 8036 87948 8876 88004
rect 8932 87948 8942 88004
rect 17602 87948 17612 88004
rect 17668 87948 17836 88004
rect 17892 87948 17902 88004
rect 17042 87836 17052 87892
rect 17108 87836 18620 87892
rect 18676 87836 20412 87892
rect 20468 87836 20478 87892
rect 8006 87780 8016 87836
rect 8072 87780 8120 87836
rect 8176 87780 8224 87836
rect 8280 87780 8290 87836
rect 14810 87780 14820 87836
rect 14876 87780 14924 87836
rect 14980 87780 15028 87836
rect 15084 87780 15094 87836
rect 21614 87780 21624 87836
rect 21680 87780 21728 87836
rect 21784 87780 21832 87836
rect 21888 87780 21898 87836
rect 28418 87780 28428 87836
rect 28484 87780 28532 87836
rect 28588 87780 28636 87836
rect 28692 87780 28702 87836
rect 16604 87724 18844 87780
rect 18900 87724 18910 87780
rect 16604 87668 16660 87724
rect 14690 87612 14700 87668
rect 14756 87612 14766 87668
rect 15474 87612 15484 87668
rect 15540 87612 15596 87668
rect 15652 87612 16604 87668
rect 16660 87612 16670 87668
rect 17490 87612 17500 87668
rect 17556 87612 19404 87668
rect 19460 87612 19470 87668
rect 14700 87556 14756 87612
rect 2034 87500 2044 87556
rect 2100 87500 5292 87556
rect 5348 87500 5358 87556
rect 13010 87500 13020 87556
rect 13076 87500 13804 87556
rect 13860 87500 15036 87556
rect 15092 87500 15102 87556
rect 17500 87444 17556 87612
rect 3042 87388 3052 87444
rect 3108 87388 5068 87444
rect 5124 87388 5134 87444
rect 6738 87388 6748 87444
rect 6804 87388 17556 87444
rect 25778 87388 25788 87444
rect 25844 87388 26460 87444
rect 26516 87388 26526 87444
rect 7858 87276 7868 87332
rect 7924 87276 9660 87332
rect 9716 87276 10108 87332
rect 10164 87276 10174 87332
rect 13906 87276 13916 87332
rect 13972 87276 14252 87332
rect 14308 87276 14318 87332
rect 17266 87276 17276 87332
rect 17332 87276 17836 87332
rect 17892 87276 17902 87332
rect 24434 87276 24444 87332
rect 24500 87276 25564 87332
rect 25620 87276 25630 87332
rect 26338 87276 26348 87332
rect 26404 87276 27468 87332
rect 27524 87276 27534 87332
rect 13234 87164 13244 87220
rect 13300 87164 15036 87220
rect 15092 87164 18676 87220
rect 24882 87164 24892 87220
rect 24948 87164 26908 87220
rect 26964 87164 26974 87220
rect 18620 87108 18676 87164
rect 18620 87052 20300 87108
rect 20356 87052 20366 87108
rect 26002 87052 26012 87108
rect 26068 87052 26796 87108
rect 26852 87052 26862 87108
rect 4604 86996 4614 87052
rect 4670 86996 4718 87052
rect 4774 86996 4822 87052
rect 4878 86996 4888 87052
rect 11408 86996 11418 87052
rect 11474 86996 11522 87052
rect 11578 86996 11626 87052
rect 11682 86996 11692 87052
rect 18212 86996 18222 87052
rect 18278 86996 18326 87052
rect 18382 86996 18430 87052
rect 18486 86996 18496 87052
rect 25016 86996 25026 87052
rect 25082 86996 25130 87052
rect 25186 86996 25234 87052
rect 25290 86996 25300 87052
rect 15362 86828 15372 86884
rect 15428 86828 15438 86884
rect 16482 86828 16492 86884
rect 16548 86828 17948 86884
rect 18004 86828 18956 86884
rect 19012 86828 19022 86884
rect 22754 86828 22764 86884
rect 22820 86828 23996 86884
rect 24052 86828 24062 86884
rect 15372 86772 15428 86828
rect 6514 86716 6524 86772
rect 6580 86716 8988 86772
rect 9044 86716 9054 86772
rect 10098 86716 10108 86772
rect 10164 86716 11228 86772
rect 11284 86716 11294 86772
rect 15026 86716 15036 86772
rect 15092 86716 15428 86772
rect 24322 86716 24332 86772
rect 24388 86716 27692 86772
rect 27748 86716 27758 86772
rect 7522 86604 7532 86660
rect 7588 86604 12236 86660
rect 12292 86604 12302 86660
rect 18610 86604 18620 86660
rect 18676 86604 19180 86660
rect 19236 86604 21084 86660
rect 21140 86604 21150 86660
rect 23538 86604 23548 86660
rect 23604 86604 27244 86660
rect 27300 86604 27310 86660
rect 9202 86492 9212 86548
rect 9268 86492 10892 86548
rect 10948 86492 10958 86548
rect 20188 86492 21196 86548
rect 21252 86492 21980 86548
rect 22036 86492 22876 86548
rect 22932 86492 22942 86548
rect 20188 86436 20244 86492
rect 8642 86380 8652 86436
rect 8708 86380 8988 86436
rect 9044 86380 9548 86436
rect 9604 86380 10780 86436
rect 10836 86380 10846 86436
rect 15026 86380 15036 86436
rect 15092 86380 20188 86436
rect 20244 86380 20254 86436
rect 21522 86380 21532 86436
rect 21588 86380 23884 86436
rect 23940 86380 23950 86436
rect 15446 86268 15484 86324
rect 15540 86268 15550 86324
rect 19954 86268 19964 86324
rect 20020 86268 20748 86324
rect 20804 86268 20814 86324
rect 8006 86212 8016 86268
rect 8072 86212 8120 86268
rect 8176 86212 8224 86268
rect 8280 86212 8290 86268
rect 14810 86212 14820 86268
rect 14876 86212 14924 86268
rect 14980 86212 15028 86268
rect 15084 86212 15094 86268
rect 21614 86212 21624 86268
rect 21680 86212 21728 86268
rect 21784 86212 21832 86268
rect 21888 86212 21898 86268
rect 28418 86212 28428 86268
rect 28484 86212 28532 86268
rect 28588 86212 28636 86268
rect 28692 86212 28702 86268
rect 7298 86044 7308 86100
rect 7364 86044 9772 86100
rect 9828 86044 9838 86100
rect 24994 86044 25004 86100
rect 25060 86044 25788 86100
rect 25844 86044 25854 86100
rect 2034 85932 2044 85988
rect 2100 85932 7084 85988
rect 7140 85932 7150 85988
rect 8642 85932 8652 85988
rect 8708 85932 9660 85988
rect 9716 85932 9726 85988
rect 13570 85932 13580 85988
rect 13636 85932 15708 85988
rect 15764 85932 15932 85988
rect 15988 85932 17276 85988
rect 17332 85932 17342 85988
rect 7746 85820 7756 85876
rect 7812 85820 11004 85876
rect 11060 85820 13692 85876
rect 13748 85820 15036 85876
rect 15092 85820 15102 85876
rect 18722 85820 18732 85876
rect 18788 85820 19404 85876
rect 19460 85820 19470 85876
rect 24658 85820 24668 85876
rect 24724 85820 25452 85876
rect 25508 85820 25518 85876
rect 5842 85708 5852 85764
rect 5908 85708 6972 85764
rect 7028 85708 8316 85764
rect 8372 85708 8382 85764
rect 16818 85708 16828 85764
rect 16884 85708 18172 85764
rect 18228 85708 19068 85764
rect 19124 85708 19628 85764
rect 19684 85708 19964 85764
rect 20020 85708 20030 85764
rect 24546 85708 24556 85764
rect 24612 85708 26348 85764
rect 26404 85708 26414 85764
rect 8866 85596 8876 85652
rect 8932 85596 12012 85652
rect 12068 85596 12078 85652
rect 16706 85596 16716 85652
rect 16772 85596 17052 85652
rect 17108 85596 17118 85652
rect 23986 85596 23996 85652
rect 24052 85596 25956 85652
rect 26450 85596 26460 85652
rect 26516 85596 27468 85652
rect 27524 85596 27534 85652
rect 25900 85540 25956 85596
rect 25900 85484 26796 85540
rect 26852 85484 27356 85540
rect 27412 85484 27692 85540
rect 27748 85484 27758 85540
rect 0 85428 400 85456
rect 4604 85428 4614 85484
rect 4670 85428 4718 85484
rect 4774 85428 4822 85484
rect 4878 85428 4888 85484
rect 11408 85428 11418 85484
rect 11474 85428 11522 85484
rect 11578 85428 11626 85484
rect 11682 85428 11692 85484
rect 18212 85428 18222 85484
rect 18278 85428 18326 85484
rect 18382 85428 18430 85484
rect 18486 85428 18496 85484
rect 25016 85428 25026 85484
rect 25082 85428 25130 85484
rect 25186 85428 25234 85484
rect 25290 85428 25300 85484
rect 0 85372 1708 85428
rect 1764 85372 2492 85428
rect 2548 85372 2558 85428
rect 0 85344 400 85372
rect 15474 85260 15484 85316
rect 15540 85260 16380 85316
rect 16436 85260 19180 85316
rect 19236 85260 19246 85316
rect 25442 85260 25452 85316
rect 25508 85260 26572 85316
rect 26628 85260 26638 85316
rect 24210 85148 24220 85204
rect 24276 85148 25564 85204
rect 25620 85148 28140 85204
rect 28196 85148 28206 85204
rect 3042 85036 3052 85092
rect 3108 85036 4956 85092
rect 5012 85036 5022 85092
rect 16594 85036 16604 85092
rect 16660 85036 18620 85092
rect 18676 85036 18686 85092
rect 25666 85036 25676 85092
rect 25732 85036 26124 85092
rect 26180 85036 26190 85092
rect 12786 84924 12796 84980
rect 12852 84924 14028 84980
rect 14084 84924 16156 84980
rect 16212 84924 16222 84980
rect 20514 84924 20524 84980
rect 20580 84924 21308 84980
rect 21364 84924 21374 84980
rect 26562 84924 26572 84980
rect 26628 84924 27916 84980
rect 27972 84924 27982 84980
rect 19506 84812 19516 84868
rect 19572 84812 20636 84868
rect 20692 84812 22876 84868
rect 22932 84812 22942 84868
rect 24658 84812 24668 84868
rect 24724 84812 27692 84868
rect 27748 84812 27758 84868
rect 8006 84644 8016 84700
rect 8072 84644 8120 84700
rect 8176 84644 8224 84700
rect 8280 84644 8290 84700
rect 14810 84644 14820 84700
rect 14876 84644 14924 84700
rect 14980 84644 15028 84700
rect 15084 84644 15094 84700
rect 21614 84644 21624 84700
rect 21680 84644 21728 84700
rect 21784 84644 21832 84700
rect 21888 84644 21898 84700
rect 4946 84476 4956 84532
rect 5012 84476 5740 84532
rect 5796 84476 5806 84532
rect 8978 84476 8988 84532
rect 9044 84476 10332 84532
rect 10388 84476 10398 84532
rect 10210 84364 10220 84420
rect 10276 84364 11452 84420
rect 11508 84364 14364 84420
rect 14420 84364 14430 84420
rect 14802 84364 14812 84420
rect 14868 84364 15484 84420
rect 15540 84364 15550 84420
rect 17042 84364 17052 84420
rect 17108 84364 20076 84420
rect 20132 84364 20142 84420
rect 20738 84364 20748 84420
rect 20804 84364 21308 84420
rect 21364 84364 21374 84420
rect 26012 84308 26068 84812
rect 28418 84644 28428 84700
rect 28484 84644 28532 84700
rect 28588 84644 28636 84700
rect 28692 84644 28702 84700
rect 26898 84588 26908 84644
rect 26964 84588 28140 84644
rect 28196 84588 28206 84644
rect 26226 84364 26236 84420
rect 26292 84364 27132 84420
rect 27188 84364 27198 84420
rect 9874 84252 9884 84308
rect 9940 84252 10668 84308
rect 10724 84252 11116 84308
rect 11172 84252 13804 84308
rect 13860 84252 13870 84308
rect 16258 84252 16268 84308
rect 16324 84252 17612 84308
rect 17668 84252 17678 84308
rect 20962 84252 20972 84308
rect 21028 84252 21038 84308
rect 24434 84252 24444 84308
rect 24500 84252 25564 84308
rect 25620 84252 25630 84308
rect 26012 84252 26124 84308
rect 26180 84252 26190 84308
rect 26338 84252 26348 84308
rect 26404 84252 27580 84308
rect 27636 84252 27646 84308
rect 19394 84140 19404 84196
rect 19460 84140 20748 84196
rect 20804 84140 20814 84196
rect 8754 84028 8764 84084
rect 8820 84028 10108 84084
rect 10164 84028 10174 84084
rect 18722 84028 18732 84084
rect 18788 84028 20412 84084
rect 20468 84028 20478 84084
rect 18610 83916 18620 83972
rect 18676 83916 19068 83972
rect 19124 83916 19134 83972
rect 20150 83916 20188 83972
rect 20244 83916 20254 83972
rect 4604 83860 4614 83916
rect 4670 83860 4718 83916
rect 4774 83860 4822 83916
rect 4878 83860 4888 83916
rect 11408 83860 11418 83916
rect 11474 83860 11522 83916
rect 11578 83860 11626 83916
rect 11682 83860 11692 83916
rect 18212 83860 18222 83916
rect 18278 83860 18326 83916
rect 18382 83860 18430 83916
rect 18486 83860 18496 83916
rect 20972 83748 21028 84252
rect 21756 84140 23660 84196
rect 23716 84140 23726 84196
rect 21186 84028 21196 84084
rect 21252 84028 21532 84084
rect 21588 84028 21598 84084
rect 21756 83972 21812 84140
rect 24770 84028 24780 84084
rect 24836 84028 26460 84084
rect 26516 84028 26526 84084
rect 21634 83916 21644 83972
rect 21700 83916 21812 83972
rect 22754 83916 22764 83972
rect 22820 83916 23660 83972
rect 23716 83916 23726 83972
rect 25554 83916 25564 83972
rect 25620 83916 26684 83972
rect 26740 83916 26750 83972
rect 25016 83860 25026 83916
rect 25082 83860 25130 83916
rect 25186 83860 25234 83916
rect 25290 83860 25300 83916
rect 22642 83804 22652 83860
rect 22708 83804 24220 83860
rect 24276 83804 24286 83860
rect 14924 83692 15260 83748
rect 15316 83692 15932 83748
rect 15988 83692 15998 83748
rect 20710 83692 20748 83748
rect 20804 83692 20814 83748
rect 20972 83692 23212 83748
rect 23268 83692 23278 83748
rect 14924 83524 14980 83692
rect 15586 83580 15596 83636
rect 15652 83580 16604 83636
rect 16660 83580 16670 83636
rect 18946 83580 18956 83636
rect 19012 83580 22652 83636
rect 22708 83580 22718 83636
rect 23538 83580 23548 83636
rect 23604 83580 24332 83636
rect 24388 83580 24398 83636
rect 14466 83468 14476 83524
rect 14532 83468 14542 83524
rect 14914 83468 14924 83524
rect 14980 83468 14990 83524
rect 15092 83468 15708 83524
rect 15764 83468 15774 83524
rect 18386 83468 18396 83524
rect 18452 83468 19292 83524
rect 19348 83468 19358 83524
rect 19954 83468 19964 83524
rect 20020 83468 21980 83524
rect 22036 83468 22046 83524
rect 22418 83468 22428 83524
rect 22484 83468 23772 83524
rect 23828 83468 24444 83524
rect 24500 83468 24510 83524
rect 14476 83412 14532 83468
rect 15092 83412 15148 83468
rect 1698 83356 1708 83412
rect 1764 83356 2492 83412
rect 2548 83356 2558 83412
rect 3266 83356 3276 83412
rect 3332 83356 4172 83412
rect 4228 83356 5740 83412
rect 5796 83356 5806 83412
rect 6178 83356 6188 83412
rect 6244 83356 6748 83412
rect 6804 83356 6814 83412
rect 14476 83356 15148 83412
rect 18834 83356 18844 83412
rect 18900 83356 20300 83412
rect 20356 83356 20366 83412
rect 4050 83244 4060 83300
rect 4116 83244 4620 83300
rect 4676 83244 6524 83300
rect 6580 83244 6590 83300
rect 11554 83244 11564 83300
rect 11620 83244 12572 83300
rect 12628 83244 12638 83300
rect 12786 83244 12796 83300
rect 12852 83244 13468 83300
rect 13524 83244 13534 83300
rect 16818 83244 16828 83300
rect 16884 83244 17612 83300
rect 17668 83244 17678 83300
rect 19618 83244 19628 83300
rect 19684 83244 21308 83300
rect 21364 83244 21374 83300
rect 8006 83076 8016 83132
rect 8072 83076 8120 83132
rect 8176 83076 8224 83132
rect 8280 83076 8290 83132
rect 14810 83076 14820 83132
rect 14876 83076 14924 83132
rect 14980 83076 15028 83132
rect 15084 83076 15094 83132
rect 21614 83076 21624 83132
rect 21680 83076 21728 83132
rect 21784 83076 21832 83132
rect 21888 83076 21898 83132
rect 28418 83076 28428 83132
rect 28484 83076 28532 83132
rect 28588 83076 28636 83132
rect 28692 83076 28702 83132
rect 10210 83020 10220 83076
rect 10276 83020 11228 83076
rect 11284 83020 11294 83076
rect 20822 83020 20860 83076
rect 20916 83020 20926 83076
rect 10322 82908 10332 82964
rect 10388 82908 10780 82964
rect 10836 82908 11116 82964
rect 11172 82908 12908 82964
rect 12964 82908 12974 82964
rect 15362 82908 15372 82964
rect 15428 82908 15932 82964
rect 15988 82908 17500 82964
rect 17556 82908 17566 82964
rect 4834 82796 4844 82852
rect 4900 82796 5628 82852
rect 5684 82796 5694 82852
rect 21074 82796 21084 82852
rect 21140 82796 22092 82852
rect 22148 82796 22158 82852
rect 24546 82796 24556 82852
rect 24612 82796 26236 82852
rect 26292 82796 26302 82852
rect 27990 82796 28028 82852
rect 28084 82796 28094 82852
rect 0 82740 400 82768
rect 0 82684 1708 82740
rect 1764 82684 1774 82740
rect 2034 82684 2044 82740
rect 2100 82684 3276 82740
rect 3332 82684 3342 82740
rect 15586 82684 15596 82740
rect 15652 82684 15708 82740
rect 15764 82684 16044 82740
rect 16100 82684 16716 82740
rect 16772 82684 16782 82740
rect 24658 82684 24668 82740
rect 24724 82684 26124 82740
rect 26180 82684 26190 82740
rect 26852 82684 27244 82740
rect 27300 82684 27310 82740
rect 0 82656 400 82684
rect 26852 82516 26908 82684
rect 2818 82460 2828 82516
rect 2884 82460 3388 82516
rect 3444 82460 3454 82516
rect 4050 82460 4060 82516
rect 4116 82460 4126 82516
rect 6738 82460 6748 82516
rect 6804 82460 12124 82516
rect 12180 82460 12190 82516
rect 22978 82460 22988 82516
rect 23044 82460 26908 82516
rect 4060 82292 4116 82460
rect 15810 82348 15820 82404
rect 15876 82348 17276 82404
rect 17332 82348 17342 82404
rect 4604 82292 4614 82348
rect 4670 82292 4718 82348
rect 4774 82292 4822 82348
rect 4878 82292 4888 82348
rect 11408 82292 11418 82348
rect 11474 82292 11522 82348
rect 11578 82292 11626 82348
rect 11682 82292 11692 82348
rect 18212 82292 18222 82348
rect 18278 82292 18326 82348
rect 18382 82292 18430 82348
rect 18486 82292 18496 82348
rect 18610 82292 18620 82348
rect 18676 82292 18686 82348
rect 25016 82292 25026 82348
rect 25082 82292 25130 82348
rect 25186 82292 25234 82348
rect 25290 82292 25300 82348
rect 1810 82236 1820 82292
rect 1876 82236 4116 82292
rect 18620 82236 19292 82292
rect 19348 82236 19358 82292
rect 26898 82236 26908 82292
rect 26964 82236 27468 82292
rect 27524 82236 27534 82292
rect 3042 82124 3052 82180
rect 3108 82124 3780 82180
rect 25218 82124 25228 82180
rect 25284 82124 25788 82180
rect 25844 82124 26236 82180
rect 26292 82124 27244 82180
rect 27300 82124 27310 82180
rect 3724 81956 3780 82124
rect 16370 82012 16380 82068
rect 16436 82012 16940 82068
rect 16996 82012 18396 82068
rect 18452 82012 18462 82068
rect 23762 82012 23772 82068
rect 23828 82012 24780 82068
rect 24836 82012 24846 82068
rect 2258 81900 2268 81956
rect 2324 81900 3388 81956
rect 3714 81900 3724 81956
rect 3780 81900 5684 81956
rect 7746 81900 7756 81956
rect 7812 81900 9548 81956
rect 9604 81900 9614 81956
rect 20178 81900 20188 81956
rect 20244 81900 21532 81956
rect 21588 81900 21598 81956
rect 22530 81900 22540 81956
rect 22596 81900 23212 81956
rect 23268 81900 23278 81956
rect 26338 81900 26348 81956
rect 26404 81900 26572 81956
rect 26628 81900 27468 81956
rect 27524 81900 27534 81956
rect 3332 81844 3388 81900
rect 5628 81844 5684 81900
rect 3332 81788 4844 81844
rect 4900 81788 4910 81844
rect 5618 81788 5628 81844
rect 5684 81788 7644 81844
rect 7700 81788 8092 81844
rect 8148 81788 8158 81844
rect 20290 81788 20300 81844
rect 20356 81788 20524 81844
rect 20580 81788 21308 81844
rect 21364 81788 22652 81844
rect 22708 81788 22718 81844
rect 24210 81788 24220 81844
rect 24276 81788 24556 81844
rect 24612 81788 24622 81844
rect 3332 81676 5068 81732
rect 5124 81676 10780 81732
rect 10836 81676 10846 81732
rect 11554 81676 11564 81732
rect 11620 81676 13692 81732
rect 13748 81676 13916 81732
rect 13972 81676 14476 81732
rect 14532 81676 14812 81732
rect 14868 81676 14878 81732
rect 16930 81676 16940 81732
rect 16996 81676 17724 81732
rect 17780 81676 17790 81732
rect 20738 81676 20748 81732
rect 20804 81676 21980 81732
rect 22036 81676 22046 81732
rect 3332 81284 3388 81676
rect 10658 81564 10668 81620
rect 10724 81564 11004 81620
rect 11060 81564 14028 81620
rect 14084 81564 14094 81620
rect 8006 81508 8016 81564
rect 8072 81508 8120 81564
rect 8176 81508 8224 81564
rect 8280 81508 8290 81564
rect 14810 81508 14820 81564
rect 14876 81508 14924 81564
rect 14980 81508 15028 81564
rect 15084 81508 15094 81564
rect 21614 81508 21624 81564
rect 21680 81508 21728 81564
rect 21784 81508 21832 81564
rect 21888 81508 21898 81564
rect 28418 81508 28428 81564
rect 28484 81508 28532 81564
rect 28588 81508 28636 81564
rect 28692 81508 28702 81564
rect 9426 81340 9436 81396
rect 9492 81340 10220 81396
rect 10276 81340 11564 81396
rect 11620 81340 11630 81396
rect 19058 81340 19068 81396
rect 19124 81340 19292 81396
rect 19348 81340 20748 81396
rect 20804 81340 22764 81396
rect 22820 81340 24668 81396
rect 24724 81340 24734 81396
rect 2594 81228 2604 81284
rect 2660 81228 3388 81284
rect 11330 81228 11340 81284
rect 11396 81228 20468 81284
rect 20626 81228 20636 81284
rect 20692 81228 23884 81284
rect 23940 81228 27020 81284
rect 27076 81228 27086 81284
rect 7298 81116 7308 81172
rect 7364 81116 9772 81172
rect 9828 81116 9838 81172
rect 16594 81116 16604 81172
rect 16660 81116 17724 81172
rect 17780 81116 17790 81172
rect 19394 81116 19404 81172
rect 19460 81116 19740 81172
rect 19796 81116 19964 81172
rect 20020 81116 20030 81172
rect 20412 81060 20468 81228
rect 21970 81116 21980 81172
rect 22036 81116 22988 81172
rect 23044 81116 26460 81172
rect 26516 81116 27132 81172
rect 27188 81116 27356 81172
rect 27412 81116 27422 81172
rect 6178 81004 6188 81060
rect 6244 81004 7756 81060
rect 7812 81004 7822 81060
rect 14130 81004 14140 81060
rect 14196 81004 19068 81060
rect 19124 81004 19134 81060
rect 20412 81004 22204 81060
rect 22260 81004 22270 81060
rect 24098 81004 24108 81060
rect 24164 81004 25228 81060
rect 25284 81004 25294 81060
rect 25778 81004 25788 81060
rect 25844 81004 26348 81060
rect 26404 81004 26414 81060
rect 5170 80892 5180 80948
rect 5236 80892 6636 80948
rect 6692 80892 6972 80948
rect 7028 80892 7038 80948
rect 11106 80892 11116 80948
rect 11172 80892 12796 80948
rect 12852 80892 12862 80948
rect 14242 80892 14252 80948
rect 14308 80892 16492 80948
rect 16548 80892 16558 80948
rect 17154 80892 17164 80948
rect 17220 80892 17612 80948
rect 17668 80892 17678 80948
rect 17938 80892 17948 80948
rect 18004 80892 18172 80948
rect 18228 80892 18238 80948
rect 24546 80892 24556 80948
rect 24612 80892 25452 80948
rect 25508 80892 25518 80948
rect 26226 80892 26236 80948
rect 26292 80892 26572 80948
rect 26628 80892 26638 80948
rect 27458 80780 27468 80836
rect 27524 80780 28028 80836
rect 28084 80780 28094 80836
rect 4604 80724 4614 80780
rect 4670 80724 4718 80780
rect 4774 80724 4822 80780
rect 4878 80724 4888 80780
rect 11408 80724 11418 80780
rect 11474 80724 11522 80780
rect 11578 80724 11626 80780
rect 11682 80724 11692 80780
rect 18212 80724 18222 80780
rect 18278 80724 18326 80780
rect 18382 80724 18430 80780
rect 18486 80724 18496 80780
rect 25016 80724 25026 80780
rect 25082 80724 25130 80780
rect 25186 80724 25234 80780
rect 25290 80724 25300 80780
rect 26562 80668 26572 80724
rect 26628 80668 26908 80724
rect 26964 80668 26974 80724
rect 14018 80556 14028 80612
rect 14084 80556 14364 80612
rect 14420 80556 14430 80612
rect 17042 80556 17052 80612
rect 17108 80556 17836 80612
rect 17892 80556 18844 80612
rect 18900 80556 19516 80612
rect 19572 80556 19582 80612
rect 19842 80556 19852 80612
rect 19908 80556 22540 80612
rect 22596 80556 22606 80612
rect 24546 80556 24556 80612
rect 24612 80556 25228 80612
rect 25284 80556 25294 80612
rect 26450 80556 26460 80612
rect 26516 80556 26908 80612
rect 26852 80500 26908 80556
rect 7858 80444 7868 80500
rect 7924 80444 22092 80500
rect 22148 80444 22158 80500
rect 23426 80444 23436 80500
rect 23492 80444 24444 80500
rect 24500 80444 24510 80500
rect 26852 80444 27020 80500
rect 27076 80444 27086 80500
rect 24770 80332 24780 80388
rect 24836 80332 25564 80388
rect 25620 80332 25630 80388
rect 17490 80220 17500 80276
rect 17556 80220 18732 80276
rect 18788 80220 18798 80276
rect 20514 80220 20524 80276
rect 20580 80220 21196 80276
rect 21252 80220 21262 80276
rect 2034 80108 2044 80164
rect 2100 80108 6076 80164
rect 6132 80108 17892 80164
rect 22642 80108 22652 80164
rect 22708 80108 23324 80164
rect 23380 80108 23390 80164
rect 26646 80108 26684 80164
rect 26740 80108 26750 80164
rect 0 80052 400 80080
rect 0 79996 1708 80052
rect 1764 79996 2492 80052
rect 2548 79996 2558 80052
rect 5030 79996 5068 80052
rect 5124 79996 5740 80052
rect 5796 79996 6524 80052
rect 6580 79996 6590 80052
rect 0 79968 400 79996
rect 8006 79940 8016 79996
rect 8072 79940 8120 79996
rect 8176 79940 8224 79996
rect 8280 79940 8290 79996
rect 14810 79940 14820 79996
rect 14876 79940 14924 79996
rect 14980 79940 15028 79996
rect 15084 79940 15094 79996
rect 17836 79940 17892 80108
rect 22082 79996 22092 80052
rect 22148 79996 27132 80052
rect 27188 79996 27198 80052
rect 21614 79940 21624 79996
rect 21680 79940 21728 79996
rect 21784 79940 21832 79996
rect 21888 79940 21898 79996
rect 28418 79940 28428 79996
rect 28484 79940 28532 79996
rect 28588 79940 28636 79996
rect 28692 79940 28702 79996
rect 17826 79884 17836 79940
rect 17892 79884 17902 79940
rect 17714 79772 17724 79828
rect 17780 79772 23996 79828
rect 24052 79772 24062 79828
rect 24546 79772 24556 79828
rect 24612 79772 26236 79828
rect 26292 79772 27916 79828
rect 27972 79772 27982 79828
rect 14578 79660 14588 79716
rect 14644 79660 14812 79716
rect 14868 79660 14878 79716
rect 17602 79660 17612 79716
rect 17668 79660 19068 79716
rect 19124 79660 19134 79716
rect 19954 79660 19964 79716
rect 20020 79660 20860 79716
rect 20916 79660 20926 79716
rect 9986 79548 9996 79604
rect 10052 79548 11676 79604
rect 11732 79548 11742 79604
rect 12002 79548 12012 79604
rect 12068 79548 12684 79604
rect 12740 79548 14924 79604
rect 14980 79548 16604 79604
rect 16660 79548 17948 79604
rect 18004 79548 18014 79604
rect 21522 79548 21532 79604
rect 21588 79548 23772 79604
rect 23828 79548 24220 79604
rect 24276 79548 25004 79604
rect 25060 79548 25788 79604
rect 25844 79548 25854 79604
rect 10546 79324 10556 79380
rect 10612 79324 12012 79380
rect 12068 79324 13132 79380
rect 13188 79324 13198 79380
rect 18162 79324 18172 79380
rect 18228 79324 19068 79380
rect 19124 79324 19134 79380
rect 4604 79156 4614 79212
rect 4670 79156 4718 79212
rect 4774 79156 4822 79212
rect 4878 79156 4888 79212
rect 11408 79156 11418 79212
rect 11474 79156 11522 79212
rect 11578 79156 11626 79212
rect 11682 79156 11692 79212
rect 18212 79156 18222 79212
rect 18278 79156 18326 79212
rect 18382 79156 18430 79212
rect 18486 79156 18496 79212
rect 25016 79156 25026 79212
rect 25082 79156 25130 79212
rect 25186 79156 25234 79212
rect 25290 79156 25300 79212
rect 14242 79100 14252 79156
rect 14308 79100 14700 79156
rect 14756 79100 14766 79156
rect 9874 78988 9884 79044
rect 9940 78988 12460 79044
rect 12516 78988 14588 79044
rect 14644 78988 14654 79044
rect 4498 78876 4508 78932
rect 4564 78876 4844 78932
rect 4900 78876 8316 78932
rect 8372 78876 8382 78932
rect 10322 78876 10332 78932
rect 10388 78876 11004 78932
rect 11060 78876 12236 78932
rect 12292 78876 12302 78932
rect 13234 78876 13244 78932
rect 13300 78876 13916 78932
rect 13972 78876 13982 78932
rect 25554 78876 25564 78932
rect 25620 78876 28140 78932
rect 28196 78876 28206 78932
rect 6178 78764 6188 78820
rect 6244 78764 7868 78820
rect 7924 78764 12572 78820
rect 12628 78764 12638 78820
rect 13010 78764 13020 78820
rect 13076 78764 13692 78820
rect 13748 78764 13758 78820
rect 14466 78764 14476 78820
rect 14532 78764 20188 78820
rect 20244 78764 23772 78820
rect 23828 78764 23838 78820
rect 4050 78652 4060 78708
rect 4116 78652 5852 78708
rect 5908 78652 6916 78708
rect 10322 78652 10332 78708
rect 10388 78652 11004 78708
rect 11060 78652 19740 78708
rect 19796 78652 21868 78708
rect 21924 78652 23324 78708
rect 23380 78652 23390 78708
rect 6860 78596 6916 78652
rect 3154 78540 3164 78596
rect 3220 78540 5068 78596
rect 5124 78540 6412 78596
rect 6468 78540 6478 78596
rect 6850 78540 6860 78596
rect 6916 78540 7868 78596
rect 7924 78540 8820 78596
rect 13010 78540 13020 78596
rect 13076 78540 16044 78596
rect 16100 78540 16110 78596
rect 19282 78540 19292 78596
rect 19348 78540 19628 78596
rect 19684 78540 21532 78596
rect 21588 78540 21598 78596
rect 22082 78540 22092 78596
rect 22148 78540 22540 78596
rect 22596 78540 22606 78596
rect 22754 78540 22764 78596
rect 22820 78540 23212 78596
rect 23268 78540 23278 78596
rect 23492 78540 24220 78596
rect 24276 78540 25116 78596
rect 25172 78540 25182 78596
rect 8764 78484 8820 78540
rect 22540 78484 22596 78540
rect 23492 78484 23548 78540
rect 8754 78428 8764 78484
rect 8820 78428 13468 78484
rect 13524 78428 14252 78484
rect 14308 78428 14318 78484
rect 14466 78428 14476 78484
rect 14532 78428 14542 78484
rect 19170 78428 19180 78484
rect 19236 78428 21308 78484
rect 21364 78428 21374 78484
rect 22540 78428 23548 78484
rect 8006 78372 8016 78428
rect 8072 78372 8120 78428
rect 8176 78372 8224 78428
rect 8280 78372 8290 78428
rect 14476 78372 14532 78428
rect 14810 78372 14820 78428
rect 14876 78372 14924 78428
rect 14980 78372 15028 78428
rect 15084 78372 15094 78428
rect 21614 78372 21624 78428
rect 21680 78372 21728 78428
rect 21784 78372 21832 78428
rect 21888 78372 21898 78428
rect 28418 78372 28428 78428
rect 28484 78372 28532 78428
rect 28588 78372 28636 78428
rect 28692 78372 28702 78428
rect 9436 78316 14532 78372
rect 16818 78316 16828 78372
rect 16884 78316 18844 78372
rect 18900 78316 18910 78372
rect 2818 78204 2828 78260
rect 2884 78204 4060 78260
rect 4116 78204 4126 78260
rect 9436 78148 9492 78316
rect 13570 78204 13580 78260
rect 13636 78204 14700 78260
rect 14756 78204 14766 78260
rect 15586 78204 15596 78260
rect 15652 78204 17500 78260
rect 17556 78204 17566 78260
rect 17714 78204 17724 78260
rect 17780 78204 18172 78260
rect 18228 78204 18508 78260
rect 18564 78204 18574 78260
rect 5954 78092 5964 78148
rect 6020 78092 9492 78148
rect 14354 78092 14364 78148
rect 14420 78092 17108 78148
rect 17052 78036 17108 78092
rect 2930 77980 2940 78036
rect 2996 77980 3500 78036
rect 3556 77980 3566 78036
rect 7858 77980 7868 78036
rect 7924 77980 9884 78036
rect 9940 77980 9950 78036
rect 17052 77980 17500 78036
rect 17556 77980 17948 78036
rect 18004 77980 19740 78036
rect 19796 77980 19806 78036
rect 13682 77868 13692 77924
rect 13748 77868 17388 77924
rect 17444 77868 17454 77924
rect 17602 77868 17612 77924
rect 17668 77868 19292 77924
rect 19348 77868 19358 77924
rect 24434 77868 24444 77924
rect 24500 77868 26012 77924
rect 26068 77868 26078 77924
rect 17826 77756 17836 77812
rect 17892 77756 18508 77812
rect 18564 77756 18574 77812
rect 18834 77756 18844 77812
rect 18900 77756 19180 77812
rect 19236 77756 20412 77812
rect 20468 77756 22092 77812
rect 22148 77756 22158 77812
rect 23202 77756 23212 77812
rect 23268 77756 24668 77812
rect 24724 77756 24734 77812
rect 6962 77644 6972 77700
rect 7028 77644 8540 77700
rect 8596 77644 9100 77700
rect 9156 77644 9166 77700
rect 4604 77588 4614 77644
rect 4670 77588 4718 77644
rect 4774 77588 4822 77644
rect 4878 77588 4888 77644
rect 11408 77588 11418 77644
rect 11474 77588 11522 77644
rect 11578 77588 11626 77644
rect 11682 77588 11692 77644
rect 18212 77588 18222 77644
rect 18278 77588 18326 77644
rect 18382 77588 18430 77644
rect 18486 77588 18496 77644
rect 25016 77588 25026 77644
rect 25082 77588 25130 77644
rect 25186 77588 25234 77644
rect 25290 77588 25300 77644
rect 17378 77420 17388 77476
rect 17444 77420 20636 77476
rect 20692 77420 20702 77476
rect 0 77364 400 77392
rect 0 77308 1708 77364
rect 1764 77308 1932 77364
rect 1988 77308 1998 77364
rect 17154 77308 17164 77364
rect 17220 77308 17612 77364
rect 17668 77308 17678 77364
rect 20514 77308 20524 77364
rect 20580 77308 21420 77364
rect 21476 77308 21486 77364
rect 0 77280 400 77308
rect 3332 77196 3500 77252
rect 3556 77196 3566 77252
rect 9650 77196 9660 77252
rect 9716 77196 10108 77252
rect 10164 77196 13468 77252
rect 13524 77196 13534 77252
rect 15026 77196 15036 77252
rect 15092 77196 17836 77252
rect 17892 77196 21084 77252
rect 21140 77196 21150 77252
rect 21410 77196 21420 77252
rect 21476 77196 21980 77252
rect 22036 77196 24780 77252
rect 24836 77196 24846 77252
rect 3332 77140 3388 77196
rect 2034 77084 2044 77140
rect 2100 77084 2716 77140
rect 2772 77084 3388 77140
rect 10770 77084 10780 77140
rect 10836 77084 11900 77140
rect 11956 77084 11966 77140
rect 13010 77084 13020 77140
rect 13076 77084 18396 77140
rect 18452 77084 20188 77140
rect 20244 77084 20254 77140
rect 22166 77084 22204 77140
rect 22260 77084 22652 77140
rect 22708 77084 23660 77140
rect 23716 77084 23726 77140
rect 24322 77084 24332 77140
rect 24388 77084 25900 77140
rect 25956 77084 25966 77140
rect 26226 77084 26236 77140
rect 26292 77084 27356 77140
rect 27412 77084 27422 77140
rect 11218 76972 11228 77028
rect 11284 76972 13580 77028
rect 13636 76972 13646 77028
rect 13906 76972 13916 77028
rect 13972 76972 19964 77028
rect 20020 76972 20030 77028
rect 24658 76972 24668 77028
rect 24724 76972 25564 77028
rect 25620 76972 25630 77028
rect 25900 76916 25956 77084
rect 27122 76972 27132 77028
rect 27188 76972 28140 77028
rect 28196 76972 28206 77028
rect 9538 76860 9548 76916
rect 9604 76860 12796 76916
rect 12852 76860 13132 76916
rect 13188 76860 13198 76916
rect 25900 76860 26684 76916
rect 26740 76860 27020 76916
rect 27076 76860 27086 76916
rect 8006 76804 8016 76860
rect 8072 76804 8120 76860
rect 8176 76804 8224 76860
rect 8280 76804 8290 76860
rect 14810 76804 14820 76860
rect 14876 76804 14924 76860
rect 14980 76804 15028 76860
rect 15084 76804 15094 76860
rect 21614 76804 21624 76860
rect 21680 76804 21728 76860
rect 21784 76804 21832 76860
rect 21888 76804 21898 76860
rect 28418 76804 28428 76860
rect 28484 76804 28532 76860
rect 28588 76804 28636 76860
rect 28692 76804 28702 76860
rect 25330 76748 25340 76804
rect 25396 76748 26460 76804
rect 26516 76748 26526 76804
rect 4610 76636 4620 76692
rect 4676 76636 6132 76692
rect 8754 76636 8764 76692
rect 8820 76636 11116 76692
rect 11172 76636 11182 76692
rect 22866 76636 22876 76692
rect 22932 76636 23772 76692
rect 23828 76636 23838 76692
rect 24882 76636 24892 76692
rect 24948 76636 27020 76692
rect 27076 76636 27086 76692
rect 6076 76580 6132 76636
rect 3490 76524 3500 76580
rect 3556 76524 3724 76580
rect 3780 76524 5068 76580
rect 5124 76524 5134 76580
rect 6066 76524 6076 76580
rect 6132 76524 7084 76580
rect 7140 76524 7150 76580
rect 10434 76524 10444 76580
rect 10500 76524 13244 76580
rect 13300 76524 13310 76580
rect 4050 76412 4060 76468
rect 4116 76412 5292 76468
rect 5348 76412 6860 76468
rect 6916 76412 6926 76468
rect 9762 76412 9772 76468
rect 9828 76412 10108 76468
rect 10164 76412 11788 76468
rect 11844 76412 11854 76468
rect 14018 76412 14028 76468
rect 14084 76412 14140 76468
rect 14196 76412 16492 76468
rect 16548 76412 16558 76468
rect 26338 76412 26348 76468
rect 26404 76412 26796 76468
rect 26852 76412 27580 76468
rect 27636 76412 27646 76468
rect 5506 76300 5516 76356
rect 5572 76300 5740 76356
rect 5796 76300 6524 76356
rect 6580 76300 7924 76356
rect 8530 76300 8540 76356
rect 8596 76300 12124 76356
rect 12180 76300 12190 76356
rect 17602 76300 17612 76356
rect 17668 76300 18956 76356
rect 19012 76300 19022 76356
rect 20626 76300 20636 76356
rect 20692 76300 21420 76356
rect 21476 76300 21756 76356
rect 21812 76300 21822 76356
rect 22530 76300 22540 76356
rect 22596 76300 23548 76356
rect 23604 76300 23614 76356
rect 7868 76244 7924 76300
rect 6290 76188 6300 76244
rect 6356 76188 7644 76244
rect 7700 76188 7710 76244
rect 7868 76188 8988 76244
rect 9044 76188 11004 76244
rect 11060 76188 11070 76244
rect 12786 76188 12796 76244
rect 12852 76188 23884 76244
rect 23940 76188 26684 76244
rect 26740 76188 26750 76244
rect 7074 76076 7084 76132
rect 7140 76076 7756 76132
rect 7812 76076 7822 76132
rect 18946 76076 18956 76132
rect 19012 76076 21532 76132
rect 21588 76076 22652 76132
rect 22708 76076 22718 76132
rect 4604 76020 4614 76076
rect 4670 76020 4718 76076
rect 4774 76020 4822 76076
rect 4878 76020 4888 76076
rect 11408 76020 11418 76076
rect 11474 76020 11522 76076
rect 11578 76020 11626 76076
rect 11682 76020 11692 76076
rect 18212 76020 18222 76076
rect 18278 76020 18326 76076
rect 18382 76020 18430 76076
rect 18486 76020 18496 76076
rect 25016 76020 25026 76076
rect 25082 76020 25130 76076
rect 25186 76020 25234 76076
rect 25290 76020 25300 76076
rect 15222 75964 15260 76020
rect 15316 75964 15326 76020
rect 6850 75852 6860 75908
rect 6916 75852 23884 75908
rect 23940 75852 24556 75908
rect 24612 75852 24622 75908
rect 9762 75740 9772 75796
rect 9828 75740 10220 75796
rect 10276 75740 10286 75796
rect 13458 75740 13468 75796
rect 13524 75740 16828 75796
rect 16884 75740 16894 75796
rect 20188 75740 20748 75796
rect 20804 75740 22316 75796
rect 22372 75740 22540 75796
rect 22596 75740 22606 75796
rect 24770 75740 24780 75796
rect 24836 75740 25676 75796
rect 25732 75740 25742 75796
rect 20188 75684 20244 75740
rect 2930 75628 2940 75684
rect 2996 75628 4956 75684
rect 5012 75628 5022 75684
rect 12114 75628 12124 75684
rect 12180 75628 15764 75684
rect 17490 75628 17500 75684
rect 17556 75628 18284 75684
rect 18340 75628 20188 75684
rect 20244 75628 20254 75684
rect 20412 75628 23100 75684
rect 23156 75628 23166 75684
rect 25218 75628 25228 75684
rect 25284 75628 26572 75684
rect 26628 75628 27020 75684
rect 27076 75628 27356 75684
rect 27412 75628 27422 75684
rect 8642 75516 8652 75572
rect 8708 75516 10444 75572
rect 10500 75516 10510 75572
rect 10994 75516 11004 75572
rect 11060 75516 15652 75572
rect 6962 75404 6972 75460
rect 7028 75404 8540 75460
rect 8596 75404 9772 75460
rect 9828 75404 9838 75460
rect 13570 75404 13580 75460
rect 13636 75404 13692 75460
rect 13748 75404 13758 75460
rect 15596 75348 15652 75516
rect 15708 75460 15764 75628
rect 17378 75516 17388 75572
rect 17444 75516 17724 75572
rect 17780 75516 19628 75572
rect 19684 75516 19694 75572
rect 20412 75460 20468 75628
rect 23650 75516 23660 75572
rect 23716 75516 27132 75572
rect 27188 75516 27198 75572
rect 15708 75404 17276 75460
rect 17332 75404 17948 75460
rect 18004 75404 18014 75460
rect 20402 75404 20412 75460
rect 20468 75404 20478 75460
rect 20636 75404 25228 75460
rect 25284 75404 25294 75460
rect 26898 75404 26908 75460
rect 26964 75404 27804 75460
rect 27860 75404 27870 75460
rect 20636 75348 20692 75404
rect 15586 75292 15596 75348
rect 15652 75292 15932 75348
rect 15988 75292 20692 75348
rect 8006 75236 8016 75292
rect 8072 75236 8120 75292
rect 8176 75236 8224 75292
rect 8280 75236 8290 75292
rect 14810 75236 14820 75292
rect 14876 75236 14924 75292
rect 14980 75236 15028 75292
rect 15084 75236 15094 75292
rect 21614 75236 21624 75292
rect 21680 75236 21728 75292
rect 21784 75236 21832 75292
rect 21888 75236 21898 75292
rect 26236 75180 26796 75236
rect 26852 75180 26862 75236
rect 26236 75124 26292 75180
rect 27020 75124 27076 75404
rect 28418 75236 28428 75292
rect 28484 75236 28532 75292
rect 28588 75236 28636 75292
rect 28692 75236 28702 75292
rect 7970 75068 7980 75124
rect 8036 75068 8764 75124
rect 8820 75068 9996 75124
rect 10052 75068 10062 75124
rect 11190 75068 11228 75124
rect 11284 75068 12348 75124
rect 12404 75068 13860 75124
rect 15138 75068 15148 75124
rect 15204 75068 16380 75124
rect 16436 75068 16446 75124
rect 17714 75068 17724 75124
rect 17780 75068 18060 75124
rect 18116 75068 18126 75124
rect 18610 75068 18620 75124
rect 18676 75068 20860 75124
rect 20916 75068 26292 75124
rect 26348 75068 27076 75124
rect 13804 75012 13860 75068
rect 12562 74956 12572 75012
rect 12628 74956 13580 75012
rect 13636 74956 13646 75012
rect 13804 74956 24108 75012
rect 24164 74956 24556 75012
rect 24612 74956 24622 75012
rect 26348 74900 26404 75068
rect 2034 74844 2044 74900
rect 2100 74844 2828 74900
rect 2884 74844 3612 74900
rect 3668 74844 3678 74900
rect 6066 74844 6076 74900
rect 6132 74844 6860 74900
rect 6916 74844 6926 74900
rect 11442 74844 11452 74900
rect 11508 74844 11900 74900
rect 11956 74844 12460 74900
rect 12516 74844 12526 74900
rect 13234 74844 13244 74900
rect 13300 74844 14028 74900
rect 14084 74844 14094 74900
rect 14578 74844 14588 74900
rect 14644 74844 15036 74900
rect 15092 74844 15102 74900
rect 16818 74844 16828 74900
rect 16884 74844 26348 74900
rect 26404 74844 26414 74900
rect 16828 74788 16884 74844
rect 4162 74732 4172 74788
rect 4228 74732 5292 74788
rect 5348 74732 5964 74788
rect 6020 74732 6030 74788
rect 14354 74732 14364 74788
rect 14420 74732 14924 74788
rect 14980 74732 16884 74788
rect 19926 74732 19964 74788
rect 20020 74732 20030 74788
rect 22530 74732 22540 74788
rect 22596 74732 23212 74788
rect 23268 74732 23278 74788
rect 23426 74732 23436 74788
rect 23492 74732 26124 74788
rect 26180 74732 26190 74788
rect 0 74676 400 74704
rect 0 74620 1708 74676
rect 1764 74620 2268 74676
rect 2324 74620 2334 74676
rect 13990 74620 14028 74676
rect 14084 74620 16044 74676
rect 16100 74620 16110 74676
rect 16482 74620 16492 74676
rect 16548 74620 17276 74676
rect 17332 74620 17342 74676
rect 18060 74620 24892 74676
rect 24948 74620 24958 74676
rect 0 74592 400 74620
rect 18060 74564 18116 74620
rect 11890 74508 11900 74564
rect 11956 74508 12796 74564
rect 12852 74508 14252 74564
rect 14308 74508 14318 74564
rect 15092 74508 18116 74564
rect 18610 74508 18620 74564
rect 18676 74508 19180 74564
rect 19236 74508 19246 74564
rect 4604 74452 4614 74508
rect 4670 74452 4718 74508
rect 4774 74452 4822 74508
rect 4878 74452 4888 74508
rect 11408 74452 11418 74508
rect 11474 74452 11522 74508
rect 11578 74452 11626 74508
rect 11682 74452 11692 74508
rect 15092 74452 15148 74508
rect 18212 74452 18222 74508
rect 18278 74452 18326 74508
rect 18382 74452 18430 74508
rect 18486 74452 18496 74508
rect 25016 74452 25026 74508
rect 25082 74452 25130 74508
rect 25186 74452 25234 74508
rect 25290 74452 25300 74508
rect 11778 74396 11788 74452
rect 11844 74396 12124 74452
rect 12180 74396 12348 74452
rect 12404 74396 15148 74452
rect 23538 74396 23548 74452
rect 23604 74396 23642 74452
rect 26572 74396 26796 74452
rect 26852 74396 26862 74452
rect 26572 74340 26628 74396
rect 3154 74284 3164 74340
rect 3220 74284 4060 74340
rect 4116 74284 4126 74340
rect 5954 74284 5964 74340
rect 6020 74284 26572 74340
rect 26628 74284 26638 74340
rect 26786 74284 26796 74340
rect 26852 74284 27580 74340
rect 27636 74284 27646 74340
rect 2482 74172 2492 74228
rect 2548 74172 2940 74228
rect 2996 74172 3612 74228
rect 3668 74172 3678 74228
rect 11218 74172 11228 74228
rect 11284 74172 11788 74228
rect 11844 74172 11854 74228
rect 13794 74172 13804 74228
rect 13860 74172 18508 74228
rect 18564 74172 18574 74228
rect 18946 74172 18956 74228
rect 19012 74172 19292 74228
rect 19348 74172 19358 74228
rect 22530 74172 22540 74228
rect 22596 74172 24220 74228
rect 24276 74172 24286 74228
rect 24994 74172 25004 74228
rect 25060 74172 25676 74228
rect 25732 74172 28028 74228
rect 28084 74172 28094 74228
rect 8988 74060 9996 74116
rect 10052 74060 10062 74116
rect 12534 74060 12572 74116
rect 12628 74060 12638 74116
rect 15698 74060 15708 74116
rect 15764 74060 19852 74116
rect 19908 74060 20300 74116
rect 20356 74060 20366 74116
rect 26562 74060 26572 74116
rect 26628 74060 27020 74116
rect 27076 74060 27086 74116
rect 8988 74004 9044 74060
rect 6514 73948 6524 74004
rect 6580 73948 7196 74004
rect 7252 73948 7262 74004
rect 8978 73948 8988 74004
rect 9044 73948 9054 74004
rect 9314 73948 9324 74004
rect 9380 73948 11676 74004
rect 11732 73948 11742 74004
rect 13682 73948 13692 74004
rect 13748 73948 13804 74004
rect 13860 73948 13870 74004
rect 18956 73948 19516 74004
rect 19572 73948 19582 74004
rect 25666 73948 25676 74004
rect 25732 73948 27132 74004
rect 27188 73948 28140 74004
rect 28196 73948 28206 74004
rect 4834 73836 4844 73892
rect 4900 73836 5740 73892
rect 5796 73836 5806 73892
rect 8754 73836 8764 73892
rect 8820 73836 9772 73892
rect 9828 73836 9838 73892
rect 13122 73836 13132 73892
rect 13188 73836 14588 73892
rect 14644 73836 15372 73892
rect 15428 73836 15438 73892
rect 18956 73780 19012 73948
rect 23202 73836 23212 73892
rect 23268 73836 23660 73892
rect 23716 73836 23726 73892
rect 23874 73836 23884 73892
rect 23940 73836 23978 73892
rect 24518 73836 24556 73892
rect 24612 73836 24892 73892
rect 24948 73836 24958 73892
rect 25330 73836 25340 73892
rect 25396 73836 28252 73892
rect 28308 73836 28318 73892
rect 18722 73724 18732 73780
rect 18788 73724 19012 73780
rect 22754 73724 22764 73780
rect 22820 73724 24332 73780
rect 24388 73724 24398 73780
rect 8006 73668 8016 73724
rect 8072 73668 8120 73724
rect 8176 73668 8224 73724
rect 8280 73668 8290 73724
rect 14810 73668 14820 73724
rect 14876 73668 14924 73724
rect 14980 73668 15028 73724
rect 15084 73668 15094 73724
rect 21614 73668 21624 73724
rect 21680 73668 21728 73724
rect 21784 73668 21832 73724
rect 21888 73668 21898 73724
rect 28418 73668 28428 73724
rect 28484 73668 28532 73724
rect 28588 73668 28636 73724
rect 28692 73668 28702 73724
rect 18834 73612 18844 73668
rect 18900 73612 19964 73668
rect 20020 73612 20030 73668
rect 23538 73612 23548 73668
rect 23604 73612 23642 73668
rect 26674 73612 26684 73668
rect 26740 73612 27244 73668
rect 27300 73612 27310 73668
rect 2930 73500 2940 73556
rect 2996 73500 3006 73556
rect 8418 73500 8428 73556
rect 8484 73500 9548 73556
rect 9604 73500 10892 73556
rect 10948 73500 15596 73556
rect 15652 73500 15662 73556
rect 16604 73500 20300 73556
rect 20356 73500 20366 73556
rect 23650 73500 23660 73556
rect 23716 73500 25452 73556
rect 25508 73500 26460 73556
rect 26516 73500 26526 73556
rect 2034 73388 2044 73444
rect 2100 73388 2716 73444
rect 2772 73388 2782 73444
rect 2940 73332 2996 73500
rect 16604 73444 16660 73500
rect 14018 73388 14028 73444
rect 14084 73388 14700 73444
rect 14756 73388 14766 73444
rect 15250 73388 15260 73444
rect 15316 73388 15820 73444
rect 15876 73388 16660 73444
rect 18022 73388 18060 73444
rect 18116 73388 20748 73444
rect 20804 73388 20814 73444
rect 22978 73388 22988 73444
rect 23044 73388 23604 73444
rect 23986 73388 23996 73444
rect 24052 73388 24332 73444
rect 24388 73388 24398 73444
rect 23548 73332 23604 73388
rect 2370 73276 2380 73332
rect 2436 73276 2996 73332
rect 13794 73276 13804 73332
rect 13860 73276 13916 73332
rect 13972 73276 13982 73332
rect 14242 73276 14252 73332
rect 14308 73276 17948 73332
rect 18004 73276 18014 73332
rect 18274 73276 18284 73332
rect 18340 73276 23268 73332
rect 23538 73276 23548 73332
rect 23604 73276 23614 73332
rect 13682 73164 13692 73220
rect 13748 73164 15148 73220
rect 15204 73164 15260 73220
rect 15316 73164 15326 73220
rect 15782 73164 15820 73220
rect 15876 73164 17500 73220
rect 17556 73164 17566 73220
rect 21858 73164 21868 73220
rect 21924 73164 22428 73220
rect 22484 73164 22988 73220
rect 23044 73164 23054 73220
rect 23212 73108 23268 73276
rect 15474 73052 15484 73108
rect 15540 73052 21308 73108
rect 21364 73052 21374 73108
rect 21634 73052 21644 73108
rect 21700 73052 22316 73108
rect 22372 73052 22382 73108
rect 23202 73052 23212 73108
rect 23268 73052 23278 73108
rect 21074 72940 21084 72996
rect 21140 72940 21868 72996
rect 21924 72940 21934 72996
rect 22194 72940 22204 72996
rect 22260 72940 22764 72996
rect 22820 72940 24668 72996
rect 24724 72940 24734 72996
rect 4604 72884 4614 72940
rect 4670 72884 4718 72940
rect 4774 72884 4822 72940
rect 4878 72884 4888 72940
rect 11408 72884 11418 72940
rect 11474 72884 11522 72940
rect 11578 72884 11626 72940
rect 11682 72884 11692 72940
rect 18212 72884 18222 72940
rect 18278 72884 18326 72940
rect 18382 72884 18430 72940
rect 18486 72884 18496 72940
rect 25016 72884 25026 72940
rect 25082 72884 25130 72940
rect 25186 72884 25234 72940
rect 25290 72884 25300 72940
rect 12226 72828 12236 72884
rect 12292 72828 12684 72884
rect 12740 72828 12750 72884
rect 15586 72828 15596 72884
rect 15652 72828 16492 72884
rect 16548 72828 16558 72884
rect 25778 72828 25788 72884
rect 25844 72828 26460 72884
rect 26516 72828 26526 72884
rect 7186 72716 7196 72772
rect 7252 72716 7868 72772
rect 7924 72716 8540 72772
rect 8596 72716 8606 72772
rect 12786 72716 12796 72772
rect 12852 72716 14028 72772
rect 14084 72716 14094 72772
rect 15092 72716 16324 72772
rect 23398 72716 23436 72772
rect 23492 72716 23502 72772
rect 15092 72660 15148 72716
rect 16268 72660 16324 72716
rect 6178 72604 6188 72660
rect 6244 72604 6972 72660
rect 7028 72604 7038 72660
rect 7970 72604 7980 72660
rect 8036 72604 9324 72660
rect 9380 72604 9390 72660
rect 10098 72604 10108 72660
rect 10164 72604 11116 72660
rect 11172 72604 12908 72660
rect 12964 72604 14476 72660
rect 14532 72604 15148 72660
rect 16258 72604 16268 72660
rect 16324 72604 16334 72660
rect 16706 72604 16716 72660
rect 16772 72604 17836 72660
rect 17892 72604 17902 72660
rect 1810 72492 1820 72548
rect 1876 72492 4396 72548
rect 4452 72492 4956 72548
rect 5012 72492 7644 72548
rect 7700 72492 8092 72548
rect 8148 72492 8158 72548
rect 8866 72492 8876 72548
rect 8932 72492 13580 72548
rect 13636 72492 13646 72548
rect 13804 72492 14588 72548
rect 14644 72492 16380 72548
rect 16436 72492 16446 72548
rect 17266 72492 17276 72548
rect 17332 72492 19180 72548
rect 19236 72492 19246 72548
rect 19506 72492 19516 72548
rect 19572 72492 19582 72548
rect 21158 72492 21196 72548
rect 21252 72492 21262 72548
rect 22530 72492 22540 72548
rect 22596 72492 22988 72548
rect 23044 72492 23054 72548
rect 23202 72492 23212 72548
rect 23268 72492 23548 72548
rect 13804 72436 13860 72492
rect 19516 72436 19572 72492
rect 23492 72436 23548 72492
rect 3490 72380 3500 72436
rect 3556 72380 5068 72436
rect 5124 72380 6076 72436
rect 6132 72380 6636 72436
rect 6692 72380 6702 72436
rect 9996 72380 13860 72436
rect 15138 72380 15148 72436
rect 15204 72380 15932 72436
rect 15988 72380 15998 72436
rect 18946 72380 18956 72436
rect 19012 72380 19572 72436
rect 21858 72380 21868 72436
rect 21924 72380 22540 72436
rect 22596 72380 22606 72436
rect 23492 72380 24388 72436
rect 9996 72324 10052 72380
rect 24332 72324 24388 72380
rect 9062 72268 9100 72324
rect 9156 72268 9166 72324
rect 9986 72268 9996 72324
rect 10052 72268 10062 72324
rect 12786 72268 12796 72324
rect 12852 72268 14140 72324
rect 14196 72268 14206 72324
rect 15250 72268 15260 72324
rect 15316 72268 15372 72324
rect 15428 72268 15438 72324
rect 15586 72268 15596 72324
rect 15652 72268 15690 72324
rect 19506 72268 19516 72324
rect 19572 72268 20524 72324
rect 20580 72268 21084 72324
rect 21140 72268 21150 72324
rect 22082 72268 22092 72324
rect 22148 72268 23772 72324
rect 23828 72268 24108 72324
rect 24164 72268 24174 72324
rect 24332 72268 24556 72324
rect 24612 72268 24622 72324
rect 3042 72156 3052 72212
rect 3108 72156 3612 72212
rect 3668 72156 3678 72212
rect 10434 72156 10444 72212
rect 10500 72156 11228 72212
rect 11284 72156 12012 72212
rect 12068 72156 12078 72212
rect 12226 72156 12236 72212
rect 12292 72156 12302 72212
rect 15362 72156 15372 72212
rect 15428 72156 16716 72212
rect 16772 72156 16782 72212
rect 21970 72156 21980 72212
rect 22036 72156 25004 72212
rect 25060 72156 25070 72212
rect 8006 72100 8016 72156
rect 8072 72100 8120 72156
rect 8176 72100 8224 72156
rect 8280 72100 8290 72156
rect 12236 72100 12292 72156
rect 14810 72100 14820 72156
rect 14876 72100 14924 72156
rect 14980 72100 15028 72156
rect 15084 72100 15094 72156
rect 21614 72100 21624 72156
rect 21680 72100 21728 72156
rect 21784 72100 21832 72156
rect 21888 72100 21898 72156
rect 28418 72100 28428 72156
rect 28484 72100 28532 72156
rect 28588 72100 28636 72156
rect 28692 72100 28702 72156
rect 11666 72044 11676 72100
rect 11732 72044 14252 72100
rect 14308 72044 14318 72100
rect 16370 72044 16380 72100
rect 16436 72044 21028 72100
rect 22306 72044 22316 72100
rect 22372 72044 24556 72100
rect 24612 72044 24622 72100
rect 25666 72044 25676 72100
rect 25732 72044 26684 72100
rect 26740 72044 26750 72100
rect 0 71988 400 72016
rect 0 71932 1708 71988
rect 1764 71932 1774 71988
rect 10098 71932 10108 71988
rect 10164 71932 10556 71988
rect 10612 71932 10622 71988
rect 11778 71932 11788 71988
rect 11844 71932 12908 71988
rect 12964 71932 12974 71988
rect 14354 71932 14364 71988
rect 14420 71932 15036 71988
rect 15092 71932 15102 71988
rect 16482 71932 16492 71988
rect 16548 71932 17500 71988
rect 17556 71932 17566 71988
rect 18610 71932 18620 71988
rect 18676 71932 19068 71988
rect 19124 71932 19134 71988
rect 0 71904 400 71932
rect 20972 71876 21028 72044
rect 21522 71932 21532 71988
rect 21588 71932 27468 71988
rect 27524 71932 27534 71988
rect 2258 71820 2268 71876
rect 2324 71820 3276 71876
rect 3332 71820 3342 71876
rect 4162 71820 4172 71876
rect 4228 71820 4508 71876
rect 4564 71820 4574 71876
rect 10994 71820 11004 71876
rect 11060 71820 11564 71876
rect 11620 71820 11630 71876
rect 12002 71820 12012 71876
rect 12068 71820 15484 71876
rect 15540 71820 15550 71876
rect 18050 71820 18060 71876
rect 18116 71820 20748 71876
rect 20804 71820 20814 71876
rect 20972 71820 25564 71876
rect 25620 71820 25630 71876
rect 2594 71708 2604 71764
rect 2660 71708 3388 71764
rect 3444 71708 3454 71764
rect 8418 71708 8428 71764
rect 8484 71708 8764 71764
rect 8820 71708 8830 71764
rect 10770 71708 10780 71764
rect 10836 71708 15484 71764
rect 15540 71708 15550 71764
rect 15698 71708 15708 71764
rect 15764 71708 24668 71764
rect 24724 71708 24734 71764
rect 3938 71596 3948 71652
rect 4004 71596 4508 71652
rect 4564 71596 4574 71652
rect 5170 71596 5180 71652
rect 5236 71596 5740 71652
rect 5796 71596 5806 71652
rect 8978 71596 8988 71652
rect 9044 71596 9436 71652
rect 9492 71596 9502 71652
rect 9650 71596 9660 71652
rect 9716 71596 16212 71652
rect 16454 71596 16492 71652
rect 16548 71596 16558 71652
rect 18274 71596 18284 71652
rect 18340 71596 23660 71652
rect 23716 71596 23726 71652
rect 16156 71540 16212 71596
rect 9538 71484 9548 71540
rect 9604 71484 13468 71540
rect 13524 71484 13534 71540
rect 13906 71484 13916 71540
rect 13972 71484 13982 71540
rect 14214 71484 14252 71540
rect 14308 71484 14318 71540
rect 14914 71484 14924 71540
rect 14980 71484 15372 71540
rect 15428 71484 15438 71540
rect 16146 71484 16156 71540
rect 16212 71484 16222 71540
rect 17266 71484 17276 71540
rect 17332 71484 19292 71540
rect 19348 71484 19358 71540
rect 21382 71484 21420 71540
rect 21476 71484 21486 71540
rect 22502 71484 22540 71540
rect 22596 71484 22606 71540
rect 23314 71484 23324 71540
rect 23380 71484 23436 71540
rect 23492 71484 25340 71540
rect 25396 71484 25406 71540
rect 13916 71428 13972 71484
rect 13916 71372 17948 71428
rect 18004 71372 18014 71428
rect 4604 71316 4614 71372
rect 4670 71316 4718 71372
rect 4774 71316 4822 71372
rect 4878 71316 4888 71372
rect 11408 71316 11418 71372
rect 11474 71316 11522 71372
rect 11578 71316 11626 71372
rect 11682 71316 11692 71372
rect 18212 71316 18222 71372
rect 18278 71316 18326 71372
rect 18382 71316 18430 71372
rect 18486 71316 18496 71372
rect 25016 71316 25026 71372
rect 25082 71316 25130 71372
rect 25186 71316 25234 71372
rect 25290 71316 25300 71372
rect 11788 71260 17276 71316
rect 17332 71260 17342 71316
rect 23202 71260 23212 71316
rect 23268 71260 23436 71316
rect 23492 71260 23502 71316
rect 11788 71204 11844 71260
rect 10658 71148 10668 71204
rect 10724 71148 11844 71204
rect 13010 71148 13020 71204
rect 13076 71148 13468 71204
rect 13524 71148 13534 71204
rect 13906 71148 13916 71204
rect 13972 71148 14140 71204
rect 14196 71148 14206 71204
rect 14466 71148 14476 71204
rect 14532 71148 16716 71204
rect 16772 71148 16782 71204
rect 17938 71148 17948 71204
rect 18004 71148 18844 71204
rect 18900 71148 18910 71204
rect 3826 71036 3836 71092
rect 3892 71036 7700 71092
rect 7970 71036 7980 71092
rect 8036 71036 8876 71092
rect 8932 71036 13244 71092
rect 13300 71036 13310 71092
rect 13468 71036 26012 71092
rect 26068 71036 26684 71092
rect 26740 71036 26750 71092
rect 27010 71036 27020 71092
rect 27076 71036 28140 71092
rect 28196 71036 28206 71092
rect 6066 70924 6076 70980
rect 6132 70924 6860 70980
rect 6916 70924 6926 70980
rect 7644 70868 7700 71036
rect 10434 70924 10444 70980
rect 10500 70924 11228 70980
rect 11284 70924 11294 70980
rect 13468 70868 13524 71036
rect 13654 70924 13692 70980
rect 13748 70924 13758 70980
rect 13906 70924 13916 70980
rect 13972 70924 14924 70980
rect 14980 70924 14990 70980
rect 15092 70924 15260 70980
rect 15316 70924 15326 70980
rect 15474 70924 15484 70980
rect 15540 70924 15876 70980
rect 16006 70924 16044 70980
rect 16100 70924 16110 70980
rect 16370 70924 16380 70980
rect 16436 70924 16828 70980
rect 16884 70924 16894 70980
rect 19058 70924 19068 70980
rect 19124 70924 19740 70980
rect 19796 70924 20188 70980
rect 20244 70924 20254 70980
rect 20514 70924 20524 70980
rect 20580 70924 21532 70980
rect 21588 70924 21598 70980
rect 23314 70924 23324 70980
rect 23380 70924 23418 70980
rect 15092 70868 15148 70924
rect 15820 70868 15876 70924
rect 6738 70812 6748 70868
rect 6804 70812 7420 70868
rect 7476 70812 7486 70868
rect 7644 70812 13524 70868
rect 13766 70812 13804 70868
rect 13860 70812 13870 70868
rect 14102 70812 14140 70868
rect 14196 70812 15148 70868
rect 15362 70812 15372 70868
rect 15428 70812 15484 70868
rect 15540 70812 15550 70868
rect 15820 70812 23100 70868
rect 23156 70812 23436 70868
rect 23492 70812 23502 70868
rect 1922 70700 1932 70756
rect 1988 70700 2604 70756
rect 2660 70700 2670 70756
rect 3266 70700 3276 70756
rect 3332 70700 3948 70756
rect 4004 70700 4014 70756
rect 4162 70700 4172 70756
rect 4228 70700 4508 70756
rect 4564 70700 5964 70756
rect 6020 70700 6030 70756
rect 7308 70700 7980 70756
rect 8036 70700 8046 70756
rect 10770 70700 10780 70756
rect 10836 70700 12460 70756
rect 12516 70700 14028 70756
rect 14084 70700 14094 70756
rect 14242 70700 14252 70756
rect 14308 70700 14644 70756
rect 16706 70700 16716 70756
rect 16772 70700 18284 70756
rect 18340 70700 18350 70756
rect 19506 70700 19516 70756
rect 19572 70700 20188 70756
rect 20244 70700 24780 70756
rect 24836 70700 24846 70756
rect 7308 70644 7364 70700
rect 5058 70588 5068 70644
rect 5124 70588 5628 70644
rect 5684 70588 7364 70644
rect 8530 70588 8540 70644
rect 8596 70588 9772 70644
rect 9828 70588 9838 70644
rect 10434 70588 10444 70644
rect 10500 70588 11788 70644
rect 11844 70588 11854 70644
rect 12898 70588 12908 70644
rect 12964 70588 13244 70644
rect 13300 70588 13580 70644
rect 13636 70588 13646 70644
rect 14130 70588 14140 70644
rect 14196 70588 14364 70644
rect 14420 70588 14430 70644
rect 8006 70532 8016 70588
rect 8072 70532 8120 70588
rect 8176 70532 8224 70588
rect 8280 70532 8290 70588
rect 14588 70532 14644 70700
rect 15250 70588 15260 70644
rect 15316 70588 15596 70644
rect 15652 70588 15662 70644
rect 16034 70588 16044 70644
rect 16100 70588 17500 70644
rect 17556 70588 17566 70644
rect 18162 70588 18172 70644
rect 18228 70588 19068 70644
rect 19124 70588 19134 70644
rect 20822 70588 20860 70644
rect 20916 70588 20926 70644
rect 21970 70588 21980 70644
rect 22036 70588 22074 70644
rect 14810 70532 14820 70588
rect 14876 70532 14924 70588
rect 14980 70532 15028 70588
rect 15084 70532 15094 70588
rect 21614 70532 21624 70588
rect 21680 70532 21728 70588
rect 21784 70532 21832 70588
rect 21888 70532 21898 70588
rect 28418 70532 28428 70588
rect 28484 70532 28532 70588
rect 28588 70532 28636 70588
rect 28692 70532 28702 70588
rect 1810 70476 1820 70532
rect 1876 70476 3052 70532
rect 3108 70476 3118 70532
rect 3332 70476 5180 70532
rect 5236 70476 5852 70532
rect 5908 70476 5918 70532
rect 14578 70476 14588 70532
rect 14644 70476 14654 70532
rect 3332 70084 3388 70476
rect 7074 70364 7084 70420
rect 7140 70364 9772 70420
rect 9828 70364 9838 70420
rect 9986 70364 9996 70420
rect 10052 70364 10220 70420
rect 10276 70364 10286 70420
rect 10658 70364 10668 70420
rect 10724 70364 11340 70420
rect 11396 70364 11406 70420
rect 14140 70364 19740 70420
rect 19796 70364 21308 70420
rect 21364 70364 21644 70420
rect 21700 70364 21710 70420
rect 27122 70364 27132 70420
rect 27188 70364 27916 70420
rect 27972 70364 27982 70420
rect 14140 70308 14196 70364
rect 9538 70252 9548 70308
rect 9604 70252 10892 70308
rect 10948 70252 10958 70308
rect 11116 70252 14196 70308
rect 18386 70252 18396 70308
rect 18452 70252 19516 70308
rect 19572 70252 20300 70308
rect 20356 70252 20366 70308
rect 11116 70196 11172 70252
rect 5506 70140 5516 70196
rect 5572 70140 11172 70196
rect 12898 70140 12908 70196
rect 12964 70140 13356 70196
rect 13412 70140 13422 70196
rect 14018 70140 14028 70196
rect 14084 70140 15148 70196
rect 15204 70140 15214 70196
rect 3042 70028 3052 70084
rect 3108 70028 3388 70084
rect 11890 70028 11900 70084
rect 11956 70028 12684 70084
rect 12740 70028 13468 70084
rect 13524 70028 13534 70084
rect 15026 70028 15036 70084
rect 15092 70028 20748 70084
rect 20804 70028 20814 70084
rect 21746 70028 21756 70084
rect 21812 70028 23324 70084
rect 23380 70028 23390 70084
rect 25778 70028 25788 70084
rect 25844 70028 26796 70084
rect 26852 70028 27468 70084
rect 27524 70028 27534 70084
rect 15446 69916 15484 69972
rect 15540 69916 15550 69972
rect 15810 69916 15820 69972
rect 15876 69916 26908 69972
rect 26964 69916 26974 69972
rect 9398 69804 9436 69860
rect 9492 69804 9502 69860
rect 12684 69804 13132 69860
rect 13188 69804 13198 69860
rect 4604 69748 4614 69804
rect 4670 69748 4718 69804
rect 4774 69748 4822 69804
rect 4878 69748 4888 69804
rect 11408 69748 11418 69804
rect 11474 69748 11522 69804
rect 11578 69748 11626 69804
rect 11682 69748 11692 69804
rect 12684 69636 12740 69804
rect 18212 69748 18222 69804
rect 18278 69748 18326 69804
rect 18382 69748 18430 69804
rect 18486 69748 18496 69804
rect 25016 69748 25026 69804
rect 25082 69748 25130 69804
rect 25186 69748 25234 69804
rect 25290 69748 25300 69804
rect 12674 69580 12684 69636
rect 12740 69580 12750 69636
rect 13458 69468 13468 69524
rect 13524 69468 14140 69524
rect 14196 69468 15036 69524
rect 15092 69468 15102 69524
rect 15596 69468 15932 69524
rect 15988 69468 16716 69524
rect 16772 69468 16782 69524
rect 18946 69468 18956 69524
rect 19012 69468 19404 69524
rect 19460 69468 19470 69524
rect 15596 69412 15652 69468
rect 13206 69356 13244 69412
rect 13300 69356 13310 69412
rect 14018 69356 14028 69412
rect 14084 69356 14812 69412
rect 14868 69356 15652 69412
rect 16902 69356 16940 69412
rect 16996 69356 17006 69412
rect 17826 69356 17836 69412
rect 17892 69356 17902 69412
rect 0 69300 400 69328
rect 0 69244 1820 69300
rect 1876 69244 1886 69300
rect 9314 69244 9324 69300
rect 9380 69244 15260 69300
rect 15316 69244 15326 69300
rect 16146 69244 16156 69300
rect 16212 69244 16828 69300
rect 16884 69244 16894 69300
rect 0 69216 400 69244
rect 17836 69188 17892 69356
rect 18722 69244 18732 69300
rect 18788 69244 20132 69300
rect 25778 69244 25788 69300
rect 25844 69244 26348 69300
rect 26404 69244 27804 69300
rect 27860 69244 27870 69300
rect 20076 69188 20132 69244
rect 8418 69132 8428 69188
rect 8484 69132 9212 69188
rect 9268 69132 9278 69188
rect 9426 69132 9436 69188
rect 9492 69132 9530 69188
rect 9986 69132 9996 69188
rect 10052 69132 10444 69188
rect 10500 69132 11228 69188
rect 11284 69132 11294 69188
rect 11778 69132 11788 69188
rect 11844 69132 13916 69188
rect 13972 69132 14028 69188
rect 14084 69132 14094 69188
rect 14690 69132 14700 69188
rect 14756 69132 15316 69188
rect 15586 69132 15596 69188
rect 15652 69132 16268 69188
rect 16324 69132 17388 69188
rect 17444 69132 17454 69188
rect 17836 69132 19516 69188
rect 19572 69132 19582 69188
rect 20066 69132 20076 69188
rect 20132 69132 20412 69188
rect 20468 69132 20478 69188
rect 15260 69076 15316 69132
rect 3378 69020 3388 69076
rect 3444 69020 3836 69076
rect 3892 69020 3902 69076
rect 15260 69020 18284 69076
rect 18340 69020 20748 69076
rect 20804 69020 20814 69076
rect 8006 68964 8016 69020
rect 8072 68964 8120 69020
rect 8176 68964 8224 69020
rect 8280 68964 8290 69020
rect 14810 68964 14820 69020
rect 14876 68964 14924 69020
rect 14980 68964 15028 69020
rect 15084 68964 15094 69020
rect 15260 68964 15316 69020
rect 21614 68964 21624 69020
rect 21680 68964 21728 69020
rect 21784 68964 21832 69020
rect 21888 68964 21898 69020
rect 28418 68964 28428 69020
rect 28484 68964 28532 69020
rect 28588 68964 28636 69020
rect 28692 68964 28702 69020
rect 15250 68908 15260 68964
rect 15316 68908 15326 68964
rect 15586 68908 15596 68964
rect 15652 68908 17164 68964
rect 17220 68908 17836 68964
rect 17892 68908 17902 68964
rect 3490 68796 3500 68852
rect 3556 68796 3668 68852
rect 16706 68796 16716 68852
rect 16772 68796 17948 68852
rect 18004 68796 18014 68852
rect 18610 68796 18620 68852
rect 18676 68796 19068 68852
rect 19124 68796 19134 68852
rect 19394 68796 19404 68852
rect 19460 68796 19852 68852
rect 19908 68796 20748 68852
rect 20804 68796 23548 68852
rect 23604 68796 23614 68852
rect 2454 68572 2492 68628
rect 2548 68572 2558 68628
rect 2818 68572 2828 68628
rect 2884 68572 3388 68628
rect 3444 68572 3454 68628
rect 2492 68516 2548 68572
rect 3612 68516 3668 68796
rect 19404 68740 19460 68796
rect 12002 68684 12012 68740
rect 12068 68684 12236 68740
rect 12292 68684 15820 68740
rect 15876 68684 17836 68740
rect 17892 68684 19460 68740
rect 24210 68684 24220 68740
rect 24276 68684 25340 68740
rect 25396 68684 26012 68740
rect 26068 68684 26078 68740
rect 14018 68572 14028 68628
rect 14084 68572 14252 68628
rect 14308 68572 14588 68628
rect 14644 68572 14654 68628
rect 16034 68572 16044 68628
rect 16100 68572 17612 68628
rect 17668 68572 17678 68628
rect 2492 68460 4396 68516
rect 4452 68460 4462 68516
rect 13468 68460 14588 68516
rect 14644 68460 14654 68516
rect 17378 68460 17388 68516
rect 17444 68460 19292 68516
rect 19348 68460 19358 68516
rect 21746 68460 21756 68516
rect 21812 68460 22988 68516
rect 23044 68460 23436 68516
rect 23492 68460 23502 68516
rect 24434 68460 24444 68516
rect 24500 68460 25228 68516
rect 25284 68460 25294 68516
rect 13468 68404 13524 68460
rect 17388 68404 17444 68460
rect 3490 68348 3500 68404
rect 3556 68348 3948 68404
rect 4004 68348 4014 68404
rect 4162 68348 4172 68404
rect 4228 68348 4396 68404
rect 4452 68348 4462 68404
rect 13458 68348 13468 68404
rect 13524 68348 13534 68404
rect 16930 68348 16940 68404
rect 16996 68348 17444 68404
rect 24546 68348 24556 68404
rect 24612 68348 27244 68404
rect 27300 68348 27310 68404
rect 13682 68236 13692 68292
rect 13748 68236 14476 68292
rect 14532 68236 14542 68292
rect 4604 68180 4614 68236
rect 4670 68180 4718 68236
rect 4774 68180 4822 68236
rect 4878 68180 4888 68236
rect 11408 68180 11418 68236
rect 11474 68180 11522 68236
rect 11578 68180 11626 68236
rect 11682 68180 11692 68236
rect 18212 68180 18222 68236
rect 18278 68180 18326 68236
rect 18382 68180 18430 68236
rect 18486 68180 18496 68236
rect 25016 68180 25026 68236
rect 25082 68180 25130 68236
rect 25186 68180 25234 68236
rect 25290 68180 25300 68236
rect 20150 68124 20188 68180
rect 20244 68124 20254 68180
rect 21382 68124 21420 68180
rect 21476 68124 21486 68180
rect 22838 68012 22876 68068
rect 22932 68012 22942 68068
rect 4946 67900 4956 67956
rect 5012 67900 7756 67956
rect 7812 67900 7822 67956
rect 12898 67900 12908 67956
rect 12964 67900 13468 67956
rect 13524 67900 13534 67956
rect 18722 67900 18732 67956
rect 18788 67900 19292 67956
rect 19348 67900 19358 67956
rect 9622 67788 9660 67844
rect 9716 67788 9726 67844
rect 11666 67788 11676 67844
rect 11732 67788 12460 67844
rect 12516 67788 12526 67844
rect 18946 67788 18956 67844
rect 19012 67788 20300 67844
rect 20356 67788 20366 67844
rect 21858 67788 21868 67844
rect 21924 67788 22876 67844
rect 22932 67788 22942 67844
rect 26002 67788 26012 67844
rect 26068 67788 27356 67844
rect 27412 67788 27422 67844
rect 5170 67676 5180 67732
rect 5236 67676 6300 67732
rect 6356 67676 10668 67732
rect 10724 67676 10892 67732
rect 10948 67676 10958 67732
rect 19058 67676 19068 67732
rect 19124 67676 19852 67732
rect 19908 67676 20188 67732
rect 20244 67676 20254 67732
rect 21522 67676 21532 67732
rect 21588 67676 22204 67732
rect 22260 67676 22270 67732
rect 23202 67676 23212 67732
rect 23268 67676 24444 67732
rect 24500 67676 24510 67732
rect 9660 67620 9716 67676
rect 5954 67564 5964 67620
rect 6020 67564 7084 67620
rect 7140 67564 7150 67620
rect 9650 67564 9660 67620
rect 9716 67564 9726 67620
rect 11442 67564 11452 67620
rect 11508 67564 12460 67620
rect 12516 67564 12526 67620
rect 13878 67564 13916 67620
rect 13972 67564 13982 67620
rect 19366 67564 19404 67620
rect 19460 67564 19470 67620
rect 19730 67564 19740 67620
rect 19796 67564 23100 67620
rect 23156 67564 23166 67620
rect 23314 67564 23324 67620
rect 23380 67564 23418 67620
rect 8006 67396 8016 67452
rect 8072 67396 8120 67452
rect 8176 67396 8224 67452
rect 8280 67396 8290 67452
rect 14810 67396 14820 67452
rect 14876 67396 14924 67452
rect 14980 67396 15028 67452
rect 15084 67396 15094 67452
rect 21614 67396 21624 67452
rect 21680 67396 21728 67452
rect 21784 67396 21832 67452
rect 21888 67396 21898 67452
rect 28418 67396 28428 67452
rect 28484 67396 28532 67452
rect 28588 67396 28636 67452
rect 28692 67396 28702 67452
rect 12450 67340 12460 67396
rect 12516 67340 14028 67396
rect 14084 67340 14094 67396
rect 16482 67340 16492 67396
rect 16548 67340 18060 67396
rect 18116 67340 18126 67396
rect 26562 67340 26572 67396
rect 26628 67340 27356 67396
rect 27412 67340 27422 67396
rect 2034 67116 2044 67172
rect 2100 67116 2716 67172
rect 2772 67116 2782 67172
rect 13458 67116 13468 67172
rect 13524 67116 17948 67172
rect 18004 67116 18620 67172
rect 18676 67116 18686 67172
rect 24658 67116 24668 67172
rect 24724 67116 25340 67172
rect 25396 67116 26796 67172
rect 26852 67116 26862 67172
rect 1586 67004 1596 67060
rect 1652 67004 4732 67060
rect 4788 67004 4798 67060
rect 10742 67004 10780 67060
rect 10836 67004 10846 67060
rect 11554 67004 11564 67060
rect 11620 67004 12572 67060
rect 12628 67004 12638 67060
rect 17574 67004 17612 67060
rect 17668 67004 18396 67060
rect 18452 67004 18462 67060
rect 3332 66892 3836 66948
rect 3892 66892 3902 66948
rect 6402 66892 6412 66948
rect 6468 66892 7980 66948
rect 8036 66892 8046 66948
rect 9650 66892 9660 66948
rect 9716 66892 9726 66948
rect 10994 66892 11004 66948
rect 11060 66892 12012 66948
rect 12068 66892 12078 66948
rect 17826 66892 17836 66948
rect 17892 66892 21084 66948
rect 21140 66892 21150 66948
rect 3332 66836 3388 66892
rect 9660 66836 9716 66892
rect 2370 66780 2380 66836
rect 2436 66780 3388 66836
rect 7858 66780 7868 66836
rect 7924 66780 8876 66836
rect 8932 66780 9716 66836
rect 12758 66780 12796 66836
rect 12852 66780 15484 66836
rect 15540 66780 16380 66836
rect 16436 66780 16446 66836
rect 23314 66780 23324 66836
rect 23380 66780 25228 66836
rect 25284 66780 27132 66836
rect 27188 66780 27198 66836
rect 0 66612 400 66640
rect 4604 66612 4614 66668
rect 4670 66612 4718 66668
rect 4774 66612 4822 66668
rect 4878 66612 4888 66668
rect 11408 66612 11418 66668
rect 11474 66612 11522 66668
rect 11578 66612 11626 66668
rect 11682 66612 11692 66668
rect 18212 66612 18222 66668
rect 18278 66612 18326 66668
rect 18382 66612 18430 66668
rect 18486 66612 18496 66668
rect 25016 66612 25026 66668
rect 25082 66612 25130 66668
rect 25186 66612 25234 66668
rect 25290 66612 25300 66668
rect 0 66556 1708 66612
rect 1764 66556 1774 66612
rect 20738 66556 20748 66612
rect 20804 66556 21196 66612
rect 21252 66556 21262 66612
rect 0 66528 400 66556
rect 8978 66444 8988 66500
rect 9044 66444 9548 66500
rect 9604 66444 9614 66500
rect 13542 66444 13580 66500
rect 13636 66444 13646 66500
rect 8306 66332 8316 66388
rect 8372 66332 12908 66388
rect 12964 66332 15148 66388
rect 15250 66332 15260 66388
rect 15316 66332 16380 66388
rect 16436 66332 16446 66388
rect 15092 66276 15148 66332
rect 13458 66220 13468 66276
rect 13524 66220 13534 66276
rect 13794 66220 13804 66276
rect 13860 66220 14252 66276
rect 14308 66220 14318 66276
rect 15092 66220 21084 66276
rect 21140 66220 22876 66276
rect 22932 66220 23436 66276
rect 23492 66220 23502 66276
rect 13468 66164 13524 66220
rect 5170 66108 5180 66164
rect 5236 66108 6076 66164
rect 6132 66108 6142 66164
rect 13468 66108 16828 66164
rect 16884 66108 16894 66164
rect 17500 66108 18956 66164
rect 19012 66108 19022 66164
rect 22082 66108 22092 66164
rect 22148 66108 22540 66164
rect 22596 66108 22606 66164
rect 13692 66052 13748 66108
rect 17500 66052 17556 66108
rect 5842 65996 5852 66052
rect 5908 65996 6860 66052
rect 6916 65996 6926 66052
rect 13682 65996 13692 66052
rect 13748 65996 13758 66052
rect 16370 65996 16380 66052
rect 16436 65996 17500 66052
rect 17556 65996 17566 66052
rect 18946 65996 18956 66052
rect 19012 65996 19068 66052
rect 19124 65996 19404 66052
rect 19460 65996 19470 66052
rect 20514 65996 20524 66052
rect 20580 65996 20748 66052
rect 20804 65996 21532 66052
rect 21588 65996 21598 66052
rect 8006 65828 8016 65884
rect 8072 65828 8120 65884
rect 8176 65828 8224 65884
rect 8280 65828 8290 65884
rect 14810 65828 14820 65884
rect 14876 65828 14924 65884
rect 14980 65828 15028 65884
rect 15084 65828 15094 65884
rect 21614 65828 21624 65884
rect 21680 65828 21728 65884
rect 21784 65828 21832 65884
rect 21888 65828 21898 65884
rect 28418 65828 28428 65884
rect 28484 65828 28532 65884
rect 28588 65828 28636 65884
rect 28692 65828 28702 65884
rect 2818 65772 2828 65828
rect 2884 65772 3500 65828
rect 3556 65772 3566 65828
rect 14354 65772 14364 65828
rect 14420 65772 14476 65828
rect 14532 65772 14542 65828
rect 22390 65772 22428 65828
rect 22484 65772 22494 65828
rect 23986 65772 23996 65828
rect 24052 65772 24668 65828
rect 24724 65772 24734 65828
rect 6514 65660 6524 65716
rect 6580 65660 7420 65716
rect 7476 65660 7486 65716
rect 12450 65660 12460 65716
rect 12516 65660 15540 65716
rect 21298 65660 21308 65716
rect 21364 65660 21980 65716
rect 22036 65660 22764 65716
rect 22820 65660 22830 65716
rect 14588 65604 14644 65660
rect 3042 65548 3052 65604
rect 3108 65548 3276 65604
rect 3332 65548 4172 65604
rect 4228 65548 4396 65604
rect 4452 65548 4462 65604
rect 13430 65548 13468 65604
rect 13524 65548 13534 65604
rect 14466 65548 14476 65604
rect 14532 65548 14644 65604
rect 15484 65492 15540 65660
rect 17938 65548 17948 65604
rect 18004 65548 18060 65604
rect 18116 65548 18732 65604
rect 18788 65548 18798 65604
rect 19170 65548 19180 65604
rect 19236 65548 19516 65604
rect 19572 65548 19964 65604
rect 20020 65548 20030 65604
rect 22306 65548 22316 65604
rect 22372 65548 23100 65604
rect 23156 65548 23166 65604
rect 25442 65548 25452 65604
rect 25508 65548 27916 65604
rect 27972 65548 27982 65604
rect 2454 65436 2492 65492
rect 2548 65436 2558 65492
rect 7186 65436 7196 65492
rect 7252 65436 7644 65492
rect 7700 65436 8428 65492
rect 8484 65436 8494 65492
rect 12674 65436 12684 65492
rect 12740 65436 14364 65492
rect 14420 65436 14430 65492
rect 15474 65436 15484 65492
rect 15540 65436 15550 65492
rect 17266 65436 17276 65492
rect 17332 65436 18508 65492
rect 18564 65436 18574 65492
rect 22418 65436 22428 65492
rect 22484 65436 23996 65492
rect 24052 65436 24444 65492
rect 24500 65436 24510 65492
rect 24770 65436 24780 65492
rect 24836 65436 25788 65492
rect 25844 65436 26908 65492
rect 26964 65436 27804 65492
rect 27860 65436 27870 65492
rect 3826 65324 3836 65380
rect 3892 65324 4620 65380
rect 4676 65324 4686 65380
rect 13122 65324 13132 65380
rect 13188 65324 13804 65380
rect 13860 65324 13870 65380
rect 14018 65324 14028 65380
rect 14084 65324 14812 65380
rect 14868 65324 14878 65380
rect 18274 65324 18284 65380
rect 18340 65324 23268 65380
rect 25554 65324 25564 65380
rect 25620 65324 26124 65380
rect 26180 65324 27356 65380
rect 27412 65324 27422 65380
rect 23212 65268 23268 65324
rect 4274 65212 4284 65268
rect 4340 65212 4350 65268
rect 23202 65212 23212 65268
rect 23268 65212 23278 65268
rect 23538 65212 23548 65268
rect 23604 65212 24444 65268
rect 24500 65212 24510 65268
rect 4284 64820 4340 65212
rect 23548 65156 23604 65212
rect 21858 65100 21868 65156
rect 21924 65100 23324 65156
rect 23380 65100 23604 65156
rect 4604 65044 4614 65100
rect 4670 65044 4718 65100
rect 4774 65044 4822 65100
rect 4878 65044 4888 65100
rect 11408 65044 11418 65100
rect 11474 65044 11522 65100
rect 11578 65044 11626 65100
rect 11682 65044 11692 65100
rect 18212 65044 18222 65100
rect 18278 65044 18326 65100
rect 18382 65044 18430 65100
rect 18486 65044 18496 65100
rect 25016 65044 25026 65100
rect 25082 65044 25130 65100
rect 25186 65044 25234 65100
rect 25290 65044 25300 65100
rect 20290 64876 20300 64932
rect 20356 64876 21308 64932
rect 21364 64876 21374 64932
rect 21522 64876 21532 64932
rect 21588 64876 27020 64932
rect 27076 64876 27086 64932
rect 4274 64764 4284 64820
rect 4340 64764 4350 64820
rect 5730 64764 5740 64820
rect 5796 64764 6636 64820
rect 6692 64764 8988 64820
rect 9044 64764 9436 64820
rect 9492 64764 9502 64820
rect 12236 64764 13748 64820
rect 15586 64764 15596 64820
rect 15652 64764 22316 64820
rect 22372 64764 22382 64820
rect 22866 64764 22876 64820
rect 22932 64764 24220 64820
rect 24276 64764 24286 64820
rect 12236 64708 12292 64764
rect 4134 64652 4172 64708
rect 4228 64652 4238 64708
rect 7186 64652 7196 64708
rect 7252 64652 12292 64708
rect 13692 64596 13748 64764
rect 17238 64652 17276 64708
rect 17332 64652 17342 64708
rect 19618 64652 19628 64708
rect 19684 64652 20524 64708
rect 20580 64652 20590 64708
rect 22754 64652 22764 64708
rect 22820 64652 26348 64708
rect 26404 64652 26414 64708
rect 1698 64540 1708 64596
rect 1764 64540 1932 64596
rect 1988 64540 1998 64596
rect 2258 64540 2268 64596
rect 2324 64540 3052 64596
rect 3108 64540 4620 64596
rect 4676 64540 4686 64596
rect 10322 64540 10332 64596
rect 10388 64540 11228 64596
rect 11284 64540 11788 64596
rect 13692 64540 19964 64596
rect 20020 64540 20030 64596
rect 20738 64540 20748 64596
rect 20804 64540 22092 64596
rect 22148 64540 22158 64596
rect 11732 64484 11788 64540
rect 19964 64484 20020 64540
rect 2034 64428 2044 64484
rect 2100 64428 2828 64484
rect 2884 64428 3948 64484
rect 4004 64428 4014 64484
rect 6066 64428 6076 64484
rect 6132 64428 9884 64484
rect 9940 64428 10444 64484
rect 10500 64428 10510 64484
rect 11732 64428 13468 64484
rect 13524 64428 14252 64484
rect 14308 64428 14318 64484
rect 16594 64428 16604 64484
rect 16660 64428 17388 64484
rect 17444 64428 17454 64484
rect 19964 64428 20972 64484
rect 21028 64428 21038 64484
rect 21420 64428 25564 64484
rect 25620 64428 25900 64484
rect 25956 64428 25966 64484
rect 9202 64316 9212 64372
rect 9268 64316 13356 64372
rect 13412 64316 13422 64372
rect 19170 64316 19180 64372
rect 19236 64316 19246 64372
rect 8006 64260 8016 64316
rect 8072 64260 8120 64316
rect 8176 64260 8224 64316
rect 8280 64260 8290 64316
rect 14810 64260 14820 64316
rect 14876 64260 14924 64316
rect 14980 64260 15028 64316
rect 15084 64260 15094 64316
rect 19180 64260 19236 64316
rect 13122 64204 13132 64260
rect 13188 64204 13198 64260
rect 19180 64204 19404 64260
rect 19460 64204 20748 64260
rect 20804 64204 20814 64260
rect 13132 64148 13188 64204
rect 21420 64148 21476 64428
rect 21614 64260 21624 64316
rect 21680 64260 21728 64316
rect 21784 64260 21832 64316
rect 21888 64260 21898 64316
rect 28418 64260 28428 64316
rect 28484 64260 28532 64316
rect 28588 64260 28636 64316
rect 28692 64260 28702 64316
rect 22306 64204 22316 64260
rect 22372 64204 23436 64260
rect 23492 64204 23502 64260
rect 3266 64092 3276 64148
rect 3332 64092 4172 64148
rect 4228 64092 4238 64148
rect 6402 64092 6412 64148
rect 6468 64092 13188 64148
rect 15092 64092 21476 64148
rect 21858 64092 21868 64148
rect 21924 64092 22876 64148
rect 22932 64092 22942 64148
rect 23492 64092 24668 64148
rect 24724 64092 25116 64148
rect 25172 64092 25182 64148
rect 25666 64092 25676 64148
rect 25732 64092 26012 64148
rect 26068 64092 26078 64148
rect 26562 64092 26572 64148
rect 26628 64092 26684 64148
rect 26740 64092 26750 64148
rect 15092 64036 15148 64092
rect 23492 64036 23548 64092
rect 6178 63980 6188 64036
rect 6244 63980 15148 64036
rect 16482 63980 16492 64036
rect 16548 63980 17724 64036
rect 17780 63980 17790 64036
rect 21298 63980 21308 64036
rect 21364 63980 22428 64036
rect 22484 63980 22494 64036
rect 23100 63980 23548 64036
rect 25116 64036 25172 64092
rect 25116 63980 27468 64036
rect 27524 63980 28028 64036
rect 28084 63980 28094 64036
rect 0 63924 400 63952
rect 23100 63924 23156 63980
rect 0 63868 1820 63924
rect 1876 63868 1886 63924
rect 2706 63868 2716 63924
rect 2772 63868 3724 63924
rect 3780 63868 3790 63924
rect 4498 63868 4508 63924
rect 4564 63868 5180 63924
rect 5236 63868 5246 63924
rect 6066 63868 6076 63924
rect 6132 63868 7084 63924
rect 7140 63868 7150 63924
rect 7410 63868 7420 63924
rect 7476 63868 8820 63924
rect 8978 63868 8988 63924
rect 9044 63868 9660 63924
rect 9716 63868 10108 63924
rect 10164 63868 12012 63924
rect 12068 63868 12684 63924
rect 12740 63868 13356 63924
rect 13412 63868 13422 63924
rect 17378 63868 17388 63924
rect 17444 63868 23100 63924
rect 23156 63868 23166 63924
rect 23762 63868 23772 63924
rect 23828 63868 24220 63924
rect 24276 63868 25788 63924
rect 25844 63868 25854 63924
rect 0 63840 400 63868
rect 8764 63812 8820 63868
rect 26012 63812 26068 63980
rect 3042 63756 3052 63812
rect 3108 63756 3500 63812
rect 3556 63756 3566 63812
rect 6626 63756 6636 63812
rect 6692 63756 7532 63812
rect 7588 63756 7598 63812
rect 8764 63756 8876 63812
rect 8932 63756 9996 63812
rect 10052 63756 10062 63812
rect 17836 63756 20356 63812
rect 20514 63756 20524 63812
rect 20580 63756 21756 63812
rect 21812 63756 21822 63812
rect 23426 63756 23436 63812
rect 23492 63756 24108 63812
rect 24164 63756 24174 63812
rect 25666 63756 25676 63812
rect 25732 63756 26068 63812
rect 26852 63756 27132 63812
rect 27188 63756 27198 63812
rect 17836 63700 17892 63756
rect 9622 63644 9660 63700
rect 9716 63644 9726 63700
rect 13570 63644 13580 63700
rect 13636 63644 13916 63700
rect 13972 63644 13982 63700
rect 14924 63644 15260 63700
rect 15316 63644 17892 63700
rect 14924 63588 14980 63644
rect 20300 63588 20356 63756
rect 26852 63700 26908 63756
rect 20738 63644 20748 63700
rect 20804 63644 20972 63700
rect 21028 63644 21644 63700
rect 21700 63644 22092 63700
rect 22148 63644 22876 63700
rect 22932 63644 22942 63700
rect 26450 63644 26460 63700
rect 26516 63644 26908 63700
rect 27234 63644 27244 63700
rect 27300 63644 28140 63700
rect 28196 63644 28206 63700
rect 14914 63532 14924 63588
rect 14980 63532 14990 63588
rect 18722 63532 18732 63588
rect 18788 63532 19292 63588
rect 19348 63532 19358 63588
rect 20300 63532 22316 63588
rect 22372 63532 24780 63588
rect 24836 63532 24846 63588
rect 26674 63532 26684 63588
rect 26740 63532 26796 63588
rect 26852 63532 26862 63588
rect 4604 63476 4614 63532
rect 4670 63476 4718 63532
rect 4774 63476 4822 63532
rect 4878 63476 4888 63532
rect 11408 63476 11418 63532
rect 11474 63476 11522 63532
rect 11578 63476 11626 63532
rect 11682 63476 11692 63532
rect 18212 63476 18222 63532
rect 18278 63476 18326 63532
rect 18382 63476 18430 63532
rect 18486 63476 18496 63532
rect 25016 63476 25026 63532
rect 25082 63476 25130 63532
rect 25186 63476 25234 63532
rect 25290 63476 25300 63532
rect 5058 63420 5068 63476
rect 5124 63420 5852 63476
rect 5908 63420 5918 63476
rect 15810 63420 15820 63476
rect 15876 63420 16268 63476
rect 16324 63420 16334 63476
rect 22866 63420 22876 63476
rect 22932 63420 23100 63476
rect 23156 63420 23166 63476
rect 6626 63308 6636 63364
rect 6692 63308 14476 63364
rect 14532 63308 15260 63364
rect 15316 63308 15484 63364
rect 15540 63308 15550 63364
rect 16370 63308 16380 63364
rect 16436 63308 16828 63364
rect 16884 63308 16894 63364
rect 18162 63308 18172 63364
rect 18228 63308 18956 63364
rect 19012 63308 19022 63364
rect 3714 63196 3724 63252
rect 3780 63196 4620 63252
rect 4676 63196 4686 63252
rect 9650 63196 9660 63252
rect 9716 63196 10220 63252
rect 10276 63196 10286 63252
rect 11554 63196 11564 63252
rect 11620 63196 17612 63252
rect 17668 63196 17678 63252
rect 25890 63196 25900 63252
rect 25956 63196 26348 63252
rect 26404 63196 27020 63252
rect 27076 63196 27086 63252
rect 11778 63084 11788 63140
rect 11844 63084 12236 63140
rect 12292 63084 12302 63140
rect 12450 63084 12460 63140
rect 12516 63084 13020 63140
rect 13076 63084 13468 63140
rect 13524 63084 13534 63140
rect 13906 63084 13916 63140
rect 13972 63084 16268 63140
rect 16324 63084 16334 63140
rect 17126 63084 17164 63140
rect 17220 63084 17230 63140
rect 19058 63084 19068 63140
rect 19124 63084 19180 63140
rect 19236 63084 19628 63140
rect 19684 63084 19694 63140
rect 20066 63084 20076 63140
rect 20132 63084 26796 63140
rect 26852 63084 26862 63140
rect 20076 63028 20132 63084
rect 3154 62972 3164 63028
rect 3220 62972 18620 63028
rect 18676 62972 20132 63028
rect 22866 62972 22876 63028
rect 22932 62972 23660 63028
rect 23716 62972 23726 63028
rect 24322 62972 24332 63028
rect 24388 62972 27244 63028
rect 27300 62972 27310 63028
rect 3938 62860 3948 62916
rect 4004 62860 4956 62916
rect 5012 62860 5022 62916
rect 8418 62860 8428 62916
rect 8484 62860 12684 62916
rect 12740 62860 14028 62916
rect 14084 62860 16100 62916
rect 16230 62860 16268 62916
rect 16324 62860 16334 62916
rect 16492 62860 23436 62916
rect 23492 62860 23502 62916
rect 26562 62860 26572 62916
rect 26628 62860 27356 62916
rect 27412 62860 27422 62916
rect 16044 62804 16100 62860
rect 16492 62804 16548 62860
rect 8754 62748 8764 62804
rect 8820 62748 11228 62804
rect 11284 62748 12460 62804
rect 12516 62748 12526 62804
rect 16044 62748 16548 62804
rect 16818 62748 16828 62804
rect 16884 62748 17500 62804
rect 17556 62748 17566 62804
rect 8006 62692 8016 62748
rect 8072 62692 8120 62748
rect 8176 62692 8224 62748
rect 8280 62692 8290 62748
rect 14810 62692 14820 62748
rect 14876 62692 14924 62748
rect 14980 62692 15028 62748
rect 15084 62692 15094 62748
rect 21614 62692 21624 62748
rect 21680 62692 21728 62748
rect 21784 62692 21832 62748
rect 21888 62692 21898 62748
rect 28418 62692 28428 62748
rect 28484 62692 28532 62748
rect 28588 62692 28636 62748
rect 28692 62692 28702 62748
rect 9212 62636 10108 62692
rect 10164 62636 10174 62692
rect 11218 62636 11228 62692
rect 11284 62636 13916 62692
rect 13972 62636 13982 62692
rect 17154 62636 17164 62692
rect 17220 62636 17724 62692
rect 17780 62636 17790 62692
rect 19702 62636 19740 62692
rect 19796 62636 19806 62692
rect 6738 62524 6748 62580
rect 6804 62524 7980 62580
rect 8036 62524 8428 62580
rect 8484 62524 8494 62580
rect 9212 62468 9268 62636
rect 9986 62524 9996 62580
rect 10052 62524 11004 62580
rect 11060 62524 12236 62580
rect 12292 62524 13020 62580
rect 13076 62524 13086 62580
rect 14242 62524 14252 62580
rect 14308 62524 19292 62580
rect 19348 62524 19358 62580
rect 20626 62524 20636 62580
rect 20692 62524 23100 62580
rect 23156 62524 23166 62580
rect 20636 62468 20692 62524
rect 8306 62412 8316 62468
rect 8372 62412 9268 62468
rect 9324 62412 18396 62468
rect 18452 62412 19180 62468
rect 19236 62412 20692 62468
rect 6514 62300 6524 62356
rect 6580 62300 7084 62356
rect 7140 62300 7756 62356
rect 7812 62300 8764 62356
rect 8820 62300 8830 62356
rect 9324 62244 9380 62412
rect 12674 62300 12684 62356
rect 12740 62300 14364 62356
rect 14420 62300 14430 62356
rect 14588 62300 15372 62356
rect 15428 62300 15438 62356
rect 15586 62300 15596 62356
rect 15652 62300 16044 62356
rect 16100 62300 16110 62356
rect 16818 62300 16828 62356
rect 16884 62300 18620 62356
rect 18676 62300 18686 62356
rect 14588 62244 14644 62300
rect 5842 62188 5852 62244
rect 5908 62188 6636 62244
rect 6692 62188 9380 62244
rect 14466 62188 14476 62244
rect 14532 62188 14644 62244
rect 17462 62188 17500 62244
rect 17556 62188 17566 62244
rect 22082 62188 22092 62244
rect 22148 62188 22428 62244
rect 22484 62188 22494 62244
rect 23202 62188 23212 62244
rect 23268 62188 23548 62244
rect 23604 62188 24220 62244
rect 24276 62188 24286 62244
rect 24658 62188 24668 62244
rect 24724 62188 25228 62244
rect 25284 62188 25294 62244
rect 5170 62076 5180 62132
rect 5236 62076 5964 62132
rect 6020 62076 15148 62132
rect 15362 62076 15372 62132
rect 15428 62076 15820 62132
rect 15876 62076 15886 62132
rect 17602 62076 17612 62132
rect 17668 62076 19572 62132
rect 15092 62020 15148 62076
rect 19516 62020 19572 62076
rect 15092 61964 18116 62020
rect 19506 61964 19516 62020
rect 19572 61964 19582 62020
rect 4604 61908 4614 61964
rect 4670 61908 4718 61964
rect 4774 61908 4822 61964
rect 4878 61908 4888 61964
rect 11408 61908 11418 61964
rect 11474 61908 11522 61964
rect 11578 61908 11626 61964
rect 11682 61908 11692 61964
rect 14354 61852 14364 61908
rect 14420 61852 14476 61908
rect 14532 61852 14542 61908
rect 14700 61852 15932 61908
rect 15988 61852 16828 61908
rect 16884 61852 16894 61908
rect 14700 61796 14756 61852
rect 18060 61796 18116 61964
rect 18212 61908 18222 61964
rect 18278 61908 18326 61964
rect 18382 61908 18430 61964
rect 18486 61908 18496 61964
rect 25016 61908 25026 61964
rect 25082 61908 25130 61964
rect 25186 61908 25234 61964
rect 25290 61908 25300 61964
rect 3490 61740 3500 61796
rect 3556 61740 5292 61796
rect 5348 61740 12124 61796
rect 12180 61740 12190 61796
rect 12338 61740 12348 61796
rect 12404 61740 13580 61796
rect 13636 61740 14756 61796
rect 15558 61740 15596 61796
rect 15652 61740 15662 61796
rect 16930 61740 16940 61796
rect 16996 61740 17724 61796
rect 17780 61740 17790 61796
rect 18060 61740 25340 61796
rect 25396 61740 26236 61796
rect 26292 61740 26302 61796
rect 26852 61684 26908 61796
rect 26964 61740 26974 61796
rect 4386 61628 4396 61684
rect 4452 61628 4620 61684
rect 4676 61628 6188 61684
rect 6244 61628 6254 61684
rect 10546 61628 10556 61684
rect 10612 61628 24108 61684
rect 24164 61628 26908 61684
rect 6066 61516 6076 61572
rect 6132 61516 6860 61572
rect 6916 61516 6926 61572
rect 9986 61516 9996 61572
rect 10052 61516 14924 61572
rect 14980 61516 14990 61572
rect 15250 61516 15260 61572
rect 15316 61516 15372 61572
rect 15428 61516 15438 61572
rect 15586 61516 15596 61572
rect 15652 61516 16604 61572
rect 16660 61516 16670 61572
rect 21410 61516 21420 61572
rect 21476 61516 22652 61572
rect 22708 61516 23324 61572
rect 23380 61516 23390 61572
rect 15596 61460 15652 61516
rect 2034 61404 2044 61460
rect 2100 61404 3276 61460
rect 3332 61404 3342 61460
rect 7074 61404 7084 61460
rect 7140 61404 12124 61460
rect 12180 61404 12190 61460
rect 13346 61404 13356 61460
rect 13412 61404 13916 61460
rect 13972 61404 13982 61460
rect 14140 61404 15652 61460
rect 16258 61404 16268 61460
rect 16324 61404 16828 61460
rect 16884 61404 16894 61460
rect 19506 61404 19516 61460
rect 19572 61404 23996 61460
rect 24052 61404 24062 61460
rect 14140 61348 14196 61404
rect 2370 61292 2380 61348
rect 2436 61292 2716 61348
rect 2772 61292 4172 61348
rect 4228 61292 4238 61348
rect 6738 61292 6748 61348
rect 6804 61292 7532 61348
rect 7588 61292 7598 61348
rect 11778 61292 11788 61348
rect 11844 61292 12348 61348
rect 12404 61292 12414 61348
rect 12674 61292 12684 61348
rect 12740 61292 12796 61348
rect 12852 61292 13132 61348
rect 13188 61292 13198 61348
rect 14130 61292 14140 61348
rect 14196 61292 14206 61348
rect 15260 61292 24332 61348
rect 24388 61292 24398 61348
rect 0 61236 400 61264
rect 0 61180 1708 61236
rect 1764 61180 2492 61236
rect 2548 61180 2558 61236
rect 0 61152 400 61180
rect 8006 61124 8016 61180
rect 8072 61124 8120 61180
rect 8176 61124 8224 61180
rect 8280 61124 8290 61180
rect 14810 61124 14820 61180
rect 14876 61124 14924 61180
rect 14980 61124 15028 61180
rect 15084 61124 15094 61180
rect 5170 61068 5180 61124
rect 5236 61068 5740 61124
rect 5796 61068 5806 61124
rect 15260 61012 15316 61292
rect 16146 61180 16156 61236
rect 16212 61180 17836 61236
rect 17892 61180 20412 61236
rect 20468 61180 20478 61236
rect 22306 61180 22316 61236
rect 22372 61180 25116 61236
rect 25172 61180 25182 61236
rect 21614 61124 21624 61180
rect 21680 61124 21728 61180
rect 21784 61124 21832 61180
rect 21888 61124 21898 61180
rect 28418 61124 28428 61180
rect 28484 61124 28532 61180
rect 28588 61124 28636 61180
rect 28692 61124 28702 61180
rect 16146 61068 16156 61124
rect 16212 61068 16940 61124
rect 16996 61068 18172 61124
rect 18228 61068 18238 61124
rect 9650 60956 9660 61012
rect 9716 60956 10332 61012
rect 10388 60956 10398 61012
rect 14466 60956 14476 61012
rect 14532 60956 15316 61012
rect 15810 60956 15820 61012
rect 15876 60956 17164 61012
rect 17220 60956 17230 61012
rect 11218 60844 11228 60900
rect 11284 60844 11452 60900
rect 11508 60844 11518 60900
rect 19394 60844 19404 60900
rect 19460 60844 20188 60900
rect 20244 60844 20972 60900
rect 21028 60844 21038 60900
rect 25666 60844 25676 60900
rect 25732 60844 26684 60900
rect 26740 60844 26750 60900
rect 7522 60732 7532 60788
rect 7588 60732 8316 60788
rect 8372 60732 8382 60788
rect 8978 60732 8988 60788
rect 9044 60732 10332 60788
rect 10388 60732 10398 60788
rect 12338 60732 12348 60788
rect 12404 60732 13804 60788
rect 13860 60732 14028 60788
rect 14084 60732 14094 60788
rect 14354 60732 14364 60788
rect 14420 60732 17948 60788
rect 18004 60732 18014 60788
rect 18722 60732 18732 60788
rect 18788 60732 19404 60788
rect 19460 60732 19470 60788
rect 19618 60732 19628 60788
rect 19684 60732 19964 60788
rect 20020 60732 20030 60788
rect 20178 60732 20188 60788
rect 20244 60732 21308 60788
rect 21364 60732 21374 60788
rect 2146 60620 2156 60676
rect 2212 60620 3724 60676
rect 3780 60620 3790 60676
rect 9762 60620 9772 60676
rect 9828 60620 10108 60676
rect 10164 60620 10174 60676
rect 12898 60620 12908 60676
rect 12964 60620 16380 60676
rect 16436 60620 17164 60676
rect 17220 60620 21196 60676
rect 21252 60620 21262 60676
rect 22082 60620 22092 60676
rect 22148 60620 22428 60676
rect 22484 60620 23100 60676
rect 23156 60620 23166 60676
rect 2594 60508 2604 60564
rect 2660 60508 3388 60564
rect 3444 60508 3454 60564
rect 3798 60508 3836 60564
rect 3892 60508 3902 60564
rect 4386 60508 4396 60564
rect 4452 60508 5740 60564
rect 5796 60508 5806 60564
rect 10434 60508 10444 60564
rect 10500 60508 10780 60564
rect 10836 60508 10846 60564
rect 14242 60508 14252 60564
rect 14308 60508 14924 60564
rect 14980 60508 14990 60564
rect 15222 60508 15260 60564
rect 15316 60508 15326 60564
rect 16594 60508 16604 60564
rect 16660 60508 17836 60564
rect 17892 60508 17902 60564
rect 18582 60508 18620 60564
rect 18676 60508 18686 60564
rect 19618 60508 19628 60564
rect 19684 60508 20300 60564
rect 20356 60508 20366 60564
rect 20626 60508 20636 60564
rect 20692 60508 21420 60564
rect 21476 60508 21868 60564
rect 21924 60508 21934 60564
rect 20636 60452 20692 60508
rect 6738 60396 6748 60452
rect 6804 60396 11228 60452
rect 11284 60396 11294 60452
rect 14242 60396 14252 60452
rect 14308 60396 17388 60452
rect 17444 60396 17454 60452
rect 17602 60396 17612 60452
rect 17668 60396 17948 60452
rect 18004 60396 18014 60452
rect 20402 60396 20412 60452
rect 20468 60396 20692 60452
rect 22418 60396 22428 60452
rect 22484 60396 23100 60452
rect 23156 60396 23166 60452
rect 4604 60340 4614 60396
rect 4670 60340 4718 60396
rect 4774 60340 4822 60396
rect 4878 60340 4888 60396
rect 11408 60340 11418 60396
rect 11474 60340 11522 60396
rect 11578 60340 11626 60396
rect 11682 60340 11692 60396
rect 18212 60340 18222 60396
rect 18278 60340 18326 60396
rect 18382 60340 18430 60396
rect 18486 60340 18496 60396
rect 25016 60340 25026 60396
rect 25082 60340 25130 60396
rect 25186 60340 25234 60396
rect 25290 60340 25300 60396
rect 12898 60284 12908 60340
rect 12964 60284 15372 60340
rect 15428 60284 16268 60340
rect 16324 60284 16334 60340
rect 19506 60284 19516 60340
rect 19572 60284 20076 60340
rect 20132 60284 20142 60340
rect 22726 60284 22764 60340
rect 22820 60284 22830 60340
rect 5730 60172 5740 60228
rect 5796 60172 8428 60228
rect 8484 60172 8988 60228
rect 9044 60172 9054 60228
rect 13682 60172 13692 60228
rect 13748 60172 15484 60228
rect 15540 60172 15550 60228
rect 17238 60172 17276 60228
rect 17332 60172 17342 60228
rect 23762 60172 23772 60228
rect 23828 60172 24780 60228
rect 24836 60172 24846 60228
rect 26674 60172 26684 60228
rect 26740 60172 28028 60228
rect 28084 60172 28094 60228
rect 7858 60060 7868 60116
rect 7924 60060 8540 60116
rect 8596 60060 8606 60116
rect 14242 60060 14252 60116
rect 14308 60060 21644 60116
rect 21700 60060 23660 60116
rect 23716 60060 23726 60116
rect 26338 60060 26348 60116
rect 26404 60060 26796 60116
rect 26852 60060 28140 60116
rect 28196 60060 28206 60116
rect 11732 59948 11900 60004
rect 11956 59948 11966 60004
rect 14326 59948 14364 60004
rect 14420 59948 14430 60004
rect 18162 59948 18172 60004
rect 18228 59948 20076 60004
rect 20132 59948 20142 60004
rect 24546 59948 24556 60004
rect 24612 59948 25340 60004
rect 25396 59948 25406 60004
rect 3266 59836 3276 59892
rect 3332 59836 4620 59892
rect 4676 59836 4686 59892
rect 11732 59780 11788 59948
rect 13906 59836 13916 59892
rect 13972 59836 17500 59892
rect 17556 59836 17566 59892
rect 19170 59836 19180 59892
rect 19236 59836 20636 59892
rect 20692 59836 20702 59892
rect 22754 59836 22764 59892
rect 22820 59836 23772 59892
rect 23828 59836 23838 59892
rect 10434 59724 10444 59780
rect 10500 59724 11788 59780
rect 11844 59724 11854 59780
rect 13794 59724 13804 59780
rect 13860 59724 14028 59780
rect 14084 59724 14140 59780
rect 14196 59724 14206 59780
rect 16118 59724 16156 59780
rect 16212 59724 16222 59780
rect 18498 59724 18508 59780
rect 18564 59724 22428 59780
rect 22484 59724 22494 59780
rect 19058 59612 19068 59668
rect 19124 59612 19180 59668
rect 19236 59612 19246 59668
rect 8006 59556 8016 59612
rect 8072 59556 8120 59612
rect 8176 59556 8224 59612
rect 8280 59556 8290 59612
rect 14810 59556 14820 59612
rect 14876 59556 14924 59612
rect 14980 59556 15028 59612
rect 15084 59556 15094 59612
rect 21614 59556 21624 59612
rect 21680 59556 21728 59612
rect 21784 59556 21832 59612
rect 21888 59556 21898 59612
rect 28418 59556 28428 59612
rect 28484 59556 28532 59612
rect 28588 59556 28636 59612
rect 28692 59556 28702 59612
rect 5170 59388 5180 59444
rect 5236 59388 5740 59444
rect 5796 59388 7420 59444
rect 7476 59388 7486 59444
rect 8530 59388 8540 59444
rect 8596 59388 9884 59444
rect 9940 59388 9950 59444
rect 14802 59388 14812 59444
rect 14868 59388 16156 59444
rect 16212 59388 16222 59444
rect 22642 59388 22652 59444
rect 22708 59388 23436 59444
rect 23492 59388 23502 59444
rect 24546 59388 24556 59444
rect 24612 59388 26236 59444
rect 26292 59388 26302 59444
rect 26572 59388 26908 59444
rect 26964 59388 26974 59444
rect 7420 59332 7476 59388
rect 7420 59276 8932 59332
rect 9090 59276 9100 59332
rect 9156 59276 10444 59332
rect 10500 59276 10510 59332
rect 14690 59276 14700 59332
rect 14756 59276 17500 59332
rect 17556 59276 17566 59332
rect 18946 59276 18956 59332
rect 19012 59276 20300 59332
rect 20356 59276 20366 59332
rect 8876 59220 8932 59276
rect 26572 59220 26628 59388
rect 26852 59276 27356 59332
rect 27412 59276 27422 59332
rect 6514 59164 6524 59220
rect 6580 59164 6860 59220
rect 6916 59164 7756 59220
rect 7812 59164 7822 59220
rect 8876 59164 9660 59220
rect 9716 59164 9726 59220
rect 14018 59164 14028 59220
rect 14084 59164 15036 59220
rect 15092 59164 15102 59220
rect 16818 59164 16828 59220
rect 16884 59164 18172 59220
rect 18228 59164 18238 59220
rect 22978 59164 22988 59220
rect 23044 59164 23548 59220
rect 23604 59164 23614 59220
rect 26226 59164 26236 59220
rect 26292 59164 26572 59220
rect 26628 59164 26638 59220
rect 26852 59108 26908 59276
rect 6178 59052 6188 59108
rect 6244 59052 6748 59108
rect 6804 59052 6814 59108
rect 15820 59052 15932 59108
rect 15988 59052 15998 59108
rect 23426 59052 23436 59108
rect 23492 59052 24444 59108
rect 24500 59052 24510 59108
rect 25890 59052 25900 59108
rect 25956 59052 26908 59108
rect 15820 58996 15876 59052
rect 4610 58940 4620 58996
rect 4676 58940 11900 58996
rect 11956 58940 11966 58996
rect 12898 58940 12908 58996
rect 12964 58940 13356 58996
rect 13412 58940 13422 58996
rect 15810 58940 15820 58996
rect 15876 58940 15886 58996
rect 10434 58828 10444 58884
rect 10500 58828 10780 58884
rect 10836 58828 10846 58884
rect 14466 58828 14476 58884
rect 14532 58828 15260 58884
rect 15316 58828 15596 58884
rect 15652 58828 15662 58884
rect 19506 58828 19516 58884
rect 19572 58828 21532 58884
rect 21588 58828 22092 58884
rect 22148 58828 22158 58884
rect 25442 58828 25452 58884
rect 25508 58828 26684 58884
rect 26740 58828 26750 58884
rect 4604 58772 4614 58828
rect 4670 58772 4718 58828
rect 4774 58772 4822 58828
rect 4878 58772 4888 58828
rect 11408 58772 11418 58828
rect 11474 58772 11522 58828
rect 11578 58772 11626 58828
rect 11682 58772 11692 58828
rect 18212 58772 18222 58828
rect 18278 58772 18326 58828
rect 18382 58772 18430 58828
rect 18486 58772 18496 58828
rect 25016 58772 25026 58828
rect 25082 58772 25130 58828
rect 25186 58772 25234 58828
rect 25290 58772 25300 58828
rect 4134 58716 4172 58772
rect 4228 58716 4238 58772
rect 13570 58716 13580 58772
rect 13636 58716 15484 58772
rect 15540 58716 15932 58772
rect 15988 58716 15998 58772
rect 2370 58604 2380 58660
rect 2436 58604 2772 58660
rect 2930 58604 2940 58660
rect 2996 58604 3724 58660
rect 3780 58604 3790 58660
rect 11778 58604 11788 58660
rect 11844 58604 12572 58660
rect 12628 58604 12638 58660
rect 14466 58604 14476 58660
rect 14532 58604 15036 58660
rect 15092 58604 16380 58660
rect 16436 58604 16446 58660
rect 20626 58604 20636 58660
rect 20692 58604 25676 58660
rect 25732 58604 25742 58660
rect 0 58548 400 58576
rect 2716 58548 2772 58604
rect 0 58492 1708 58548
rect 1764 58492 2492 58548
rect 2548 58492 2558 58548
rect 2716 58492 2828 58548
rect 2884 58492 4620 58548
rect 4676 58492 4686 58548
rect 7746 58492 7756 58548
rect 7812 58492 10556 58548
rect 10612 58492 11396 58548
rect 13010 58492 13020 58548
rect 13076 58492 13356 58548
rect 13412 58492 13422 58548
rect 13794 58492 13804 58548
rect 13860 58492 22316 58548
rect 22372 58492 22382 58548
rect 22866 58492 22876 58548
rect 22932 58492 23772 58548
rect 23828 58492 24892 58548
rect 24948 58492 25900 58548
rect 25956 58492 25966 58548
rect 0 58464 400 58492
rect 2034 58380 2044 58436
rect 2100 58380 5628 58436
rect 5684 58380 5694 58436
rect 9090 58380 9100 58436
rect 9156 58380 10892 58436
rect 10948 58380 10958 58436
rect 2716 58268 4060 58324
rect 4116 58268 4126 58324
rect 2716 58212 2772 58268
rect 4284 58212 4340 58380
rect 11340 58324 11396 58492
rect 14578 58380 14588 58436
rect 14644 58380 15148 58436
rect 15204 58380 15214 58436
rect 16342 58380 16380 58436
rect 16436 58380 16446 58436
rect 8838 58268 8876 58324
rect 8932 58268 8942 58324
rect 9202 58268 9212 58324
rect 9268 58268 9548 58324
rect 9604 58268 9614 58324
rect 10518 58268 10556 58324
rect 10612 58268 10622 58324
rect 11330 58268 11340 58324
rect 11396 58268 11406 58324
rect 12562 58268 12572 58324
rect 12628 58268 12638 58324
rect 14018 58268 14028 58324
rect 14084 58268 14364 58324
rect 14420 58268 17052 58324
rect 17108 58268 18396 58324
rect 18452 58268 18462 58324
rect 24434 58268 24444 58324
rect 24500 58268 27244 58324
rect 27300 58268 27310 58324
rect 12572 58212 12628 58268
rect 2258 58156 2268 58212
rect 2324 58156 2716 58212
rect 2772 58156 2782 58212
rect 3826 58156 3836 58212
rect 3892 58156 4340 58212
rect 7522 58156 7532 58212
rect 7588 58156 11004 58212
rect 11060 58156 20188 58212
rect 20244 58156 20254 58212
rect 21074 58156 21084 58212
rect 21140 58156 22316 58212
rect 22372 58156 22382 58212
rect 24098 58156 24108 58212
rect 24164 58156 24892 58212
rect 24948 58156 24958 58212
rect 9650 58044 9660 58100
rect 9716 58044 12012 58100
rect 12068 58044 14364 58100
rect 14420 58044 14430 58100
rect 8006 57988 8016 58044
rect 8072 57988 8120 58044
rect 8176 57988 8224 58044
rect 8280 57988 8290 58044
rect 14810 57988 14820 58044
rect 14876 57988 14924 58044
rect 14980 57988 15028 58044
rect 15084 57988 15094 58044
rect 21614 57988 21624 58044
rect 21680 57988 21728 58044
rect 21784 57988 21832 58044
rect 21888 57988 21898 58044
rect 28418 57988 28428 58044
rect 28484 57988 28532 58044
rect 28588 57988 28636 58044
rect 28692 57988 28702 58044
rect 5814 57932 5852 57988
rect 5908 57932 5918 57988
rect 8978 57932 8988 57988
rect 9044 57932 12236 57988
rect 12292 57932 12302 57988
rect 12450 57932 12460 57988
rect 12516 57932 12554 57988
rect 13244 57932 14644 57988
rect 15250 57932 15260 57988
rect 15316 57932 15354 57988
rect 23398 57932 23436 57988
rect 23492 57932 23502 57988
rect 13244 57876 13300 57932
rect 14588 57876 14644 57932
rect 1810 57820 1820 57876
rect 1876 57820 5068 57876
rect 5124 57820 5134 57876
rect 6290 57820 6300 57876
rect 6356 57820 6636 57876
rect 6692 57820 7084 57876
rect 7140 57820 7150 57876
rect 8530 57820 8540 57876
rect 8596 57820 10108 57876
rect 10164 57820 13300 57876
rect 13458 57820 13468 57876
rect 13524 57820 13692 57876
rect 13748 57820 13758 57876
rect 14588 57820 23996 57876
rect 24052 57820 24444 57876
rect 24500 57820 24510 57876
rect 6066 57708 6076 57764
rect 6132 57708 6300 57764
rect 6356 57708 12180 57764
rect 13122 57708 13132 57764
rect 13188 57708 17500 57764
rect 17556 57708 17566 57764
rect 19394 57708 19404 57764
rect 19460 57708 19964 57764
rect 20020 57708 20030 57764
rect 20178 57708 20188 57764
rect 20244 57708 20748 57764
rect 20804 57708 21644 57764
rect 21700 57708 21710 57764
rect 23492 57708 23884 57764
rect 23940 57708 23950 57764
rect 25554 57708 25564 57764
rect 25620 57708 26236 57764
rect 26292 57708 26302 57764
rect 10658 57596 10668 57652
rect 10724 57596 11340 57652
rect 11396 57596 11406 57652
rect 12124 57540 12180 57708
rect 16482 57596 16492 57652
rect 16548 57596 16828 57652
rect 16884 57596 17836 57652
rect 17892 57596 17902 57652
rect 23426 57596 23436 57652
rect 23492 57596 23548 57708
rect 26450 57596 26460 57652
rect 26516 57596 26908 57652
rect 26964 57596 26974 57652
rect 10322 57484 10332 57540
rect 10388 57484 11116 57540
rect 11172 57484 11900 57540
rect 11956 57484 11966 57540
rect 12124 57484 19852 57540
rect 19908 57484 19918 57540
rect 22530 57484 22540 57540
rect 22596 57484 23212 57540
rect 23268 57484 23278 57540
rect 10780 57372 13580 57428
rect 13636 57372 13646 57428
rect 14140 57372 14588 57428
rect 14644 57372 14654 57428
rect 23762 57372 23772 57428
rect 23828 57372 24444 57428
rect 24500 57372 25340 57428
rect 25396 57372 26460 57428
rect 26516 57372 26796 57428
rect 26852 57372 26862 57428
rect 3602 57260 3612 57316
rect 3668 57260 3724 57316
rect 3780 57260 3790 57316
rect 5618 57260 5628 57316
rect 5684 57260 7532 57316
rect 7588 57260 7598 57316
rect 4604 57204 4614 57260
rect 4670 57204 4718 57260
rect 4774 57204 4822 57260
rect 4878 57204 4888 57260
rect 10780 57204 10836 57372
rect 14140 57316 14196 57372
rect 13682 57260 13692 57316
rect 13748 57260 14196 57316
rect 14354 57260 14364 57316
rect 14420 57260 18116 57316
rect 24070 57260 24108 57316
rect 24164 57260 24174 57316
rect 11408 57204 11418 57260
rect 11474 57204 11522 57260
rect 11578 57204 11626 57260
rect 11682 57204 11692 57260
rect 6066 57148 6076 57204
rect 6132 57148 6142 57204
rect 10770 57148 10780 57204
rect 10836 57148 10846 57204
rect 12226 57148 12236 57204
rect 12292 57148 12684 57204
rect 12740 57148 12750 57204
rect 14130 57148 14140 57204
rect 14196 57148 15484 57204
rect 15540 57148 15550 57204
rect 6076 57092 6132 57148
rect 18060 57092 18116 57260
rect 18212 57204 18222 57260
rect 18278 57204 18326 57260
rect 18382 57204 18430 57260
rect 18486 57204 18496 57260
rect 25016 57204 25026 57260
rect 25082 57204 25130 57260
rect 25186 57204 25234 57260
rect 25290 57204 25300 57260
rect 18620 57148 19180 57204
rect 19236 57148 19852 57204
rect 19908 57148 19918 57204
rect 21970 57148 21980 57204
rect 22036 57148 22204 57204
rect 22260 57148 22270 57204
rect 23202 57148 23212 57204
rect 23268 57148 24332 57204
rect 24388 57148 24668 57204
rect 24724 57148 24734 57204
rect 18620 57092 18676 57148
rect 3154 57036 3164 57092
rect 3220 57036 3500 57092
rect 3556 57036 3566 57092
rect 6076 57036 6468 57092
rect 12786 57036 12796 57092
rect 12852 57036 13916 57092
rect 13972 57036 16492 57092
rect 16548 57036 16558 57092
rect 18060 57036 18676 57092
rect 26338 57036 26348 57092
rect 26404 57036 26796 57092
rect 26852 57036 26862 57092
rect 27010 57036 27020 57092
rect 27076 57036 27916 57092
rect 27972 57036 27982 57092
rect 6412 56980 6468 57036
rect 5366 56924 5404 56980
rect 5460 56924 5470 56980
rect 6402 56924 6412 56980
rect 6468 56924 6478 56980
rect 10770 56924 10780 56980
rect 10836 56924 12012 56980
rect 12068 56924 12078 56980
rect 12450 56924 12460 56980
rect 12516 56924 13580 56980
rect 13636 56924 13646 56980
rect 13794 56924 13804 56980
rect 13860 56924 14588 56980
rect 14644 56924 16604 56980
rect 16660 56924 16670 56980
rect 23986 56924 23996 56980
rect 24052 56924 24556 56980
rect 24612 56924 24622 56980
rect 25526 56924 25564 56980
rect 25620 56924 25630 56980
rect 26674 56924 26684 56980
rect 26740 56924 27692 56980
rect 27748 56924 28140 56980
rect 28196 56924 28206 56980
rect 4610 56812 4620 56868
rect 4676 56812 6860 56868
rect 6916 56812 6926 56868
rect 15362 56812 15372 56868
rect 15428 56812 15932 56868
rect 15988 56812 15998 56868
rect 17014 56812 17052 56868
rect 17108 56812 17118 56868
rect 21970 56812 21980 56868
rect 22036 56812 22316 56868
rect 22372 56812 22382 56868
rect 3574 56700 3612 56756
rect 3668 56700 4060 56756
rect 4116 56700 4396 56756
rect 4452 56700 4462 56756
rect 5254 56700 5292 56756
rect 5348 56700 5358 56756
rect 5506 56700 5516 56756
rect 5572 56700 5610 56756
rect 5814 56700 5852 56756
rect 5908 56700 5918 56756
rect 7522 56700 7532 56756
rect 7588 56700 8428 56756
rect 8484 56700 8494 56756
rect 15026 56700 15036 56756
rect 15092 56700 16492 56756
rect 16548 56700 16558 56756
rect 19478 56700 19516 56756
rect 19572 56700 21420 56756
rect 21476 56700 21486 56756
rect 25890 56700 25900 56756
rect 25956 56700 26908 56756
rect 26964 56700 26974 56756
rect 3490 56588 3500 56644
rect 3556 56588 5628 56644
rect 5684 56588 5694 56644
rect 9650 56588 9660 56644
rect 9716 56588 10220 56644
rect 10276 56588 10286 56644
rect 11890 56588 11900 56644
rect 11956 56588 19068 56644
rect 19124 56588 19134 56644
rect 24322 56588 24332 56644
rect 24388 56588 26012 56644
rect 26068 56588 27468 56644
rect 27524 56588 27534 56644
rect 4246 56476 4284 56532
rect 4340 56476 4350 56532
rect 5170 56476 5180 56532
rect 5236 56476 6188 56532
rect 6244 56476 6636 56532
rect 6692 56476 6702 56532
rect 9762 56476 9772 56532
rect 9828 56476 10108 56532
rect 10164 56476 10174 56532
rect 12226 56476 12236 56532
rect 12292 56476 12908 56532
rect 12964 56476 13692 56532
rect 13748 56476 13758 56532
rect 5180 56420 5236 56476
rect 8006 56420 8016 56476
rect 8072 56420 8120 56476
rect 8176 56420 8224 56476
rect 8280 56420 8290 56476
rect 14810 56420 14820 56476
rect 14876 56420 14924 56476
rect 14980 56420 15028 56476
rect 15084 56420 15094 56476
rect 21614 56420 21624 56476
rect 21680 56420 21728 56476
rect 21784 56420 21832 56476
rect 21888 56420 21898 56476
rect 28418 56420 28428 56476
rect 28484 56420 28532 56476
rect 28588 56420 28636 56476
rect 28692 56420 28702 56476
rect 3378 56364 3388 56420
rect 3444 56364 5236 56420
rect 8642 56364 8652 56420
rect 8708 56364 13916 56420
rect 13972 56364 13982 56420
rect 16146 56364 16156 56420
rect 16212 56364 16940 56420
rect 16996 56364 17006 56420
rect 17378 56364 17388 56420
rect 17444 56364 19068 56420
rect 19124 56364 19134 56420
rect 8978 56252 8988 56308
rect 9044 56252 10892 56308
rect 10948 56252 11116 56308
rect 11172 56252 11182 56308
rect 16594 56252 16604 56308
rect 16660 56252 20636 56308
rect 20692 56252 20702 56308
rect 21522 56252 21532 56308
rect 21588 56252 22204 56308
rect 22260 56252 22270 56308
rect 22502 56252 22540 56308
rect 22596 56252 22606 56308
rect 3602 56140 3612 56196
rect 3668 56140 3836 56196
rect 3892 56140 6748 56196
rect 6804 56140 6814 56196
rect 8866 56140 8876 56196
rect 8932 56140 9548 56196
rect 9604 56140 9614 56196
rect 10294 56140 10332 56196
rect 10388 56140 10398 56196
rect 11218 56140 11228 56196
rect 11284 56140 11452 56196
rect 11508 56140 13244 56196
rect 13300 56140 13310 56196
rect 15026 56140 15036 56196
rect 15092 56140 18004 56196
rect 19058 56140 19068 56196
rect 19124 56140 21196 56196
rect 21252 56140 22652 56196
rect 22708 56140 22718 56196
rect 25666 56140 25676 56196
rect 25732 56140 26124 56196
rect 26180 56140 26190 56196
rect 17948 56084 18004 56140
rect 4162 56028 4172 56084
rect 4228 56028 4956 56084
rect 5012 56028 12572 56084
rect 12628 56028 12638 56084
rect 12898 56028 12908 56084
rect 12964 56028 13692 56084
rect 13748 56028 13758 56084
rect 15474 56028 15484 56084
rect 15540 56028 15550 56084
rect 17938 56028 17948 56084
rect 18004 56028 18014 56084
rect 18274 56028 18284 56084
rect 18340 56028 18956 56084
rect 19012 56028 19022 56084
rect 19282 56028 19292 56084
rect 19348 56028 23436 56084
rect 23492 56028 23502 56084
rect 25778 56028 25788 56084
rect 25844 56028 26348 56084
rect 26404 56028 26414 56084
rect 15484 55972 15540 56028
rect 6626 55916 6636 55972
rect 6692 55916 7420 55972
rect 7476 55916 9772 55972
rect 9828 55916 9838 55972
rect 10322 55916 10332 55972
rect 10388 55916 15540 55972
rect 16930 55916 16940 55972
rect 16996 55916 17612 55972
rect 17668 55916 17678 55972
rect 17938 55916 17948 55972
rect 18004 55916 18172 55972
rect 18228 55916 18238 55972
rect 19618 55916 19628 55972
rect 19684 55916 19694 55972
rect 20178 55916 20188 55972
rect 20244 55916 21420 55972
rect 21476 55916 21486 55972
rect 25666 55916 25676 55972
rect 25732 55916 26012 55972
rect 26068 55916 26078 55972
rect 0 55860 400 55888
rect 19628 55860 19684 55916
rect 0 55804 1708 55860
rect 1764 55804 2492 55860
rect 2548 55804 2558 55860
rect 4274 55804 4284 55860
rect 4340 55804 5516 55860
rect 5572 55804 5582 55860
rect 8082 55804 8092 55860
rect 8148 55804 10108 55860
rect 10164 55804 10174 55860
rect 10434 55804 10444 55860
rect 10500 55804 10892 55860
rect 10948 55804 10958 55860
rect 11116 55804 11452 55860
rect 11508 55804 11518 55860
rect 13906 55804 13916 55860
rect 13972 55804 19684 55860
rect 0 55776 400 55804
rect 4604 55636 4614 55692
rect 4670 55636 4718 55692
rect 4774 55636 4822 55692
rect 4878 55636 4888 55692
rect 3826 55580 3836 55636
rect 3892 55580 4172 55636
rect 4228 55580 4238 55636
rect 11116 55412 11172 55804
rect 11778 55692 11788 55748
rect 11844 55692 12908 55748
rect 12964 55692 14140 55748
rect 14196 55692 14206 55748
rect 19506 55692 19516 55748
rect 19572 55692 20188 55748
rect 20244 55692 21868 55748
rect 21924 55692 24220 55748
rect 24276 55692 24286 55748
rect 11408 55636 11418 55692
rect 11474 55636 11522 55692
rect 11578 55636 11626 55692
rect 11682 55636 11692 55692
rect 18212 55636 18222 55692
rect 18278 55636 18326 55692
rect 18382 55636 18430 55692
rect 18486 55636 18496 55692
rect 25016 55636 25026 55692
rect 25082 55636 25130 55692
rect 25186 55636 25234 55692
rect 25290 55636 25300 55692
rect 22082 55580 22092 55636
rect 22148 55580 22158 55636
rect 11330 55468 11340 55524
rect 11396 55468 12796 55524
rect 12852 55468 12862 55524
rect 15474 55468 15484 55524
rect 15540 55468 16604 55524
rect 16660 55468 16670 55524
rect 17378 55468 17388 55524
rect 17444 55468 19964 55524
rect 20020 55468 20030 55524
rect 21270 55468 21308 55524
rect 21364 55468 21374 55524
rect 22092 55412 22148 55580
rect 22306 55468 22316 55524
rect 22372 55468 23044 55524
rect 22988 55412 23044 55468
rect 7746 55356 7756 55412
rect 7812 55356 7980 55412
rect 8036 55356 8652 55412
rect 8708 55356 8718 55412
rect 9426 55356 9436 55412
rect 9492 55356 11172 55412
rect 12562 55356 12572 55412
rect 12628 55356 13468 55412
rect 13524 55356 13534 55412
rect 20738 55356 20748 55412
rect 20804 55356 22764 55412
rect 22820 55356 22830 55412
rect 22988 55356 23212 55412
rect 23268 55356 23278 55412
rect 26002 55356 26012 55412
rect 26068 55356 26460 55412
rect 26516 55356 26526 55412
rect 27010 55356 27020 55412
rect 27076 55356 28028 55412
rect 28084 55356 28094 55412
rect 13570 55244 13580 55300
rect 13636 55244 14476 55300
rect 14532 55244 14542 55300
rect 15922 55244 15932 55300
rect 15988 55244 17612 55300
rect 17668 55244 17678 55300
rect 20962 55244 20972 55300
rect 21028 55244 25340 55300
rect 25396 55244 25564 55300
rect 25620 55244 25630 55300
rect 26786 55244 26796 55300
rect 26852 55244 27356 55300
rect 27412 55244 28140 55300
rect 28196 55244 28206 55300
rect 17612 55188 17668 55244
rect 9650 55132 9660 55188
rect 9716 55132 11564 55188
rect 11620 55132 11630 55188
rect 12002 55132 12012 55188
rect 12068 55132 12460 55188
rect 12516 55132 14028 55188
rect 14084 55132 15372 55188
rect 15428 55132 15438 55188
rect 17126 55132 17164 55188
rect 17220 55132 17230 55188
rect 17612 55132 21644 55188
rect 21700 55132 21710 55188
rect 22866 55132 22876 55188
rect 22932 55132 24108 55188
rect 24164 55132 24174 55188
rect 24546 55132 24556 55188
rect 24612 55132 25116 55188
rect 25172 55132 25182 55188
rect 25778 55132 25788 55188
rect 25844 55132 27244 55188
rect 27300 55132 27310 55188
rect 10630 55020 10668 55076
rect 10724 55020 14364 55076
rect 14420 55020 14430 55076
rect 20850 55020 20860 55076
rect 20916 55020 22036 55076
rect 22194 55020 22204 55076
rect 22260 55020 26012 55076
rect 26068 55020 26078 55076
rect 26562 55020 26572 55076
rect 26628 55020 27188 55076
rect 21980 54964 22036 55020
rect 9986 54908 9996 54964
rect 10052 54908 12012 54964
rect 12068 54908 12078 54964
rect 21980 54908 24668 54964
rect 24724 54908 24734 54964
rect 8006 54852 8016 54908
rect 8072 54852 8120 54908
rect 8176 54852 8224 54908
rect 8280 54852 8290 54908
rect 14810 54852 14820 54908
rect 14876 54852 14924 54908
rect 14980 54852 15028 54908
rect 15084 54852 15094 54908
rect 21614 54852 21624 54908
rect 21680 54852 21728 54908
rect 21784 54852 21832 54908
rect 21888 54852 21898 54908
rect 22652 54852 22708 54908
rect 27132 54852 27188 55020
rect 28418 54852 28428 54908
rect 28484 54852 28532 54908
rect 28588 54852 28636 54908
rect 28692 54852 28702 54908
rect 9202 54796 9212 54852
rect 9268 54796 10556 54852
rect 10612 54796 10622 54852
rect 19170 54796 19180 54852
rect 19236 54796 19628 54852
rect 19684 54796 19694 54852
rect 22642 54796 22652 54852
rect 22708 54796 22718 54852
rect 23090 54796 23100 54852
rect 23156 54796 23212 54852
rect 23268 54796 23278 54852
rect 23874 54796 23884 54852
rect 23940 54796 24108 54852
rect 24164 54796 25788 54852
rect 25844 54796 26908 54852
rect 27122 54796 27132 54852
rect 27188 54796 27198 54852
rect 3714 54684 3724 54740
rect 3780 54684 5292 54740
rect 5348 54684 5358 54740
rect 19730 54684 19740 54740
rect 19796 54684 23436 54740
rect 23492 54684 24108 54740
rect 24164 54684 24174 54740
rect 25330 54684 25340 54740
rect 25396 54684 25788 54740
rect 25844 54684 26348 54740
rect 26404 54684 26414 54740
rect 2594 54572 2604 54628
rect 2660 54572 2828 54628
rect 2884 54572 3500 54628
rect 3556 54572 3566 54628
rect 4386 54572 4396 54628
rect 4452 54572 5404 54628
rect 5460 54572 6076 54628
rect 6132 54572 12796 54628
rect 12852 54572 12862 54628
rect 20514 54572 20524 54628
rect 20580 54572 21084 54628
rect 21140 54572 21150 54628
rect 21634 54572 21644 54628
rect 21700 54572 23772 54628
rect 23828 54572 25676 54628
rect 25732 54572 26236 54628
rect 26292 54572 26302 54628
rect 26852 54516 26908 54796
rect 2146 54460 2156 54516
rect 2212 54460 3276 54516
rect 3332 54460 8540 54516
rect 8596 54460 8606 54516
rect 17714 54460 17724 54516
rect 17780 54460 21196 54516
rect 21252 54460 23660 54516
rect 23716 54460 23726 54516
rect 26852 54460 27692 54516
rect 27748 54460 27758 54516
rect 6178 54348 6188 54404
rect 6244 54348 6412 54404
rect 6468 54348 6478 54404
rect 13122 54348 13132 54404
rect 13188 54348 14140 54404
rect 14196 54348 20860 54404
rect 20916 54348 20926 54404
rect 21074 54348 21084 54404
rect 21140 54348 22428 54404
rect 22484 54348 22494 54404
rect 25330 54348 25340 54404
rect 25396 54348 26012 54404
rect 26068 54348 26684 54404
rect 26740 54348 26750 54404
rect 3266 54236 3276 54292
rect 3332 54236 3948 54292
rect 4004 54236 4014 54292
rect 8530 54236 8540 54292
rect 8596 54236 10444 54292
rect 10500 54236 12908 54292
rect 12964 54236 13580 54292
rect 13636 54236 13646 54292
rect 19954 54236 19964 54292
rect 20020 54236 20524 54292
rect 20580 54236 20590 54292
rect 20738 54236 20748 54292
rect 20804 54236 21196 54292
rect 21252 54236 21262 54292
rect 8194 54124 8204 54180
rect 8260 54124 10332 54180
rect 10388 54124 10556 54180
rect 10612 54124 10622 54180
rect 20066 54124 20076 54180
rect 20132 54124 21980 54180
rect 22036 54124 22046 54180
rect 23090 54124 23100 54180
rect 23156 54124 23436 54180
rect 23492 54124 23502 54180
rect 4604 54068 4614 54124
rect 4670 54068 4718 54124
rect 4774 54068 4822 54124
rect 4878 54068 4888 54124
rect 11408 54068 11418 54124
rect 11474 54068 11522 54124
rect 11578 54068 11626 54124
rect 11682 54068 11692 54124
rect 18212 54068 18222 54124
rect 18278 54068 18326 54124
rect 18382 54068 18430 54124
rect 18486 54068 18496 54124
rect 25016 54068 25026 54124
rect 25082 54068 25130 54124
rect 25186 54068 25234 54124
rect 25290 54068 25300 54124
rect 6402 54012 6412 54068
rect 6468 54012 9100 54068
rect 9156 54012 9166 54068
rect 11890 54012 11900 54068
rect 11956 54012 12348 54068
rect 12404 54012 12414 54068
rect 20290 54012 20300 54068
rect 20356 54012 23772 54068
rect 23828 54012 23838 54068
rect 4050 53900 4060 53956
rect 4116 53900 4508 53956
rect 4564 53900 4574 53956
rect 4722 53900 4732 53956
rect 4788 53900 18340 53956
rect 20850 53900 20860 53956
rect 20916 53900 26460 53956
rect 26516 53900 26526 53956
rect 18284 53844 18340 53900
rect 4610 53788 4620 53844
rect 4676 53788 5292 53844
rect 5348 53788 5358 53844
rect 5842 53788 5852 53844
rect 5908 53788 6300 53844
rect 6356 53788 6366 53844
rect 6598 53788 6636 53844
rect 6692 53788 6702 53844
rect 7298 53788 7308 53844
rect 7364 53788 8540 53844
rect 8596 53788 8606 53844
rect 9650 53788 9660 53844
rect 9716 53788 10220 53844
rect 10276 53788 10286 53844
rect 11106 53788 11116 53844
rect 11172 53788 11788 53844
rect 11844 53788 11854 53844
rect 12870 53788 12908 53844
rect 12964 53788 12974 53844
rect 18284 53788 20692 53844
rect 23314 53788 23324 53844
rect 23380 53788 24108 53844
rect 24164 53788 24174 53844
rect 26124 53788 28028 53844
rect 28084 53788 28094 53844
rect 20636 53732 20692 53788
rect 1810 53676 1820 53732
rect 1876 53676 3836 53732
rect 3892 53676 5628 53732
rect 5684 53676 5694 53732
rect 8978 53676 8988 53732
rect 9044 53676 10444 53732
rect 10500 53676 10510 53732
rect 11218 53676 11228 53732
rect 11284 53676 13132 53732
rect 13188 53676 13198 53732
rect 13356 53676 14924 53732
rect 14980 53676 14990 53732
rect 16258 53676 16268 53732
rect 16324 53676 16716 53732
rect 16772 53676 16782 53732
rect 18386 53676 18396 53732
rect 18452 53676 19068 53732
rect 19124 53676 19134 53732
rect 20262 53676 20300 53732
rect 20356 53676 20366 53732
rect 20626 53676 20636 53732
rect 20692 53676 20702 53732
rect 21196 53676 23212 53732
rect 23268 53676 23278 53732
rect 13356 53620 13412 53676
rect 21196 53620 21252 53676
rect 26124 53620 26180 53788
rect 26338 53676 26348 53732
rect 26404 53676 26796 53732
rect 26852 53676 26862 53732
rect 1698 53564 1708 53620
rect 1764 53564 1932 53620
rect 1988 53564 1998 53620
rect 4134 53564 4172 53620
rect 4228 53564 4956 53620
rect 5012 53564 5022 53620
rect 6262 53564 6300 53620
rect 6356 53564 6366 53620
rect 6738 53564 6748 53620
rect 6804 53564 8428 53620
rect 8484 53564 8764 53620
rect 8820 53564 8830 53620
rect 9986 53564 9996 53620
rect 10052 53564 12348 53620
rect 12404 53564 12414 53620
rect 12572 53564 13412 53620
rect 15026 53564 15036 53620
rect 15092 53564 15372 53620
rect 15428 53564 15438 53620
rect 18498 53564 18508 53620
rect 18564 53564 19236 53620
rect 19842 53564 19852 53620
rect 19908 53564 20076 53620
rect 20132 53564 21252 53620
rect 21308 53564 21644 53620
rect 21700 53564 21710 53620
rect 22194 53564 22204 53620
rect 22260 53564 23996 53620
rect 24052 53564 24062 53620
rect 26086 53564 26124 53620
rect 26180 53564 26190 53620
rect 26674 53564 26684 53620
rect 26740 53564 26750 53620
rect 27234 53564 27244 53620
rect 27300 53564 27692 53620
rect 27748 53564 27758 53620
rect 12572 53508 12628 53564
rect 19180 53508 19236 53564
rect 21308 53508 21364 53564
rect 26684 53508 26740 53564
rect 2930 53452 2940 53508
rect 2996 53452 7644 53508
rect 7700 53452 10780 53508
rect 10836 53452 10846 53508
rect 10994 53452 11004 53508
rect 11060 53452 11788 53508
rect 11844 53452 11854 53508
rect 12002 53452 12012 53508
rect 12068 53452 12628 53508
rect 12908 53452 14364 53508
rect 14420 53452 14700 53508
rect 14756 53452 14766 53508
rect 14914 53452 14924 53508
rect 14980 53452 16100 53508
rect 16258 53452 16268 53508
rect 16324 53452 16380 53508
rect 16436 53452 18956 53508
rect 19012 53452 19022 53508
rect 19170 53452 19180 53508
rect 19236 53452 19404 53508
rect 19460 53452 19470 53508
rect 20290 53452 20300 53508
rect 20356 53452 21364 53508
rect 21420 53452 21980 53508
rect 22036 53452 22046 53508
rect 22978 53452 22988 53508
rect 23044 53452 23884 53508
rect 23940 53452 23950 53508
rect 24210 53452 24220 53508
rect 24276 53452 27020 53508
rect 27076 53452 27580 53508
rect 27636 53452 28140 53508
rect 28196 53452 28206 53508
rect 8642 53340 8652 53396
rect 8708 53340 12012 53396
rect 12068 53340 12124 53396
rect 12180 53340 12684 53396
rect 12740 53340 12750 53396
rect 8006 53284 8016 53340
rect 8072 53284 8120 53340
rect 8176 53284 8224 53340
rect 8280 53284 8290 53340
rect 12908 53284 12964 53452
rect 16044 53396 16100 53452
rect 21420 53396 21476 53452
rect 16044 53340 21476 53396
rect 21980 53396 22036 53452
rect 21980 53340 24556 53396
rect 24612 53340 24622 53396
rect 26646 53340 26684 53396
rect 26740 53340 26750 53396
rect 14810 53284 14820 53340
rect 14876 53284 14924 53340
rect 14980 53284 15028 53340
rect 15084 53284 15094 53340
rect 21614 53284 21624 53340
rect 21680 53284 21728 53340
rect 21784 53284 21832 53340
rect 21888 53284 21898 53340
rect 24556 53284 24612 53340
rect 28418 53284 28428 53340
rect 28484 53284 28532 53340
rect 28588 53284 28636 53340
rect 28692 53284 28702 53340
rect 3826 53228 3836 53284
rect 3892 53228 5180 53284
rect 5236 53228 6300 53284
rect 6356 53228 6366 53284
rect 9090 53228 9100 53284
rect 9156 53228 11788 53284
rect 11844 53228 12572 53284
rect 12628 53228 12964 53284
rect 15586 53228 15596 53284
rect 15652 53228 18396 53284
rect 18452 53228 18462 53284
rect 22502 53228 22540 53284
rect 22596 53228 22606 53284
rect 24556 53228 26572 53284
rect 26628 53228 27132 53284
rect 27188 53228 27198 53284
rect 0 53172 400 53200
rect 0 53116 1932 53172
rect 1988 53116 1998 53172
rect 2818 53116 2828 53172
rect 2884 53116 8876 53172
rect 8932 53116 8942 53172
rect 9510 53116 9548 53172
rect 9604 53116 9614 53172
rect 9772 53116 20300 53172
rect 20356 53116 20366 53172
rect 21298 53116 21308 53172
rect 21364 53116 22652 53172
rect 22708 53116 22718 53172
rect 23090 53116 23100 53172
rect 23156 53116 25116 53172
rect 25172 53116 25788 53172
rect 25844 53116 25854 53172
rect 0 53088 400 53116
rect 4386 53004 4396 53060
rect 4452 53004 5068 53060
rect 5124 53004 5134 53060
rect 5702 53004 5740 53060
rect 5796 53004 9212 53060
rect 9268 53004 9278 53060
rect 4396 52948 4452 53004
rect 9772 52948 9828 53116
rect 23100 53060 23156 53116
rect 10098 53004 10108 53060
rect 10164 53004 10220 53060
rect 10276 53004 10286 53060
rect 11078 53004 11116 53060
rect 11172 53004 12124 53060
rect 12180 53004 12190 53060
rect 15026 53004 15036 53060
rect 15092 53004 15260 53060
rect 15316 53004 15708 53060
rect 15764 53004 15774 53060
rect 15922 53004 15932 53060
rect 15988 53004 16492 53060
rect 16548 53004 17948 53060
rect 18004 53004 18014 53060
rect 20514 53004 20524 53060
rect 20580 53004 20860 53060
rect 20916 53004 20926 53060
rect 21634 53004 21644 53060
rect 21700 53004 22428 53060
rect 22484 53004 23156 53060
rect 3332 52892 4452 52948
rect 4610 52892 4620 52948
rect 4676 52892 9828 52948
rect 10322 52892 10332 52948
rect 10388 52892 10556 52948
rect 10612 52892 10622 52948
rect 13654 52892 13692 52948
rect 13748 52892 15372 52948
rect 15428 52892 16268 52948
rect 16324 52892 16334 52948
rect 16818 52892 16828 52948
rect 16884 52892 17388 52948
rect 17444 52892 17454 52948
rect 18582 52892 18620 52948
rect 18676 52892 18686 52948
rect 20178 52892 20188 52948
rect 20244 52892 20636 52948
rect 20692 52892 23660 52948
rect 23716 52892 23726 52948
rect 24546 52892 24556 52948
rect 24612 52892 24892 52948
rect 24948 52892 25228 52948
rect 25284 52892 25294 52948
rect 3332 52836 3388 52892
rect 2146 52780 2156 52836
rect 2212 52780 3388 52836
rect 5740 52780 19740 52836
rect 19796 52780 19806 52836
rect 20402 52780 20412 52836
rect 20468 52780 21308 52836
rect 21364 52780 21374 52836
rect 26786 52780 26796 52836
rect 26852 52780 28140 52836
rect 28196 52780 28206 52836
rect 5740 52724 5796 52780
rect 2678 52668 2716 52724
rect 2772 52668 2782 52724
rect 4722 52668 4732 52724
rect 4788 52668 5012 52724
rect 5730 52668 5740 52724
rect 5796 52668 5806 52724
rect 9202 52668 9212 52724
rect 9268 52668 10668 52724
rect 10724 52668 10734 52724
rect 10882 52668 10892 52724
rect 10948 52668 13692 52724
rect 13748 52668 16716 52724
rect 16772 52668 16782 52724
rect 17042 52668 17052 52724
rect 17108 52668 17612 52724
rect 17668 52668 17678 52724
rect 18610 52668 18620 52724
rect 18676 52668 27468 52724
rect 27524 52668 27534 52724
rect 4604 52500 4614 52556
rect 4670 52500 4718 52556
rect 4774 52500 4822 52556
rect 4878 52500 4888 52556
rect 4956 52388 5012 52668
rect 7634 52556 7644 52612
rect 7700 52556 11228 52612
rect 11284 52556 11294 52612
rect 12338 52556 12348 52612
rect 12404 52556 12796 52612
rect 12852 52556 13580 52612
rect 13636 52556 13646 52612
rect 14802 52556 14812 52612
rect 14868 52556 17052 52612
rect 17108 52556 17948 52612
rect 18004 52556 18014 52612
rect 22642 52556 22652 52612
rect 22708 52556 24780 52612
rect 24836 52556 24846 52612
rect 11408 52500 11418 52556
rect 11474 52500 11522 52556
rect 11578 52500 11626 52556
rect 11682 52500 11692 52556
rect 18212 52500 18222 52556
rect 18278 52500 18326 52556
rect 18382 52500 18430 52556
rect 18486 52500 18496 52556
rect 25016 52500 25026 52556
rect 25082 52500 25130 52556
rect 25186 52500 25234 52556
rect 25290 52500 25300 52556
rect 5730 52444 5740 52500
rect 5796 52444 5806 52500
rect 6738 52444 6748 52500
rect 6804 52444 8092 52500
rect 8148 52444 11060 52500
rect 12562 52444 12572 52500
rect 12628 52444 17724 52500
rect 17780 52444 17790 52500
rect 5740 52388 5796 52444
rect 11004 52388 11060 52444
rect 12572 52388 12628 52444
rect 3714 52332 3724 52388
rect 3780 52332 4564 52388
rect 4722 52332 4732 52388
rect 4788 52332 5796 52388
rect 7410 52332 7420 52388
rect 7476 52332 7532 52388
rect 7588 52332 10108 52388
rect 10164 52332 10174 52388
rect 10994 52332 11004 52388
rect 11060 52332 12628 52388
rect 13318 52332 13356 52388
rect 13412 52332 13422 52388
rect 18834 52332 18844 52388
rect 18900 52332 20076 52388
rect 20132 52332 24332 52388
rect 24388 52332 24398 52388
rect 2790 52220 2828 52276
rect 2884 52220 2894 52276
rect 3378 52220 3388 52276
rect 3444 52220 4284 52276
rect 4340 52220 4350 52276
rect 4508 52164 4564 52332
rect 5842 52220 5852 52276
rect 5908 52220 7084 52276
rect 7140 52220 8428 52276
rect 8484 52220 8494 52276
rect 9874 52220 9884 52276
rect 9940 52220 10332 52276
rect 10388 52220 10556 52276
rect 10612 52220 10622 52276
rect 14102 52220 14140 52276
rect 14196 52220 17500 52276
rect 17556 52220 17612 52276
rect 17668 52220 17678 52276
rect 19954 52220 19964 52276
rect 20020 52220 26236 52276
rect 26292 52220 26302 52276
rect 3490 52108 3500 52164
rect 3556 52108 3724 52164
rect 3780 52108 3790 52164
rect 4508 52108 11004 52164
rect 11060 52108 11070 52164
rect 12114 52108 12124 52164
rect 12180 52108 12908 52164
rect 12964 52108 15148 52164
rect 15204 52108 15214 52164
rect 20514 52108 20524 52164
rect 20580 52108 22428 52164
rect 22484 52108 22494 52164
rect 22652 52108 23996 52164
rect 24052 52108 25228 52164
rect 25284 52108 25294 52164
rect 25666 52108 25676 52164
rect 25732 52108 27132 52164
rect 27188 52108 27198 52164
rect 22652 52052 22708 52108
rect 26236 52052 26292 52108
rect 2258 51996 2268 52052
rect 2324 51996 4508 52052
rect 4564 51996 4574 52052
rect 5618 51996 5628 52052
rect 5684 51996 6188 52052
rect 6244 51996 7532 52052
rect 7588 51996 8428 52052
rect 8484 51996 10108 52052
rect 10164 51996 10174 52052
rect 15922 51996 15932 52052
rect 15988 51996 18172 52052
rect 18228 51996 18238 52052
rect 19170 51996 19180 52052
rect 19236 51996 19292 52052
rect 19348 51996 19358 52052
rect 20738 51996 20748 52052
rect 20804 51996 21644 52052
rect 21700 51996 21710 52052
rect 21858 51996 21868 52052
rect 21924 51996 22092 52052
rect 22148 51996 22708 52052
rect 26226 51996 26236 52052
rect 26292 51996 26302 52052
rect 26562 51996 26572 52052
rect 26628 51996 27580 52052
rect 27636 51996 27646 52052
rect 4386 51884 4396 51940
rect 4452 51884 18396 51940
rect 18452 51884 18462 51940
rect 18722 51884 18732 51940
rect 18788 51884 23436 51940
rect 23492 51884 23502 51940
rect 26002 51884 26012 51940
rect 26068 51884 26348 51940
rect 26404 51884 26414 51940
rect 8978 51772 8988 51828
rect 9044 51772 9436 51828
rect 9492 51772 9502 51828
rect 19058 51772 19068 51828
rect 19124 51772 19404 51828
rect 19460 51772 19470 51828
rect 8006 51716 8016 51772
rect 8072 51716 8120 51772
rect 8176 51716 8224 51772
rect 8280 51716 8290 51772
rect 14810 51716 14820 51772
rect 14876 51716 14924 51772
rect 14980 51716 15028 51772
rect 15084 51716 15094 51772
rect 21614 51716 21624 51772
rect 21680 51716 21728 51772
rect 21784 51716 21832 51772
rect 21888 51716 21898 51772
rect 28418 51716 28428 51772
rect 28484 51716 28532 51772
rect 28588 51716 28636 51772
rect 28692 51716 28702 51772
rect 8754 51660 8764 51716
rect 8820 51660 9548 51716
rect 9604 51660 9614 51716
rect 16258 51660 16268 51716
rect 16324 51660 16828 51716
rect 16884 51660 17500 51716
rect 17556 51660 19292 51716
rect 19348 51660 19358 51716
rect 21970 51660 21980 51716
rect 22036 51660 24220 51716
rect 24276 51660 24286 51716
rect 4722 51548 4732 51604
rect 4788 51548 5964 51604
rect 6020 51548 6030 51604
rect 7746 51548 7756 51604
rect 7812 51548 11116 51604
rect 11172 51548 11182 51604
rect 16706 51548 16716 51604
rect 16772 51548 19180 51604
rect 19236 51548 19740 51604
rect 19796 51548 19806 51604
rect 5170 51436 5180 51492
rect 5236 51436 8988 51492
rect 9044 51436 9054 51492
rect 10658 51436 10668 51492
rect 10724 51436 10780 51492
rect 10836 51436 10846 51492
rect 18694 51436 18732 51492
rect 18788 51436 18798 51492
rect 23874 51436 23884 51492
rect 23940 51436 24220 51492
rect 24276 51436 25788 51492
rect 25844 51436 25854 51492
rect 26226 51436 26236 51492
rect 26292 51436 26908 51492
rect 26964 51436 26974 51492
rect 3602 51324 3612 51380
rect 3668 51324 5852 51380
rect 5908 51324 6244 51380
rect 8754 51324 8764 51380
rect 8820 51324 9996 51380
rect 10052 51324 10062 51380
rect 13580 51324 15596 51380
rect 15652 51324 16156 51380
rect 16212 51324 19628 51380
rect 19684 51324 19694 51380
rect 22978 51324 22988 51380
rect 23044 51324 23548 51380
rect 23604 51324 24108 51380
rect 24164 51324 24174 51380
rect 26450 51324 26460 51380
rect 26516 51324 27804 51380
rect 27860 51324 27870 51380
rect 6188 51268 6244 51324
rect 5394 51212 5404 51268
rect 5460 51212 5964 51268
rect 6020 51212 6030 51268
rect 6178 51212 6188 51268
rect 6244 51212 6282 51268
rect 8194 51212 8204 51268
rect 8260 51212 9100 51268
rect 9156 51212 9166 51268
rect 13580 51156 13636 51324
rect 23174 51212 23212 51268
rect 23268 51212 23278 51268
rect 2034 51100 2044 51156
rect 2100 51100 2716 51156
rect 2772 51100 3052 51156
rect 3108 51100 3118 51156
rect 3798 51100 3836 51156
rect 3892 51100 3902 51156
rect 6402 51100 6412 51156
rect 6468 51100 7196 51156
rect 7252 51100 7262 51156
rect 10770 51100 10780 51156
rect 10836 51100 11676 51156
rect 11732 51100 11742 51156
rect 12002 51100 12012 51156
rect 12068 51100 13580 51156
rect 13636 51100 13646 51156
rect 18162 51100 18172 51156
rect 18228 51100 19964 51156
rect 20020 51100 20030 51156
rect 22194 51100 22204 51156
rect 22260 51100 24444 51156
rect 24500 51100 24510 51156
rect 24668 51100 25340 51156
rect 25396 51100 25406 51156
rect 5282 50988 5292 51044
rect 5348 50988 5628 51044
rect 5684 50988 5694 51044
rect 7858 50988 7868 51044
rect 7924 50988 8652 51044
rect 8708 50988 8718 51044
rect 13906 50988 13916 51044
rect 13972 50988 15372 51044
rect 15428 50988 15438 51044
rect 4604 50932 4614 50988
rect 4670 50932 4718 50988
rect 4774 50932 4822 50988
rect 4878 50932 4888 50988
rect 11408 50932 11418 50988
rect 11474 50932 11522 50988
rect 11578 50932 11626 50988
rect 11682 50932 11692 50988
rect 18212 50932 18222 50988
rect 18278 50932 18326 50988
rect 18382 50932 18430 50988
rect 18486 50932 18496 50988
rect 24668 50932 24724 51100
rect 26226 50988 26236 51044
rect 26292 50988 27020 51044
rect 27076 50988 27086 51044
rect 25016 50932 25026 50988
rect 25082 50932 25130 50988
rect 25186 50932 25234 50988
rect 25290 50932 25300 50988
rect 5394 50876 5404 50932
rect 5460 50876 5964 50932
rect 6020 50876 6030 50932
rect 12562 50876 12572 50932
rect 12628 50876 13244 50932
rect 13300 50876 13310 50932
rect 21298 50876 21308 50932
rect 21364 50876 23436 50932
rect 23492 50876 24724 50932
rect 4050 50764 4060 50820
rect 4116 50764 4620 50820
rect 4676 50764 7140 50820
rect 14802 50764 14812 50820
rect 14868 50764 15148 50820
rect 15204 50764 15932 50820
rect 15988 50764 16156 50820
rect 16212 50764 17948 50820
rect 18004 50764 18508 50820
rect 18564 50764 18574 50820
rect 19618 50764 19628 50820
rect 19684 50764 22652 50820
rect 22708 50764 22876 50820
rect 22932 50764 22942 50820
rect 7084 50708 7140 50764
rect 5170 50652 5180 50708
rect 5236 50652 6860 50708
rect 6916 50652 6926 50708
rect 7084 50652 10556 50708
rect 10612 50652 10622 50708
rect 13122 50652 13132 50708
rect 13188 50652 13468 50708
rect 13524 50652 13534 50708
rect 19058 50652 19068 50708
rect 19124 50652 19180 50708
rect 19236 50652 24332 50708
rect 24388 50652 24398 50708
rect 26852 50652 27244 50708
rect 27300 50652 27310 50708
rect 6178 50540 6188 50596
rect 6244 50540 7308 50596
rect 7364 50540 7420 50596
rect 7476 50540 7868 50596
rect 7924 50540 7934 50596
rect 13570 50540 13580 50596
rect 13636 50540 14252 50596
rect 14308 50540 14318 50596
rect 22278 50540 22316 50596
rect 22372 50540 22382 50596
rect 24434 50540 24444 50596
rect 24500 50540 25452 50596
rect 25508 50540 25518 50596
rect 25750 50540 25788 50596
rect 25844 50540 25854 50596
rect 0 50484 400 50512
rect 0 50428 1708 50484
rect 1764 50428 1774 50484
rect 2482 50428 2492 50484
rect 2548 50428 3164 50484
rect 3220 50428 3230 50484
rect 0 50400 400 50428
rect 6524 50260 6580 50540
rect 26852 50484 26908 50652
rect 6738 50428 6748 50484
rect 6804 50428 7532 50484
rect 7588 50428 12460 50484
rect 12516 50428 12526 50484
rect 13010 50428 13020 50484
rect 13076 50428 14476 50484
rect 14532 50428 14542 50484
rect 15026 50428 15036 50484
rect 15092 50428 16492 50484
rect 16548 50428 16558 50484
rect 17686 50428 17724 50484
rect 17780 50428 17790 50484
rect 20066 50428 20076 50484
rect 20132 50428 22428 50484
rect 22484 50428 24332 50484
rect 24388 50428 26908 50484
rect 16492 50372 16548 50428
rect 12226 50316 12236 50372
rect 12292 50316 13916 50372
rect 13972 50316 13982 50372
rect 16492 50316 17612 50372
rect 17668 50316 17678 50372
rect 19170 50316 19180 50372
rect 19236 50316 19292 50372
rect 19348 50316 20076 50372
rect 20132 50316 20142 50372
rect 6524 50204 6748 50260
rect 6804 50204 6814 50260
rect 8418 50204 8428 50260
rect 8484 50204 8522 50260
rect 8754 50204 8764 50260
rect 8820 50204 10332 50260
rect 10388 50204 13468 50260
rect 13524 50204 13534 50260
rect 8006 50148 8016 50204
rect 8072 50148 8120 50204
rect 8176 50148 8224 50204
rect 8280 50148 8290 50204
rect 14810 50148 14820 50204
rect 14876 50148 14924 50204
rect 14980 50148 15028 50204
rect 15084 50148 15094 50204
rect 21614 50148 21624 50204
rect 21680 50148 21728 50204
rect 21784 50148 21832 50204
rect 21888 50148 21898 50204
rect 28418 50148 28428 50204
rect 28484 50148 28532 50204
rect 28588 50148 28636 50204
rect 28692 50148 28702 50204
rect 2146 50092 2156 50148
rect 2212 50092 2940 50148
rect 2996 50092 3006 50148
rect 15250 50092 15260 50148
rect 15316 50092 15932 50148
rect 15988 50092 15998 50148
rect 3266 49980 3276 50036
rect 3332 49980 4284 50036
rect 4340 49980 4350 50036
rect 6290 49980 6300 50036
rect 6356 49980 6412 50036
rect 6468 49980 6478 50036
rect 10658 49980 10668 50036
rect 10724 49980 11452 50036
rect 11508 49980 11518 50036
rect 11890 49980 11900 50036
rect 11956 49980 15596 50036
rect 15652 49980 15662 50036
rect 17490 49980 17500 50036
rect 17556 49980 19516 50036
rect 19572 49980 19582 50036
rect 20962 49980 20972 50036
rect 21028 49980 24220 50036
rect 24276 49980 24286 50036
rect 2034 49868 2044 49924
rect 2100 49868 5628 49924
rect 5684 49868 5694 49924
rect 8194 49868 8204 49924
rect 8260 49868 12460 49924
rect 12516 49868 12526 49924
rect 14018 49868 14028 49924
rect 14084 49868 14364 49924
rect 14420 49868 16828 49924
rect 16884 49868 17388 49924
rect 17444 49868 17724 49924
rect 17780 49868 17790 49924
rect 18498 49868 18508 49924
rect 18564 49868 20524 49924
rect 20580 49868 20590 49924
rect 2566 49756 2604 49812
rect 2660 49756 2670 49812
rect 2818 49756 2828 49812
rect 2884 49756 3164 49812
rect 3220 49756 3230 49812
rect 6514 49756 6524 49812
rect 6580 49756 7084 49812
rect 7140 49756 8652 49812
rect 8708 49756 8718 49812
rect 10098 49756 10108 49812
rect 10164 49756 11228 49812
rect 11284 49756 11900 49812
rect 11956 49756 11966 49812
rect 17938 49756 17948 49812
rect 18004 49756 18956 49812
rect 19012 49756 19022 49812
rect 19506 49756 19516 49812
rect 19572 49756 21308 49812
rect 21364 49756 21374 49812
rect 1810 49644 1820 49700
rect 1876 49644 3388 49700
rect 10966 49644 11004 49700
rect 11060 49644 11070 49700
rect 18610 49644 18620 49700
rect 18676 49644 19068 49700
rect 19124 49644 19134 49700
rect 22530 49644 22540 49700
rect 22596 49644 23436 49700
rect 23492 49644 23502 49700
rect 25554 49644 25564 49700
rect 25620 49644 27468 49700
rect 27524 49644 27534 49700
rect 2492 49588 2548 49644
rect 3332 49588 3388 49644
rect 2482 49532 2492 49588
rect 2548 49532 2558 49588
rect 3332 49532 4620 49588
rect 4676 49532 6188 49588
rect 6244 49532 6254 49588
rect 9734 49532 9772 49588
rect 9828 49532 10780 49588
rect 10836 49532 15484 49588
rect 15540 49532 16380 49588
rect 16436 49532 16446 49588
rect 24098 49532 24108 49588
rect 24164 49532 27132 49588
rect 27188 49532 27198 49588
rect 13458 49420 13468 49476
rect 13524 49420 14140 49476
rect 14196 49420 14206 49476
rect 25554 49420 25564 49476
rect 25620 49420 26012 49476
rect 26068 49420 26078 49476
rect 4604 49364 4614 49420
rect 4670 49364 4718 49420
rect 4774 49364 4822 49420
rect 4878 49364 4888 49420
rect 11408 49364 11418 49420
rect 11474 49364 11522 49420
rect 11578 49364 11626 49420
rect 11682 49364 11692 49420
rect 18212 49364 18222 49420
rect 18278 49364 18326 49420
rect 18382 49364 18430 49420
rect 18486 49364 18496 49420
rect 25016 49364 25026 49420
rect 25082 49364 25130 49420
rect 25186 49364 25234 49420
rect 25290 49364 25300 49420
rect 1810 49308 1820 49364
rect 1876 49308 1886 49364
rect 10742 49308 10780 49364
rect 10836 49308 10846 49364
rect 25442 49308 25452 49364
rect 25508 49308 26572 49364
rect 26628 49308 26638 49364
rect 1820 48916 1876 49308
rect 4386 49196 4396 49252
rect 4452 49196 5068 49252
rect 5124 49196 5134 49252
rect 7858 49196 7868 49252
rect 7924 49196 8652 49252
rect 8708 49196 11340 49252
rect 11396 49196 14364 49252
rect 14420 49196 14430 49252
rect 22194 49196 22204 49252
rect 22260 49196 22988 49252
rect 23044 49196 23054 49252
rect 23874 49196 23884 49252
rect 23940 49196 25228 49252
rect 25284 49196 25294 49252
rect 5282 49084 5292 49140
rect 5348 49084 5628 49140
rect 5684 49084 5694 49140
rect 6850 49084 6860 49140
rect 6916 49084 8428 49140
rect 8484 49084 8494 49140
rect 11106 49084 11116 49140
rect 11172 49084 12236 49140
rect 12292 49084 12302 49140
rect 15362 49084 15372 49140
rect 15428 49084 16268 49140
rect 16324 49084 16334 49140
rect 20626 49084 20636 49140
rect 20692 49084 21420 49140
rect 21476 49084 21486 49140
rect 23996 49084 25900 49140
rect 25956 49084 25966 49140
rect 23996 49028 24052 49084
rect 3602 48972 3612 49028
rect 3668 48972 3836 49028
rect 3892 48972 3948 49028
rect 4004 48972 4014 49028
rect 4162 48972 4172 49028
rect 4228 48972 4396 49028
rect 4452 48972 4462 49028
rect 6962 48972 6972 49028
rect 7028 48972 7308 49028
rect 7364 48972 7374 49028
rect 11750 48972 11788 49028
rect 11844 48972 11854 49028
rect 12338 48972 12348 49028
rect 12404 48972 13916 49028
rect 13972 48972 13982 49028
rect 14130 48972 14140 49028
rect 14196 48972 15148 49028
rect 15204 48972 15214 49028
rect 18946 48972 18956 49028
rect 19012 48972 20076 49028
rect 20132 48972 20142 49028
rect 23650 48972 23660 49028
rect 23716 48972 23996 49028
rect 24052 48972 24062 49028
rect 24322 48972 24332 49028
rect 24388 48972 24500 49028
rect 24658 48972 24668 49028
rect 24724 48972 25228 49028
rect 25284 48972 25294 49028
rect 26310 48972 26348 49028
rect 26404 48972 26572 49028
rect 26628 48972 26638 49028
rect 24444 48916 24500 48972
rect 1810 48860 1820 48916
rect 1876 48860 1886 48916
rect 9090 48860 9100 48916
rect 9156 48860 11004 48916
rect 11060 48860 12572 48916
rect 12628 48860 12796 48916
rect 12852 48860 13804 48916
rect 13860 48860 13870 48916
rect 14438 48860 14476 48916
rect 14532 48860 14542 48916
rect 17042 48860 17052 48916
rect 17108 48860 17388 48916
rect 17444 48860 17454 48916
rect 19282 48860 19292 48916
rect 19348 48860 20188 48916
rect 20244 48860 21868 48916
rect 21924 48860 24220 48916
rect 24276 48860 24286 48916
rect 24444 48860 24892 48916
rect 24948 48860 24958 48916
rect 26674 48860 26684 48916
rect 26740 48860 26908 48916
rect 26964 48860 26974 48916
rect 3574 48748 3612 48804
rect 3668 48748 3678 48804
rect 4162 48748 4172 48804
rect 4228 48748 4620 48804
rect 4676 48748 4686 48804
rect 5730 48748 5740 48804
rect 5796 48748 6188 48804
rect 6244 48748 6412 48804
rect 6468 48748 6478 48804
rect 10546 48748 10556 48804
rect 10612 48748 12236 48804
rect 12292 48748 13020 48804
rect 13076 48748 14028 48804
rect 14084 48748 14644 48804
rect 17714 48748 17724 48804
rect 17780 48748 18956 48804
rect 19012 48748 19022 48804
rect 22194 48748 22204 48804
rect 22260 48748 24332 48804
rect 24388 48748 24398 48804
rect 9986 48636 9996 48692
rect 10052 48636 10444 48692
rect 10500 48636 11788 48692
rect 11844 48636 11854 48692
rect 14326 48636 14364 48692
rect 14420 48636 14430 48692
rect 8006 48580 8016 48636
rect 8072 48580 8120 48636
rect 8176 48580 8224 48636
rect 8280 48580 8290 48636
rect 3826 48524 3836 48580
rect 3892 48524 4284 48580
rect 4340 48524 4350 48580
rect 5842 48524 5852 48580
rect 5908 48524 6524 48580
rect 6580 48524 6590 48580
rect 14588 48468 14644 48748
rect 16706 48636 16716 48692
rect 16772 48636 19740 48692
rect 19796 48636 19806 48692
rect 22390 48636 22428 48692
rect 22484 48636 22494 48692
rect 24322 48636 24332 48692
rect 24388 48636 24892 48692
rect 24948 48636 24958 48692
rect 14810 48580 14820 48636
rect 14876 48580 14924 48636
rect 14980 48580 15028 48636
rect 15084 48580 15094 48636
rect 21614 48580 21624 48636
rect 21680 48580 21728 48636
rect 21784 48580 21832 48636
rect 21888 48580 21898 48636
rect 28418 48580 28428 48636
rect 28484 48580 28532 48636
rect 28588 48580 28636 48636
rect 28692 48580 28702 48636
rect 17462 48524 17500 48580
rect 17556 48524 17566 48580
rect 3714 48412 3724 48468
rect 3780 48412 4172 48468
rect 4228 48412 4238 48468
rect 7494 48412 7532 48468
rect 7588 48412 9436 48468
rect 9492 48412 9996 48468
rect 10052 48412 10062 48468
rect 10406 48412 10444 48468
rect 10500 48412 10510 48468
rect 11190 48412 11228 48468
rect 11284 48412 11294 48468
rect 12674 48412 12684 48468
rect 12740 48412 13132 48468
rect 13188 48412 13198 48468
rect 14588 48412 15036 48468
rect 15092 48412 15102 48468
rect 15922 48412 15932 48468
rect 15988 48412 22092 48468
rect 22148 48412 22158 48468
rect 2930 48300 2940 48356
rect 2996 48300 4956 48356
rect 5012 48300 5022 48356
rect 5842 48300 5852 48356
rect 5908 48300 6860 48356
rect 6916 48300 6926 48356
rect 8502 48300 8540 48356
rect 8596 48300 8606 48356
rect 14130 48300 14140 48356
rect 14196 48300 15204 48356
rect 15148 48244 15204 48300
rect 8306 48188 8316 48244
rect 8372 48188 10892 48244
rect 10948 48188 10958 48244
rect 15138 48188 15148 48244
rect 15204 48188 15214 48244
rect 15932 48132 15988 48412
rect 16258 48300 16268 48356
rect 16324 48300 17500 48356
rect 17556 48300 17948 48356
rect 18004 48300 18014 48356
rect 21298 48188 21308 48244
rect 21364 48188 21644 48244
rect 21700 48188 21710 48244
rect 2482 48076 2492 48132
rect 2548 48076 3052 48132
rect 3108 48076 3118 48132
rect 7410 48076 7420 48132
rect 7476 48076 8428 48132
rect 8484 48076 8494 48132
rect 9202 48076 9212 48132
rect 9268 48076 9660 48132
rect 9716 48076 9726 48132
rect 10742 48076 10780 48132
rect 10836 48076 10846 48132
rect 14130 48076 14140 48132
rect 14196 48076 15988 48132
rect 16044 48076 19292 48132
rect 19348 48076 19358 48132
rect 26086 48076 26124 48132
rect 26180 48076 26190 48132
rect 16044 48020 16100 48076
rect 4610 47964 4620 48020
rect 4676 47964 9996 48020
rect 10052 47964 10062 48020
rect 13794 47964 13804 48020
rect 13860 47964 14700 48020
rect 14756 47964 16100 48020
rect 16818 47964 16828 48020
rect 16884 47964 16894 48020
rect 17154 47964 17164 48020
rect 17220 47964 17612 48020
rect 17668 47964 17678 48020
rect 16828 47908 16884 47964
rect 4946 47852 4956 47908
rect 5012 47852 5022 47908
rect 7074 47852 7084 47908
rect 7140 47852 9212 47908
rect 9268 47852 9548 47908
rect 9604 47852 9614 47908
rect 10098 47852 10108 47908
rect 10164 47852 10612 47908
rect 16828 47852 17556 47908
rect 19730 47852 19740 47908
rect 19796 47852 20860 47908
rect 20916 47852 20926 47908
rect 0 47796 400 47824
rect 4604 47796 4614 47852
rect 4670 47796 4718 47852
rect 4774 47796 4822 47852
rect 4878 47796 4888 47852
rect 0 47740 1428 47796
rect 0 47712 400 47740
rect 1372 47460 1428 47740
rect 3154 47628 3164 47684
rect 3220 47628 3230 47684
rect 3490 47628 3500 47684
rect 3556 47628 4060 47684
rect 4116 47628 4126 47684
rect 3164 47572 3220 47628
rect 1698 47516 1708 47572
rect 1764 47516 2492 47572
rect 2548 47516 2558 47572
rect 3164 47516 3948 47572
rect 4004 47516 4732 47572
rect 4788 47516 4798 47572
rect 4956 47460 5012 47852
rect 10556 47796 10612 47852
rect 11408 47796 11418 47852
rect 11474 47796 11522 47852
rect 11578 47796 11626 47852
rect 11682 47796 11692 47852
rect 10210 47740 10220 47796
rect 10276 47740 10332 47796
rect 10388 47740 10398 47796
rect 10546 47740 10556 47796
rect 10612 47740 10622 47796
rect 16818 47740 16828 47796
rect 16884 47740 17276 47796
rect 17332 47740 17342 47796
rect 17500 47684 17556 47852
rect 18212 47796 18222 47852
rect 18278 47796 18326 47852
rect 18382 47796 18430 47852
rect 18486 47796 18496 47852
rect 25016 47796 25026 47852
rect 25082 47796 25130 47852
rect 25186 47796 25234 47852
rect 25290 47796 25300 47852
rect 20514 47740 20524 47796
rect 20580 47740 20590 47796
rect 20524 47684 20580 47740
rect 5478 47628 5516 47684
rect 5572 47628 5582 47684
rect 8194 47628 8204 47684
rect 8260 47628 9100 47684
rect 9156 47628 9772 47684
rect 9828 47628 10220 47684
rect 10276 47628 10286 47684
rect 10546 47628 10556 47684
rect 10612 47628 11452 47684
rect 11508 47628 11518 47684
rect 12422 47628 12460 47684
rect 12516 47628 15260 47684
rect 15316 47628 15326 47684
rect 17500 47628 18396 47684
rect 18452 47628 19180 47684
rect 19236 47628 20580 47684
rect 20850 47628 20860 47684
rect 20916 47628 21532 47684
rect 21588 47628 21598 47684
rect 10770 47516 10780 47572
rect 10836 47516 13916 47572
rect 13972 47516 20524 47572
rect 20580 47516 20590 47572
rect 21420 47516 22764 47572
rect 22820 47516 22830 47572
rect 23398 47516 23436 47572
rect 23492 47516 23502 47572
rect 21420 47460 21476 47516
rect 1372 47404 1764 47460
rect 2146 47404 2156 47460
rect 2212 47404 3164 47460
rect 3220 47404 3230 47460
rect 3826 47404 3836 47460
rect 3892 47404 4508 47460
rect 4564 47404 4574 47460
rect 4946 47404 4956 47460
rect 5012 47404 5022 47460
rect 9538 47404 9548 47460
rect 9604 47404 10388 47460
rect 11974 47404 12012 47460
rect 12068 47404 12078 47460
rect 12226 47404 12236 47460
rect 12292 47404 14140 47460
rect 14196 47404 17500 47460
rect 17556 47404 17566 47460
rect 18610 47404 18620 47460
rect 18676 47404 19516 47460
rect 19572 47404 19582 47460
rect 21410 47404 21420 47460
rect 21476 47404 21486 47460
rect 21970 47404 21980 47460
rect 22036 47404 23548 47460
rect 23604 47404 25564 47460
rect 25620 47404 25630 47460
rect 1708 47348 1764 47404
rect 10332 47348 10388 47404
rect 19516 47348 19572 47404
rect 1698 47292 1708 47348
rect 1764 47292 2604 47348
rect 2660 47292 2670 47348
rect 3490 47292 3500 47348
rect 3556 47292 4284 47348
rect 4340 47292 4350 47348
rect 6738 47292 6748 47348
rect 6804 47292 10108 47348
rect 10164 47292 10174 47348
rect 10332 47292 10444 47348
rect 10500 47292 10510 47348
rect 10770 47292 10780 47348
rect 10836 47292 10948 47348
rect 11330 47292 11340 47348
rect 11396 47292 14364 47348
rect 14420 47292 15932 47348
rect 15988 47292 15998 47348
rect 19516 47292 22316 47348
rect 22372 47292 23324 47348
rect 23380 47292 23390 47348
rect 10892 47236 10948 47292
rect 2034 47180 2044 47236
rect 2100 47180 5068 47236
rect 5124 47180 5740 47236
rect 5796 47180 5806 47236
rect 10434 47180 10444 47236
rect 10500 47180 10668 47236
rect 10724 47180 10734 47236
rect 10892 47180 12012 47236
rect 12068 47180 12078 47236
rect 12898 47180 12908 47236
rect 12964 47180 14364 47236
rect 14420 47180 14700 47236
rect 14756 47180 14766 47236
rect 17938 47180 17948 47236
rect 18004 47180 18042 47236
rect 19954 47180 19964 47236
rect 20020 47180 20188 47236
rect 20244 47180 20254 47236
rect 20514 47180 20524 47236
rect 20580 47180 25452 47236
rect 25508 47180 26348 47236
rect 26404 47180 26414 47236
rect 5842 47068 5852 47124
rect 5908 47068 7084 47124
rect 7140 47068 7150 47124
rect 10210 47068 10220 47124
rect 10276 47068 10332 47124
rect 10388 47068 10398 47124
rect 10546 47068 10556 47124
rect 10612 47068 11788 47124
rect 11844 47068 11854 47124
rect 14018 47068 14028 47124
rect 14084 47068 14364 47124
rect 14420 47068 14430 47124
rect 17154 47068 17164 47124
rect 17220 47068 17332 47124
rect 17490 47068 17500 47124
rect 17556 47068 17566 47124
rect 19730 47068 19740 47124
rect 19796 47068 20300 47124
rect 20356 47068 20366 47124
rect 20738 47068 20748 47124
rect 20804 47068 21476 47124
rect 23202 47068 23212 47124
rect 23268 47068 23278 47124
rect 25666 47068 25676 47124
rect 25732 47068 26012 47124
rect 26068 47068 26078 47124
rect 4834 47012 4844 47068
rect 4900 47012 4910 47068
rect 8006 47012 8016 47068
rect 8072 47012 8120 47068
rect 8176 47012 8224 47068
rect 8280 47012 8290 47068
rect 9958 47012 9996 47068
rect 10052 47012 10062 47068
rect 14810 47012 14820 47068
rect 14876 47012 14924 47068
rect 14980 47012 15028 47068
rect 15084 47012 15094 47068
rect 17266 47012 17276 47068
rect 17332 47012 17342 47068
rect 17500 47012 17556 47068
rect 4844 46956 5908 47012
rect 10882 46956 10892 47012
rect 10948 46956 11004 47012
rect 11060 46956 11070 47012
rect 17500 46956 17836 47012
rect 17892 46956 17902 47012
rect 5852 46900 5908 46956
rect 21420 46900 21476 47068
rect 21614 47012 21624 47068
rect 21680 47012 21728 47068
rect 21784 47012 21832 47068
rect 21888 47012 21898 47068
rect 23212 47012 23268 47068
rect 28418 47012 28428 47068
rect 28484 47012 28532 47068
rect 28588 47012 28636 47068
rect 28692 47012 28702 47068
rect 22092 46956 26684 47012
rect 26740 46956 26750 47012
rect 27234 46956 27244 47012
rect 27300 46956 27804 47012
rect 27860 46956 27870 47012
rect 1810 46844 1820 46900
rect 1876 46844 4060 46900
rect 4116 46844 5516 46900
rect 5572 46844 5582 46900
rect 5842 46844 5852 46900
rect 5908 46844 5918 46900
rect 20738 46844 20748 46900
rect 20804 46844 20860 46900
rect 20916 46844 20926 46900
rect 21420 46844 21644 46900
rect 21700 46844 21710 46900
rect 22092 46788 22148 46956
rect 22978 46844 22988 46900
rect 23044 46844 23100 46900
rect 23156 46844 23166 46900
rect 23986 46844 23996 46900
rect 24052 46844 24332 46900
rect 24388 46844 27132 46900
rect 27188 46844 27198 46900
rect 3602 46732 3612 46788
rect 3668 46732 4060 46788
rect 4116 46732 4126 46788
rect 5142 46732 5180 46788
rect 5236 46732 5246 46788
rect 10322 46732 10332 46788
rect 10388 46732 10892 46788
rect 10948 46732 10958 46788
rect 13206 46732 13244 46788
rect 13300 46732 13310 46788
rect 15026 46732 15036 46788
rect 15092 46732 20076 46788
rect 20132 46732 22092 46788
rect 22148 46732 22158 46788
rect 22978 46732 22988 46788
rect 23044 46732 24444 46788
rect 24500 46732 25732 46788
rect 25676 46676 25732 46732
rect 4162 46620 4172 46676
rect 4228 46620 5404 46676
rect 5460 46620 5470 46676
rect 15474 46620 15484 46676
rect 15540 46620 15932 46676
rect 15988 46620 15998 46676
rect 20290 46620 20300 46676
rect 20356 46620 20366 46676
rect 21410 46620 21420 46676
rect 21476 46620 23100 46676
rect 23156 46620 24220 46676
rect 24276 46620 24286 46676
rect 24546 46620 24556 46676
rect 24612 46620 25340 46676
rect 25396 46620 25406 46676
rect 25676 46620 25788 46676
rect 25844 46620 25854 46676
rect 3126 46508 3164 46564
rect 3220 46508 3230 46564
rect 4498 46508 4508 46564
rect 4564 46508 5852 46564
rect 5908 46508 5918 46564
rect 6290 46508 6300 46564
rect 6356 46508 6860 46564
rect 6916 46508 6926 46564
rect 8978 46508 8988 46564
rect 9044 46508 10108 46564
rect 10164 46508 10332 46564
rect 10388 46508 10398 46564
rect 11218 46508 11228 46564
rect 11284 46508 11452 46564
rect 11508 46508 11518 46564
rect 19170 46508 19180 46564
rect 19236 46508 19516 46564
rect 19572 46508 19582 46564
rect 20300 46452 20356 46620
rect 23314 46508 23324 46564
rect 23380 46508 23548 46564
rect 23604 46508 25228 46564
rect 25284 46508 25294 46564
rect 3602 46396 3612 46452
rect 3668 46396 4284 46452
rect 4340 46396 4844 46452
rect 4900 46396 4910 46452
rect 20300 46396 26572 46452
rect 26628 46396 26638 46452
rect 4604 46228 4614 46284
rect 4670 46228 4718 46284
rect 4774 46228 4822 46284
rect 4878 46228 4888 46284
rect 11408 46228 11418 46284
rect 11474 46228 11522 46284
rect 11578 46228 11626 46284
rect 11682 46228 11692 46284
rect 18212 46228 18222 46284
rect 18278 46228 18326 46284
rect 18382 46228 18430 46284
rect 18486 46228 18496 46284
rect 25016 46228 25026 46284
rect 25082 46228 25130 46284
rect 25186 46228 25234 46284
rect 25290 46228 25300 46284
rect 6402 46172 6412 46228
rect 6468 46172 7868 46228
rect 7924 46172 7934 46228
rect 22642 46172 22652 46228
rect 22708 46172 22764 46228
rect 22820 46172 22830 46228
rect 7046 46060 7084 46116
rect 7140 46060 7150 46116
rect 7298 46060 7308 46116
rect 7364 46060 7374 46116
rect 22754 46060 22764 46116
rect 22820 46060 22830 46116
rect 7308 45780 7364 46060
rect 12450 45948 12460 46004
rect 12516 45948 12796 46004
rect 12852 45948 12862 46004
rect 17014 45948 17052 46004
rect 17108 45948 17118 46004
rect 7970 45836 7980 45892
rect 8036 45836 8204 45892
rect 8260 45836 8270 45892
rect 9202 45836 9212 45892
rect 9268 45836 9436 45892
rect 9492 45836 11508 45892
rect 11890 45836 11900 45892
rect 11956 45836 13804 45892
rect 13860 45836 13870 45892
rect 14690 45836 14700 45892
rect 14756 45836 15260 45892
rect 15316 45836 15326 45892
rect 15810 45836 15820 45892
rect 15876 45836 17388 45892
rect 17444 45836 17454 45892
rect 2342 45724 2380 45780
rect 2436 45724 2446 45780
rect 6402 45724 6412 45780
rect 6468 45724 8428 45780
rect 8484 45724 8494 45780
rect 10994 45724 11004 45780
rect 11060 45724 11116 45780
rect 11172 45724 11182 45780
rect 11452 45668 11508 45836
rect 22764 45780 22820 46060
rect 25106 45948 25116 46004
rect 25172 45948 27244 46004
rect 27300 45948 27310 46004
rect 26226 45836 26236 45892
rect 26292 45836 27356 45892
rect 27412 45836 27804 45892
rect 27860 45836 27870 45892
rect 11666 45724 11676 45780
rect 11732 45724 12236 45780
rect 12292 45724 12302 45780
rect 17490 45724 17500 45780
rect 17556 45724 17836 45780
rect 17892 45724 17902 45780
rect 20412 45724 23156 45780
rect 20412 45668 20468 45724
rect 23100 45668 23156 45724
rect 5170 45612 5180 45668
rect 5236 45612 6524 45668
rect 6580 45612 6748 45668
rect 6804 45612 6814 45668
rect 8194 45612 8204 45668
rect 8260 45612 10444 45668
rect 10500 45612 10510 45668
rect 11452 45612 12124 45668
rect 12180 45612 12190 45668
rect 14466 45612 14476 45668
rect 14532 45612 14700 45668
rect 14756 45612 14766 45668
rect 19618 45612 19628 45668
rect 19684 45612 20412 45668
rect 20468 45612 20478 45668
rect 23090 45612 23100 45668
rect 23156 45612 23166 45668
rect 24322 45612 24332 45668
rect 24388 45612 24668 45668
rect 24724 45612 24780 45668
rect 24836 45612 24846 45668
rect 6150 45500 6188 45556
rect 6244 45500 6254 45556
rect 6748 45500 7756 45556
rect 7812 45500 7822 45556
rect 8418 45500 8428 45556
rect 8484 45500 9436 45556
rect 9492 45500 9502 45556
rect 9650 45500 9660 45556
rect 9716 45500 11228 45556
rect 11284 45500 11452 45556
rect 11508 45500 11518 45556
rect 6748 45444 6804 45500
rect 8006 45444 8016 45500
rect 8072 45444 8120 45500
rect 8176 45444 8224 45500
rect 8280 45444 8290 45500
rect 14810 45444 14820 45500
rect 14876 45444 14924 45500
rect 14980 45444 15028 45500
rect 15084 45444 15094 45500
rect 21614 45444 21624 45500
rect 21680 45444 21728 45500
rect 21784 45444 21832 45500
rect 21888 45444 21898 45500
rect 28418 45444 28428 45500
rect 28484 45444 28532 45500
rect 28588 45444 28636 45500
rect 28692 45444 28702 45500
rect 4050 45388 4060 45444
rect 4116 45388 5180 45444
rect 5236 45388 5246 45444
rect 6066 45388 6076 45444
rect 6132 45388 6748 45444
rect 6804 45388 6814 45444
rect 6962 45388 6972 45444
rect 7028 45388 7066 45444
rect 7186 45388 7196 45444
rect 7252 45388 7644 45444
rect 7700 45388 7710 45444
rect 9202 45388 9212 45444
rect 9268 45388 9772 45444
rect 9828 45388 9838 45444
rect 19730 45388 19740 45444
rect 19796 45388 20860 45444
rect 20916 45388 20926 45444
rect 22082 45388 22092 45444
rect 22148 45388 23548 45444
rect 23604 45388 23884 45444
rect 23940 45388 23950 45444
rect 25778 45388 25788 45444
rect 25844 45388 26236 45444
rect 26292 45388 26302 45444
rect 2370 45276 2380 45332
rect 2436 45276 2828 45332
rect 2884 45276 2894 45332
rect 5730 45276 5740 45332
rect 5796 45276 6636 45332
rect 6692 45276 7084 45332
rect 7140 45276 7150 45332
rect 8418 45276 8428 45332
rect 8484 45276 13468 45332
rect 13524 45276 13534 45332
rect 13682 45276 13692 45332
rect 13748 45276 14588 45332
rect 14644 45276 14654 45332
rect 14914 45276 14924 45332
rect 14980 45276 15708 45332
rect 15764 45276 16156 45332
rect 16212 45276 16222 45332
rect 17154 45276 17164 45332
rect 17220 45276 17612 45332
rect 17668 45276 17678 45332
rect 20738 45276 20748 45332
rect 20804 45276 23996 45332
rect 24052 45276 24062 45332
rect 3602 45164 3612 45220
rect 3668 45164 4620 45220
rect 4676 45164 9548 45220
rect 9604 45164 9614 45220
rect 12338 45164 12348 45220
rect 12404 45164 13244 45220
rect 13300 45164 18004 45220
rect 18386 45164 18396 45220
rect 18452 45164 18844 45220
rect 18900 45164 20524 45220
rect 20580 45164 20590 45220
rect 0 45108 400 45136
rect 0 45052 1708 45108
rect 1764 45052 1774 45108
rect 2818 45052 2828 45108
rect 2884 45052 3388 45108
rect 5954 45052 5964 45108
rect 6020 45052 9100 45108
rect 9156 45052 12740 45108
rect 12898 45052 12908 45108
rect 12964 45052 13468 45108
rect 13524 45052 13534 45108
rect 0 45024 400 45052
rect 3332 44940 3388 45052
rect 12684 44996 12740 45052
rect 3444 44940 3454 44996
rect 4834 44940 4844 44996
rect 4900 44940 6300 44996
rect 6356 44940 6366 44996
rect 7186 44940 7196 44996
rect 7252 44940 7532 44996
rect 7588 44940 7598 44996
rect 7970 44940 7980 44996
rect 8036 44940 8652 44996
rect 8708 44940 8718 44996
rect 8978 44940 8988 44996
rect 9044 44940 10108 44996
rect 10164 44940 11788 44996
rect 11844 44940 11854 44996
rect 12684 44940 13692 44996
rect 13748 44940 13758 44996
rect 8988 44884 9044 44940
rect 1922 44828 1932 44884
rect 1988 44828 2828 44884
rect 2884 44828 2894 44884
rect 6738 44828 6748 44884
rect 6804 44828 9044 44884
rect 10770 44828 10780 44884
rect 10836 44828 15372 44884
rect 15428 44828 15438 44884
rect 3686 44716 3724 44772
rect 3780 44716 3790 44772
rect 9650 44716 9660 44772
rect 9716 44716 11004 44772
rect 11060 44716 11070 44772
rect 12114 44716 12124 44772
rect 12180 44716 12190 44772
rect 13794 44716 13804 44772
rect 13860 44716 14812 44772
rect 14868 44716 14878 44772
rect 4604 44660 4614 44716
rect 4670 44660 4718 44716
rect 4774 44660 4822 44716
rect 4878 44660 4888 44716
rect 11408 44660 11418 44716
rect 11474 44660 11522 44716
rect 11578 44660 11626 44716
rect 11682 44660 11692 44716
rect 12124 44660 12180 44716
rect 17948 44660 18004 45164
rect 21186 45052 21196 45108
rect 21252 45052 25564 45108
rect 25620 45052 26796 45108
rect 26852 45052 27468 45108
rect 27524 45052 28140 45108
rect 28196 45052 28206 45108
rect 21746 44940 21756 44996
rect 21812 44940 21980 44996
rect 22036 44940 24444 44996
rect 24500 44940 24510 44996
rect 26450 44940 26460 44996
rect 26516 44940 27356 44996
rect 27412 44940 27422 44996
rect 22306 44828 22316 44884
rect 22372 44828 25228 44884
rect 25284 44828 27132 44884
rect 27188 44828 27198 44884
rect 18212 44660 18222 44716
rect 18278 44660 18326 44716
rect 18382 44660 18430 44716
rect 18486 44660 18496 44716
rect 25016 44660 25026 44716
rect 25082 44660 25130 44716
rect 25186 44660 25234 44716
rect 25290 44660 25300 44716
rect 3798 44604 3836 44660
rect 3892 44604 3902 44660
rect 6738 44604 6748 44660
rect 6804 44604 7532 44660
rect 7588 44604 7598 44660
rect 12086 44604 12124 44660
rect 12180 44604 13468 44660
rect 13524 44604 13534 44660
rect 17938 44604 17948 44660
rect 18004 44604 18014 44660
rect 3602 44492 3612 44548
rect 3668 44492 3948 44548
rect 4004 44492 4014 44548
rect 6178 44492 6188 44548
rect 6244 44492 6860 44548
rect 6916 44492 6926 44548
rect 7858 44492 7868 44548
rect 7924 44492 9436 44548
rect 9492 44492 9502 44548
rect 10434 44492 10444 44548
rect 10500 44492 10668 44548
rect 10724 44492 10734 44548
rect 13542 44492 13580 44548
rect 13636 44492 13646 44548
rect 14578 44492 14588 44548
rect 14644 44492 14654 44548
rect 15092 44492 17500 44548
rect 17556 44492 17836 44548
rect 17892 44492 17902 44548
rect 14588 44436 14644 44492
rect 15092 44436 15148 44492
rect 2818 44380 2828 44436
rect 2884 44380 3724 44436
rect 3780 44380 3790 44436
rect 7186 44380 7196 44436
rect 7252 44380 7980 44436
rect 8036 44380 8046 44436
rect 8866 44380 8876 44436
rect 8932 44380 8942 44436
rect 10770 44380 10780 44436
rect 10836 44380 11340 44436
rect 11396 44380 11406 44436
rect 12562 44380 12572 44436
rect 12628 44380 13692 44436
rect 13748 44380 13758 44436
rect 13906 44380 13916 44436
rect 13972 44380 14010 44436
rect 14578 44380 14588 44436
rect 14644 44380 15148 44436
rect 16930 44380 16940 44436
rect 16996 44380 17500 44436
rect 17556 44380 17566 44436
rect 8876 44324 8932 44380
rect 5842 44268 5852 44324
rect 5908 44268 6748 44324
rect 6804 44268 7308 44324
rect 7364 44268 7374 44324
rect 7634 44268 7644 44324
rect 7700 44268 9156 44324
rect 10882 44268 10892 44324
rect 10948 44268 11676 44324
rect 11732 44268 12236 44324
rect 12292 44268 12302 44324
rect 12898 44268 12908 44324
rect 12964 44268 17612 44324
rect 17668 44268 21420 44324
rect 21476 44268 22988 44324
rect 23044 44268 23054 44324
rect 23734 44268 23772 44324
rect 23828 44268 23838 44324
rect 9100 44212 9156 44268
rect 2482 44156 2492 44212
rect 2548 44156 3388 44212
rect 3444 44156 5628 44212
rect 5684 44156 5694 44212
rect 5842 44156 5852 44212
rect 5908 44156 5964 44212
rect 6020 44156 6030 44212
rect 6290 44156 6300 44212
rect 6356 44156 7868 44212
rect 7924 44156 7934 44212
rect 9100 44156 9772 44212
rect 9828 44156 9838 44212
rect 10994 44156 11004 44212
rect 11060 44156 12012 44212
rect 12068 44156 12796 44212
rect 12852 44156 12862 44212
rect 13458 44156 13468 44212
rect 13524 44156 19180 44212
rect 19236 44156 19292 44212
rect 19348 44156 21700 44212
rect 21858 44156 21868 44212
rect 21924 44156 22764 44212
rect 22820 44156 22830 44212
rect 3042 44044 3052 44100
rect 3108 44044 3836 44100
rect 3892 44044 3902 44100
rect 5170 44044 5180 44100
rect 5236 44044 6188 44100
rect 6244 44044 8652 44100
rect 8708 44044 8718 44100
rect 9100 43988 9156 44156
rect 21644 44100 21700 44156
rect 12450 44044 12460 44100
rect 12516 44044 13916 44100
rect 13972 44044 14644 44100
rect 16146 44044 16156 44100
rect 16212 44044 17500 44100
rect 17556 44044 17566 44100
rect 20178 44044 20188 44100
rect 20244 44044 20524 44100
rect 20580 44044 20590 44100
rect 21644 44044 22092 44100
rect 22148 44044 22158 44100
rect 6738 43932 6748 43988
rect 6804 43932 6842 43988
rect 8652 43932 9156 43988
rect 13682 43932 13692 43988
rect 13748 43932 14252 43988
rect 14308 43932 14318 43988
rect 8006 43876 8016 43932
rect 8072 43876 8120 43932
rect 8176 43876 8224 43932
rect 8280 43876 8290 43932
rect 8652 43876 8708 43932
rect 14588 43876 14644 44044
rect 14810 43876 14820 43932
rect 14876 43876 14924 43932
rect 14980 43876 15028 43932
rect 15084 43876 15094 43932
rect 21614 43876 21624 43932
rect 21680 43876 21728 43932
rect 21784 43876 21832 43932
rect 21888 43876 21898 43932
rect 28418 43876 28428 43932
rect 28484 43876 28532 43932
rect 28588 43876 28636 43932
rect 28692 43876 28702 43932
rect 8642 43820 8652 43876
rect 8708 43820 8718 43876
rect 10518 43820 10556 43876
rect 10612 43820 10622 43876
rect 10994 43820 11004 43876
rect 11060 43820 11228 43876
rect 11284 43820 14364 43876
rect 14420 43820 14430 43876
rect 14578 43820 14588 43876
rect 14644 43820 14654 43876
rect 15250 43820 15260 43876
rect 15316 43820 21476 43876
rect 23398 43820 23436 43876
rect 23492 43820 23502 43876
rect 25554 43820 25564 43876
rect 25620 43820 26684 43876
rect 26740 43820 26750 43876
rect 21420 43764 21476 43820
rect 1810 43708 1820 43764
rect 1876 43708 2156 43764
rect 2212 43708 2222 43764
rect 2370 43708 2380 43764
rect 2436 43708 3164 43764
rect 3220 43708 5796 43764
rect 13906 43708 13916 43764
rect 13972 43708 16604 43764
rect 16660 43708 16670 43764
rect 20178 43708 20188 43764
rect 20244 43708 20748 43764
rect 20804 43708 20814 43764
rect 21420 43708 25452 43764
rect 25508 43708 25788 43764
rect 25844 43708 25854 43764
rect 26002 43708 26012 43764
rect 26068 43708 26078 43764
rect 2482 43596 2492 43652
rect 2548 43596 3164 43652
rect 3220 43596 4172 43652
rect 4228 43596 4238 43652
rect 5740 43540 5796 43708
rect 26012 43652 26068 43708
rect 10994 43596 11004 43652
rect 11060 43596 16156 43652
rect 16212 43596 16222 43652
rect 16370 43596 16380 43652
rect 16436 43596 17948 43652
rect 18004 43596 19404 43652
rect 19460 43596 19470 43652
rect 21270 43596 21308 43652
rect 21364 43596 21374 43652
rect 22082 43596 22092 43652
rect 22148 43596 25564 43652
rect 25620 43596 25630 43652
rect 26012 43596 28140 43652
rect 28196 43596 28206 43652
rect 26460 43540 26516 43596
rect 3042 43484 3052 43540
rect 3108 43484 4396 43540
rect 4452 43484 4462 43540
rect 5730 43484 5740 43540
rect 5796 43484 6412 43540
rect 6468 43484 6478 43540
rect 8530 43484 8540 43540
rect 8596 43484 10892 43540
rect 10948 43484 11340 43540
rect 11396 43484 11406 43540
rect 11778 43484 11788 43540
rect 11844 43484 13804 43540
rect 13860 43484 13870 43540
rect 14578 43484 14588 43540
rect 14644 43484 14700 43540
rect 14756 43484 14766 43540
rect 15026 43484 15036 43540
rect 15092 43484 15260 43540
rect 15316 43484 15326 43540
rect 16146 43484 16156 43540
rect 16212 43484 19292 43540
rect 19348 43484 19358 43540
rect 20850 43484 20860 43540
rect 20916 43484 26292 43540
rect 26450 43484 26460 43540
rect 26516 43484 26526 43540
rect 26786 43484 26796 43540
rect 26852 43484 27244 43540
rect 27300 43484 27310 43540
rect 26236 43428 26292 43484
rect 3826 43372 3836 43428
rect 3892 43372 5964 43428
rect 6020 43372 9660 43428
rect 9716 43372 9726 43428
rect 13794 43372 13804 43428
rect 13860 43372 18172 43428
rect 18228 43372 18238 43428
rect 18498 43372 18508 43428
rect 18564 43372 18620 43428
rect 18676 43372 18686 43428
rect 26226 43372 26236 43428
rect 26292 43372 27356 43428
rect 27412 43372 27692 43428
rect 27748 43372 27758 43428
rect 14354 43260 14364 43316
rect 14420 43260 16044 43316
rect 16100 43260 16110 43316
rect 16706 43260 16716 43316
rect 16772 43260 20300 43316
rect 20356 43260 22540 43316
rect 22596 43260 22606 43316
rect 25890 43260 25900 43316
rect 25956 43260 26348 43316
rect 26404 43260 26414 43316
rect 26534 43260 26572 43316
rect 26628 43260 26638 43316
rect 9650 43148 9660 43204
rect 9716 43148 10892 43204
rect 10948 43148 10958 43204
rect 20962 43148 20972 43204
rect 21028 43148 21644 43204
rect 21700 43148 21710 43204
rect 4604 43092 4614 43148
rect 4670 43092 4718 43148
rect 4774 43092 4822 43148
rect 4878 43092 4888 43148
rect 11408 43092 11418 43148
rect 11474 43092 11522 43148
rect 11578 43092 11626 43148
rect 11682 43092 11692 43148
rect 18212 43092 18222 43148
rect 18278 43092 18326 43148
rect 18382 43092 18430 43148
rect 18486 43092 18496 43148
rect 25016 43092 25026 43148
rect 25082 43092 25130 43148
rect 25186 43092 25234 43148
rect 25290 43092 25300 43148
rect 10294 43036 10332 43092
rect 10388 43036 10398 43092
rect 7186 42924 7196 42980
rect 7252 42924 8540 42980
rect 8596 42924 8606 42980
rect 9314 42924 9324 42980
rect 9380 42924 9660 42980
rect 9716 42924 9726 42980
rect 12086 42924 12124 42980
rect 12180 42924 12190 42980
rect 4946 42812 4956 42868
rect 5012 42812 6076 42868
rect 6132 42812 12684 42868
rect 12740 42812 12750 42868
rect 13794 42812 13804 42868
rect 13860 42812 16492 42868
rect 16548 42812 20804 42868
rect 20748 42756 20804 42812
rect 7746 42700 7756 42756
rect 7812 42700 16716 42756
rect 16772 42700 16782 42756
rect 20066 42700 20076 42756
rect 20132 42700 20142 42756
rect 20738 42700 20748 42756
rect 20804 42700 22540 42756
rect 22596 42700 23436 42756
rect 23492 42700 25564 42756
rect 25620 42700 27692 42756
rect 27748 42700 27758 42756
rect 20076 42644 20132 42700
rect 4610 42588 4620 42644
rect 4676 42588 10780 42644
rect 10836 42588 10846 42644
rect 11106 42588 11116 42644
rect 11172 42588 20132 42644
rect 23874 42588 23884 42644
rect 23940 42588 26684 42644
rect 26740 42588 26750 42644
rect 6962 42476 6972 42532
rect 7028 42476 10444 42532
rect 10500 42476 10510 42532
rect 10994 42476 11004 42532
rect 11060 42476 11070 42532
rect 11554 42476 11564 42532
rect 11620 42476 12012 42532
rect 12068 42476 14140 42532
rect 14196 42476 14206 42532
rect 14354 42476 14364 42532
rect 14420 42476 15260 42532
rect 15316 42476 18284 42532
rect 18340 42476 18350 42532
rect 19170 42476 19180 42532
rect 19236 42476 21308 42532
rect 21364 42476 22204 42532
rect 22260 42476 22270 42532
rect 23650 42476 23660 42532
rect 23716 42476 24444 42532
rect 24500 42476 24510 42532
rect 0 42420 400 42448
rect 11004 42420 11060 42476
rect 0 42364 1708 42420
rect 1764 42364 1774 42420
rect 9874 42364 9884 42420
rect 9940 42364 10556 42420
rect 10612 42364 11060 42420
rect 12422 42364 12460 42420
rect 12516 42364 13916 42420
rect 13972 42364 13982 42420
rect 0 42336 400 42364
rect 8006 42308 8016 42364
rect 8072 42308 8120 42364
rect 8176 42308 8224 42364
rect 8280 42308 8290 42364
rect 14810 42308 14820 42364
rect 14876 42308 14924 42364
rect 14980 42308 15028 42364
rect 15084 42308 15094 42364
rect 21614 42308 21624 42364
rect 21680 42308 21728 42364
rect 21784 42308 21832 42364
rect 21888 42308 21898 42364
rect 28418 42308 28428 42364
rect 28484 42308 28532 42364
rect 28588 42308 28636 42364
rect 28692 42308 28702 42364
rect 9538 42252 9548 42308
rect 9604 42252 9996 42308
rect 10052 42252 10062 42308
rect 16818 42252 16828 42308
rect 16884 42252 17612 42308
rect 17668 42252 18732 42308
rect 18788 42252 18798 42308
rect 8306 42140 8316 42196
rect 8372 42140 9884 42196
rect 9940 42140 9950 42196
rect 11218 42140 11228 42196
rect 11284 42140 12236 42196
rect 12292 42140 12302 42196
rect 20290 42140 20300 42196
rect 20356 42140 20860 42196
rect 20916 42140 20926 42196
rect 21858 42140 21868 42196
rect 21924 42140 23436 42196
rect 23492 42140 23502 42196
rect 23986 42140 23996 42196
rect 24052 42140 24108 42196
rect 24164 42140 24174 42196
rect 24630 42140 24668 42196
rect 24724 42140 24734 42196
rect 4834 42028 4844 42084
rect 4900 42028 5740 42084
rect 5796 42028 5806 42084
rect 10994 42028 11004 42084
rect 11060 42028 11676 42084
rect 11732 42028 11742 42084
rect 15698 42028 15708 42084
rect 15764 42028 16828 42084
rect 16884 42028 16894 42084
rect 18498 42028 18508 42084
rect 18564 42028 18620 42084
rect 18676 42028 19404 42084
rect 19460 42028 20972 42084
rect 21028 42028 21038 42084
rect 22082 42028 22092 42084
rect 22148 42028 24108 42084
rect 24164 42028 24174 42084
rect 24322 42028 24332 42084
rect 24388 42028 26124 42084
rect 26180 42028 26190 42084
rect 2706 41916 2716 41972
rect 2772 41916 3724 41972
rect 3780 41916 3790 41972
rect 4162 41916 4172 41972
rect 4228 41916 5068 41972
rect 5124 41916 5134 41972
rect 7858 41916 7868 41972
rect 7924 41916 8092 41972
rect 8148 41916 8158 41972
rect 10434 41916 10444 41972
rect 10500 41916 12124 41972
rect 12180 41916 12190 41972
rect 12338 41916 12348 41972
rect 12404 41916 14812 41972
rect 14868 41916 14878 41972
rect 15092 41916 17612 41972
rect 17668 41916 17678 41972
rect 18050 41916 18060 41972
rect 18116 41916 18396 41972
rect 18452 41916 18462 41972
rect 18834 41916 18844 41972
rect 18900 41916 19068 41972
rect 19124 41916 19134 41972
rect 19954 41916 19964 41972
rect 20020 41916 20300 41972
rect 20356 41916 20366 41972
rect 21046 41916 21084 41972
rect 21140 41916 21150 41972
rect 21410 41916 21420 41972
rect 21476 41916 23884 41972
rect 23940 41916 23950 41972
rect 24658 41916 24668 41972
rect 24724 41916 24780 41972
rect 24836 41916 25564 41972
rect 25620 41916 25630 41972
rect 27458 41916 27468 41972
rect 27524 41916 28028 41972
rect 28084 41916 28094 41972
rect 7868 41860 7924 41916
rect 6850 41804 6860 41860
rect 6916 41804 7924 41860
rect 9846 41804 9884 41860
rect 9940 41804 9950 41860
rect 10322 41804 10332 41860
rect 10388 41804 10398 41860
rect 10770 41804 10780 41860
rect 10836 41804 12236 41860
rect 12292 41804 12302 41860
rect 13010 41804 13020 41860
rect 13076 41804 13580 41860
rect 13636 41804 13646 41860
rect 10332 41748 10388 41804
rect 15092 41748 15148 41916
rect 19068 41860 19124 41916
rect 15362 41804 15372 41860
rect 15428 41804 19124 41860
rect 20626 41804 20636 41860
rect 20692 41804 24556 41860
rect 24612 41804 24622 41860
rect 25218 41804 25228 41860
rect 25284 41804 25452 41860
rect 25508 41804 25518 41860
rect 27010 41804 27020 41860
rect 27076 41804 27356 41860
rect 27412 41804 27422 41860
rect 19068 41748 19124 41804
rect 3378 41692 3388 41748
rect 3444 41692 3556 41748
rect 7522 41692 7532 41748
rect 7588 41692 9548 41748
rect 9604 41692 9614 41748
rect 10332 41692 15148 41748
rect 15922 41692 15932 41748
rect 15988 41692 16716 41748
rect 16772 41692 16782 41748
rect 19068 41692 20412 41748
rect 20468 41692 20478 41748
rect 21634 41692 21644 41748
rect 21700 41692 22204 41748
rect 22260 41692 22270 41748
rect 3500 41300 3556 41692
rect 14578 41580 14588 41636
rect 14644 41580 14924 41636
rect 14980 41580 14990 41636
rect 20962 41580 20972 41636
rect 21028 41580 22316 41636
rect 22372 41580 22382 41636
rect 23986 41580 23996 41636
rect 24052 41580 24668 41636
rect 24724 41580 24734 41636
rect 25554 41580 25564 41636
rect 25620 41580 26012 41636
rect 26068 41580 26078 41636
rect 4604 41524 4614 41580
rect 4670 41524 4718 41580
rect 4774 41524 4822 41580
rect 4878 41524 4888 41580
rect 11408 41524 11418 41580
rect 11474 41524 11522 41580
rect 11578 41524 11626 41580
rect 11682 41524 11692 41580
rect 18212 41524 18222 41580
rect 18278 41524 18326 41580
rect 18382 41524 18430 41580
rect 18486 41524 18496 41580
rect 25016 41524 25026 41580
rect 25082 41524 25130 41580
rect 25186 41524 25234 41580
rect 25290 41524 25300 41580
rect 15586 41468 15596 41524
rect 15652 41468 15662 41524
rect 17686 41468 17724 41524
rect 17780 41468 17790 41524
rect 15596 41412 15652 41468
rect 15250 41356 15260 41412
rect 15316 41356 18284 41412
rect 18340 41356 18350 41412
rect 19282 41356 19292 41412
rect 19348 41356 19404 41412
rect 19460 41356 21420 41412
rect 21476 41356 21486 41412
rect 3490 41244 3500 41300
rect 3556 41244 3566 41300
rect 4946 41244 4956 41300
rect 5012 41244 5628 41300
rect 5684 41244 5694 41300
rect 9986 41244 9996 41300
rect 10052 41244 10556 41300
rect 10612 41244 10622 41300
rect 10882 41244 10892 41300
rect 10948 41244 11788 41300
rect 11844 41244 12012 41300
rect 12068 41244 12078 41300
rect 12226 41244 12236 41300
rect 12292 41244 15372 41300
rect 15428 41244 15438 41300
rect 18834 41244 18844 41300
rect 18900 41244 19516 41300
rect 19572 41244 19582 41300
rect 22866 41244 22876 41300
rect 22932 41244 25116 41300
rect 25172 41244 25182 41300
rect 25340 41244 27580 41300
rect 27636 41244 27646 41300
rect 3826 41132 3836 41188
rect 3892 41132 3902 41188
rect 6514 41132 6524 41188
rect 6580 41132 7644 41188
rect 7700 41132 7710 41188
rect 8082 41132 8092 41188
rect 8148 41132 13244 41188
rect 13300 41132 13748 41188
rect 3836 40964 3892 41132
rect 13692 41076 13748 41132
rect 14028 41132 16044 41188
rect 16100 41132 16110 41188
rect 21858 41132 21868 41188
rect 21924 41132 23212 41188
rect 23268 41132 23278 41188
rect 23538 41132 23548 41188
rect 23604 41132 23772 41188
rect 23828 41132 23838 41188
rect 6290 41020 6300 41076
rect 6356 41020 7196 41076
rect 7252 41020 7262 41076
rect 13010 41020 13020 41076
rect 13076 41020 13244 41076
rect 13300 41020 13310 41076
rect 13692 41020 13804 41076
rect 13860 41020 13870 41076
rect 14028 40964 14084 41132
rect 25340 41076 25396 41244
rect 26226 41132 26236 41188
rect 26292 41132 26572 41188
rect 26628 41132 26638 41188
rect 26786 41132 26796 41188
rect 26852 41132 26862 41188
rect 26796 41076 26852 41132
rect 16706 41020 16716 41076
rect 16772 41020 18620 41076
rect 18676 41020 18686 41076
rect 22428 41020 25396 41076
rect 26012 41020 27580 41076
rect 27636 41020 27646 41076
rect 22428 40964 22484 41020
rect 26012 40964 26068 41020
rect 2034 40908 2044 40964
rect 2100 40908 3052 40964
rect 3108 40908 3118 40964
rect 3836 40908 4396 40964
rect 4452 40908 4462 40964
rect 5068 40908 14084 40964
rect 15138 40908 15148 40964
rect 15204 40908 17948 40964
rect 18004 40908 19740 40964
rect 19796 40908 19964 40964
rect 20020 40908 22316 40964
rect 22372 40908 22484 40964
rect 23538 40908 23548 40964
rect 23604 40908 23642 40964
rect 24210 40908 24220 40964
rect 24276 40908 25788 40964
rect 25844 40908 26068 40964
rect 26786 40908 26796 40964
rect 26852 40908 27020 40964
rect 27076 40908 27086 40964
rect 5068 40852 5124 40908
rect 23548 40852 23604 40908
rect 2370 40796 2380 40852
rect 2436 40796 3164 40852
rect 3220 40796 3500 40852
rect 3556 40796 3566 40852
rect 4162 40796 4172 40852
rect 4228 40796 5124 40852
rect 7298 40796 7308 40852
rect 7364 40796 7868 40852
rect 7924 40796 7934 40852
rect 10322 40796 10332 40852
rect 10388 40796 10780 40852
rect 10836 40796 10846 40852
rect 11190 40796 11228 40852
rect 11284 40796 11294 40852
rect 11778 40796 11788 40852
rect 11844 40796 12236 40852
rect 12292 40796 12302 40852
rect 19366 40796 19404 40852
rect 19460 40796 19470 40852
rect 20066 40796 20076 40852
rect 20132 40796 21420 40852
rect 21476 40796 21486 40852
rect 23548 40796 25340 40852
rect 25396 40796 25452 40852
rect 25508 40796 25518 40852
rect 8006 40740 8016 40796
rect 8072 40740 8120 40796
rect 8176 40740 8224 40796
rect 8280 40740 8290 40796
rect 14810 40740 14820 40796
rect 14876 40740 14924 40796
rect 14980 40740 15028 40796
rect 15084 40740 15094 40796
rect 21614 40740 21624 40796
rect 21680 40740 21728 40796
rect 21784 40740 21832 40796
rect 21888 40740 21898 40796
rect 28418 40740 28428 40796
rect 28484 40740 28532 40796
rect 28588 40740 28636 40796
rect 28692 40740 28702 40796
rect 7746 40684 7756 40740
rect 7812 40684 7822 40740
rect 10882 40684 10892 40740
rect 10948 40684 11564 40740
rect 11620 40684 11630 40740
rect 16706 40684 16716 40740
rect 16772 40684 21084 40740
rect 21140 40684 21150 40740
rect 7756 40628 7812 40684
rect 2930 40572 2940 40628
rect 2996 40572 3006 40628
rect 4274 40572 4284 40628
rect 4340 40572 5516 40628
rect 5572 40572 5582 40628
rect 7756 40572 8260 40628
rect 9650 40572 9660 40628
rect 9716 40572 11228 40628
rect 11284 40572 11294 40628
rect 12898 40572 12908 40628
rect 12964 40572 13468 40628
rect 13524 40572 14028 40628
rect 14084 40572 15260 40628
rect 15316 40572 15326 40628
rect 20290 40572 20300 40628
rect 20356 40572 23324 40628
rect 23380 40572 23390 40628
rect 26226 40572 26236 40628
rect 26292 40572 26908 40628
rect 26964 40572 26974 40628
rect 28130 40572 28140 40628
rect 28196 40572 28206 40628
rect 2940 40516 2996 40572
rect 8204 40516 8260 40572
rect 2482 40460 2492 40516
rect 2548 40460 2996 40516
rect 6514 40460 6524 40516
rect 6580 40460 7756 40516
rect 7812 40460 7822 40516
rect 8194 40460 8204 40516
rect 8260 40460 11116 40516
rect 11172 40460 12796 40516
rect 12852 40460 12862 40516
rect 19954 40460 19964 40516
rect 20020 40460 20412 40516
rect 20468 40460 21980 40516
rect 22036 40460 22046 40516
rect 22866 40460 22876 40516
rect 22932 40460 23660 40516
rect 23716 40460 23726 40516
rect 24070 40460 24108 40516
rect 24164 40460 24174 40516
rect 26338 40460 26348 40516
rect 26404 40460 27132 40516
rect 27188 40460 27198 40516
rect 28140 40404 28196 40572
rect 2034 40348 2044 40404
rect 2100 40348 2828 40404
rect 2884 40348 3612 40404
rect 3668 40348 3678 40404
rect 8530 40348 8540 40404
rect 8596 40348 8988 40404
rect 9044 40348 11788 40404
rect 11844 40348 12460 40404
rect 12516 40348 12526 40404
rect 18274 40348 18284 40404
rect 18340 40348 20300 40404
rect 20356 40348 20748 40404
rect 20804 40348 20814 40404
rect 26786 40348 26796 40404
rect 26852 40348 28196 40404
rect 7074 40236 7084 40292
rect 7140 40236 8428 40292
rect 8484 40236 8494 40292
rect 9538 40236 9548 40292
rect 9604 40236 12236 40292
rect 12292 40236 13580 40292
rect 13636 40236 13646 40292
rect 16146 40236 16156 40292
rect 16212 40236 18844 40292
rect 18900 40236 18910 40292
rect 19618 40236 19628 40292
rect 19684 40236 20636 40292
rect 20692 40236 20702 40292
rect 23426 40236 23436 40292
rect 23492 40236 23548 40292
rect 23604 40236 23614 40292
rect 25890 40236 25900 40292
rect 25956 40236 26460 40292
rect 26516 40236 26526 40292
rect 3714 40124 3724 40180
rect 3780 40124 4172 40180
rect 4228 40124 4238 40180
rect 10108 40068 10164 40236
rect 16370 40124 16380 40180
rect 16436 40124 16828 40180
rect 16884 40124 16894 40180
rect 23202 40124 23212 40180
rect 23268 40124 26572 40180
rect 26628 40124 26908 40180
rect 26964 40124 26974 40180
rect 3154 40012 3164 40068
rect 3220 40012 3388 40068
rect 5506 40012 5516 40068
rect 5572 40012 7196 40068
rect 7252 40012 7262 40068
rect 7746 40012 7756 40068
rect 7812 40012 9548 40068
rect 9604 40012 9614 40068
rect 10098 40012 10108 40068
rect 10164 40012 10174 40068
rect 11778 40012 11788 40068
rect 11844 40012 12348 40068
rect 12404 40012 12414 40068
rect 3332 39956 3388 40012
rect 4604 39956 4614 40012
rect 4670 39956 4718 40012
rect 4774 39956 4822 40012
rect 4878 39956 4888 40012
rect 11408 39956 11418 40012
rect 11474 39956 11522 40012
rect 11578 39956 11626 40012
rect 11682 39956 11692 40012
rect 18212 39956 18222 40012
rect 18278 39956 18326 40012
rect 18382 39956 18430 40012
rect 18486 39956 18496 40012
rect 25016 39956 25026 40012
rect 25082 39956 25130 40012
rect 25186 39956 25234 40012
rect 25290 39956 25300 40012
rect 3332 39900 3892 39956
rect 4386 39900 4396 39956
rect 4452 39900 4462 39956
rect 2034 39788 2044 39844
rect 2100 39788 3388 39844
rect 0 39732 400 39760
rect 0 39676 1708 39732
rect 1764 39676 1774 39732
rect 0 39648 400 39676
rect 3332 39620 3388 39788
rect 3836 39732 3892 39900
rect 4396 39844 4452 39900
rect 4050 39788 4060 39844
rect 4116 39788 5628 39844
rect 5684 39788 5694 39844
rect 10658 39788 10668 39844
rect 10724 39788 11116 39844
rect 11172 39788 11182 39844
rect 11666 39788 11676 39844
rect 11732 39788 11788 39844
rect 11844 39788 11854 39844
rect 14018 39788 14028 39844
rect 14084 39788 14700 39844
rect 14756 39788 16380 39844
rect 16436 39788 16446 39844
rect 22978 39788 22988 39844
rect 23044 39788 24444 39844
rect 24500 39788 24510 39844
rect 26786 39788 26796 39844
rect 26852 39788 27356 39844
rect 27412 39788 27422 39844
rect 27682 39788 27692 39844
rect 27748 39788 28140 39844
rect 28196 39788 28206 39844
rect 3836 39676 4396 39732
rect 4452 39676 5068 39732
rect 5124 39676 6412 39732
rect 6468 39676 6478 39732
rect 13570 39676 13580 39732
rect 13636 39676 20412 39732
rect 20468 39676 20478 39732
rect 3332 39564 13692 39620
rect 13748 39564 14140 39620
rect 14196 39564 15148 39620
rect 15204 39564 15214 39620
rect 17490 39564 17500 39620
rect 17556 39564 18620 39620
rect 18676 39564 18686 39620
rect 14914 39452 14924 39508
rect 14980 39452 15260 39508
rect 15316 39452 15326 39508
rect 15474 39452 15484 39508
rect 15540 39452 17388 39508
rect 17444 39452 17454 39508
rect 24098 39452 24108 39508
rect 24164 39452 25116 39508
rect 25172 39452 25182 39508
rect 6066 39340 6076 39396
rect 6132 39340 10164 39396
rect 17714 39340 17724 39396
rect 17780 39340 18172 39396
rect 18228 39340 19852 39396
rect 19908 39340 19918 39396
rect 21270 39340 21308 39396
rect 21364 39340 21868 39396
rect 21924 39340 21934 39396
rect 27010 39340 27020 39396
rect 27076 39340 27356 39396
rect 27412 39340 27422 39396
rect 10108 39284 10164 39340
rect 5170 39228 5180 39284
rect 5236 39228 5628 39284
rect 5684 39228 5694 39284
rect 10108 39228 11788 39284
rect 11844 39228 11854 39284
rect 16034 39228 16044 39284
rect 16100 39228 17052 39284
rect 17108 39228 17118 39284
rect 20290 39228 20300 39284
rect 20356 39228 21420 39284
rect 21476 39228 21486 39284
rect 8006 39172 8016 39228
rect 8072 39172 8120 39228
rect 8176 39172 8224 39228
rect 8280 39172 8290 39228
rect 14810 39172 14820 39228
rect 14876 39172 14924 39228
rect 14980 39172 15028 39228
rect 15084 39172 15094 39228
rect 21614 39172 21624 39228
rect 21680 39172 21728 39228
rect 21784 39172 21832 39228
rect 21888 39172 21898 39228
rect 28418 39172 28428 39228
rect 28484 39172 28532 39228
rect 28588 39172 28636 39228
rect 28692 39172 28702 39228
rect 9538 39116 9548 39172
rect 9604 39116 9996 39172
rect 10052 39116 10892 39172
rect 10948 39116 13580 39172
rect 13636 39116 13646 39172
rect 20738 39116 20748 39172
rect 20804 39116 20860 39172
rect 20916 39116 20926 39172
rect 22082 39116 22092 39172
rect 22148 39116 24668 39172
rect 24724 39116 24734 39172
rect 1810 39004 1820 39060
rect 1876 39004 2268 39060
rect 2324 39004 2334 39060
rect 3490 39004 3500 39060
rect 3556 39004 4620 39060
rect 4676 39004 15372 39060
rect 15428 39004 15438 39060
rect 16818 39004 16828 39060
rect 16884 39004 16940 39060
rect 16996 39004 23212 39060
rect 23268 39004 23278 39060
rect 24098 39004 24108 39060
rect 24164 39004 26572 39060
rect 26628 39004 26638 39060
rect 3602 38892 3612 38948
rect 3668 38892 3724 38948
rect 3780 38892 3790 38948
rect 3938 38892 3948 38948
rect 4004 38892 5068 38948
rect 5124 38892 5134 38948
rect 5282 38892 5292 38948
rect 5348 38892 6076 38948
rect 6132 38892 6142 38948
rect 7746 38892 7756 38948
rect 7812 38892 8540 38948
rect 8596 38892 17836 38948
rect 17892 38892 17902 38948
rect 19842 38892 19852 38948
rect 19908 38892 25228 38948
rect 25284 38892 27468 38948
rect 27524 38892 27534 38948
rect 7606 38780 7644 38836
rect 7700 38780 7710 38836
rect 12338 38780 12348 38836
rect 12404 38780 16828 38836
rect 16884 38780 16894 38836
rect 18498 38780 18508 38836
rect 18564 38780 19740 38836
rect 19796 38780 19806 38836
rect 20038 38780 20076 38836
rect 20132 38780 20142 38836
rect 21746 38780 21756 38836
rect 21812 38780 22764 38836
rect 22820 38780 22830 38836
rect 23650 38780 23660 38836
rect 23716 38780 23996 38836
rect 24052 38780 24062 38836
rect 26898 38780 26908 38836
rect 26964 38780 26974 38836
rect 26908 38724 26964 38780
rect 11218 38668 11228 38724
rect 11284 38668 11676 38724
rect 11732 38668 11742 38724
rect 16818 38668 16828 38724
rect 16884 38668 17612 38724
rect 17668 38668 19404 38724
rect 19460 38668 19470 38724
rect 20626 38668 20636 38724
rect 20692 38668 21980 38724
rect 22036 38668 25172 38724
rect 26226 38668 26236 38724
rect 26292 38668 26964 38724
rect 25116 38612 25284 38668
rect 11228 38556 11788 38612
rect 11844 38556 11854 38612
rect 17910 38556 17948 38612
rect 18004 38556 18014 38612
rect 21410 38556 21420 38612
rect 21476 38556 22652 38612
rect 22708 38556 22718 38612
rect 25228 38556 25676 38612
rect 25732 38556 25742 38612
rect 11228 38500 11284 38556
rect 5702 38444 5740 38500
rect 5796 38444 5806 38500
rect 11218 38444 11228 38500
rect 11284 38444 11294 38500
rect 20178 38444 20188 38500
rect 20244 38444 20748 38500
rect 20804 38444 20814 38500
rect 21158 38444 21196 38500
rect 21252 38444 21262 38500
rect 22082 38444 22092 38500
rect 22148 38444 22158 38500
rect 4604 38388 4614 38444
rect 4670 38388 4718 38444
rect 4774 38388 4822 38444
rect 4878 38388 4888 38444
rect 11408 38388 11418 38444
rect 11474 38388 11522 38444
rect 11578 38388 11626 38444
rect 11682 38388 11692 38444
rect 18212 38388 18222 38444
rect 18278 38388 18326 38444
rect 18382 38388 18430 38444
rect 18486 38388 18496 38444
rect 22092 38388 22148 38444
rect 25016 38388 25026 38444
rect 25082 38388 25130 38444
rect 25186 38388 25234 38444
rect 25290 38388 25300 38444
rect 6738 38332 6748 38388
rect 6804 38332 7420 38388
rect 7476 38332 7486 38388
rect 12758 38332 12796 38388
rect 12852 38332 12862 38388
rect 19068 38332 22148 38388
rect 19068 38276 19124 38332
rect 2342 38220 2380 38276
rect 2436 38220 2446 38276
rect 9650 38220 9660 38276
rect 9716 38220 12236 38276
rect 12292 38220 13580 38276
rect 13636 38220 19124 38276
rect 24658 38220 24668 38276
rect 24724 38220 25228 38276
rect 25284 38220 25294 38276
rect 8418 38108 8428 38164
rect 8484 38108 9100 38164
rect 9156 38108 10108 38164
rect 10164 38108 10174 38164
rect 11106 38108 11116 38164
rect 11172 38108 11228 38164
rect 11284 38108 11788 38164
rect 16482 38108 16492 38164
rect 16548 38108 16828 38164
rect 16884 38108 17500 38164
rect 17556 38108 17566 38164
rect 19282 38108 19292 38164
rect 19348 38108 20076 38164
rect 20132 38108 20142 38164
rect 23986 38108 23996 38164
rect 24052 38108 26348 38164
rect 26404 38108 26414 38164
rect 2370 37996 2380 38052
rect 2436 37996 3388 38052
rect 3444 37996 3948 38052
rect 4004 37996 4014 38052
rect 4162 37996 4172 38052
rect 4228 37996 4266 38052
rect 10770 37996 10780 38052
rect 10836 37996 11228 38052
rect 11284 37996 11294 38052
rect 11732 37940 11788 38108
rect 12674 37996 12684 38052
rect 12740 37996 15932 38052
rect 15988 37996 15998 38052
rect 21746 37996 21756 38052
rect 21812 37996 22204 38052
rect 22260 37996 22270 38052
rect 22754 37996 22764 38052
rect 22820 37996 23436 38052
rect 23492 37996 23502 38052
rect 23650 37996 23660 38052
rect 23716 37996 26460 38052
rect 26516 37996 26526 38052
rect 23660 37940 23716 37996
rect 2930 37884 2940 37940
rect 2996 37884 3388 37940
rect 11732 37884 12348 37940
rect 12404 37884 16044 37940
rect 16100 37884 16110 37940
rect 19842 37884 19852 37940
rect 19908 37884 20860 37940
rect 20916 37884 20926 37940
rect 21074 37884 21084 37940
rect 21140 37884 21420 37940
rect 21476 37884 23716 37940
rect 24098 37884 24108 37940
rect 24164 37884 24174 37940
rect 24780 37884 27356 37940
rect 27412 37884 27422 37940
rect 3332 37828 3388 37884
rect 24108 37828 24164 37884
rect 24780 37828 24836 37884
rect 3332 37772 3836 37828
rect 3892 37772 4396 37828
rect 4452 37772 4462 37828
rect 7522 37772 7532 37828
rect 7588 37772 21308 37828
rect 21364 37772 21980 37828
rect 22036 37772 22046 37828
rect 23650 37772 23660 37828
rect 23716 37772 24780 37828
rect 24836 37772 24846 37828
rect 25666 37772 25676 37828
rect 25732 37772 28140 37828
rect 28196 37772 28206 37828
rect 7158 37660 7196 37716
rect 7252 37660 7262 37716
rect 18834 37660 18844 37716
rect 18900 37660 21084 37716
rect 21140 37660 21150 37716
rect 23426 37660 23436 37716
rect 23492 37660 27692 37716
rect 27748 37660 27758 37716
rect 8006 37604 8016 37660
rect 8072 37604 8120 37660
rect 8176 37604 8224 37660
rect 8280 37604 8290 37660
rect 14810 37604 14820 37660
rect 14876 37604 14924 37660
rect 14980 37604 15028 37660
rect 15084 37604 15094 37660
rect 21614 37604 21624 37660
rect 21680 37604 21728 37660
rect 21784 37604 21832 37660
rect 21888 37604 21898 37660
rect 28418 37604 28428 37660
rect 28484 37604 28532 37660
rect 28588 37604 28636 37660
rect 28692 37604 28702 37660
rect 10322 37548 10332 37604
rect 10388 37548 11228 37604
rect 11284 37548 12236 37604
rect 12292 37548 12302 37604
rect 15922 37548 15932 37604
rect 15988 37548 20300 37604
rect 20356 37548 20366 37604
rect 20514 37548 20524 37604
rect 20580 37548 20972 37604
rect 21028 37548 21038 37604
rect 24294 37548 24332 37604
rect 24388 37548 24398 37604
rect 24770 37548 24780 37604
rect 24836 37548 25116 37604
rect 25172 37548 25676 37604
rect 25732 37548 25742 37604
rect 5170 37436 5180 37492
rect 5236 37436 6412 37492
rect 6468 37436 6478 37492
rect 7410 37436 7420 37492
rect 7476 37436 8204 37492
rect 8260 37436 8270 37492
rect 8754 37436 8764 37492
rect 8820 37436 9660 37492
rect 9716 37436 9726 37492
rect 13542 37436 13580 37492
rect 13636 37436 13646 37492
rect 13906 37436 13916 37492
rect 13972 37436 14364 37492
rect 14420 37436 14430 37492
rect 15250 37436 15260 37492
rect 15316 37436 15484 37492
rect 15540 37436 15550 37492
rect 18386 37436 18396 37492
rect 18452 37436 19292 37492
rect 19348 37436 19358 37492
rect 22082 37436 22092 37492
rect 22148 37436 22988 37492
rect 23044 37436 23212 37492
rect 23268 37436 23278 37492
rect 25218 37436 25228 37492
rect 25284 37436 25452 37492
rect 25508 37436 25518 37492
rect 25778 37436 25788 37492
rect 25844 37436 26348 37492
rect 26404 37436 26414 37492
rect 6412 37380 6468 37436
rect 4386 37324 4396 37380
rect 4452 37324 4956 37380
rect 5012 37324 5022 37380
rect 6412 37324 7532 37380
rect 7588 37324 7598 37380
rect 8642 37324 8652 37380
rect 8708 37324 10108 37380
rect 10164 37324 10174 37380
rect 10994 37324 11004 37380
rect 11060 37324 18956 37380
rect 19012 37324 19022 37380
rect 20066 37324 20076 37380
rect 20132 37324 20412 37380
rect 20468 37324 22764 37380
rect 22820 37324 22830 37380
rect 26758 37324 26796 37380
rect 26852 37324 26862 37380
rect 5068 37212 5516 37268
rect 5572 37212 5852 37268
rect 5908 37212 7420 37268
rect 7476 37212 7486 37268
rect 7970 37212 7980 37268
rect 8036 37212 8316 37268
rect 8372 37212 8382 37268
rect 9986 37212 9996 37268
rect 10052 37212 11564 37268
rect 11620 37212 11630 37268
rect 14578 37212 14588 37268
rect 14644 37212 14654 37268
rect 15026 37212 15036 37268
rect 15092 37212 22876 37268
rect 22932 37212 22942 37268
rect 24546 37212 24556 37268
rect 24612 37212 25340 37268
rect 25396 37212 25406 37268
rect 5068 37156 5124 37212
rect 14588 37156 14644 37212
rect 4050 37100 4060 37156
rect 4116 37100 5068 37156
rect 5124 37100 5134 37156
rect 5954 37100 5964 37156
rect 6020 37100 11452 37156
rect 11508 37100 11518 37156
rect 14588 37100 15596 37156
rect 15652 37100 15662 37156
rect 17378 37100 17388 37156
rect 17444 37100 18396 37156
rect 18452 37100 18844 37156
rect 18900 37100 18910 37156
rect 19506 37100 19516 37156
rect 19572 37100 21756 37156
rect 21812 37100 21822 37156
rect 21970 37100 21980 37156
rect 22036 37100 22652 37156
rect 22708 37100 24332 37156
rect 24388 37100 24398 37156
rect 0 37044 400 37072
rect 0 36988 1708 37044
rect 1764 36988 2492 37044
rect 2548 36988 2558 37044
rect 4722 36988 4732 37044
rect 4788 36988 5012 37044
rect 0 36960 400 36988
rect 4604 36820 4614 36876
rect 4670 36820 4718 36876
rect 4774 36820 4822 36876
rect 4878 36820 4888 36876
rect 4956 36820 5012 36988
rect 6972 36932 7028 37100
rect 8194 36988 8204 37044
rect 8260 36988 9324 37044
rect 9380 36988 12796 37044
rect 12852 36988 12862 37044
rect 13570 36988 13580 37044
rect 13636 36988 15484 37044
rect 15540 36988 15550 37044
rect 17938 36988 17948 37044
rect 18004 36988 18788 37044
rect 18946 36988 18956 37044
rect 19012 36988 24780 37044
rect 24836 36988 24846 37044
rect 18732 36932 18788 36988
rect 6962 36876 6972 36932
rect 7028 36876 7038 36932
rect 10406 36876 10444 36932
rect 10500 36876 10510 36932
rect 10966 36876 11004 36932
rect 11060 36876 11070 36932
rect 12898 36876 12908 36932
rect 12964 36876 13692 36932
rect 13748 36876 13758 36932
rect 18732 36876 19404 36932
rect 19460 36876 19964 36932
rect 20020 36876 20030 36932
rect 26226 36876 26236 36932
rect 26292 36876 26628 36932
rect 11408 36820 11418 36876
rect 11474 36820 11522 36876
rect 11578 36820 11626 36876
rect 11682 36820 11692 36876
rect 18212 36820 18222 36876
rect 18278 36820 18326 36876
rect 18382 36820 18430 36876
rect 18486 36820 18496 36876
rect 25016 36820 25026 36876
rect 25082 36820 25130 36876
rect 25186 36820 25234 36876
rect 25290 36820 25300 36876
rect 26572 36820 26628 36876
rect 4956 36764 8204 36820
rect 8260 36764 8270 36820
rect 9874 36764 9884 36820
rect 9940 36764 10556 36820
rect 10612 36764 10622 36820
rect 12758 36764 12796 36820
rect 12852 36764 12862 36820
rect 15138 36764 15148 36820
rect 15204 36764 16044 36820
rect 16100 36764 16110 36820
rect 18610 36764 18620 36820
rect 18676 36764 19180 36820
rect 19236 36764 23212 36820
rect 23268 36764 23278 36820
rect 26562 36764 26572 36820
rect 26628 36764 26638 36820
rect 4956 36708 5012 36764
rect 3266 36652 3276 36708
rect 3332 36652 5012 36708
rect 6850 36652 6860 36708
rect 6916 36652 6972 36708
rect 7028 36652 7038 36708
rect 11778 36652 11788 36708
rect 11844 36652 14028 36708
rect 14084 36652 14094 36708
rect 14326 36652 14364 36708
rect 14420 36652 14430 36708
rect 15698 36652 15708 36708
rect 15764 36652 25452 36708
rect 25508 36652 26236 36708
rect 26292 36652 26302 36708
rect 3938 36540 3948 36596
rect 4004 36540 5180 36596
rect 5236 36540 5628 36596
rect 5684 36540 5694 36596
rect 12114 36540 12124 36596
rect 12180 36540 13972 36596
rect 18386 36540 18396 36596
rect 18452 36540 18620 36596
rect 18676 36540 18686 36596
rect 24770 36540 24780 36596
rect 24836 36540 25228 36596
rect 25284 36540 26908 36596
rect 26964 36540 26974 36596
rect 13916 36484 13972 36540
rect 3714 36428 3724 36484
rect 3780 36428 4732 36484
rect 4788 36428 4798 36484
rect 5058 36428 5068 36484
rect 5124 36428 5964 36484
rect 6020 36428 6030 36484
rect 12674 36428 12684 36484
rect 12740 36428 13188 36484
rect 13654 36428 13692 36484
rect 13748 36428 13758 36484
rect 13906 36428 13916 36484
rect 13972 36428 13982 36484
rect 14690 36428 14700 36484
rect 14756 36428 16156 36484
rect 16212 36428 16492 36484
rect 16548 36428 16558 36484
rect 18722 36428 18732 36484
rect 18788 36428 18956 36484
rect 19012 36428 19022 36484
rect 21522 36428 21532 36484
rect 21588 36428 22988 36484
rect 23044 36428 23054 36484
rect 24210 36428 24220 36484
rect 24276 36428 27020 36484
rect 27076 36428 27086 36484
rect 13132 36372 13188 36428
rect 3332 36316 4956 36372
rect 5012 36316 6748 36372
rect 6804 36316 6814 36372
rect 9986 36316 9996 36372
rect 10052 36316 12124 36372
rect 12180 36316 12572 36372
rect 12628 36316 12638 36372
rect 13132 36316 13468 36372
rect 13524 36316 13534 36372
rect 13766 36316 13804 36372
rect 13860 36316 13870 36372
rect 15092 36316 16604 36372
rect 16660 36316 17612 36372
rect 17668 36316 17678 36372
rect 26758 36316 26796 36372
rect 26852 36316 26862 36372
rect 3332 36260 3388 36316
rect 15092 36260 15148 36316
rect 2034 36204 2044 36260
rect 2100 36204 3388 36260
rect 3938 36204 3948 36260
rect 4004 36204 4396 36260
rect 4452 36204 6412 36260
rect 6468 36204 6478 36260
rect 11218 36204 11228 36260
rect 11284 36204 15148 36260
rect 15362 36204 15372 36260
rect 15428 36204 15708 36260
rect 15764 36204 15774 36260
rect 16258 36204 16268 36260
rect 16324 36204 17164 36260
rect 17220 36204 19852 36260
rect 19908 36204 19918 36260
rect 21420 36204 21644 36260
rect 21700 36204 21710 36260
rect 3826 36092 3836 36148
rect 3892 36092 4956 36148
rect 5012 36092 5022 36148
rect 6178 36092 6188 36148
rect 6244 36092 6748 36148
rect 6804 36092 6814 36148
rect 8006 36036 8016 36092
rect 8072 36036 8120 36092
rect 8176 36036 8224 36092
rect 8280 36036 8290 36092
rect 12572 36036 12628 36204
rect 21420 36148 21476 36204
rect 17462 36092 17500 36148
rect 17556 36092 17566 36148
rect 21410 36092 21420 36148
rect 21476 36092 21486 36148
rect 14810 36036 14820 36092
rect 14876 36036 14924 36092
rect 14980 36036 15028 36092
rect 15084 36036 15094 36092
rect 21614 36036 21624 36092
rect 21680 36036 21728 36092
rect 21784 36036 21832 36092
rect 21888 36036 21898 36092
rect 28418 36036 28428 36092
rect 28484 36036 28532 36092
rect 28588 36036 28636 36092
rect 28692 36036 28702 36092
rect 3826 35980 3836 36036
rect 3892 35980 4060 36036
rect 4116 35980 4126 36036
rect 12562 35980 12572 36036
rect 12628 35980 12638 36036
rect 8530 35868 8540 35924
rect 8596 35868 10108 35924
rect 10164 35868 10174 35924
rect 15250 35868 15260 35924
rect 15316 35868 16044 35924
rect 16100 35868 16110 35924
rect 21298 35868 21308 35924
rect 21364 35868 22316 35924
rect 22372 35868 22382 35924
rect 4834 35756 4844 35812
rect 4900 35756 5628 35812
rect 5684 35756 5694 35812
rect 8754 35756 8764 35812
rect 8820 35756 9660 35812
rect 9716 35756 9726 35812
rect 12898 35756 12908 35812
rect 12964 35756 13356 35812
rect 13412 35756 13422 35812
rect 15474 35756 15484 35812
rect 15540 35756 16604 35812
rect 16660 35756 16670 35812
rect 7830 35644 7868 35700
rect 7924 35644 7934 35700
rect 12450 35644 12460 35700
rect 12516 35644 16044 35700
rect 16100 35644 16110 35700
rect 16706 35644 16716 35700
rect 16772 35644 17388 35700
rect 17444 35644 17454 35700
rect 10322 35532 10332 35588
rect 10388 35532 10780 35588
rect 10836 35532 11228 35588
rect 11284 35532 11294 35588
rect 11666 35532 11676 35588
rect 11732 35532 12572 35588
rect 12628 35532 12638 35588
rect 14130 35532 14140 35588
rect 14196 35532 14812 35588
rect 14868 35532 14878 35588
rect 19170 35532 19180 35588
rect 19236 35532 19516 35588
rect 19572 35532 20300 35588
rect 20356 35532 20366 35588
rect 22754 35532 22764 35588
rect 22820 35532 22988 35588
rect 23044 35532 23054 35588
rect 24658 35532 24668 35588
rect 24724 35532 25676 35588
rect 25732 35532 26572 35588
rect 26628 35532 26638 35588
rect 11106 35420 11116 35476
rect 11172 35420 11788 35476
rect 11844 35420 11854 35476
rect 14466 35420 14476 35476
rect 14532 35420 14644 35476
rect 15698 35420 15708 35476
rect 15764 35420 16380 35476
rect 16436 35420 16446 35476
rect 17714 35420 17724 35476
rect 17780 35420 17836 35476
rect 17892 35420 17902 35476
rect 18732 35420 18956 35476
rect 19012 35420 19022 35476
rect 23650 35420 23660 35476
rect 23716 35420 24108 35476
rect 24164 35420 24174 35476
rect 24322 35420 24332 35476
rect 24388 35420 25452 35476
rect 25508 35420 25518 35476
rect 14326 35308 14364 35364
rect 14420 35308 14430 35364
rect 14588 35308 14644 35420
rect 18732 35308 18788 35420
rect 18946 35308 18956 35364
rect 19012 35308 19348 35364
rect 20822 35308 20860 35364
rect 20916 35308 20926 35364
rect 22978 35308 22988 35364
rect 23044 35308 23212 35364
rect 23268 35308 23278 35364
rect 23538 35308 23548 35364
rect 23604 35308 24220 35364
rect 24276 35308 24286 35364
rect 4604 35252 4614 35308
rect 4670 35252 4718 35308
rect 4774 35252 4822 35308
rect 4878 35252 4888 35308
rect 11408 35252 11418 35308
rect 11474 35252 11522 35308
rect 11578 35252 11626 35308
rect 11682 35252 11692 35308
rect 14578 35252 14588 35308
rect 14644 35252 14654 35308
rect 18212 35252 18222 35308
rect 18278 35252 18326 35308
rect 18382 35252 18430 35308
rect 18486 35252 18496 35308
rect 18722 35252 18732 35308
rect 18788 35252 18798 35308
rect 19292 35252 19348 35308
rect 25016 35252 25026 35308
rect 25082 35252 25130 35308
rect 25186 35252 25234 35308
rect 25290 35252 25300 35308
rect 1922 35196 1932 35252
rect 1988 35196 4060 35252
rect 4116 35196 4126 35252
rect 10966 35196 11004 35252
rect 11060 35196 11070 35252
rect 19292 35196 20636 35252
rect 20692 35196 20702 35252
rect 22082 35196 22092 35252
rect 22148 35196 22764 35252
rect 22820 35196 22830 35252
rect 23986 35196 23996 35252
rect 24052 35196 24668 35252
rect 24724 35196 24734 35252
rect 4060 35140 4116 35196
rect 4060 35084 4844 35140
rect 4900 35084 4910 35140
rect 11666 35084 11676 35140
rect 11732 35084 15820 35140
rect 15876 35084 15886 35140
rect 16342 35084 16380 35140
rect 16436 35084 16446 35140
rect 19142 35084 19180 35140
rect 19236 35084 19246 35140
rect 23762 35084 23772 35140
rect 23828 35084 25004 35140
rect 25060 35084 25900 35140
rect 25956 35084 25966 35140
rect 2930 34972 2940 35028
rect 2996 34972 7084 35028
rect 7140 34972 7150 35028
rect 8642 34972 8652 35028
rect 8708 34972 10780 35028
rect 10836 34972 10846 35028
rect 12674 34972 12684 35028
rect 12740 34972 13692 35028
rect 13748 34972 14924 35028
rect 14980 34972 14990 35028
rect 19702 34972 19740 35028
rect 19796 34972 19806 35028
rect 19964 34972 20300 35028
rect 20356 34972 20366 35028
rect 23986 34972 23996 35028
rect 24052 34972 26236 35028
rect 26292 34972 26684 35028
rect 26740 34972 26750 35028
rect 14924 34916 14980 34972
rect 19964 34916 20020 34972
rect 3490 34860 3500 34916
rect 3556 34860 4620 34916
rect 4676 34860 10108 34916
rect 10164 34860 10174 34916
rect 10406 34860 10444 34916
rect 10500 34860 10510 34916
rect 11330 34860 11340 34916
rect 11396 34860 12348 34916
rect 12404 34860 12414 34916
rect 13906 34860 13916 34916
rect 13972 34860 14700 34916
rect 14756 34860 14766 34916
rect 14924 34860 15596 34916
rect 15652 34860 15662 34916
rect 17938 34860 17948 34916
rect 18004 34860 18956 34916
rect 19012 34860 20020 34916
rect 20178 34860 20188 34916
rect 20244 34860 22092 34916
rect 22148 34860 22158 34916
rect 22754 34860 22764 34916
rect 22820 34860 26460 34916
rect 26516 34860 27356 34916
rect 27412 34860 27422 34916
rect 7746 34748 7756 34804
rect 7812 34748 8652 34804
rect 8708 34748 8988 34804
rect 9044 34748 9054 34804
rect 9762 34748 9772 34804
rect 9828 34748 11788 34804
rect 11844 34748 11854 34804
rect 12012 34748 17612 34804
rect 17668 34748 18172 34804
rect 18228 34748 18238 34804
rect 20626 34748 20636 34804
rect 20692 34748 21868 34804
rect 21924 34748 21934 34804
rect 24098 34748 24108 34804
rect 24164 34748 24668 34804
rect 24724 34748 25340 34804
rect 25396 34748 25406 34804
rect 26562 34748 26572 34804
rect 26628 34748 28028 34804
rect 28084 34748 28094 34804
rect 12012 34692 12068 34748
rect 3602 34636 3612 34692
rect 3668 34636 12068 34692
rect 18610 34636 18620 34692
rect 18676 34636 19852 34692
rect 19908 34636 20188 34692
rect 20244 34636 20254 34692
rect 20738 34636 20748 34692
rect 20804 34636 22092 34692
rect 22148 34636 22158 34692
rect 24658 34636 24668 34692
rect 24724 34636 25116 34692
rect 25172 34636 25182 34692
rect 25890 34636 25900 34692
rect 25956 34636 27132 34692
rect 27188 34636 27804 34692
rect 27860 34636 27870 34692
rect 10098 34524 10108 34580
rect 10164 34524 10668 34580
rect 10724 34524 10734 34580
rect 19730 34524 19740 34580
rect 19796 34524 19964 34580
rect 20020 34524 20030 34580
rect 22166 34524 22204 34580
rect 22260 34524 22270 34580
rect 8006 34468 8016 34524
rect 8072 34468 8120 34524
rect 8176 34468 8224 34524
rect 8280 34468 8290 34524
rect 14810 34468 14820 34524
rect 14876 34468 14924 34524
rect 14980 34468 15028 34524
rect 15084 34468 15094 34524
rect 21614 34468 21624 34524
rect 21680 34468 21728 34524
rect 21784 34468 21832 34524
rect 21888 34468 21898 34524
rect 28418 34468 28428 34524
rect 28484 34468 28532 34524
rect 28588 34468 28636 34524
rect 28692 34468 28702 34524
rect 9090 34412 9100 34468
rect 9156 34412 12404 34468
rect 21970 34412 21980 34468
rect 22036 34412 23324 34468
rect 23380 34412 23390 34468
rect 25442 34412 25452 34468
rect 25508 34412 26124 34468
rect 26180 34412 26190 34468
rect 26852 34412 27692 34468
rect 27748 34412 28140 34468
rect 28196 34412 28206 34468
rect 0 34356 400 34384
rect 12348 34356 12404 34412
rect 0 34300 1708 34356
rect 1764 34300 1774 34356
rect 3826 34300 3836 34356
rect 3892 34300 7196 34356
rect 7252 34300 7262 34356
rect 8418 34300 8428 34356
rect 8484 34300 8494 34356
rect 11106 34300 11116 34356
rect 11172 34300 11228 34356
rect 11284 34300 11294 34356
rect 11778 34300 11788 34356
rect 11844 34300 12124 34356
rect 12180 34300 12190 34356
rect 12348 34300 19068 34356
rect 19124 34300 20076 34356
rect 20132 34300 20142 34356
rect 20738 34300 20748 34356
rect 20804 34300 21196 34356
rect 21252 34300 21262 34356
rect 21746 34300 21756 34356
rect 21812 34300 22540 34356
rect 22596 34300 22606 34356
rect 25666 34300 25676 34356
rect 25732 34300 26348 34356
rect 26404 34300 26414 34356
rect 0 34272 400 34300
rect 7196 34132 7252 34300
rect 8428 34132 8484 34300
rect 11788 34132 11844 34300
rect 20748 34132 20804 34300
rect 26852 34244 26908 34412
rect 21970 34188 21980 34244
rect 22036 34188 24220 34244
rect 24276 34188 26908 34244
rect 7196 34076 7868 34132
rect 7924 34076 7934 34132
rect 8082 34076 8092 34132
rect 8148 34076 9100 34132
rect 9156 34076 9772 34132
rect 9828 34076 9838 34132
rect 11106 34076 11116 34132
rect 11172 34076 11844 34132
rect 19842 34076 19852 34132
rect 19908 34076 20804 34132
rect 23426 34076 23436 34132
rect 23492 34076 25900 34132
rect 25956 34076 25966 34132
rect 7522 33964 7532 34020
rect 7588 33964 8316 34020
rect 8372 33964 8382 34020
rect 9986 33964 9996 34020
rect 10052 33964 12460 34020
rect 12516 33964 12526 34020
rect 14130 33964 14140 34020
rect 14196 33964 15372 34020
rect 15428 33964 18060 34020
rect 18116 33964 18126 34020
rect 23650 33964 23660 34020
rect 23716 33964 25676 34020
rect 25732 33964 25742 34020
rect 8418 33852 8428 33908
rect 8484 33852 8988 33908
rect 9044 33852 10108 33908
rect 10164 33852 10174 33908
rect 10322 33852 10332 33908
rect 10388 33852 10556 33908
rect 10612 33852 11228 33908
rect 11284 33852 11294 33908
rect 12338 33852 12348 33908
rect 12404 33852 12796 33908
rect 12852 33852 22428 33908
rect 22484 33852 22494 33908
rect 26450 33852 26460 33908
rect 26516 33852 27020 33908
rect 27076 33852 27086 33908
rect 6514 33740 6524 33796
rect 6580 33740 8652 33796
rect 8708 33740 9548 33796
rect 9604 33740 9614 33796
rect 19618 33740 19628 33796
rect 19684 33740 20524 33796
rect 20580 33740 20590 33796
rect 4604 33684 4614 33740
rect 4670 33684 4718 33740
rect 4774 33684 4822 33740
rect 4878 33684 4888 33740
rect 11408 33684 11418 33740
rect 11474 33684 11522 33740
rect 11578 33684 11626 33740
rect 11682 33684 11692 33740
rect 18212 33684 18222 33740
rect 18278 33684 18326 33740
rect 18382 33684 18430 33740
rect 18486 33684 18496 33740
rect 25016 33684 25026 33740
rect 25082 33684 25130 33740
rect 25186 33684 25234 33740
rect 25290 33684 25300 33740
rect 5954 33628 5964 33684
rect 6020 33628 6030 33684
rect 7074 33628 7084 33684
rect 7140 33628 7756 33684
rect 7812 33628 7822 33684
rect 8502 33628 8540 33684
rect 8596 33628 8606 33684
rect 17042 33628 17052 33684
rect 17108 33628 17612 33684
rect 17668 33628 17678 33684
rect 19954 33628 19964 33684
rect 20020 33628 20636 33684
rect 20692 33628 20702 33684
rect 23286 33628 23324 33684
rect 23380 33628 23390 33684
rect 23622 33628 23660 33684
rect 23716 33628 23726 33684
rect 2370 33516 2380 33572
rect 2436 33516 3388 33572
rect 3444 33516 5180 33572
rect 5236 33516 5246 33572
rect 2594 33404 2604 33460
rect 2660 33404 3500 33460
rect 3556 33404 3566 33460
rect 2034 33292 2044 33348
rect 2100 33292 2716 33348
rect 2772 33292 3388 33348
rect 3444 33292 3454 33348
rect 4396 33124 4452 33516
rect 5964 33460 6020 33628
rect 10546 33516 10556 33572
rect 10612 33516 10668 33572
rect 10724 33516 10734 33572
rect 12002 33516 12012 33572
rect 12068 33516 13244 33572
rect 13300 33516 13310 33572
rect 16594 33516 16604 33572
rect 16660 33516 16940 33572
rect 16996 33516 18060 33572
rect 18116 33516 18126 33572
rect 20178 33516 20188 33572
rect 20244 33516 25340 33572
rect 25396 33516 25406 33572
rect 4834 33404 4844 33460
rect 4900 33404 6020 33460
rect 6738 33404 6748 33460
rect 6804 33404 6814 33460
rect 8194 33404 8204 33460
rect 8260 33404 21364 33460
rect 22306 33404 22316 33460
rect 22372 33404 23324 33460
rect 23380 33404 23390 33460
rect 24406 33404 24444 33460
rect 24500 33404 24510 33460
rect 26674 33404 26684 33460
rect 26740 33404 27356 33460
rect 27412 33404 27422 33460
rect 6748 33348 6804 33404
rect 21308 33348 21364 33404
rect 5142 33292 5180 33348
rect 5236 33292 5246 33348
rect 5394 33292 5404 33348
rect 5460 33292 6804 33348
rect 10434 33292 10444 33348
rect 10500 33292 10556 33348
rect 10612 33292 10622 33348
rect 11106 33292 11116 33348
rect 11172 33292 12012 33348
rect 12068 33292 12078 33348
rect 14578 33292 14588 33348
rect 14644 33292 15932 33348
rect 15988 33292 15998 33348
rect 20178 33292 20188 33348
rect 20244 33292 20748 33348
rect 20804 33292 20814 33348
rect 21298 33292 21308 33348
rect 21364 33292 21374 33348
rect 22418 33292 22428 33348
rect 22484 33292 25228 33348
rect 25284 33292 27020 33348
rect 27076 33292 27086 33348
rect 9874 33180 9884 33236
rect 9940 33180 10556 33236
rect 10612 33180 10622 33236
rect 12674 33180 12684 33236
rect 12740 33180 14364 33236
rect 14420 33180 14812 33236
rect 14868 33180 15596 33236
rect 15652 33180 15662 33236
rect 19058 33180 19068 33236
rect 19124 33180 22316 33236
rect 22372 33180 22382 33236
rect 22642 33180 22652 33236
rect 22708 33180 23940 33236
rect 23884 33124 23940 33180
rect 4386 33068 4396 33124
rect 4452 33068 4462 33124
rect 11330 33068 11340 33124
rect 11396 33068 16044 33124
rect 16100 33068 16110 33124
rect 19954 33068 19964 33124
rect 20020 33068 20188 33124
rect 20244 33068 20254 33124
rect 21410 33068 21420 33124
rect 21476 33068 22540 33124
rect 22596 33068 22606 33124
rect 22866 33068 22876 33124
rect 22932 33068 23660 33124
rect 23716 33068 23726 33124
rect 23884 33068 24444 33124
rect 24500 33068 24510 33124
rect 12338 32956 12348 33012
rect 12404 32956 13468 33012
rect 13524 32956 13534 33012
rect 19954 32956 19964 33012
rect 20020 32956 20748 33012
rect 20804 32956 20814 33012
rect 8006 32900 8016 32956
rect 8072 32900 8120 32956
rect 8176 32900 8224 32956
rect 8280 32900 8290 32956
rect 14810 32900 14820 32956
rect 14876 32900 14924 32956
rect 14980 32900 15028 32956
rect 15084 32900 15094 32956
rect 21614 32900 21624 32956
rect 21680 32900 21728 32956
rect 21784 32900 21832 32956
rect 21888 32900 21898 32956
rect 28418 32900 28428 32956
rect 28484 32900 28532 32956
rect 28588 32900 28636 32956
rect 28692 32900 28702 32956
rect 10854 32844 10892 32900
rect 10948 32844 10958 32900
rect 12002 32844 12012 32900
rect 12068 32844 12796 32900
rect 12852 32844 12862 32900
rect 23090 32844 23100 32900
rect 23156 32844 23436 32900
rect 23492 32844 23502 32900
rect 2594 32732 2604 32788
rect 2660 32732 3052 32788
rect 3108 32732 3724 32788
rect 3780 32732 3790 32788
rect 8754 32732 8764 32788
rect 8820 32732 9212 32788
rect 9268 32732 9278 32788
rect 10966 32732 11004 32788
rect 11060 32732 11070 32788
rect 11218 32732 11228 32788
rect 11284 32732 11452 32788
rect 11508 32732 11518 32788
rect 16566 32732 16604 32788
rect 16660 32732 16670 32788
rect 17462 32732 17500 32788
rect 17556 32732 17566 32788
rect 17714 32732 17724 32788
rect 17780 32732 17818 32788
rect 18498 32732 18508 32788
rect 18564 32732 18574 32788
rect 18834 32732 18844 32788
rect 18900 32732 19404 32788
rect 19460 32732 19470 32788
rect 25442 32732 25452 32788
rect 25508 32732 26348 32788
rect 26404 32732 26414 32788
rect 18508 32676 18564 32732
rect 6962 32620 6972 32676
rect 7028 32620 17388 32676
rect 17444 32620 23884 32676
rect 23940 32620 23950 32676
rect 25526 32620 25564 32676
rect 25620 32620 25630 32676
rect 18050 32508 18060 32564
rect 18116 32508 18844 32564
rect 18900 32508 19516 32564
rect 19572 32508 20300 32564
rect 20356 32508 20366 32564
rect 3938 32396 3948 32452
rect 4004 32396 4844 32452
rect 4900 32396 4910 32452
rect 6290 32396 6300 32452
rect 6356 32396 8764 32452
rect 8820 32396 8830 32452
rect 15138 32396 15148 32452
rect 15204 32396 15820 32452
rect 15876 32396 15886 32452
rect 16818 32396 16828 32452
rect 16884 32396 17500 32452
rect 17556 32396 17724 32452
rect 17780 32396 17790 32452
rect 18386 32396 18396 32452
rect 18452 32396 19964 32452
rect 20020 32396 20076 32452
rect 20132 32396 20972 32452
rect 21028 32396 21420 32452
rect 21476 32396 21486 32452
rect 23650 32396 23660 32452
rect 23716 32396 24668 32452
rect 24724 32396 24734 32452
rect 26114 32396 26124 32452
rect 26180 32396 26460 32452
rect 26516 32396 26526 32452
rect 26852 32396 27916 32452
rect 27972 32396 27982 32452
rect 26852 32340 26908 32396
rect 11228 32284 11676 32340
rect 11732 32284 11742 32340
rect 26674 32284 26684 32340
rect 26740 32284 26908 32340
rect 8754 32172 8764 32228
rect 8820 32172 9996 32228
rect 10052 32172 10062 32228
rect 4604 32116 4614 32172
rect 4670 32116 4718 32172
rect 4774 32116 4822 32172
rect 4878 32116 4888 32172
rect 11228 32116 11284 32284
rect 19058 32172 19068 32228
rect 19124 32172 24780 32228
rect 24836 32172 24846 32228
rect 11408 32116 11418 32172
rect 11474 32116 11522 32172
rect 11578 32116 11626 32172
rect 11682 32116 11692 32172
rect 18212 32116 18222 32172
rect 18278 32116 18326 32172
rect 18382 32116 18430 32172
rect 18486 32116 18496 32172
rect 25016 32116 25026 32172
rect 25082 32116 25130 32172
rect 25186 32116 25234 32172
rect 25290 32116 25300 32172
rect 6300 32060 10780 32116
rect 10836 32060 10846 32116
rect 11218 32060 11228 32116
rect 11284 32060 11294 32116
rect 12114 32060 12124 32116
rect 12180 32060 12908 32116
rect 12964 32060 12974 32116
rect 20486 32060 20524 32116
rect 20580 32060 20590 32116
rect 22978 32060 22988 32116
rect 23044 32060 23884 32116
rect 23940 32060 23950 32116
rect 26236 32060 26796 32116
rect 26852 32060 26862 32116
rect 6300 32004 6356 32060
rect 3378 31948 3388 32004
rect 3444 31948 4620 32004
rect 4676 31948 6356 32004
rect 9762 31948 9772 32004
rect 9828 31948 10668 32004
rect 10724 31948 10734 32004
rect 2146 31836 2156 31892
rect 2212 31836 4060 31892
rect 4116 31836 4126 31892
rect 9772 31836 10332 31892
rect 10388 31836 11228 31892
rect 11284 31836 11294 31892
rect 9772 31780 9828 31836
rect 2034 31724 2044 31780
rect 2100 31724 2828 31780
rect 2884 31724 4732 31780
rect 4788 31724 4798 31780
rect 9762 31724 9772 31780
rect 9828 31724 9838 31780
rect 10994 31724 11004 31780
rect 11060 31724 11564 31780
rect 11620 31724 11630 31780
rect 0 31668 400 31696
rect 11004 31668 11060 31724
rect 12124 31668 12180 32060
rect 26236 32004 26292 32060
rect 13458 31948 13468 32004
rect 13524 31948 18732 32004
rect 18788 31948 18798 32004
rect 20290 31948 20300 32004
rect 20356 31948 20412 32004
rect 20468 31948 20478 32004
rect 20626 31948 20636 32004
rect 20692 31948 20804 32004
rect 22306 31948 22316 32004
rect 22372 31948 22876 32004
rect 22932 31948 22942 32004
rect 26226 31948 26236 32004
rect 26292 31948 26302 32004
rect 20748 31892 20804 31948
rect 20748 31836 21084 31892
rect 21140 31836 21150 31892
rect 23314 31836 23324 31892
rect 23380 31836 23548 31892
rect 23604 31836 24220 31892
rect 24276 31836 24286 31892
rect 19058 31724 19068 31780
rect 19124 31724 19404 31780
rect 19460 31724 19470 31780
rect 20738 31724 20748 31780
rect 20804 31724 21308 31780
rect 21364 31724 21374 31780
rect 0 31612 1708 31668
rect 1764 31612 1774 31668
rect 7186 31612 7196 31668
rect 7252 31612 11060 31668
rect 12114 31612 12124 31668
rect 12180 31612 12190 31668
rect 12562 31612 12572 31668
rect 12628 31612 13468 31668
rect 13524 31612 13534 31668
rect 19506 31612 19516 31668
rect 19572 31612 21196 31668
rect 21252 31612 21262 31668
rect 23314 31612 23324 31668
rect 23380 31612 24668 31668
rect 24724 31612 25788 31668
rect 25844 31612 26124 31668
rect 26180 31612 26190 31668
rect 26674 31612 26684 31668
rect 26740 31612 27356 31668
rect 27412 31612 27422 31668
rect 0 31584 400 31612
rect 5170 31500 5180 31556
rect 5236 31500 5404 31556
rect 5460 31500 5470 31556
rect 10994 31500 11004 31556
rect 11060 31500 11340 31556
rect 11396 31500 11406 31556
rect 16034 31500 16044 31556
rect 16100 31500 20636 31556
rect 20692 31500 20702 31556
rect 20850 31500 20860 31556
rect 20916 31500 21532 31556
rect 21588 31500 21598 31556
rect 9874 31388 9884 31444
rect 9940 31388 10220 31444
rect 10276 31388 10286 31444
rect 16258 31388 16268 31444
rect 16324 31388 17500 31444
rect 17556 31388 17566 31444
rect 19730 31388 19740 31444
rect 19796 31388 20188 31444
rect 20244 31388 20254 31444
rect 8006 31332 8016 31388
rect 8072 31332 8120 31388
rect 8176 31332 8224 31388
rect 8280 31332 8290 31388
rect 14810 31332 14820 31388
rect 14876 31332 14924 31388
rect 14980 31332 15028 31388
rect 15084 31332 15094 31388
rect 21614 31332 21624 31388
rect 21680 31332 21728 31388
rect 21784 31332 21832 31388
rect 21888 31332 21898 31388
rect 28418 31332 28428 31388
rect 28484 31332 28532 31388
rect 28588 31332 28636 31388
rect 28692 31332 28702 31388
rect 5058 31276 5068 31332
rect 5124 31276 5852 31332
rect 5908 31276 5918 31332
rect 7606 31276 7644 31332
rect 7700 31276 7710 31332
rect 19170 31276 19180 31332
rect 19236 31276 19852 31332
rect 19908 31276 19918 31332
rect 4162 31164 4172 31220
rect 4228 31164 6300 31220
rect 6356 31164 7196 31220
rect 7252 31164 7262 31220
rect 14578 31164 14588 31220
rect 14644 31164 14812 31220
rect 14868 31164 14878 31220
rect 15474 31164 15484 31220
rect 15540 31164 16492 31220
rect 16548 31164 16558 31220
rect 17266 31164 17276 31220
rect 17332 31164 19516 31220
rect 19572 31164 19582 31220
rect 21634 31164 21644 31220
rect 21700 31164 21980 31220
rect 22036 31164 22046 31220
rect 24098 31164 24108 31220
rect 24164 31164 24892 31220
rect 24948 31164 24958 31220
rect 7634 31052 7644 31108
rect 7700 31052 7980 31108
rect 8036 31052 8046 31108
rect 14588 31052 15372 31108
rect 15428 31052 15438 31108
rect 17378 31052 17388 31108
rect 17444 31052 18172 31108
rect 18228 31052 18238 31108
rect 18946 31052 18956 31108
rect 19012 31052 19740 31108
rect 19796 31052 19806 31108
rect 21186 31052 21196 31108
rect 21252 31052 24332 31108
rect 24388 31052 24398 31108
rect 26086 31052 26124 31108
rect 26180 31052 26190 31108
rect 14588 30996 14644 31052
rect 5618 30940 5628 30996
rect 5684 30940 7532 30996
rect 7588 30940 7598 30996
rect 8418 30940 8428 30996
rect 8484 30940 9100 30996
rect 9156 30940 9548 30996
rect 9604 30940 9614 30996
rect 12898 30940 12908 30996
rect 12964 30940 14140 30996
rect 14196 30940 14588 30996
rect 14644 30940 14654 30996
rect 16930 30940 16940 30996
rect 16996 30940 17836 30996
rect 17892 30940 17902 30996
rect 18610 30940 18620 30996
rect 18676 30940 19068 30996
rect 19124 30940 19134 30996
rect 21074 30940 21084 30996
rect 21140 30940 21980 30996
rect 22036 30940 22046 30996
rect 25890 30940 25900 30996
rect 25956 30940 26908 30996
rect 5506 30828 5516 30884
rect 5572 30828 6412 30884
rect 6468 30828 6636 30884
rect 6692 30828 6702 30884
rect 7532 30660 7588 30940
rect 26852 30884 26908 30940
rect 8082 30828 8092 30884
rect 8148 30828 8876 30884
rect 8932 30828 8942 30884
rect 14242 30828 14252 30884
rect 14308 30828 16828 30884
rect 16884 30828 16894 30884
rect 23986 30828 23996 30884
rect 24052 30828 24668 30884
rect 24724 30828 25340 30884
rect 25396 30828 25788 30884
rect 25844 30828 25854 30884
rect 26852 30828 27580 30884
rect 27636 30828 27646 30884
rect 19618 30716 19628 30772
rect 19684 30716 23548 30772
rect 23604 30716 23614 30772
rect 7532 30604 7924 30660
rect 4604 30548 4614 30604
rect 4670 30548 4718 30604
rect 4774 30548 4822 30604
rect 4878 30548 4888 30604
rect 7868 30548 7924 30604
rect 11408 30548 11418 30604
rect 11474 30548 11522 30604
rect 11578 30548 11626 30604
rect 11682 30548 11692 30604
rect 18212 30548 18222 30604
rect 18278 30548 18326 30604
rect 18382 30548 18430 30604
rect 18486 30548 18496 30604
rect 25016 30548 25026 30604
rect 25082 30548 25130 30604
rect 25186 30548 25234 30604
rect 25290 30548 25300 30604
rect 7858 30492 7868 30548
rect 7924 30492 7934 30548
rect 4722 30380 4732 30436
rect 4788 30380 8092 30436
rect 8148 30380 8158 30436
rect 8418 30380 8428 30436
rect 8484 30380 8494 30436
rect 21382 30380 21420 30436
rect 21476 30380 21486 30436
rect 8428 30324 8484 30380
rect 5170 30268 5180 30324
rect 5236 30268 5852 30324
rect 5908 30268 5918 30324
rect 6738 30268 6748 30324
rect 6804 30268 7308 30324
rect 7364 30268 7374 30324
rect 7634 30268 7644 30324
rect 7700 30268 8484 30324
rect 9538 30268 9548 30324
rect 9604 30268 10556 30324
rect 10612 30268 11452 30324
rect 11508 30268 11518 30324
rect 12562 30268 12572 30324
rect 12628 30268 14252 30324
rect 14308 30268 14318 30324
rect 15372 30268 15708 30324
rect 15764 30268 15774 30324
rect 17602 30268 17612 30324
rect 17668 30268 18396 30324
rect 18452 30268 18462 30324
rect 15372 30212 15428 30268
rect 3938 30156 3948 30212
rect 4004 30156 4014 30212
rect 5058 30156 5068 30212
rect 5124 30156 5740 30212
rect 5796 30156 10332 30212
rect 10388 30156 10398 30212
rect 10658 30156 10668 30212
rect 10724 30156 12012 30212
rect 12068 30156 12796 30212
rect 12852 30156 12862 30212
rect 14476 30156 15428 30212
rect 15586 30156 15596 30212
rect 15652 30156 16380 30212
rect 16436 30156 19852 30212
rect 19908 30156 19918 30212
rect 20178 30156 20188 30212
rect 20244 30156 20748 30212
rect 20804 30156 20814 30212
rect 23650 30156 23660 30212
rect 23716 30156 26236 30212
rect 26292 30156 26302 30212
rect 3948 30100 4004 30156
rect 3948 30044 6188 30100
rect 6244 30044 6254 30100
rect 8978 30044 8988 30100
rect 9044 30044 9324 30100
rect 9380 30044 9390 30100
rect 9874 30044 9884 30100
rect 9940 30044 10444 30100
rect 10500 30044 10892 30100
rect 10948 30044 11900 30100
rect 11956 30044 11966 30100
rect 3948 29988 4004 30044
rect 14476 29988 14532 30156
rect 15362 30044 15372 30100
rect 15428 30044 16716 30100
rect 16772 30044 20300 30100
rect 20356 30044 23996 30100
rect 24052 30044 24062 30100
rect 24658 30044 24668 30100
rect 24724 30044 27132 30100
rect 27188 30044 27916 30100
rect 27972 30044 27982 30100
rect 3602 29932 3612 29988
rect 3668 29932 4004 29988
rect 4386 29932 4396 29988
rect 4452 29932 5180 29988
rect 5236 29932 5516 29988
rect 5572 29932 5582 29988
rect 8306 29932 8316 29988
rect 8372 29932 9660 29988
rect 9716 29932 9726 29988
rect 10210 29932 10220 29988
rect 10276 29932 10780 29988
rect 10836 29932 10846 29988
rect 12674 29932 12684 29988
rect 12740 29932 12908 29988
rect 12964 29932 14532 29988
rect 14914 29932 14924 29988
rect 14980 29932 15260 29988
rect 15316 29932 17388 29988
rect 17444 29932 19292 29988
rect 19348 29932 20188 29988
rect 20244 29932 20254 29988
rect 21858 29932 21868 29988
rect 21924 29932 23660 29988
rect 23716 29932 23726 29988
rect 3938 29820 3948 29876
rect 4004 29820 4732 29876
rect 4788 29820 4798 29876
rect 6850 29820 6860 29876
rect 6916 29820 7196 29876
rect 7252 29820 7262 29876
rect 8530 29820 8540 29876
rect 8596 29820 8988 29876
rect 9044 29820 9054 29876
rect 20738 29820 20748 29876
rect 20804 29820 21420 29876
rect 21476 29820 21486 29876
rect 22530 29820 22540 29876
rect 22596 29820 22988 29876
rect 23044 29820 23054 29876
rect 24770 29820 24780 29876
rect 24836 29820 25340 29876
rect 25396 29820 25406 29876
rect 8006 29764 8016 29820
rect 8072 29764 8120 29820
rect 8176 29764 8224 29820
rect 8280 29764 8290 29820
rect 14810 29764 14820 29820
rect 14876 29764 14924 29820
rect 14980 29764 15028 29820
rect 15084 29764 15094 29820
rect 21614 29764 21624 29820
rect 21680 29764 21728 29820
rect 21784 29764 21832 29820
rect 21888 29764 21898 29820
rect 28418 29764 28428 29820
rect 28484 29764 28532 29820
rect 28588 29764 28636 29820
rect 28692 29764 28702 29820
rect 19282 29708 19292 29764
rect 19348 29708 19628 29764
rect 19684 29708 19694 29764
rect 7084 29596 11788 29652
rect 12338 29596 12348 29652
rect 12404 29596 14588 29652
rect 14644 29596 14654 29652
rect 14802 29596 14812 29652
rect 14868 29596 21868 29652
rect 21924 29596 21934 29652
rect 22530 29596 22540 29652
rect 22596 29596 23212 29652
rect 23268 29596 23278 29652
rect 7084 29540 7140 29596
rect 11732 29540 11788 29596
rect 3602 29484 3612 29540
rect 3668 29484 5628 29540
rect 5684 29484 5694 29540
rect 7074 29484 7084 29540
rect 7140 29484 7150 29540
rect 10546 29484 10556 29540
rect 10612 29484 11172 29540
rect 11732 29484 22316 29540
rect 22372 29484 22382 29540
rect 11116 29428 11172 29484
rect 4274 29372 4284 29428
rect 4340 29372 10892 29428
rect 10948 29372 10958 29428
rect 11116 29372 19852 29428
rect 19908 29372 19918 29428
rect 20290 29372 20300 29428
rect 20356 29372 21308 29428
rect 21364 29372 21374 29428
rect 2482 29260 2492 29316
rect 2548 29260 3164 29316
rect 3220 29260 3230 29316
rect 9650 29260 9660 29316
rect 9716 29260 14812 29316
rect 14868 29260 14878 29316
rect 17826 29260 17836 29316
rect 17892 29260 19292 29316
rect 19348 29260 19358 29316
rect 23874 29260 23884 29316
rect 23940 29260 24556 29316
rect 24612 29260 24622 29316
rect 24770 29260 24780 29316
rect 24836 29260 25228 29316
rect 25284 29260 25294 29316
rect 11106 29148 11116 29204
rect 11172 29148 12012 29204
rect 12068 29148 12078 29204
rect 15138 29148 15148 29204
rect 15204 29148 15596 29204
rect 15652 29148 15662 29204
rect 18498 29148 18508 29204
rect 18564 29148 19348 29204
rect 19292 29092 19348 29148
rect 8502 29036 8540 29092
rect 8596 29036 8606 29092
rect 13346 29036 13356 29092
rect 13412 29036 14028 29092
rect 14084 29036 14094 29092
rect 19282 29036 19292 29092
rect 19348 29036 19358 29092
rect 0 28980 400 29008
rect 4604 28980 4614 29036
rect 4670 28980 4718 29036
rect 4774 28980 4822 29036
rect 4878 28980 4888 29036
rect 11408 28980 11418 29036
rect 11474 28980 11522 29036
rect 11578 28980 11626 29036
rect 11682 28980 11692 29036
rect 18212 28980 18222 29036
rect 18278 28980 18326 29036
rect 18382 28980 18430 29036
rect 18486 28980 18496 29036
rect 25016 28980 25026 29036
rect 25082 28980 25130 29036
rect 25186 28980 25234 29036
rect 25290 28980 25300 29036
rect 0 28924 1708 28980
rect 1764 28924 1774 28980
rect 12460 28924 14252 28980
rect 14308 28924 14318 28980
rect 0 28896 400 28924
rect 12460 28868 12516 28924
rect 5170 28812 5180 28868
rect 5236 28812 12460 28868
rect 12516 28812 12526 28868
rect 14130 28812 14140 28868
rect 14196 28812 15036 28868
rect 15092 28812 15102 28868
rect 24434 28812 24444 28868
rect 24500 28812 25564 28868
rect 25620 28812 25630 28868
rect 2706 28700 2716 28756
rect 2772 28700 3500 28756
rect 3556 28700 3566 28756
rect 4274 28700 4284 28756
rect 4340 28700 4620 28756
rect 4676 28700 4686 28756
rect 6850 28700 6860 28756
rect 6916 28700 7756 28756
rect 7812 28700 7822 28756
rect 10434 28700 10444 28756
rect 10500 28700 10556 28756
rect 10612 28700 11116 28756
rect 11172 28700 11182 28756
rect 11778 28700 11788 28756
rect 11844 28700 12908 28756
rect 12964 28700 13356 28756
rect 13412 28700 13422 28756
rect 13906 28700 13916 28756
rect 13972 28700 14812 28756
rect 14868 28700 15148 28756
rect 15250 28700 15260 28756
rect 15316 28700 15708 28756
rect 15764 28700 15774 28756
rect 18386 28700 18396 28756
rect 18452 28700 18844 28756
rect 18900 28700 18910 28756
rect 25330 28700 25340 28756
rect 25396 28700 27356 28756
rect 27412 28700 27422 28756
rect 15092 28644 15148 28700
rect 1698 28588 1708 28644
rect 1764 28588 2604 28644
rect 2660 28588 2670 28644
rect 2930 28588 2940 28644
rect 2996 28588 4172 28644
rect 4228 28588 4238 28644
rect 14130 28588 14140 28644
rect 14196 28588 14924 28644
rect 14980 28588 14990 28644
rect 15092 28588 16044 28644
rect 16100 28588 19068 28644
rect 19124 28588 19134 28644
rect 22978 28588 22988 28644
rect 23044 28588 24780 28644
rect 24836 28588 25004 28644
rect 25060 28588 25070 28644
rect 25666 28588 25676 28644
rect 25732 28588 26460 28644
rect 26516 28588 26526 28644
rect 4274 28476 4284 28532
rect 4340 28476 5068 28532
rect 5124 28476 5134 28532
rect 13654 28476 13692 28532
rect 13748 28476 15708 28532
rect 15764 28476 15774 28532
rect 20514 28476 20524 28532
rect 20580 28476 23548 28532
rect 23604 28476 23614 28532
rect 24770 28476 24780 28532
rect 24836 28476 26348 28532
rect 26404 28476 26414 28532
rect 13346 28364 13356 28420
rect 13412 28364 17836 28420
rect 17892 28364 17902 28420
rect 20514 28364 20524 28420
rect 20580 28364 21980 28420
rect 22036 28364 22540 28420
rect 22596 28364 22606 28420
rect 25750 28364 25788 28420
rect 25844 28364 26236 28420
rect 26292 28364 26302 28420
rect 25554 28252 25564 28308
rect 25620 28252 26124 28308
rect 26180 28252 26190 28308
rect 26646 28252 26684 28308
rect 26740 28252 26750 28308
rect 8006 28196 8016 28252
rect 8072 28196 8120 28252
rect 8176 28196 8224 28252
rect 8280 28196 8290 28252
rect 14810 28196 14820 28252
rect 14876 28196 14924 28252
rect 14980 28196 15028 28252
rect 15084 28196 15094 28252
rect 21614 28196 21624 28252
rect 21680 28196 21728 28252
rect 21784 28196 21832 28252
rect 21888 28196 21898 28252
rect 28418 28196 28428 28252
rect 28484 28196 28532 28252
rect 28588 28196 28636 28252
rect 28692 28196 28702 28252
rect 9874 28140 9884 28196
rect 9940 28140 10332 28196
rect 10388 28140 10398 28196
rect 10770 28140 10780 28196
rect 10836 28140 10846 28196
rect 12562 28140 12572 28196
rect 12628 28140 12740 28196
rect 14242 28140 14252 28196
rect 14308 28140 14588 28196
rect 14644 28140 14654 28196
rect 23538 28140 23548 28196
rect 23604 28140 23772 28196
rect 23828 28140 23838 28196
rect 26562 28140 26572 28196
rect 26628 28140 27804 28196
rect 27860 28140 27870 28196
rect 10780 28084 10836 28140
rect 12684 28084 12740 28140
rect 1810 28028 1820 28084
rect 1876 28028 2940 28084
rect 2996 28028 5068 28084
rect 5124 28028 5964 28084
rect 6020 28028 6030 28084
rect 9996 28028 10836 28084
rect 11554 28028 11564 28084
rect 11620 28028 12460 28084
rect 12516 28028 12526 28084
rect 12684 28028 15260 28084
rect 15316 28028 15326 28084
rect 16716 28028 17052 28084
rect 17108 28028 17836 28084
rect 17892 28028 17902 28084
rect 22082 28028 22092 28084
rect 22148 28028 22988 28084
rect 23044 28028 23054 28084
rect 9996 27860 10052 28028
rect 16716 27972 16772 28028
rect 10210 27916 10220 27972
rect 10276 27916 10780 27972
rect 10836 27916 16772 27972
rect 16930 27916 16940 27972
rect 16996 27916 19628 27972
rect 19684 27916 19694 27972
rect 25890 27916 25900 27972
rect 25956 27916 27804 27972
rect 27860 27916 27870 27972
rect 2146 27804 2156 27860
rect 2212 27804 5852 27860
rect 5908 27804 5918 27860
rect 8082 27804 8092 27860
rect 8148 27804 8988 27860
rect 9044 27804 13692 27860
rect 13748 27804 14028 27860
rect 14084 27804 14094 27860
rect 14914 27804 14924 27860
rect 14980 27804 16380 27860
rect 16436 27804 16446 27860
rect 23538 27804 23548 27860
rect 23604 27804 24276 27860
rect 26450 27804 26460 27860
rect 26516 27804 26684 27860
rect 26740 27804 26750 27860
rect 8866 27692 8876 27748
rect 8932 27692 9660 27748
rect 9716 27692 15036 27748
rect 15092 27692 15102 27748
rect 15250 27692 15260 27748
rect 15316 27692 16156 27748
rect 16212 27692 19292 27748
rect 19348 27692 19358 27748
rect 9202 27580 9212 27636
rect 9268 27580 11004 27636
rect 11060 27580 11340 27636
rect 11396 27580 12180 27636
rect 12338 27580 12348 27636
rect 12404 27580 17388 27636
rect 17444 27580 18844 27636
rect 18900 27580 18910 27636
rect 12124 27524 12180 27580
rect 24220 27524 24276 27804
rect 26338 27580 26348 27636
rect 26404 27580 27020 27636
rect 27076 27580 27086 27636
rect 12124 27468 12796 27524
rect 12852 27468 13356 27524
rect 13412 27468 13422 27524
rect 13682 27468 13692 27524
rect 13748 27468 14364 27524
rect 14420 27468 14430 27524
rect 17686 27468 17724 27524
rect 17780 27468 17790 27524
rect 20738 27468 20748 27524
rect 20804 27468 21196 27524
rect 21252 27468 21262 27524
rect 24210 27468 24220 27524
rect 24276 27468 24286 27524
rect 4604 27412 4614 27468
rect 4670 27412 4718 27468
rect 4774 27412 4822 27468
rect 4878 27412 4888 27468
rect 11408 27412 11418 27468
rect 11474 27412 11522 27468
rect 11578 27412 11626 27468
rect 11682 27412 11692 27468
rect 18212 27412 18222 27468
rect 18278 27412 18326 27468
rect 18382 27412 18430 27468
rect 18486 27412 18496 27468
rect 25016 27412 25026 27468
rect 25082 27412 25130 27468
rect 25186 27412 25234 27468
rect 25290 27412 25300 27468
rect 8530 27356 8540 27412
rect 8596 27356 9548 27412
rect 9604 27356 9614 27412
rect 10518 27356 10556 27412
rect 10612 27356 10622 27412
rect 13122 27356 13132 27412
rect 13188 27356 15596 27412
rect 15652 27356 15662 27412
rect 19954 27356 19964 27412
rect 20020 27356 20076 27412
rect 20132 27356 20142 27412
rect 20514 27356 20524 27412
rect 20580 27356 21308 27412
rect 21364 27356 21374 27412
rect 26086 27356 26124 27412
rect 26180 27356 26190 27412
rect 6850 27244 6860 27300
rect 6916 27244 7644 27300
rect 7700 27244 9212 27300
rect 9268 27244 9278 27300
rect 20738 27244 20748 27300
rect 20804 27244 20972 27300
rect 21028 27244 21038 27300
rect 23090 27244 23100 27300
rect 23156 27244 25228 27300
rect 25284 27244 27020 27300
rect 27076 27244 27086 27300
rect 2818 27132 2828 27188
rect 2884 27132 3612 27188
rect 3668 27132 3836 27188
rect 3892 27132 5068 27188
rect 5124 27132 5628 27188
rect 5684 27132 5694 27188
rect 6402 27132 6412 27188
rect 6468 27132 7308 27188
rect 7364 27132 7374 27188
rect 7746 27132 7756 27188
rect 7812 27132 8316 27188
rect 8372 27132 9772 27188
rect 9828 27132 9838 27188
rect 15092 27132 16716 27188
rect 16772 27132 16782 27188
rect 16940 27132 18172 27188
rect 18228 27132 19068 27188
rect 19124 27132 24444 27188
rect 24500 27132 26460 27188
rect 26516 27132 26526 27188
rect 26674 27132 26684 27188
rect 26740 27132 27356 27188
rect 27412 27132 27422 27188
rect 15092 27076 15148 27132
rect 16940 27076 16996 27132
rect 5842 27020 5852 27076
rect 5908 27020 6748 27076
rect 6804 27020 6814 27076
rect 9650 27020 9660 27076
rect 9716 27020 12908 27076
rect 12964 27020 13580 27076
rect 13636 27020 15148 27076
rect 15250 27020 15260 27076
rect 15316 27020 16996 27076
rect 17378 27020 17388 27076
rect 17444 27020 18620 27076
rect 18676 27020 18686 27076
rect 19254 27020 19292 27076
rect 19348 27020 19358 27076
rect 19506 27020 19516 27076
rect 19572 27020 20076 27076
rect 20132 27020 20412 27076
rect 20468 27020 20478 27076
rect 20738 27020 20748 27076
rect 20804 27020 21308 27076
rect 21364 27020 21374 27076
rect 23202 27020 23212 27076
rect 23268 27020 23660 27076
rect 23716 27020 23726 27076
rect 25330 27020 25340 27076
rect 25396 27020 26236 27076
rect 26292 27020 27244 27076
rect 27300 27020 27310 27076
rect 13692 26852 13748 27020
rect 18274 26908 18284 26964
rect 18340 26908 24556 26964
rect 24612 26908 24622 26964
rect 1698 26796 1708 26852
rect 1764 26796 2940 26852
rect 2996 26796 3006 26852
rect 13682 26796 13692 26852
rect 13748 26796 13758 26852
rect 14130 26796 14140 26852
rect 14196 26796 16380 26852
rect 16436 26796 18172 26852
rect 18228 26796 18238 26852
rect 20374 26796 20412 26852
rect 20468 26796 20478 26852
rect 20636 26796 22652 26852
rect 22708 26796 22718 26852
rect 24882 26796 24892 26852
rect 24948 26796 25900 26852
rect 25956 26796 25966 26852
rect 20636 26740 20692 26796
rect 19142 26684 19180 26740
rect 19236 26684 19246 26740
rect 20188 26684 20692 26740
rect 23090 26684 23100 26740
rect 23156 26684 23324 26740
rect 23380 26684 23390 26740
rect 8006 26628 8016 26684
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8280 26628 8290 26684
rect 14810 26628 14820 26684
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 15084 26628 15094 26684
rect 13356 26460 14364 26516
rect 14420 26460 14430 26516
rect 13356 26404 13412 26460
rect 1922 26348 1932 26404
rect 1988 26348 3388 26404
rect 3444 26348 4284 26404
rect 4340 26348 4350 26404
rect 6178 26348 6188 26404
rect 6244 26348 12460 26404
rect 12516 26348 13412 26404
rect 15698 26348 15708 26404
rect 15764 26348 17388 26404
rect 17444 26348 18620 26404
rect 18676 26348 19740 26404
rect 19796 26348 19806 26404
rect 19926 26348 19964 26404
rect 20020 26348 20030 26404
rect 0 26292 400 26320
rect 0 26236 1708 26292
rect 1764 26236 1774 26292
rect 4946 26236 4956 26292
rect 5012 26236 10780 26292
rect 10836 26236 11116 26292
rect 11172 26236 15372 26292
rect 15428 26236 15438 26292
rect 16492 26236 17780 26292
rect 19170 26236 19180 26292
rect 19236 26236 19628 26292
rect 19684 26236 19694 26292
rect 0 26208 400 26236
rect 16492 26180 16548 26236
rect 17724 26180 17780 26236
rect 20188 26180 20244 26684
rect 21614 26628 21624 26684
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21888 26628 21898 26684
rect 28418 26628 28428 26684
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28692 26628 28702 26684
rect 21298 26460 21308 26516
rect 21364 26460 22204 26516
rect 22260 26460 22270 26516
rect 22866 26460 22876 26516
rect 22932 26460 23660 26516
rect 23716 26460 23884 26516
rect 23940 26460 23950 26516
rect 27346 26460 27356 26516
rect 27412 26460 28140 26516
rect 28196 26460 28206 26516
rect 20626 26236 20636 26292
rect 20692 26236 21644 26292
rect 21700 26236 22652 26292
rect 22708 26236 22718 26292
rect 23538 26236 23548 26292
rect 23604 26236 24892 26292
rect 24948 26236 25452 26292
rect 25508 26236 25518 26292
rect 12114 26124 12124 26180
rect 12180 26124 13132 26180
rect 13188 26124 13198 26180
rect 14578 26124 14588 26180
rect 14644 26124 16548 26180
rect 16706 26124 16716 26180
rect 16772 26124 17500 26180
rect 17556 26124 17566 26180
rect 17724 26124 20244 26180
rect 22306 26124 22316 26180
rect 22372 26124 23212 26180
rect 23268 26124 23278 26180
rect 23492 26124 25900 26180
rect 25956 26124 25966 26180
rect 23492 26068 23548 26124
rect 9538 26012 9548 26068
rect 9604 26012 10332 26068
rect 10388 26012 10398 26068
rect 12674 26012 12684 26068
rect 12740 26012 12908 26068
rect 12964 26012 13356 26068
rect 13412 26012 15148 26068
rect 15204 26012 15214 26068
rect 17826 26012 17836 26068
rect 17892 26012 18508 26068
rect 18564 26012 18574 26068
rect 19170 26012 19180 26068
rect 19236 26012 19404 26068
rect 19460 26012 19470 26068
rect 20748 26012 21980 26068
rect 22036 26012 23548 26068
rect 20748 25956 20804 26012
rect 10770 25900 10780 25956
rect 10836 25900 10892 25956
rect 10948 25900 10958 25956
rect 18722 25900 18732 25956
rect 18788 25900 20748 25956
rect 20804 25900 20814 25956
rect 20962 25900 20972 25956
rect 21028 25900 21038 25956
rect 23510 25900 23548 25956
rect 23604 25900 23614 25956
rect 4604 25844 4614 25900
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4878 25844 4888 25900
rect 11408 25844 11418 25900
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11682 25844 11692 25900
rect 18212 25844 18222 25900
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18486 25844 18496 25900
rect 18834 25788 18844 25844
rect 18900 25788 19180 25844
rect 19236 25788 19292 25844
rect 19348 25788 19358 25844
rect 20290 25788 20300 25844
rect 20356 25788 20366 25844
rect 20300 25732 20356 25788
rect 20972 25732 21028 25900
rect 25016 25844 25026 25900
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25290 25844 25300 25900
rect 15362 25676 15372 25732
rect 15428 25676 21028 25732
rect 3266 25564 3276 25620
rect 3332 25564 5068 25620
rect 5124 25564 6412 25620
rect 6468 25564 6478 25620
rect 12786 25564 12796 25620
rect 12852 25564 13356 25620
rect 13412 25564 13804 25620
rect 13860 25564 13870 25620
rect 20962 25564 20972 25620
rect 21028 25564 22204 25620
rect 22260 25564 22270 25620
rect 2034 25452 2044 25508
rect 2100 25452 2716 25508
rect 2772 25452 3500 25508
rect 3556 25452 3566 25508
rect 4050 25452 4060 25508
rect 4116 25452 6636 25508
rect 6692 25452 14588 25508
rect 14644 25452 14654 25508
rect 19282 25452 19292 25508
rect 19348 25452 23100 25508
rect 23156 25452 23166 25508
rect 2258 25340 2268 25396
rect 2324 25340 4620 25396
rect 4676 25340 5740 25396
rect 5796 25340 5806 25396
rect 18582 25340 18620 25396
rect 18676 25340 18686 25396
rect 20738 25340 20748 25396
rect 20804 25340 21420 25396
rect 21476 25340 21486 25396
rect 22978 25340 22988 25396
rect 23044 25340 23772 25396
rect 23828 25340 23838 25396
rect 25666 25340 25676 25396
rect 25732 25340 27020 25396
rect 27076 25340 27086 25396
rect 7186 25228 7196 25284
rect 7252 25228 8988 25284
rect 9044 25228 9660 25284
rect 9716 25228 10444 25284
rect 10500 25228 10510 25284
rect 11890 25228 11900 25284
rect 11956 25228 12460 25284
rect 12516 25228 14364 25284
rect 14420 25228 14430 25284
rect 16034 25228 16044 25284
rect 16100 25228 19740 25284
rect 19796 25228 19806 25284
rect 21084 25228 22316 25284
rect 22372 25228 22382 25284
rect 21084 25172 21140 25228
rect 16930 25116 16940 25172
rect 16996 25116 19516 25172
rect 19572 25116 19582 25172
rect 21074 25116 21084 25172
rect 21140 25116 21150 25172
rect 23762 25116 23772 25172
rect 23828 25116 24444 25172
rect 24500 25116 24510 25172
rect 8006 25060 8016 25116
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8280 25060 8290 25116
rect 14810 25060 14820 25116
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 15084 25060 15094 25116
rect 21614 25060 21624 25116
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21888 25060 21898 25116
rect 28418 25060 28428 25116
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28692 25060 28702 25116
rect 24098 25004 24108 25060
rect 24164 25004 24444 25060
rect 24500 25004 24510 25060
rect 4498 24892 4508 24948
rect 4564 24892 4956 24948
rect 5012 24892 5740 24948
rect 5796 24892 6076 24948
rect 6132 24892 7756 24948
rect 7812 24892 7822 24948
rect 11750 24892 11788 24948
rect 11844 24892 11854 24948
rect 15698 24892 15708 24948
rect 15764 24892 16268 24948
rect 16324 24892 16334 24948
rect 18722 24892 18732 24948
rect 18788 24892 19068 24948
rect 19124 24892 19134 24948
rect 20178 24892 20188 24948
rect 20244 24892 20860 24948
rect 20916 24892 20926 24948
rect 21158 24892 21196 24948
rect 21252 24892 21262 24948
rect 25414 24892 25452 24948
rect 25508 24892 25518 24948
rect 3602 24780 3612 24836
rect 3668 24780 12348 24836
rect 12404 24780 12414 24836
rect 19590 24780 19628 24836
rect 19684 24780 19694 24836
rect 4060 24724 4116 24780
rect 2930 24668 2940 24724
rect 2996 24668 3500 24724
rect 3556 24668 3566 24724
rect 4050 24668 4060 24724
rect 4116 24668 4126 24724
rect 9090 24668 9100 24724
rect 9156 24668 9772 24724
rect 9828 24668 9838 24724
rect 20738 24668 20748 24724
rect 20804 24668 20972 24724
rect 21028 24668 21038 24724
rect 24220 24668 24780 24724
rect 24836 24668 25900 24724
rect 25956 24668 27356 24724
rect 27412 24668 27422 24724
rect 24220 24612 24276 24668
rect 15138 24556 15148 24612
rect 15204 24556 16268 24612
rect 16324 24556 16334 24612
rect 17042 24556 17052 24612
rect 17108 24556 18396 24612
rect 18452 24556 19852 24612
rect 19908 24556 19918 24612
rect 24210 24556 24220 24612
rect 24276 24556 24286 24612
rect 24658 24556 24668 24612
rect 24724 24556 25564 24612
rect 25620 24556 26124 24612
rect 26180 24556 26190 24612
rect 16268 24500 16324 24556
rect 16268 24444 17948 24500
rect 18004 24444 20076 24500
rect 20132 24444 20142 24500
rect 24220 24444 27244 24500
rect 27300 24444 27310 24500
rect 24220 24388 24276 24444
rect 9734 24332 9772 24388
rect 9828 24332 10444 24388
rect 10500 24332 10510 24388
rect 19618 24332 19628 24388
rect 19684 24332 19852 24388
rect 19908 24332 21420 24388
rect 21476 24332 21486 24388
rect 24210 24332 24220 24388
rect 24276 24332 24286 24388
rect 26226 24332 26236 24388
rect 26292 24332 26302 24388
rect 4604 24276 4614 24332
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4878 24276 4888 24332
rect 11408 24276 11418 24332
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11682 24276 11692 24332
rect 18212 24276 18222 24332
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18486 24276 18496 24332
rect 25016 24276 25026 24332
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25290 24276 25300 24332
rect 12786 24220 12796 24276
rect 12852 24220 13468 24276
rect 13524 24220 13534 24276
rect 18946 24220 18956 24276
rect 19012 24220 19740 24276
rect 19796 24220 19806 24276
rect 26236 24164 26292 24332
rect 26562 24220 26572 24276
rect 26628 24220 26684 24276
rect 26740 24220 26750 24276
rect 4050 24108 4060 24164
rect 4116 24108 4620 24164
rect 4676 24108 4686 24164
rect 10098 24108 10108 24164
rect 10164 24108 10780 24164
rect 10836 24108 13916 24164
rect 13972 24108 14476 24164
rect 14532 24108 15372 24164
rect 15428 24108 15438 24164
rect 16146 24108 16156 24164
rect 16212 24108 16940 24164
rect 16996 24108 17006 24164
rect 18498 24108 18508 24164
rect 18564 24108 18844 24164
rect 18900 24108 18910 24164
rect 24546 24108 24556 24164
rect 24612 24108 26292 24164
rect 10434 23996 10444 24052
rect 10500 23996 11564 24052
rect 11620 23996 11630 24052
rect 14018 23996 14028 24052
rect 14084 23996 19852 24052
rect 19908 23996 19918 24052
rect 20178 23996 20188 24052
rect 20244 23996 20636 24052
rect 20692 23996 20860 24052
rect 20916 23996 20926 24052
rect 25330 23996 25340 24052
rect 25396 23996 26236 24052
rect 26292 23996 26302 24052
rect 11218 23884 11228 23940
rect 11284 23884 12012 23940
rect 12068 23884 12078 23940
rect 16706 23884 16716 23940
rect 16772 23884 17612 23940
rect 17668 23884 20412 23940
rect 20468 23884 20478 23940
rect 24994 23884 25004 23940
rect 25060 23884 26348 23940
rect 26404 23884 26414 23940
rect 10658 23772 10668 23828
rect 10724 23772 11676 23828
rect 11732 23772 11742 23828
rect 12786 23772 12796 23828
rect 12852 23772 13692 23828
rect 13748 23772 13758 23828
rect 14802 23772 14812 23828
rect 14868 23772 15708 23828
rect 15764 23772 15774 23828
rect 16566 23772 16604 23828
rect 16660 23772 16670 23828
rect 17378 23772 17388 23828
rect 17444 23772 18060 23828
rect 18116 23772 18126 23828
rect 25442 23772 25452 23828
rect 25508 23772 26572 23828
rect 26628 23772 26638 23828
rect 9174 23660 9212 23716
rect 9268 23660 9278 23716
rect 11554 23660 11564 23716
rect 11620 23660 13020 23716
rect 13076 23660 13086 23716
rect 13234 23660 13244 23716
rect 13300 23660 17052 23716
rect 17108 23660 18844 23716
rect 18900 23660 19292 23716
rect 19348 23660 20076 23716
rect 20132 23660 21196 23716
rect 21252 23660 22764 23716
rect 22820 23660 22830 23716
rect 23426 23660 23436 23716
rect 23492 23660 23996 23716
rect 24052 23660 24062 23716
rect 24322 23660 24332 23716
rect 24388 23660 25004 23716
rect 25060 23660 25070 23716
rect 26002 23660 26012 23716
rect 26068 23660 27692 23716
rect 27748 23660 27758 23716
rect 0 23604 400 23632
rect 13244 23604 13300 23660
rect 23996 23604 24052 23660
rect 0 23548 1652 23604
rect 1810 23548 1820 23604
rect 1876 23548 4956 23604
rect 5012 23548 5022 23604
rect 12646 23548 12684 23604
rect 12740 23548 12750 23604
rect 12898 23548 12908 23604
rect 12964 23548 13300 23604
rect 22194 23548 22204 23604
rect 22260 23548 22316 23604
rect 22372 23548 22382 23604
rect 23996 23548 26796 23604
rect 26852 23548 26862 23604
rect 0 23520 400 23548
rect 1596 23492 1652 23548
rect 8006 23492 8016 23548
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8280 23492 8290 23548
rect 14810 23492 14820 23548
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 15084 23492 15094 23548
rect 21614 23492 21624 23548
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21888 23492 21898 23548
rect 28418 23492 28428 23548
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28692 23492 28702 23548
rect 1596 23436 1764 23492
rect 8642 23436 8652 23492
rect 8708 23436 9324 23492
rect 9380 23436 9390 23492
rect 23734 23436 23772 23492
rect 23828 23436 23838 23492
rect 23986 23436 23996 23492
rect 24052 23436 25676 23492
rect 25732 23436 25742 23492
rect 1708 23380 1764 23436
rect 1698 23324 1708 23380
rect 1764 23324 1774 23380
rect 2034 23324 2044 23380
rect 2100 23324 3164 23380
rect 3220 23324 3388 23380
rect 4610 23324 4620 23380
rect 4676 23324 11788 23380
rect 11844 23324 11854 23380
rect 13010 23324 13020 23380
rect 13076 23324 15148 23380
rect 15204 23324 15214 23380
rect 19842 23324 19852 23380
rect 19908 23324 20300 23380
rect 20356 23324 20366 23380
rect 21410 23324 21420 23380
rect 21476 23324 22204 23380
rect 22260 23324 22428 23380
rect 22484 23324 23100 23380
rect 23156 23324 23166 23380
rect 26674 23324 26684 23380
rect 26740 23324 26796 23380
rect 26852 23324 26862 23380
rect 3332 23156 3388 23324
rect 11788 23268 11844 23324
rect 6626 23212 6636 23268
rect 6692 23212 7532 23268
rect 7588 23212 7598 23268
rect 11788 23212 14532 23268
rect 21970 23212 21980 23268
rect 22036 23212 22652 23268
rect 22708 23212 22718 23268
rect 23762 23212 23772 23268
rect 23828 23212 25228 23268
rect 25284 23212 25294 23268
rect 14476 23156 14532 23212
rect 3332 23100 4508 23156
rect 4564 23100 4574 23156
rect 14466 23100 14476 23156
rect 14532 23100 14542 23156
rect 15810 23100 15820 23156
rect 15876 23100 16380 23156
rect 16436 23100 16446 23156
rect 20626 23100 20636 23156
rect 20692 23100 20702 23156
rect 26674 23100 26684 23156
rect 26740 23100 27356 23156
rect 27412 23100 27422 23156
rect 20636 23044 20692 23100
rect 6290 22988 6300 23044
rect 6356 22988 7196 23044
rect 7252 22988 7262 23044
rect 12226 22988 12236 23044
rect 12292 22988 13356 23044
rect 13412 22988 13692 23044
rect 13748 22988 16828 23044
rect 16884 22988 17612 23044
rect 17668 22988 17948 23044
rect 18004 22988 19068 23044
rect 19124 22988 19516 23044
rect 19572 22988 19740 23044
rect 19796 22988 19806 23044
rect 20636 22988 23716 23044
rect 24658 22988 24668 23044
rect 24724 22988 28028 23044
rect 28084 22988 28094 23044
rect 7298 22876 7308 22932
rect 7364 22876 8316 22932
rect 8372 22876 8382 22932
rect 11890 22876 11900 22932
rect 11956 22876 12460 22932
rect 12516 22876 12526 22932
rect 15446 22876 15484 22932
rect 15540 22876 15550 22932
rect 20402 22876 20412 22932
rect 20468 22876 21196 22932
rect 21252 22876 21262 22932
rect 22194 22876 22204 22932
rect 22260 22876 22652 22932
rect 22708 22876 22718 22932
rect 15250 22764 15260 22820
rect 15316 22764 15596 22820
rect 15652 22764 15662 22820
rect 17350 22764 17388 22820
rect 17444 22764 17454 22820
rect 4604 22708 4614 22764
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4878 22708 4888 22764
rect 11408 22708 11418 22764
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11682 22708 11692 22764
rect 18212 22708 18222 22764
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18486 22708 18496 22764
rect 23660 22708 23716 22988
rect 25016 22708 25026 22764
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25290 22708 25300 22764
rect 15698 22652 15708 22708
rect 15764 22652 16380 22708
rect 16436 22652 16446 22708
rect 19282 22652 19292 22708
rect 19348 22652 22988 22708
rect 23044 22652 23054 22708
rect 23660 22652 23884 22708
rect 23940 22652 23950 22708
rect 3826 22540 3836 22596
rect 3892 22540 4620 22596
rect 4676 22540 5516 22596
rect 5572 22540 5582 22596
rect 8194 22540 8204 22596
rect 8260 22540 8652 22596
rect 8708 22540 8876 22596
rect 8932 22540 9660 22596
rect 9716 22540 10108 22596
rect 10164 22540 11004 22596
rect 11060 22540 12012 22596
rect 12068 22540 19292 22596
rect 19348 22540 25116 22596
rect 25172 22540 25182 22596
rect 13570 22428 13580 22484
rect 13636 22428 14700 22484
rect 14756 22428 16604 22484
rect 16660 22428 16670 22484
rect 17826 22428 17836 22484
rect 17892 22428 18620 22484
rect 18676 22428 20300 22484
rect 20356 22428 22092 22484
rect 22148 22428 22316 22484
rect 22372 22428 22382 22484
rect 22866 22428 22876 22484
rect 22932 22428 23436 22484
rect 23492 22428 23996 22484
rect 24052 22428 24062 22484
rect 11778 22316 11788 22372
rect 11844 22316 12684 22372
rect 12740 22316 16044 22372
rect 16100 22316 17052 22372
rect 17108 22316 17118 22372
rect 19058 22316 19068 22372
rect 19124 22316 19852 22372
rect 19908 22316 19918 22372
rect 23734 22316 23772 22372
rect 23828 22316 23838 22372
rect 3266 22204 3276 22260
rect 3332 22204 3724 22260
rect 3780 22204 3790 22260
rect 25106 22204 25116 22260
rect 25172 22204 27020 22260
rect 27076 22204 27086 22260
rect 1810 22092 1820 22148
rect 1876 22092 4396 22148
rect 4452 22092 4462 22148
rect 15138 22092 15148 22148
rect 15204 22092 15596 22148
rect 15652 22092 17500 22148
rect 17556 22092 17566 22148
rect 17714 22092 17724 22148
rect 17780 22092 17818 22148
rect 18162 22092 18172 22148
rect 18228 22092 22820 22148
rect 2706 21980 2716 22036
rect 2772 21980 3500 22036
rect 3556 21980 3566 22036
rect 8006 21924 8016 21980
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8280 21924 8290 21980
rect 14810 21924 14820 21980
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 15084 21924 15094 21980
rect 21614 21924 21624 21980
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21888 21924 21898 21980
rect 22764 21924 22820 22092
rect 28418 21924 28428 21980
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28692 21924 28702 21980
rect 22754 21868 22764 21924
rect 22820 21868 23548 21924
rect 23604 21868 23614 21924
rect 9650 21756 9660 21812
rect 9716 21756 12348 21812
rect 12404 21756 12908 21812
rect 12964 21756 13580 21812
rect 13636 21756 13646 21812
rect 19058 21756 19068 21812
rect 19124 21756 19628 21812
rect 19684 21756 21420 21812
rect 21476 21756 21486 21812
rect 23090 21756 23100 21812
rect 23156 21756 24332 21812
rect 24388 21756 24398 21812
rect 7970 21644 7980 21700
rect 8036 21644 8428 21700
rect 8484 21644 9884 21700
rect 9940 21644 9950 21700
rect 14466 21644 14476 21700
rect 14532 21644 15148 21700
rect 15204 21644 16492 21700
rect 16548 21644 16558 21700
rect 20962 21644 20972 21700
rect 21028 21644 23268 21700
rect 23426 21644 23436 21700
rect 23492 21644 26236 21700
rect 26292 21644 26302 21700
rect 23212 21588 23268 21644
rect 17602 21532 17612 21588
rect 17668 21532 17948 21588
rect 18004 21532 18956 21588
rect 19012 21532 22652 21588
rect 22708 21532 22718 21588
rect 23212 21532 24220 21588
rect 24276 21532 25452 21588
rect 25508 21532 25518 21588
rect 10434 21420 10444 21476
rect 10500 21420 12460 21476
rect 12516 21420 12526 21476
rect 14242 21420 14252 21476
rect 14308 21420 15036 21476
rect 15092 21420 18060 21476
rect 18116 21420 18126 21476
rect 20738 21420 20748 21476
rect 20804 21420 21868 21476
rect 21924 21420 21934 21476
rect 6850 21308 6860 21364
rect 6916 21308 8316 21364
rect 8372 21308 8382 21364
rect 16940 21308 17724 21364
rect 17780 21308 18396 21364
rect 18452 21308 19180 21364
rect 19236 21308 19246 21364
rect 25778 21308 25788 21364
rect 25844 21308 26908 21364
rect 26964 21308 26974 21364
rect 16940 21252 16996 21308
rect 2370 21196 2380 21252
rect 2436 21196 3052 21252
rect 3108 21196 3612 21252
rect 3668 21196 3678 21252
rect 16930 21196 16940 21252
rect 16996 21196 17006 21252
rect 4604 21140 4614 21196
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4878 21140 4888 21196
rect 11408 21140 11418 21196
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11682 21140 11692 21196
rect 18212 21140 18222 21196
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18486 21140 18496 21196
rect 25016 21140 25026 21196
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25290 21140 25300 21196
rect 7186 21084 7196 21140
rect 7252 21084 10556 21140
rect 10612 21084 10622 21140
rect 7410 20972 7420 21028
rect 7476 20972 9100 21028
rect 9156 20972 10780 21028
rect 10836 20972 10846 21028
rect 10994 20972 11004 21028
rect 11060 20972 11676 21028
rect 11732 20972 11742 21028
rect 19506 20972 19516 21028
rect 19572 20972 20076 21028
rect 20132 20972 20142 21028
rect 26338 20972 26348 21028
rect 26404 20972 27132 21028
rect 27188 20972 27198 21028
rect 0 20916 400 20944
rect 0 20860 1820 20916
rect 1876 20860 1886 20916
rect 5058 20860 5068 20916
rect 5124 20860 8204 20916
rect 8260 20860 8270 20916
rect 9426 20860 9436 20916
rect 9492 20860 9502 20916
rect 10210 20860 10220 20916
rect 10276 20860 11340 20916
rect 11396 20860 12908 20916
rect 12964 20860 14252 20916
rect 14308 20860 15708 20916
rect 15764 20860 16604 20916
rect 16660 20860 17836 20916
rect 17892 20860 19572 20916
rect 0 20832 400 20860
rect 9436 20804 9492 20860
rect 19516 20804 19572 20860
rect 2034 20748 2044 20804
rect 2100 20748 2716 20804
rect 2772 20748 2782 20804
rect 8642 20748 8652 20804
rect 8708 20748 9772 20804
rect 9828 20748 9838 20804
rect 11778 20748 11788 20804
rect 11844 20748 13132 20804
rect 13188 20748 13198 20804
rect 19506 20748 19516 20804
rect 19572 20748 19582 20804
rect 22642 20748 22652 20804
rect 22708 20748 22876 20804
rect 22932 20748 22942 20804
rect 23986 20748 23996 20804
rect 24052 20748 27132 20804
rect 27188 20748 28140 20804
rect 28196 20748 28206 20804
rect 6178 20636 6188 20692
rect 6244 20636 7084 20692
rect 7140 20636 7150 20692
rect 7298 20636 7308 20692
rect 7364 20636 7756 20692
rect 7812 20636 9436 20692
rect 9492 20636 10556 20692
rect 10612 20636 10622 20692
rect 12450 20636 12460 20692
rect 12516 20636 13692 20692
rect 13748 20636 13758 20692
rect 18050 20636 18060 20692
rect 18116 20636 20412 20692
rect 20468 20636 20478 20692
rect 24434 20636 24444 20692
rect 24500 20636 25788 20692
rect 25844 20636 25854 20692
rect 26114 20636 26124 20692
rect 26180 20636 27468 20692
rect 27524 20636 27534 20692
rect 9762 20524 9772 20580
rect 9828 20524 10668 20580
rect 10724 20524 10734 20580
rect 13458 20524 13468 20580
rect 13524 20524 13534 20580
rect 21410 20524 21420 20580
rect 21476 20524 22204 20580
rect 22260 20524 22270 20580
rect 22418 20524 22428 20580
rect 22484 20524 22876 20580
rect 22932 20524 22942 20580
rect 8006 20356 8016 20412
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8280 20356 8290 20412
rect 3042 20300 3052 20356
rect 3108 20300 3388 20356
rect 3444 20300 3454 20356
rect 13468 20244 13524 20524
rect 14810 20356 14820 20412
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 15084 20356 15094 20412
rect 21614 20356 21624 20412
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21888 20356 21898 20412
rect 28418 20356 28428 20412
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28692 20356 28702 20412
rect 25442 20300 25452 20356
rect 25508 20300 27916 20356
rect 27972 20300 27982 20356
rect 6626 20188 6636 20244
rect 6692 20188 8876 20244
rect 8932 20188 9996 20244
rect 10052 20188 10062 20244
rect 10546 20188 10556 20244
rect 10612 20188 11452 20244
rect 11508 20188 15148 20244
rect 15092 20132 15148 20188
rect 17052 20188 18956 20244
rect 19012 20188 19022 20244
rect 22082 20188 22092 20244
rect 22148 20188 23100 20244
rect 23156 20188 23166 20244
rect 23436 20188 23548 20244
rect 23604 20188 23772 20244
rect 23828 20188 23838 20244
rect 17052 20132 17108 20188
rect 23436 20132 23492 20188
rect 3266 20076 3276 20132
rect 3332 20076 3500 20132
rect 3556 20076 4396 20132
rect 4452 20076 5404 20132
rect 5460 20076 5470 20132
rect 12898 20076 12908 20132
rect 12964 20076 13916 20132
rect 13972 20076 13982 20132
rect 15092 20076 15484 20132
rect 15540 20076 16044 20132
rect 16100 20076 17052 20132
rect 17108 20076 17118 20132
rect 22306 20076 22316 20132
rect 22372 20076 23492 20132
rect 24658 20076 24668 20132
rect 24724 20076 26572 20132
rect 26628 20076 27020 20132
rect 27076 20076 27086 20132
rect 2706 19964 2716 20020
rect 2772 19964 3948 20020
rect 4004 19964 4014 20020
rect 10770 19964 10780 20020
rect 10836 19964 12460 20020
rect 12516 19964 12526 20020
rect 15372 19964 16268 20020
rect 16324 19964 16334 20020
rect 25330 19964 25340 20020
rect 25396 19964 28028 20020
rect 28084 19964 28094 20020
rect 15372 19908 15428 19964
rect 3826 19852 3836 19908
rect 3892 19852 4956 19908
rect 5012 19852 5022 19908
rect 9090 19852 9100 19908
rect 9156 19852 15372 19908
rect 15428 19852 15438 19908
rect 20066 19852 20076 19908
rect 20132 19852 21308 19908
rect 21364 19852 21374 19908
rect 4498 19740 4508 19796
rect 4564 19740 12460 19796
rect 12516 19740 12526 19796
rect 4604 19572 4614 19628
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4878 19572 4888 19628
rect 11408 19572 11418 19628
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11682 19572 11692 19628
rect 18212 19572 18222 19628
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18486 19572 18496 19628
rect 25016 19572 25026 19628
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25290 19572 25300 19628
rect 16594 19404 16604 19460
rect 16660 19404 18284 19460
rect 18340 19404 18350 19460
rect 19506 19404 19516 19460
rect 19572 19404 20300 19460
rect 20356 19404 21644 19460
rect 21700 19404 22540 19460
rect 22596 19404 22606 19460
rect 6402 19292 6412 19348
rect 6468 19292 7196 19348
rect 7252 19292 7262 19348
rect 15334 19292 15372 19348
rect 15428 19292 15438 19348
rect 20514 19292 20524 19348
rect 20580 19292 22652 19348
rect 22708 19292 24444 19348
rect 24500 19292 24668 19348
rect 24724 19292 24734 19348
rect 6066 19180 6076 19236
rect 6132 19180 6636 19236
rect 6692 19180 6702 19236
rect 7746 19180 7756 19236
rect 7812 19180 8540 19236
rect 8596 19180 8606 19236
rect 12450 19180 12460 19236
rect 12516 19180 13804 19236
rect 13860 19180 22428 19236
rect 22484 19180 25452 19236
rect 25508 19180 25518 19236
rect 14018 19068 14028 19124
rect 14084 19068 15596 19124
rect 15652 19068 15662 19124
rect 16034 19068 16044 19124
rect 16100 19068 16268 19124
rect 16324 19068 16492 19124
rect 16548 19068 16558 19124
rect 21522 19068 21532 19124
rect 21588 19068 21756 19124
rect 21812 19068 21822 19124
rect 5954 18956 5964 19012
rect 6020 18956 6524 19012
rect 6580 18956 6590 19012
rect 6962 18956 6972 19012
rect 7028 18956 7644 19012
rect 7700 18956 7710 19012
rect 12786 18956 12796 19012
rect 12852 18956 13580 19012
rect 13636 18956 13646 19012
rect 15810 18956 15820 19012
rect 15876 18956 18620 19012
rect 18676 18956 18956 19012
rect 19012 18956 19404 19012
rect 19460 18956 19470 19012
rect 20066 18956 20076 19012
rect 20132 18956 20636 19012
rect 20692 18956 22316 19012
rect 22372 18956 22382 19012
rect 24434 18956 24444 19012
rect 24500 18956 26348 19012
rect 26404 18956 26414 19012
rect 8006 18788 8016 18844
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8280 18788 8290 18844
rect 14810 18788 14820 18844
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 15084 18788 15094 18844
rect 21614 18788 21624 18844
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21888 18788 21898 18844
rect 28418 18788 28428 18844
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28692 18788 28702 18844
rect 26114 18732 26124 18788
rect 26180 18732 27020 18788
rect 27076 18732 27804 18788
rect 27860 18732 27870 18788
rect 23090 18620 23100 18676
rect 23156 18620 24332 18676
rect 24388 18620 26348 18676
rect 26404 18620 26414 18676
rect 2594 18508 2604 18564
rect 2660 18508 3836 18564
rect 3892 18508 3902 18564
rect 6626 18508 6636 18564
rect 6692 18508 10108 18564
rect 10164 18508 10780 18564
rect 10836 18508 10846 18564
rect 24658 18508 24668 18564
rect 24724 18508 27580 18564
rect 27636 18508 27646 18564
rect 3714 18396 3724 18452
rect 3780 18396 4396 18452
rect 4452 18396 4462 18452
rect 7522 18396 7532 18452
rect 7588 18396 8540 18452
rect 8596 18396 9660 18452
rect 9716 18396 9726 18452
rect 11554 18396 11564 18452
rect 11620 18396 11630 18452
rect 12338 18396 12348 18452
rect 12404 18396 13580 18452
rect 13636 18396 13646 18452
rect 15092 18396 17612 18452
rect 17668 18396 17948 18452
rect 18004 18396 18014 18452
rect 19730 18396 19740 18452
rect 19796 18396 20748 18452
rect 20804 18396 20814 18452
rect 23426 18396 23436 18452
rect 23492 18396 25228 18452
rect 25284 18396 25294 18452
rect 25666 18396 25676 18452
rect 25732 18396 26236 18452
rect 26292 18396 26302 18452
rect 11564 18340 11620 18396
rect 15092 18340 15148 18396
rect 4946 18284 4956 18340
rect 5012 18284 9100 18340
rect 9156 18284 9166 18340
rect 10322 18284 10332 18340
rect 10388 18284 15148 18340
rect 16258 18284 16268 18340
rect 16324 18284 16828 18340
rect 16884 18284 16894 18340
rect 0 18228 400 18256
rect 0 18172 1708 18228
rect 1764 18172 2492 18228
rect 2548 18172 2558 18228
rect 15810 18172 15820 18228
rect 15876 18172 17500 18228
rect 17556 18172 22092 18228
rect 22148 18172 22158 18228
rect 0 18144 400 18172
rect 7858 18060 7868 18116
rect 7924 18060 8540 18116
rect 8596 18060 9212 18116
rect 9268 18060 9278 18116
rect 4604 18004 4614 18060
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4878 18004 4888 18060
rect 11408 18004 11418 18060
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11682 18004 11692 18060
rect 18212 18004 18222 18060
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18486 18004 18496 18060
rect 25016 18004 25026 18060
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25290 18004 25300 18060
rect 13682 17948 13692 18004
rect 13748 17948 14588 18004
rect 14644 17948 14654 18004
rect 16930 17948 16940 18004
rect 16996 17948 17006 18004
rect 10434 17836 10444 17892
rect 10500 17836 11228 17892
rect 11284 17836 15932 17892
rect 15988 17836 15998 17892
rect 5170 17724 5180 17780
rect 5236 17724 5740 17780
rect 5796 17724 6636 17780
rect 6692 17724 8988 17780
rect 9044 17724 9054 17780
rect 15250 17724 15260 17780
rect 15316 17724 15484 17780
rect 15540 17724 15550 17780
rect 2034 17612 2044 17668
rect 2100 17612 2940 17668
rect 2996 17612 4172 17668
rect 4228 17612 4238 17668
rect 11666 17612 11676 17668
rect 11732 17612 12572 17668
rect 12628 17612 12638 17668
rect 14018 17612 14028 17668
rect 14084 17612 14588 17668
rect 14644 17612 14654 17668
rect 14914 17612 14924 17668
rect 14980 17612 15708 17668
rect 15764 17612 15774 17668
rect 16940 17556 16996 17948
rect 22978 17612 22988 17668
rect 23044 17612 24108 17668
rect 24164 17612 25900 17668
rect 25956 17612 25966 17668
rect 12338 17500 12348 17556
rect 12404 17500 14700 17556
rect 14756 17500 14766 17556
rect 15474 17500 15484 17556
rect 15540 17500 16268 17556
rect 16324 17500 16334 17556
rect 16930 17500 16940 17556
rect 16996 17500 17006 17556
rect 18610 17500 18620 17556
rect 18676 17500 18956 17556
rect 19012 17500 19022 17556
rect 21298 17500 21308 17556
rect 21364 17500 23436 17556
rect 23492 17500 23502 17556
rect 25900 17444 25956 17612
rect 3042 17388 3052 17444
rect 3108 17388 3388 17444
rect 3444 17388 3454 17444
rect 8418 17388 8428 17444
rect 8484 17388 9436 17444
rect 9492 17388 10220 17444
rect 10276 17388 10286 17444
rect 12002 17388 12012 17444
rect 12068 17388 12460 17444
rect 12516 17388 17276 17444
rect 17332 17388 17342 17444
rect 21196 17388 25228 17444
rect 25284 17388 25294 17444
rect 25900 17388 28028 17444
rect 28084 17388 28094 17444
rect 21196 17332 21252 17388
rect 12898 17276 12908 17332
rect 12964 17276 14252 17332
rect 14308 17276 14318 17332
rect 15922 17276 15932 17332
rect 15988 17276 16716 17332
rect 16772 17276 18844 17332
rect 18900 17276 19068 17332
rect 19124 17276 19740 17332
rect 19796 17276 21196 17332
rect 21252 17276 21262 17332
rect 8006 17220 8016 17276
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8280 17220 8290 17276
rect 14810 17220 14820 17276
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 15084 17220 15094 17276
rect 21614 17220 21624 17276
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21888 17220 21898 17276
rect 28418 17220 28428 17276
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28692 17220 28702 17276
rect 15362 17164 15372 17220
rect 15428 17164 16268 17220
rect 16324 17164 16334 17220
rect 22754 17164 22764 17220
rect 22820 17164 23996 17220
rect 24052 17164 24668 17220
rect 24724 17164 26012 17220
rect 26068 17164 27020 17220
rect 27076 17164 27086 17220
rect 7410 17052 7420 17108
rect 7476 17052 8204 17108
rect 8260 17052 10332 17108
rect 10388 17052 10398 17108
rect 11666 17052 11676 17108
rect 11732 17052 16884 17108
rect 17266 17052 17276 17108
rect 17332 17052 18060 17108
rect 18116 17052 20524 17108
rect 20580 17052 20590 17108
rect 20962 17052 20972 17108
rect 21028 17052 21756 17108
rect 21812 17052 21822 17108
rect 7186 16940 7196 16996
rect 7252 16940 7756 16996
rect 7812 16940 7822 16996
rect 16230 16940 16268 16996
rect 16324 16940 16334 16996
rect 16828 16884 16884 17052
rect 18610 16940 18620 16996
rect 18676 16940 19180 16996
rect 19236 16940 19246 16996
rect 19964 16940 20300 16996
rect 20356 16940 22652 16996
rect 22708 16940 26348 16996
rect 26404 16940 26414 16996
rect 19964 16884 20020 16940
rect 5170 16828 5180 16884
rect 5236 16828 6076 16884
rect 6132 16828 6142 16884
rect 10210 16828 10220 16884
rect 10276 16828 10780 16884
rect 10836 16828 10846 16884
rect 14242 16828 14252 16884
rect 14308 16828 15204 16884
rect 16818 16828 16828 16884
rect 16884 16828 17612 16884
rect 17668 16828 20020 16884
rect 20178 16828 20188 16884
rect 20244 16828 22204 16884
rect 22260 16828 22270 16884
rect 26562 16828 26572 16884
rect 26628 16828 27580 16884
rect 27636 16828 27646 16884
rect 15148 16772 15204 16828
rect 5618 16716 5628 16772
rect 5684 16716 5852 16772
rect 5908 16716 6748 16772
rect 6804 16716 6814 16772
rect 15148 16716 15596 16772
rect 15652 16716 15662 16772
rect 4604 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4888 16492
rect 11408 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11692 16492
rect 18212 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18496 16492
rect 25016 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25300 16492
rect 9762 16268 9772 16324
rect 9828 16268 12124 16324
rect 12180 16268 12190 16324
rect 13794 16156 13804 16212
rect 13860 16156 14588 16212
rect 14644 16156 14654 16212
rect 15138 16156 15148 16212
rect 15204 16156 17052 16212
rect 17108 16156 18396 16212
rect 18452 16156 18732 16212
rect 18788 16156 20076 16212
rect 20132 16156 20142 16212
rect 10210 16044 10220 16100
rect 10276 16044 12796 16100
rect 12852 16044 12862 16100
rect 18050 16044 18060 16100
rect 18116 16044 20300 16100
rect 20356 16044 21308 16100
rect 21364 16044 21374 16100
rect 11106 15820 11116 15876
rect 11172 15820 12460 15876
rect 12516 15820 12526 15876
rect 12786 15820 12796 15876
rect 12852 15820 13692 15876
rect 13748 15820 19292 15876
rect 19348 15820 19358 15876
rect 11218 15708 11228 15764
rect 11284 15708 12348 15764
rect 12404 15708 13020 15764
rect 13076 15708 13086 15764
rect 22642 15708 22652 15764
rect 22708 15708 22718 15764
rect 8006 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8290 15708
rect 14810 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15094 15708
rect 21614 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21898 15708
rect 22652 15652 22708 15708
rect 28418 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28702 15708
rect 22652 15596 24724 15652
rect 0 15540 400 15568
rect 0 15484 1820 15540
rect 1876 15484 1886 15540
rect 6514 15484 6524 15540
rect 6580 15484 7756 15540
rect 7812 15484 8540 15540
rect 8596 15484 8606 15540
rect 13346 15484 13356 15540
rect 13412 15484 18788 15540
rect 18946 15484 18956 15540
rect 19012 15484 19964 15540
rect 20020 15484 20636 15540
rect 20692 15484 20702 15540
rect 0 15456 400 15484
rect 6066 15372 6076 15428
rect 6132 15372 7084 15428
rect 7140 15372 7150 15428
rect 7410 15372 7420 15428
rect 7476 15372 10668 15428
rect 10724 15372 10734 15428
rect 15138 15372 15148 15428
rect 15204 15372 16604 15428
rect 16660 15372 16670 15428
rect 18732 15316 18788 15484
rect 22652 15428 22708 15596
rect 24668 15540 24724 15596
rect 24658 15484 24668 15540
rect 24724 15484 26796 15540
rect 26852 15484 26862 15540
rect 19282 15372 19292 15428
rect 19348 15372 19740 15428
rect 19796 15372 22708 15428
rect 6178 15260 6188 15316
rect 6244 15260 7868 15316
rect 7924 15260 7934 15316
rect 14802 15260 14812 15316
rect 14868 15260 15260 15316
rect 15316 15260 15326 15316
rect 18722 15260 18732 15316
rect 18788 15260 20188 15316
rect 20244 15260 24108 15316
rect 24164 15260 24556 15316
rect 24612 15260 26348 15316
rect 26404 15260 26414 15316
rect 2034 15148 2044 15204
rect 2100 15148 2604 15204
rect 2660 15148 3500 15204
rect 3556 15148 3566 15204
rect 3826 15148 3836 15204
rect 3892 15148 5628 15204
rect 5684 15148 6860 15204
rect 6916 15148 6926 15204
rect 7410 15148 7420 15204
rect 7476 15148 7980 15204
rect 8036 15148 8046 15204
rect 14578 15148 14588 15204
rect 14644 15148 21196 15204
rect 21252 15148 22204 15204
rect 22260 15148 23548 15204
rect 23604 15148 23614 15204
rect 16706 15036 16716 15092
rect 16772 15036 22876 15092
rect 22932 15036 22942 15092
rect 2034 14924 2044 14980
rect 2100 14924 2380 14980
rect 2436 14924 2716 14980
rect 2772 14924 2782 14980
rect 16902 14924 16940 14980
rect 16996 14924 17006 14980
rect 4604 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4888 14924
rect 11408 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11692 14924
rect 18212 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18496 14924
rect 25016 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25300 14924
rect 2258 14700 2268 14756
rect 2324 14700 2334 14756
rect 9846 14700 9884 14756
rect 9940 14700 9950 14756
rect 10108 14700 19180 14756
rect 19236 14700 19246 14756
rect 24322 14700 24332 14756
rect 24388 14700 25676 14756
rect 25732 14700 25742 14756
rect 2268 14532 2324 14700
rect 10108 14644 10164 14700
rect 5058 14588 5068 14644
rect 5124 14588 5516 14644
rect 5572 14588 5582 14644
rect 8754 14588 8764 14644
rect 8820 14588 10164 14644
rect 14578 14588 14588 14644
rect 14644 14588 20748 14644
rect 20804 14588 21532 14644
rect 21588 14588 21598 14644
rect 2268 14476 2492 14532
rect 2548 14476 2558 14532
rect 2818 14364 2828 14420
rect 2884 14364 3276 14420
rect 3332 14364 3342 14420
rect 4610 14364 4620 14420
rect 4676 14364 4956 14420
rect 5012 14364 5964 14420
rect 6020 14364 6030 14420
rect 7298 14364 7308 14420
rect 7364 14364 8540 14420
rect 8596 14364 8606 14420
rect 19058 14364 19068 14420
rect 19124 14364 21196 14420
rect 21252 14364 23212 14420
rect 23268 14364 24444 14420
rect 24500 14364 24510 14420
rect 22092 14308 22148 14364
rect 5814 14252 5852 14308
rect 5908 14252 5918 14308
rect 12002 14252 12012 14308
rect 12068 14252 14140 14308
rect 14196 14252 15708 14308
rect 15764 14252 15774 14308
rect 22082 14252 22092 14308
rect 22148 14252 22158 14308
rect 8006 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8290 14140
rect 14810 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15094 14140
rect 21614 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21898 14140
rect 28418 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28702 14140
rect 2258 13916 2268 13972
rect 2324 13916 3388 13972
rect 3444 13916 3500 13972
rect 3556 13916 3566 13972
rect 9874 13916 9884 13972
rect 9940 13916 11564 13972
rect 11620 13916 11630 13972
rect 14242 13916 14252 13972
rect 14308 13916 15036 13972
rect 15092 13916 15260 13972
rect 15316 13916 16716 13972
rect 16772 13916 16782 13972
rect 2482 13804 2492 13860
rect 2548 13804 2716 13860
rect 2772 13804 3612 13860
rect 3668 13804 3678 13860
rect 8306 13804 8316 13860
rect 8372 13804 10444 13860
rect 10500 13804 10510 13860
rect 14914 13804 14924 13860
rect 14980 13804 17948 13860
rect 18004 13804 19068 13860
rect 19124 13804 19134 13860
rect 26852 13804 27132 13860
rect 27188 13804 27198 13860
rect 26852 13748 26908 13804
rect 8082 13692 8092 13748
rect 8148 13692 10780 13748
rect 10836 13692 10846 13748
rect 13794 13692 13804 13748
rect 13860 13692 14812 13748
rect 14868 13692 14878 13748
rect 21970 13692 21980 13748
rect 22036 13692 23548 13748
rect 23604 13692 26908 13748
rect 3378 13580 3388 13636
rect 3444 13580 4956 13636
rect 5012 13580 5022 13636
rect 9986 13580 9996 13636
rect 10052 13580 17052 13636
rect 17108 13580 17118 13636
rect 17714 13580 17724 13636
rect 17780 13580 18396 13636
rect 18452 13580 18462 13636
rect 24210 13580 24220 13636
rect 24276 13580 25788 13636
rect 25844 13580 26460 13636
rect 26516 13580 26526 13636
rect 4162 13468 4172 13524
rect 4228 13468 5964 13524
rect 6020 13468 6030 13524
rect 9762 13468 9772 13524
rect 9828 13468 10892 13524
rect 10948 13468 10958 13524
rect 6962 13356 6972 13412
rect 7028 13356 7644 13412
rect 7700 13356 8652 13412
rect 8708 13356 9548 13412
rect 9604 13356 9614 13412
rect 9846 13356 9884 13412
rect 9940 13356 9950 13412
rect 12674 13356 12684 13412
rect 12740 13356 13804 13412
rect 13860 13356 13870 13412
rect 4604 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4888 13356
rect 11408 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11692 13356
rect 18212 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18496 13356
rect 25016 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25300 13356
rect 26226 13244 26236 13300
rect 26292 13244 26516 13300
rect 26460 13188 26516 13244
rect 7074 13132 7084 13188
rect 7140 13132 12236 13188
rect 12292 13132 13692 13188
rect 13748 13132 13758 13188
rect 26450 13132 26460 13188
rect 26516 13132 26526 13188
rect 5506 13020 5516 13076
rect 5572 13020 8092 13076
rect 8148 13020 8158 13076
rect 10322 13020 10332 13076
rect 10388 13020 11340 13076
rect 11396 13020 12124 13076
rect 12180 13020 14140 13076
rect 14196 13020 14924 13076
rect 14980 13020 14990 13076
rect 24098 13020 24108 13076
rect 24164 13020 24444 13076
rect 24500 13020 24510 13076
rect 20178 12908 20188 12964
rect 20244 12908 20524 12964
rect 20580 12908 22764 12964
rect 22820 12908 23548 12964
rect 23604 12908 26124 12964
rect 26180 12908 26572 12964
rect 26628 12908 26638 12964
rect 0 12852 400 12880
rect 0 12796 1708 12852
rect 1764 12796 1774 12852
rect 6178 12796 6188 12852
rect 6244 12796 7084 12852
rect 7140 12796 7150 12852
rect 9324 12796 10108 12852
rect 10164 12796 11452 12852
rect 11508 12796 11518 12852
rect 17938 12796 17948 12852
rect 18004 12796 18396 12852
rect 18452 12796 18462 12852
rect 0 12768 400 12796
rect 9324 12740 9380 12796
rect 7410 12684 7420 12740
rect 7476 12684 8540 12740
rect 8596 12684 9324 12740
rect 9380 12684 9390 12740
rect 9874 12684 9884 12740
rect 9940 12684 11788 12740
rect 11844 12684 11854 12740
rect 13570 12684 13580 12740
rect 13636 12684 16548 12740
rect 16706 12684 16716 12740
rect 16772 12684 17388 12740
rect 17444 12684 18172 12740
rect 18228 12684 19628 12740
rect 19684 12684 20972 12740
rect 21028 12684 22540 12740
rect 22596 12684 22988 12740
rect 23044 12684 23054 12740
rect 16492 12628 16548 12684
rect 16492 12572 18284 12628
rect 18340 12572 20188 12628
rect 20244 12572 20254 12628
rect 8006 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8290 12572
rect 14810 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15094 12572
rect 21614 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21898 12572
rect 28418 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28702 12572
rect 2370 12348 2380 12404
rect 2436 12348 4060 12404
rect 4116 12348 4126 12404
rect 5954 12348 5964 12404
rect 6020 12348 13356 12404
rect 13412 12348 13422 12404
rect 14690 12348 14700 12404
rect 14756 12348 16380 12404
rect 16436 12348 17724 12404
rect 17780 12348 18620 12404
rect 18676 12348 18686 12404
rect 18918 12348 18956 12404
rect 19012 12348 19022 12404
rect 21746 12348 21756 12404
rect 21812 12348 22204 12404
rect 22260 12348 22270 12404
rect 9538 12236 9548 12292
rect 9604 12236 10556 12292
rect 10612 12236 11004 12292
rect 11060 12236 18452 12292
rect 18610 12236 18620 12292
rect 18676 12236 19292 12292
rect 19348 12236 19358 12292
rect 18396 12180 18452 12236
rect 2706 12124 2716 12180
rect 2772 12124 3052 12180
rect 3108 12124 4284 12180
rect 4340 12124 4350 12180
rect 8978 12124 8988 12180
rect 9044 12124 9772 12180
rect 9828 12124 15484 12180
rect 15540 12124 15550 12180
rect 17378 12124 17388 12180
rect 17444 12124 17724 12180
rect 17780 12124 17790 12180
rect 18396 12124 21980 12180
rect 22036 12124 22046 12180
rect 23426 12124 23436 12180
rect 23492 12124 24668 12180
rect 24724 12124 25228 12180
rect 25284 12124 26460 12180
rect 26516 12124 26526 12180
rect 7298 12012 7308 12068
rect 7364 12012 8540 12068
rect 8596 12012 8606 12068
rect 16258 12012 16268 12068
rect 16324 12012 16828 12068
rect 16884 12012 17444 12068
rect 18498 12012 18508 12068
rect 18564 12012 19292 12068
rect 19348 12012 19358 12068
rect 17388 11956 17444 12012
rect 17388 11900 18620 11956
rect 18676 11900 18686 11956
rect 17388 11844 17444 11900
rect 17378 11788 17388 11844
rect 17444 11788 17454 11844
rect 18610 11788 18620 11844
rect 18676 11788 19740 11844
rect 19796 11788 19806 11844
rect 20178 11788 20188 11844
rect 20244 11788 22596 11844
rect 4604 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4888 11788
rect 11408 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11692 11788
rect 18212 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18496 11788
rect 18620 11732 18676 11788
rect 22540 11732 22596 11788
rect 25016 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25300 11788
rect 6402 11676 6412 11732
rect 6468 11676 6478 11732
rect 13570 11676 13580 11732
rect 13636 11676 14364 11732
rect 14420 11676 15148 11732
rect 15204 11676 15214 11732
rect 18610 11676 18620 11732
rect 18676 11676 18686 11732
rect 20402 11676 20412 11732
rect 20468 11676 20478 11732
rect 22530 11676 22540 11732
rect 22596 11676 22606 11732
rect 6412 11620 6468 11676
rect 20412 11620 20468 11676
rect 3938 11564 3948 11620
rect 4004 11564 6468 11620
rect 8754 11564 8764 11620
rect 8820 11564 11900 11620
rect 11956 11564 11966 11620
rect 15810 11564 15820 11620
rect 15876 11564 20468 11620
rect 20962 11564 20972 11620
rect 21028 11564 22316 11620
rect 22372 11564 22382 11620
rect 3332 11452 6748 11508
rect 6804 11452 6814 11508
rect 7858 11452 7868 11508
rect 7924 11452 9884 11508
rect 9940 11452 9950 11508
rect 10098 11452 10108 11508
rect 10164 11452 15148 11508
rect 19954 11452 19964 11508
rect 20020 11452 21308 11508
rect 21364 11452 22428 11508
rect 22484 11452 22494 11508
rect 3332 11396 3388 11452
rect 15092 11396 15148 11452
rect 2034 11340 2044 11396
rect 2100 11340 3388 11396
rect 3490 11340 3500 11396
rect 3556 11340 4508 11396
rect 4564 11340 4574 11396
rect 5814 11340 5852 11396
rect 5908 11340 5918 11396
rect 6066 11340 6076 11396
rect 6132 11340 11508 11396
rect 11890 11340 11900 11396
rect 11956 11340 12572 11396
rect 12628 11340 14476 11396
rect 14532 11340 14542 11396
rect 15092 11340 20076 11396
rect 20132 11340 20748 11396
rect 20804 11340 20814 11396
rect 11452 11284 11508 11340
rect 2818 11228 2828 11284
rect 2884 11228 4956 11284
rect 5012 11228 5022 11284
rect 5170 11228 5180 11284
rect 5236 11228 6300 11284
rect 6356 11228 6366 11284
rect 9202 11228 9212 11284
rect 9268 11228 10668 11284
rect 10724 11228 11228 11284
rect 11284 11228 11294 11284
rect 11452 11228 12908 11284
rect 12964 11228 13916 11284
rect 13972 11228 13982 11284
rect 14578 11228 14588 11284
rect 14644 11228 15820 11284
rect 15876 11228 15886 11284
rect 5180 11172 5236 11228
rect 2034 11116 2044 11172
rect 2100 11116 3388 11172
rect 4274 11116 4284 11172
rect 4340 11116 5236 11172
rect 5842 11116 5852 11172
rect 5908 11116 6636 11172
rect 6692 11116 10108 11172
rect 10164 11116 10174 11172
rect 11666 11116 11676 11172
rect 11732 11116 12460 11172
rect 12516 11116 13468 11172
rect 13524 11116 13534 11172
rect 15698 11116 15708 11172
rect 15764 11116 16940 11172
rect 16996 11116 17006 11172
rect 22082 11116 22092 11172
rect 22148 11116 22316 11172
rect 22372 11116 22382 11172
rect 2258 10892 2268 10948
rect 2324 10892 2604 10948
rect 2660 10892 2670 10948
rect 3332 10836 3388 11116
rect 10434 11004 10444 11060
rect 10500 11004 13580 11060
rect 13636 11004 13646 11060
rect 8006 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8290 11004
rect 14810 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15094 11004
rect 21614 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21898 11004
rect 28418 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28702 11004
rect 8372 10892 11788 10948
rect 11844 10892 11854 10948
rect 8372 10836 8428 10892
rect 1810 10780 1820 10836
rect 1876 10780 2156 10836
rect 2212 10780 2222 10836
rect 3332 10780 5068 10836
rect 5124 10780 8428 10836
rect 9874 10780 9884 10836
rect 9940 10780 10780 10836
rect 10836 10780 10846 10836
rect 12114 10780 12124 10836
rect 12180 10780 12796 10836
rect 12852 10780 14924 10836
rect 14980 10780 14990 10836
rect 17938 10780 17948 10836
rect 18004 10780 18732 10836
rect 18788 10780 18798 10836
rect 20262 10780 20300 10836
rect 20356 10780 20366 10836
rect 22530 10780 22540 10836
rect 22596 10780 24108 10836
rect 24164 10780 25788 10836
rect 25844 10780 25854 10836
rect 7746 10668 7756 10724
rect 7812 10668 8764 10724
rect 8820 10668 8830 10724
rect 14028 10612 14084 10780
rect 15362 10668 15372 10724
rect 15428 10668 16324 10724
rect 16706 10668 16716 10724
rect 16772 10668 19068 10724
rect 19124 10668 21644 10724
rect 21700 10668 22652 10724
rect 22708 10668 23212 10724
rect 23268 10668 23660 10724
rect 23716 10668 23726 10724
rect 16268 10612 16324 10668
rect 6738 10556 6748 10612
rect 6804 10556 8092 10612
rect 8148 10556 8158 10612
rect 11106 10556 11116 10612
rect 11172 10556 11788 10612
rect 11844 10556 11854 10612
rect 14018 10556 14028 10612
rect 14084 10556 14094 10612
rect 16230 10556 16268 10612
rect 16324 10556 16334 10612
rect 16482 10556 16492 10612
rect 16548 10556 16940 10612
rect 16996 10556 17612 10612
rect 17668 10556 17678 10612
rect 20178 10556 20188 10612
rect 20244 10556 21308 10612
rect 21364 10556 21374 10612
rect 13346 10444 13356 10500
rect 13412 10444 15708 10500
rect 15764 10444 15774 10500
rect 17378 10444 17388 10500
rect 17444 10444 20300 10500
rect 20356 10444 20366 10500
rect 21186 10444 21196 10500
rect 21252 10444 21980 10500
rect 22036 10444 26348 10500
rect 26404 10444 26414 10500
rect 6290 10332 6300 10388
rect 6356 10332 7644 10388
rect 7700 10332 7710 10388
rect 13794 10332 13804 10388
rect 13860 10332 16492 10388
rect 16548 10332 18508 10388
rect 18564 10332 18574 10388
rect 2034 10220 2044 10276
rect 2100 10220 2380 10276
rect 2436 10220 3388 10276
rect 3444 10220 3454 10276
rect 13570 10220 13580 10276
rect 13636 10220 14588 10276
rect 14644 10220 14654 10276
rect 14914 10220 14924 10276
rect 14980 10220 15372 10276
rect 15428 10220 16716 10276
rect 16772 10220 16782 10276
rect 0 10164 400 10192
rect 4604 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4888 10220
rect 11408 10164 11418 10220
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11682 10164 11692 10220
rect 18212 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18496 10220
rect 19516 10164 19572 10444
rect 25016 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25300 10220
rect 0 10108 2716 10164
rect 2772 10108 2782 10164
rect 4956 10108 5068 10164
rect 5124 10108 5134 10164
rect 14466 10108 14476 10164
rect 14532 10108 16268 10164
rect 16324 10108 16334 10164
rect 19506 10108 19516 10164
rect 19572 10108 19582 10164
rect 0 10080 400 10108
rect 4956 10052 5012 10108
rect 4834 9996 4844 10052
rect 4900 9996 5012 10052
rect 14690 9996 14700 10052
rect 14756 9996 15148 10052
rect 15204 9996 15214 10052
rect 16594 9996 16604 10052
rect 16660 9996 17836 10052
rect 17892 9996 20524 10052
rect 20580 9996 21532 10052
rect 21588 9996 21598 10052
rect 4498 9884 4508 9940
rect 4564 9884 6636 9940
rect 6692 9884 6702 9940
rect 15586 9884 15596 9940
rect 15652 9884 17052 9940
rect 17108 9884 17118 9940
rect 18610 9884 18620 9940
rect 18676 9884 19852 9940
rect 19908 9884 19918 9940
rect 9762 9772 9772 9828
rect 9828 9772 12796 9828
rect 12852 9772 12862 9828
rect 24882 9772 24892 9828
rect 24948 9772 25564 9828
rect 25620 9772 26012 9828
rect 26068 9772 26078 9828
rect 17378 9660 17388 9716
rect 17444 9660 18060 9716
rect 18116 9660 18126 9716
rect 16818 9436 16828 9492
rect 16884 9436 17388 9492
rect 17444 9436 17454 9492
rect 17602 9436 17612 9492
rect 17668 9436 19068 9492
rect 19124 9436 19628 9492
rect 19684 9436 19694 9492
rect 8006 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8290 9436
rect 14810 9380 14820 9436
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 15084 9380 15094 9436
rect 21614 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21898 9436
rect 28418 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28702 9436
rect 13458 9212 13468 9268
rect 13524 9212 14812 9268
rect 14868 9212 14878 9268
rect 15092 9212 15484 9268
rect 15540 9212 15550 9268
rect 1922 9100 1932 9156
rect 1988 9100 2380 9156
rect 2436 9100 3948 9156
rect 4004 9100 4014 9156
rect 13122 9100 13132 9156
rect 13188 9100 14140 9156
rect 14196 9100 14700 9156
rect 14756 9100 14766 9156
rect 14700 8932 14756 9100
rect 15092 9044 15148 9212
rect 16258 9100 16268 9156
rect 16324 9100 16828 9156
rect 16884 9100 17948 9156
rect 18004 9100 18844 9156
rect 18900 9100 21980 9156
rect 22036 9100 22046 9156
rect 14914 8988 14924 9044
rect 14980 8988 15148 9044
rect 22642 8988 22652 9044
rect 22708 8988 23436 9044
rect 23492 8988 23502 9044
rect 14700 8876 16156 8932
rect 16212 8876 16716 8932
rect 16772 8876 17836 8932
rect 17892 8876 17902 8932
rect 20934 8876 20972 8932
rect 21028 8876 21038 8932
rect 4604 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4888 8652
rect 11408 8596 11418 8652
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11682 8596 11692 8652
rect 18212 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18496 8652
rect 25016 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25300 8652
rect 2594 8428 2604 8484
rect 2660 8428 5516 8484
rect 5572 8428 6300 8484
rect 6356 8428 6366 8484
rect 3724 8372 3780 8428
rect 4732 8372 4788 8428
rect 2146 8316 2156 8372
rect 2212 8316 2828 8372
rect 2884 8316 3164 8372
rect 3220 8316 3230 8372
rect 3714 8316 3724 8372
rect 3780 8316 3790 8372
rect 4722 8316 4732 8372
rect 4788 8316 4798 8372
rect 13234 8316 13244 8372
rect 13300 8316 14252 8372
rect 14308 8316 14318 8372
rect 15026 8316 15036 8372
rect 15092 8316 18172 8372
rect 18228 8316 18238 8372
rect 20626 8316 20636 8372
rect 20692 8316 21196 8372
rect 21252 8316 21262 8372
rect 3378 8204 3388 8260
rect 3444 8204 15148 8260
rect 17378 8204 17388 8260
rect 17444 8204 18620 8260
rect 18676 8204 19292 8260
rect 19348 8204 19358 8260
rect 15092 8148 15148 8204
rect 6626 8092 6636 8148
rect 6692 8092 8092 8148
rect 8148 8092 8158 8148
rect 15092 8092 19740 8148
rect 19796 8092 19806 8148
rect 5058 7980 5068 8036
rect 5124 7980 5404 8036
rect 5460 7980 17276 8036
rect 17332 7980 17342 8036
rect 20598 7980 20636 8036
rect 20692 7980 20702 8036
rect 5170 7868 5180 7924
rect 5236 7868 6076 7924
rect 6132 7868 7420 7924
rect 7476 7868 7486 7924
rect 8006 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8290 7868
rect 14810 7812 14820 7868
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 15084 7812 15094 7868
rect 21614 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21898 7868
rect 28418 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28702 7868
rect 2930 7644 2940 7700
rect 2996 7644 5068 7700
rect 5124 7644 5134 7700
rect 6178 7644 6188 7700
rect 6244 7644 9212 7700
rect 9268 7644 9278 7700
rect 20290 7644 20300 7700
rect 20356 7644 20524 7700
rect 20580 7644 22092 7700
rect 22148 7644 23212 7700
rect 23268 7644 23278 7700
rect 2818 7532 2828 7588
rect 2884 7532 5516 7588
rect 5572 7532 5582 7588
rect 8978 7532 8988 7588
rect 9044 7532 17724 7588
rect 17780 7532 17790 7588
rect 0 7476 400 7504
rect 0 7420 1708 7476
rect 1764 7420 2492 7476
rect 2548 7420 2558 7476
rect 23874 7420 23884 7476
rect 23940 7420 24780 7476
rect 24836 7420 24846 7476
rect 0 7392 400 7420
rect 16146 7308 16156 7364
rect 16212 7308 19068 7364
rect 19124 7308 20300 7364
rect 20356 7308 20366 7364
rect 4604 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4888 7084
rect 11408 7028 11418 7084
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11682 7028 11692 7084
rect 18212 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18496 7084
rect 25016 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25300 7084
rect 4722 6636 4732 6692
rect 4788 6636 5404 6692
rect 5460 6636 5470 6692
rect 15698 6636 15708 6692
rect 15764 6636 19516 6692
rect 19572 6636 19582 6692
rect 19740 6636 20972 6692
rect 21028 6636 21644 6692
rect 21700 6636 21710 6692
rect 23762 6636 23772 6692
rect 23828 6636 24444 6692
rect 24500 6636 24510 6692
rect 19740 6580 19796 6636
rect 3378 6524 3388 6580
rect 3444 6524 4060 6580
rect 4116 6524 4396 6580
rect 4452 6524 19796 6580
rect 20514 6524 20524 6580
rect 20580 6524 21308 6580
rect 21364 6524 21374 6580
rect 2034 6300 2044 6356
rect 2100 6300 7644 6356
rect 7700 6300 7710 6356
rect 8006 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8290 6300
rect 14810 6244 14820 6300
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 15084 6244 15094 6300
rect 21614 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21898 6300
rect 28418 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28702 6300
rect 3826 6076 3836 6132
rect 3892 6076 18732 6132
rect 18788 6076 18798 6132
rect 24434 6076 24444 6132
rect 24500 6076 25452 6132
rect 25508 6076 25518 6132
rect 20066 5964 20076 6020
rect 20132 5964 22540 6020
rect 22596 5964 22606 6020
rect 23426 5964 23436 6020
rect 23492 5964 24556 6020
rect 24612 5964 24622 6020
rect 24770 5964 24780 6020
rect 24836 5964 26012 6020
rect 26068 5964 26078 6020
rect 20850 5852 20860 5908
rect 20916 5852 21868 5908
rect 21924 5852 21934 5908
rect 23650 5852 23660 5908
rect 23716 5852 25900 5908
rect 25956 5852 25966 5908
rect 19842 5740 19852 5796
rect 19908 5740 22428 5796
rect 22484 5740 22494 5796
rect 24546 5740 24556 5796
rect 24612 5740 25564 5796
rect 25620 5740 25630 5796
rect 22194 5628 22204 5684
rect 22260 5628 23884 5684
rect 23940 5628 23950 5684
rect 4604 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4888 5516
rect 11408 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11692 5516
rect 18212 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18496 5516
rect 25016 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25300 5516
rect 20402 5292 20412 5348
rect 20468 5292 25676 5348
rect 25732 5292 25742 5348
rect 21746 5180 21756 5236
rect 21812 5180 22540 5236
rect 22596 5180 22606 5236
rect 18722 5068 18732 5124
rect 18788 5068 20748 5124
rect 20804 5068 21532 5124
rect 21588 5068 21598 5124
rect 19628 4956 20412 5012
rect 20468 4956 21980 5012
rect 22036 4956 22046 5012
rect 0 4788 400 4816
rect 19628 4788 19684 4956
rect 19842 4844 19852 4900
rect 19908 4844 20636 4900
rect 20692 4844 20702 4900
rect 23986 4844 23996 4900
rect 24052 4844 26012 4900
rect 26068 4844 26078 4900
rect 0 4732 1708 4788
rect 1764 4732 2492 4788
rect 2548 4732 2558 4788
rect 19618 4732 19628 4788
rect 19684 4732 19694 4788
rect 0 4704 400 4732
rect 8006 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8290 4732
rect 14810 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15094 4732
rect 21614 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21898 4732
rect 28418 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28702 4732
rect 20066 4620 20076 4676
rect 20132 4620 20636 4676
rect 20692 4620 20702 4676
rect 23202 4396 23212 4452
rect 23268 4396 25228 4452
rect 25284 4396 25294 4452
rect 24210 4284 24220 4340
rect 24276 4284 25340 4340
rect 25396 4284 25406 4340
rect 11666 4172 11676 4228
rect 11732 4172 23212 4228
rect 23268 4172 23278 4228
rect 24882 4172 24892 4228
rect 24948 4172 26908 4228
rect 26964 4172 26974 4228
rect 11554 4060 11564 4116
rect 11620 4060 12180 4116
rect 18050 4060 18060 4116
rect 18116 4060 18284 4116
rect 18340 4060 19292 4116
rect 19348 4060 19358 4116
rect 23650 4060 23660 4116
rect 23716 4060 26460 4116
rect 26516 4060 26526 4116
rect 12124 4004 12180 4060
rect 12114 3948 12124 4004
rect 12180 3948 12190 4004
rect 20514 3948 20524 4004
rect 20580 3948 23996 4004
rect 24052 3948 24062 4004
rect 4604 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4888 3948
rect 11408 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11692 3948
rect 18212 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18496 3948
rect 25016 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25300 3948
rect 20626 3836 20636 3892
rect 20692 3836 23660 3892
rect 23716 3836 23726 3892
rect 13010 3724 13020 3780
rect 13076 3724 20300 3780
rect 20356 3724 22316 3780
rect 22372 3724 22382 3780
rect 22754 3724 22764 3780
rect 22820 3724 24892 3780
rect 24948 3724 24958 3780
rect 19730 3612 19740 3668
rect 19796 3612 21980 3668
rect 22036 3612 22046 3668
rect 23202 3612 23212 3668
rect 23268 3612 27916 3668
rect 27972 3612 27982 3668
rect 8754 3500 8764 3556
rect 8820 3500 9660 3556
rect 9716 3500 9726 3556
rect 10994 3500 11004 3556
rect 11060 3500 11788 3556
rect 11844 3500 11854 3556
rect 23202 3500 23212 3556
rect 23268 3500 24108 3556
rect 24164 3500 24174 3556
rect 25778 3500 25788 3556
rect 25844 3500 27580 3556
rect 27636 3500 27646 3556
rect 4946 3388 4956 3444
rect 5012 3388 5740 3444
rect 5796 3388 5806 3444
rect 6402 3388 6412 3444
rect 6468 3388 12124 3444
rect 12180 3388 12190 3444
rect 17500 3388 19404 3444
rect 19460 3388 19470 3444
rect 19842 3388 19852 3444
rect 19908 3388 19964 3444
rect 20020 3388 20030 3444
rect 20962 3388 20972 3444
rect 21028 3388 23324 3444
rect 23380 3388 23390 3444
rect 26114 3388 26124 3444
rect 26180 3388 27132 3444
rect 27188 3388 27198 3444
rect 17500 3220 17556 3388
rect 21410 3276 21420 3332
rect 21476 3276 23772 3332
rect 23828 3276 23838 3332
rect 8372 3164 10220 3220
rect 10276 3164 10286 3220
rect 17490 3164 17500 3220
rect 17556 3164 17566 3220
rect 19170 3164 19180 3220
rect 19236 3164 20748 3220
rect 20804 3164 20814 3220
rect 8006 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8290 3164
rect 8372 2996 8428 3164
rect 14810 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15094 3164
rect 21614 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21898 3164
rect 28418 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28702 3164
rect 17714 3052 17724 3108
rect 17780 3052 17948 3108
rect 18004 3052 19292 3108
rect 19348 3052 19358 3108
rect 8082 2940 8092 2996
rect 8148 2940 8428 2996
rect 11666 2940 11676 2996
rect 11732 2940 12572 2996
rect 12628 2940 12638 2996
rect 22642 2940 22652 2996
rect 22708 2940 23436 2996
rect 23492 2940 25340 2996
rect 25396 2940 25406 2996
rect 25666 2940 25676 2996
rect 25732 2940 26236 2996
rect 26292 2940 26302 2996
rect 18386 2828 18396 2884
rect 18452 2828 23660 2884
rect 23716 2828 23726 2884
rect 24658 2828 24668 2884
rect 24724 2828 25452 2884
rect 25508 2828 27356 2884
rect 27412 2828 27422 2884
rect 4274 2716 4284 2772
rect 4340 2716 6188 2772
rect 6244 2716 6254 2772
rect 9986 2716 9996 2772
rect 10052 2716 10556 2772
rect 10612 2716 10622 2772
rect 17378 2716 17388 2772
rect 17444 2716 19852 2772
rect 19908 2716 22876 2772
rect 22932 2716 22942 2772
rect 24098 2716 24108 2772
rect 24164 2716 25900 2772
rect 25956 2716 26684 2772
rect 26740 2716 26750 2772
rect 11228 2604 13580 2660
rect 13636 2604 13646 2660
rect 16258 2604 16268 2660
rect 16324 2604 17052 2660
rect 17108 2604 17612 2660
rect 17668 2604 17678 2660
rect 22418 2604 22428 2660
rect 22484 2604 28140 2660
rect 28196 2604 28206 2660
rect 11228 2436 11284 2604
rect 12898 2492 12908 2548
rect 12964 2492 14364 2548
rect 14420 2492 14430 2548
rect 11218 2380 11228 2436
rect 11284 2380 11294 2436
rect 4604 2324 4614 2380
rect 4670 2324 4718 2380
rect 4774 2324 4822 2380
rect 4878 2324 4888 2380
rect 11408 2324 11418 2380
rect 11474 2324 11522 2380
rect 11578 2324 11626 2380
rect 11682 2324 11692 2380
rect 18212 2324 18222 2380
rect 18278 2324 18326 2380
rect 18382 2324 18430 2380
rect 18486 2324 18496 2380
rect 25016 2324 25026 2380
rect 25082 2324 25130 2380
rect 25186 2324 25234 2380
rect 25290 2324 25300 2380
rect 3602 2156 3612 2212
rect 3668 2156 6300 2212
rect 6356 2156 6366 2212
rect 10770 2156 10780 2212
rect 10836 2156 10948 2212
rect 12338 2156 12348 2212
rect 12404 2156 12796 2212
rect 12852 2156 14140 2212
rect 14196 2156 14206 2212
rect 18050 2156 18060 2212
rect 18116 2156 18172 2212
rect 18228 2156 18238 2212
rect 20066 2156 20076 2212
rect 20132 2156 20748 2212
rect 20804 2156 20814 2212
rect 21410 2156 21420 2212
rect 21476 2156 21486 2212
rect 2380 1820 3276 1876
rect 3332 1820 3948 1876
rect 4004 1820 4014 1876
rect 4722 1820 4732 1876
rect 4788 1820 5404 1876
rect 5460 1820 5470 1876
rect 2380 1764 2436 1820
rect 10892 1764 10948 2156
rect 21420 2100 21476 2156
rect 18946 2044 18956 2100
rect 19012 2044 21476 2100
rect 24210 2044 24220 2100
rect 24276 2044 27580 2100
rect 27636 2044 27646 2100
rect 13458 1932 13468 1988
rect 13524 1932 14140 1988
rect 14196 1932 14700 1988
rect 14756 1932 14766 1988
rect 19506 1932 19516 1988
rect 19572 1932 20524 1988
rect 20580 1932 20590 1988
rect 21522 1932 21532 1988
rect 21588 1932 22428 1988
rect 22484 1932 22494 1988
rect 23538 1932 23548 1988
rect 23604 1932 25676 1988
rect 25732 1932 25742 1988
rect 16146 1820 16156 1876
rect 16212 1820 16940 1876
rect 16996 1820 17006 1876
rect 18498 1820 18508 1876
rect 18564 1820 18844 1876
rect 18900 1820 18910 1876
rect 19394 1820 19404 1876
rect 19460 1820 19628 1876
rect 19684 1820 19694 1876
rect 24322 1820 24332 1876
rect 24388 1820 27356 1876
rect 27412 1820 27422 1876
rect 2370 1708 2380 1764
rect 2436 1708 2446 1764
rect 10882 1708 10892 1764
rect 10948 1708 10958 1764
rect 24882 1708 24892 1764
rect 24948 1708 26908 1764
rect 26964 1708 26974 1764
rect 8006 1540 8016 1596
rect 8072 1540 8120 1596
rect 8176 1540 8224 1596
rect 8280 1540 8290 1596
rect 14810 1540 14820 1596
rect 14876 1540 14924 1596
rect 14980 1540 15028 1596
rect 15084 1540 15094 1596
rect 21614 1540 21624 1596
rect 21680 1540 21728 1596
rect 21784 1540 21832 1596
rect 21888 1540 21898 1596
rect 28418 1540 28428 1596
rect 28484 1540 28532 1596
rect 28588 1540 28636 1596
rect 28692 1540 28702 1596
rect 22418 476 22428 532
rect 22484 476 23212 532
rect 23268 476 23278 532
<< via3 >>
rect 4614 118356 4670 118412
rect 4718 118356 4774 118412
rect 4822 118356 4878 118412
rect 11418 118356 11474 118412
rect 11522 118356 11578 118412
rect 11626 118356 11682 118412
rect 18222 118356 18278 118412
rect 18326 118356 18382 118412
rect 18430 118356 18486 118412
rect 25026 118356 25082 118412
rect 25130 118356 25186 118412
rect 25234 118356 25290 118412
rect 8016 117572 8072 117628
rect 8120 117572 8176 117628
rect 8224 117572 8280 117628
rect 14820 117572 14876 117628
rect 14924 117572 14980 117628
rect 15028 117572 15084 117628
rect 21624 117572 21680 117628
rect 21728 117572 21784 117628
rect 21832 117572 21888 117628
rect 28428 117572 28484 117628
rect 28532 117572 28588 117628
rect 28636 117572 28692 117628
rect 4614 116788 4670 116844
rect 4718 116788 4774 116844
rect 4822 116788 4878 116844
rect 11418 116788 11474 116844
rect 11522 116788 11578 116844
rect 11626 116788 11682 116844
rect 18222 116788 18278 116844
rect 18326 116788 18382 116844
rect 18430 116788 18486 116844
rect 25026 116788 25082 116844
rect 25130 116788 25186 116844
rect 25234 116788 25290 116844
rect 8016 116004 8072 116060
rect 8120 116004 8176 116060
rect 8224 116004 8280 116060
rect 14820 116004 14876 116060
rect 14924 116004 14980 116060
rect 15028 116004 15084 116060
rect 21624 116004 21680 116060
rect 21728 116004 21784 116060
rect 21832 116004 21888 116060
rect 28428 116004 28484 116060
rect 28532 116004 28588 116060
rect 28636 116004 28692 116060
rect 4614 115220 4670 115276
rect 4718 115220 4774 115276
rect 4822 115220 4878 115276
rect 11418 115220 11474 115276
rect 11522 115220 11578 115276
rect 11626 115220 11682 115276
rect 18222 115220 18278 115276
rect 18326 115220 18382 115276
rect 18430 115220 18486 115276
rect 25026 115220 25082 115276
rect 25130 115220 25186 115276
rect 25234 115220 25290 115276
rect 8016 114436 8072 114492
rect 8120 114436 8176 114492
rect 8224 114436 8280 114492
rect 14820 114436 14876 114492
rect 14924 114436 14980 114492
rect 15028 114436 15084 114492
rect 21624 114436 21680 114492
rect 21728 114436 21784 114492
rect 21832 114436 21888 114492
rect 28428 114436 28484 114492
rect 28532 114436 28588 114492
rect 28636 114436 28692 114492
rect 4614 113652 4670 113708
rect 4718 113652 4774 113708
rect 4822 113652 4878 113708
rect 11418 113652 11474 113708
rect 11522 113652 11578 113708
rect 11626 113652 11682 113708
rect 18222 113652 18278 113708
rect 18326 113652 18382 113708
rect 18430 113652 18486 113708
rect 25026 113652 25082 113708
rect 25130 113652 25186 113708
rect 25234 113652 25290 113708
rect 8016 112868 8072 112924
rect 8120 112868 8176 112924
rect 8224 112868 8280 112924
rect 14820 112868 14876 112924
rect 14924 112868 14980 112924
rect 15028 112868 15084 112924
rect 21624 112868 21680 112924
rect 21728 112868 21784 112924
rect 21832 112868 21888 112924
rect 28428 112868 28484 112924
rect 28532 112868 28588 112924
rect 28636 112868 28692 112924
rect 4614 112084 4670 112140
rect 4718 112084 4774 112140
rect 4822 112084 4878 112140
rect 11418 112084 11474 112140
rect 11522 112084 11578 112140
rect 11626 112084 11682 112140
rect 18222 112084 18278 112140
rect 18326 112084 18382 112140
rect 18430 112084 18486 112140
rect 25026 112084 25082 112140
rect 25130 112084 25186 112140
rect 25234 112084 25290 112140
rect 8016 111300 8072 111356
rect 8120 111300 8176 111356
rect 8224 111300 8280 111356
rect 14820 111300 14876 111356
rect 14924 111300 14980 111356
rect 15028 111300 15084 111356
rect 21624 111300 21680 111356
rect 21728 111300 21784 111356
rect 21832 111300 21888 111356
rect 28428 111300 28484 111356
rect 28532 111300 28588 111356
rect 28636 111300 28692 111356
rect 4614 110516 4670 110572
rect 4718 110516 4774 110572
rect 4822 110516 4878 110572
rect 11418 110516 11474 110572
rect 11522 110516 11578 110572
rect 11626 110516 11682 110572
rect 18222 110516 18278 110572
rect 18326 110516 18382 110572
rect 18430 110516 18486 110572
rect 25026 110516 25082 110572
rect 25130 110516 25186 110572
rect 25234 110516 25290 110572
rect 8016 109732 8072 109788
rect 8120 109732 8176 109788
rect 8224 109732 8280 109788
rect 14820 109732 14876 109788
rect 14924 109732 14980 109788
rect 15028 109732 15084 109788
rect 21624 109732 21680 109788
rect 21728 109732 21784 109788
rect 21832 109732 21888 109788
rect 28428 109732 28484 109788
rect 28532 109732 28588 109788
rect 28636 109732 28692 109788
rect 4614 108948 4670 109004
rect 4718 108948 4774 109004
rect 4822 108948 4878 109004
rect 11418 108948 11474 109004
rect 11522 108948 11578 109004
rect 11626 108948 11682 109004
rect 18222 108948 18278 109004
rect 18326 108948 18382 109004
rect 18430 108948 18486 109004
rect 25026 108948 25082 109004
rect 25130 108948 25186 109004
rect 25234 108948 25290 109004
rect 8016 108164 8072 108220
rect 8120 108164 8176 108220
rect 8224 108164 8280 108220
rect 14820 108164 14876 108220
rect 14924 108164 14980 108220
rect 15028 108164 15084 108220
rect 21624 108164 21680 108220
rect 21728 108164 21784 108220
rect 21832 108164 21888 108220
rect 28428 108164 28484 108220
rect 28532 108164 28588 108220
rect 28636 108164 28692 108220
rect 4614 107380 4670 107436
rect 4718 107380 4774 107436
rect 4822 107380 4878 107436
rect 11418 107380 11474 107436
rect 11522 107380 11578 107436
rect 11626 107380 11682 107436
rect 18222 107380 18278 107436
rect 18326 107380 18382 107436
rect 18430 107380 18486 107436
rect 25026 107380 25082 107436
rect 25130 107380 25186 107436
rect 25234 107380 25290 107436
rect 8016 106596 8072 106652
rect 8120 106596 8176 106652
rect 8224 106596 8280 106652
rect 14820 106596 14876 106652
rect 14924 106596 14980 106652
rect 15028 106596 15084 106652
rect 21624 106596 21680 106652
rect 21728 106596 21784 106652
rect 21832 106596 21888 106652
rect 28428 106596 28484 106652
rect 28532 106596 28588 106652
rect 28636 106596 28692 106652
rect 4614 105812 4670 105868
rect 4718 105812 4774 105868
rect 4822 105812 4878 105868
rect 11418 105812 11474 105868
rect 11522 105812 11578 105868
rect 11626 105812 11682 105868
rect 18222 105812 18278 105868
rect 18326 105812 18382 105868
rect 18430 105812 18486 105868
rect 25026 105812 25082 105868
rect 25130 105812 25186 105868
rect 25234 105812 25290 105868
rect 24444 105644 24500 105700
rect 8016 105028 8072 105084
rect 8120 105028 8176 105084
rect 8224 105028 8280 105084
rect 14820 105028 14876 105084
rect 14924 105028 14980 105084
rect 15028 105028 15084 105084
rect 21624 105028 21680 105084
rect 21728 105028 21784 105084
rect 21832 105028 21888 105084
rect 28428 105028 28484 105084
rect 28532 105028 28588 105084
rect 28636 105028 28692 105084
rect 8540 104300 8596 104356
rect 4614 104244 4670 104300
rect 4718 104244 4774 104300
rect 4822 104244 4878 104300
rect 11418 104244 11474 104300
rect 11522 104244 11578 104300
rect 11626 104244 11682 104300
rect 18222 104244 18278 104300
rect 18326 104244 18382 104300
rect 18430 104244 18486 104300
rect 25026 104244 25082 104300
rect 25130 104244 25186 104300
rect 25234 104244 25290 104300
rect 8540 103740 8596 103796
rect 9436 103740 9492 103796
rect 8016 103460 8072 103516
rect 8120 103460 8176 103516
rect 8224 103460 8280 103516
rect 14820 103460 14876 103516
rect 14924 103460 14980 103516
rect 15028 103460 15084 103516
rect 21624 103460 21680 103516
rect 21728 103460 21784 103516
rect 21832 103460 21888 103516
rect 28428 103460 28484 103516
rect 28532 103460 28588 103516
rect 28636 103460 28692 103516
rect 9660 102732 9716 102788
rect 4614 102676 4670 102732
rect 4718 102676 4774 102732
rect 4822 102676 4878 102732
rect 11418 102676 11474 102732
rect 11522 102676 11578 102732
rect 11626 102676 11682 102732
rect 18222 102676 18278 102732
rect 18326 102676 18382 102732
rect 18430 102676 18486 102732
rect 25026 102676 25082 102732
rect 25130 102676 25186 102732
rect 25234 102676 25290 102732
rect 6524 102508 6580 102564
rect 9436 102172 9492 102228
rect 8016 101892 8072 101948
rect 8120 101892 8176 101948
rect 8224 101892 8280 101948
rect 14820 101892 14876 101948
rect 14924 101892 14980 101948
rect 15028 101892 15084 101948
rect 21624 101892 21680 101948
rect 21728 101892 21784 101948
rect 21832 101892 21888 101948
rect 28428 101892 28484 101948
rect 28532 101892 28588 101948
rect 28636 101892 28692 101948
rect 4614 101108 4670 101164
rect 4718 101108 4774 101164
rect 4822 101108 4878 101164
rect 11418 101108 11474 101164
rect 11522 101108 11578 101164
rect 11626 101108 11682 101164
rect 18222 101108 18278 101164
rect 18326 101108 18382 101164
rect 18430 101108 18486 101164
rect 25026 101108 25082 101164
rect 25130 101108 25186 101164
rect 25234 101108 25290 101164
rect 8016 100324 8072 100380
rect 8120 100324 8176 100380
rect 8224 100324 8280 100380
rect 14820 100324 14876 100380
rect 14924 100324 14980 100380
rect 15028 100324 15084 100380
rect 21624 100324 21680 100380
rect 21728 100324 21784 100380
rect 21832 100324 21888 100380
rect 28428 100324 28484 100380
rect 28532 100324 28588 100380
rect 28636 100324 28692 100380
rect 4614 99540 4670 99596
rect 4718 99540 4774 99596
rect 4822 99540 4878 99596
rect 11418 99540 11474 99596
rect 11522 99540 11578 99596
rect 11626 99540 11682 99596
rect 18222 99540 18278 99596
rect 18326 99540 18382 99596
rect 18430 99540 18486 99596
rect 25026 99540 25082 99596
rect 25130 99540 25186 99596
rect 25234 99540 25290 99596
rect 8016 98756 8072 98812
rect 8120 98756 8176 98812
rect 8224 98756 8280 98812
rect 14820 98756 14876 98812
rect 14924 98756 14980 98812
rect 15028 98756 15084 98812
rect 21624 98756 21680 98812
rect 21728 98756 21784 98812
rect 21832 98756 21888 98812
rect 28428 98756 28484 98812
rect 28532 98756 28588 98812
rect 28636 98756 28692 98812
rect 17948 98700 18004 98756
rect 18060 98476 18116 98532
rect 4614 97972 4670 98028
rect 4718 97972 4774 98028
rect 4822 97972 4878 98028
rect 11418 97972 11474 98028
rect 11522 97972 11578 98028
rect 11626 97972 11682 98028
rect 18222 97972 18278 98028
rect 18326 97972 18382 98028
rect 18430 97972 18486 98028
rect 25026 97972 25082 98028
rect 25130 97972 25186 98028
rect 25234 97972 25290 98028
rect 15260 97692 15316 97748
rect 18060 97580 18116 97636
rect 24444 97356 24500 97412
rect 14252 97244 14308 97300
rect 8016 97188 8072 97244
rect 8120 97188 8176 97244
rect 8224 97188 8280 97244
rect 14820 97188 14876 97244
rect 14924 97188 14980 97244
rect 15028 97188 15084 97244
rect 21624 97188 21680 97244
rect 21728 97188 21784 97244
rect 21832 97188 21888 97244
rect 28428 97188 28484 97244
rect 28532 97188 28588 97244
rect 28636 97188 28692 97244
rect 14028 97132 14084 97188
rect 14364 97132 14420 97188
rect 9660 97020 9716 97076
rect 13916 96908 13972 96964
rect 14252 96908 14308 96964
rect 17948 96796 18004 96852
rect 4614 96404 4670 96460
rect 4718 96404 4774 96460
rect 4822 96404 4878 96460
rect 11418 96404 11474 96460
rect 11522 96404 11578 96460
rect 11626 96404 11682 96460
rect 18222 96404 18278 96460
rect 18326 96404 18382 96460
rect 18430 96404 18486 96460
rect 25026 96404 25082 96460
rect 25130 96404 25186 96460
rect 25234 96404 25290 96460
rect 10892 96348 10948 96404
rect 14028 96348 14084 96404
rect 14588 96124 14644 96180
rect 10892 95788 10948 95844
rect 14364 95788 14420 95844
rect 8016 95620 8072 95676
rect 8120 95620 8176 95676
rect 8224 95620 8280 95676
rect 14820 95620 14876 95676
rect 14924 95620 14980 95676
rect 15028 95620 15084 95676
rect 21624 95620 21680 95676
rect 21728 95620 21784 95676
rect 21832 95620 21888 95676
rect 28428 95620 28484 95676
rect 28532 95620 28588 95676
rect 28636 95620 28692 95676
rect 14588 95228 14644 95284
rect 13916 95116 13972 95172
rect 19068 95116 19124 95172
rect 4614 94836 4670 94892
rect 4718 94836 4774 94892
rect 4822 94836 4878 94892
rect 11418 94836 11474 94892
rect 11522 94836 11578 94892
rect 11626 94836 11682 94892
rect 18222 94836 18278 94892
rect 18326 94836 18382 94892
rect 18430 94836 18486 94892
rect 25026 94836 25082 94892
rect 25130 94836 25186 94892
rect 25234 94836 25290 94892
rect 19740 94668 19796 94724
rect 6524 94556 6580 94612
rect 19068 94444 19124 94500
rect 15372 94220 15428 94276
rect 8016 94052 8072 94108
rect 8120 94052 8176 94108
rect 8224 94052 8280 94108
rect 14820 94052 14876 94108
rect 14924 94052 14980 94108
rect 15028 94052 15084 94108
rect 21624 94052 21680 94108
rect 21728 94052 21784 94108
rect 21832 94052 21888 94108
rect 15260 93996 15316 94052
rect 28428 94052 28484 94108
rect 28532 94052 28588 94108
rect 28636 94052 28692 94108
rect 15596 93884 15652 93940
rect 15260 93772 15316 93828
rect 20524 93660 20580 93716
rect 23100 93548 23156 93604
rect 4614 93268 4670 93324
rect 4718 93268 4774 93324
rect 4822 93268 4878 93324
rect 11418 93268 11474 93324
rect 11522 93268 11578 93324
rect 11626 93268 11682 93324
rect 18222 93268 18278 93324
rect 18326 93268 18382 93324
rect 18430 93268 18486 93324
rect 25026 93268 25082 93324
rect 25130 93268 25186 93324
rect 25234 93268 25290 93324
rect 15596 93212 15652 93268
rect 20860 92764 20916 92820
rect 20188 92652 20244 92708
rect 8016 92484 8072 92540
rect 8120 92484 8176 92540
rect 8224 92484 8280 92540
rect 14820 92484 14876 92540
rect 14924 92484 14980 92540
rect 15028 92484 15084 92540
rect 21624 92484 21680 92540
rect 21728 92484 21784 92540
rect 21832 92484 21888 92540
rect 28428 92484 28484 92540
rect 28532 92484 28588 92540
rect 28636 92484 28692 92540
rect 17836 92316 17892 92372
rect 4614 91700 4670 91756
rect 4718 91700 4774 91756
rect 4822 91700 4878 91756
rect 11418 91700 11474 91756
rect 11522 91700 11578 91756
rect 11626 91700 11682 91756
rect 18222 91700 18278 91756
rect 18326 91700 18382 91756
rect 18430 91700 18486 91756
rect 25026 91700 25082 91756
rect 25130 91700 25186 91756
rect 25234 91700 25290 91756
rect 22988 91644 23044 91700
rect 25564 91644 25620 91700
rect 22876 91532 22932 91588
rect 15372 91420 15428 91476
rect 8016 90916 8072 90972
rect 8120 90916 8176 90972
rect 8224 90916 8280 90972
rect 14820 90916 14876 90972
rect 14924 90916 14980 90972
rect 15028 90916 15084 90972
rect 21624 90916 21680 90972
rect 21728 90916 21784 90972
rect 21832 90916 21888 90972
rect 28428 90916 28484 90972
rect 28532 90916 28588 90972
rect 28636 90916 28692 90972
rect 10892 90636 10948 90692
rect 4614 90132 4670 90188
rect 4718 90132 4774 90188
rect 4822 90132 4878 90188
rect 11418 90132 11474 90188
rect 11522 90132 11578 90188
rect 11626 90132 11682 90188
rect 18222 90132 18278 90188
rect 18326 90132 18382 90188
rect 18430 90132 18486 90188
rect 25026 90132 25082 90188
rect 25130 90132 25186 90188
rect 25234 90132 25290 90188
rect 22876 89964 22932 90020
rect 8016 89348 8072 89404
rect 8120 89348 8176 89404
rect 8224 89348 8280 89404
rect 14820 89348 14876 89404
rect 14924 89348 14980 89404
rect 15028 89348 15084 89404
rect 21624 89348 21680 89404
rect 21728 89348 21784 89404
rect 21832 89348 21888 89404
rect 28428 89348 28484 89404
rect 28532 89348 28588 89404
rect 28636 89348 28692 89404
rect 15372 89180 15428 89236
rect 22988 89180 23044 89236
rect 15708 89068 15764 89124
rect 19740 88732 19796 88788
rect 4614 88564 4670 88620
rect 4718 88564 4774 88620
rect 4822 88564 4878 88620
rect 11418 88564 11474 88620
rect 11522 88564 11578 88620
rect 11626 88564 11682 88620
rect 18222 88564 18278 88620
rect 18326 88564 18382 88620
rect 18430 88564 18486 88620
rect 25026 88564 25082 88620
rect 25130 88564 25186 88620
rect 25234 88564 25290 88620
rect 15484 88060 15540 88116
rect 3388 87948 3444 88004
rect 17836 87948 17892 88004
rect 8016 87780 8072 87836
rect 8120 87780 8176 87836
rect 8224 87780 8280 87836
rect 14820 87780 14876 87836
rect 14924 87780 14980 87836
rect 15028 87780 15084 87836
rect 21624 87780 21680 87836
rect 21728 87780 21784 87836
rect 21832 87780 21888 87836
rect 28428 87780 28484 87836
rect 28532 87780 28588 87836
rect 28636 87780 28692 87836
rect 15596 87612 15652 87668
rect 4614 86996 4670 87052
rect 4718 86996 4774 87052
rect 4822 86996 4878 87052
rect 11418 86996 11474 87052
rect 11522 86996 11578 87052
rect 11626 86996 11682 87052
rect 18222 86996 18278 87052
rect 18326 86996 18382 87052
rect 18430 86996 18486 87052
rect 25026 86996 25082 87052
rect 25130 86996 25186 87052
rect 25234 86996 25290 87052
rect 15484 86268 15540 86324
rect 8016 86212 8072 86268
rect 8120 86212 8176 86268
rect 8224 86212 8280 86268
rect 14820 86212 14876 86268
rect 14924 86212 14980 86268
rect 15028 86212 15084 86268
rect 21624 86212 21680 86268
rect 21728 86212 21784 86268
rect 21832 86212 21888 86268
rect 28428 86212 28484 86268
rect 28532 86212 28588 86268
rect 28636 86212 28692 86268
rect 15708 85932 15764 85988
rect 4614 85428 4670 85484
rect 4718 85428 4774 85484
rect 4822 85428 4878 85484
rect 11418 85428 11474 85484
rect 11522 85428 11578 85484
rect 11626 85428 11682 85484
rect 18222 85428 18278 85484
rect 18326 85428 18382 85484
rect 18430 85428 18486 85484
rect 25026 85428 25082 85484
rect 25130 85428 25186 85484
rect 25234 85428 25290 85484
rect 8016 84644 8072 84700
rect 8120 84644 8176 84700
rect 8224 84644 8280 84700
rect 14820 84644 14876 84700
rect 14924 84644 14980 84700
rect 15028 84644 15084 84700
rect 21624 84644 21680 84700
rect 21728 84644 21784 84700
rect 21832 84644 21888 84700
rect 20748 84364 20804 84420
rect 28428 84644 28484 84700
rect 28532 84644 28588 84700
rect 28636 84644 28692 84700
rect 20188 83916 20244 83972
rect 4614 83860 4670 83916
rect 4718 83860 4774 83916
rect 4822 83860 4878 83916
rect 11418 83860 11474 83916
rect 11522 83860 11578 83916
rect 11626 83860 11682 83916
rect 18222 83860 18278 83916
rect 18326 83860 18382 83916
rect 18430 83860 18486 83916
rect 25564 83916 25620 83972
rect 25026 83860 25082 83916
rect 25130 83860 25186 83916
rect 25234 83860 25290 83916
rect 20748 83692 20804 83748
rect 8016 83076 8072 83132
rect 8120 83076 8176 83132
rect 8224 83076 8280 83132
rect 14820 83076 14876 83132
rect 14924 83076 14980 83132
rect 15028 83076 15084 83132
rect 21624 83076 21680 83132
rect 21728 83076 21784 83132
rect 21832 83076 21888 83132
rect 28428 83076 28484 83132
rect 28532 83076 28588 83132
rect 28636 83076 28692 83132
rect 20860 83020 20916 83076
rect 28028 82796 28084 82852
rect 15708 82684 15764 82740
rect 4614 82292 4670 82348
rect 4718 82292 4774 82348
rect 4822 82292 4878 82348
rect 11418 82292 11474 82348
rect 11522 82292 11578 82348
rect 11626 82292 11682 82348
rect 18222 82292 18278 82348
rect 18326 82292 18382 82348
rect 18430 82292 18486 82348
rect 25026 82292 25082 82348
rect 25130 82292 25186 82348
rect 25234 82292 25290 82348
rect 8016 81508 8072 81564
rect 8120 81508 8176 81564
rect 8224 81508 8280 81564
rect 14820 81508 14876 81564
rect 14924 81508 14980 81564
rect 15028 81508 15084 81564
rect 21624 81508 21680 81564
rect 21728 81508 21784 81564
rect 21832 81508 21888 81564
rect 28428 81508 28484 81564
rect 28532 81508 28588 81564
rect 28636 81508 28692 81564
rect 22204 81004 22260 81060
rect 12796 80892 12852 80948
rect 28028 80780 28084 80836
rect 4614 80724 4670 80780
rect 4718 80724 4774 80780
rect 4822 80724 4878 80780
rect 11418 80724 11474 80780
rect 11522 80724 11578 80780
rect 11626 80724 11682 80780
rect 18222 80724 18278 80780
rect 18326 80724 18382 80780
rect 18430 80724 18486 80780
rect 25026 80724 25082 80780
rect 25130 80724 25186 80780
rect 25234 80724 25290 80780
rect 14028 80556 14084 80612
rect 21196 80220 21252 80276
rect 26684 80108 26740 80164
rect 5068 79996 5124 80052
rect 8016 79940 8072 79996
rect 8120 79940 8176 79996
rect 8224 79940 8280 79996
rect 14820 79940 14876 79996
rect 14924 79940 14980 79996
rect 15028 79940 15084 79996
rect 21624 79940 21680 79996
rect 21728 79940 21784 79996
rect 21832 79940 21888 79996
rect 28428 79940 28484 79996
rect 28532 79940 28588 79996
rect 28636 79940 28692 79996
rect 14588 79660 14644 79716
rect 4614 79156 4670 79212
rect 4718 79156 4774 79212
rect 4822 79156 4878 79212
rect 11418 79156 11474 79212
rect 11522 79156 11578 79212
rect 11626 79156 11682 79212
rect 18222 79156 18278 79212
rect 18326 79156 18382 79212
rect 18430 79156 18486 79212
rect 25026 79156 25082 79212
rect 25130 79156 25186 79212
rect 25234 79156 25290 79212
rect 14252 79100 14308 79156
rect 14588 78988 14644 79044
rect 12572 78764 12628 78820
rect 14476 78764 14532 78820
rect 16044 78540 16100 78596
rect 14476 78428 14532 78484
rect 8016 78372 8072 78428
rect 8120 78372 8176 78428
rect 8224 78372 8280 78428
rect 14820 78372 14876 78428
rect 14924 78372 14980 78428
rect 15028 78372 15084 78428
rect 21624 78372 21680 78428
rect 21728 78372 21784 78428
rect 21832 78372 21888 78428
rect 28428 78372 28484 78428
rect 28532 78372 28588 78428
rect 28636 78372 28692 78428
rect 9100 77644 9156 77700
rect 4614 77588 4670 77644
rect 4718 77588 4774 77644
rect 4822 77588 4878 77644
rect 11418 77588 11474 77644
rect 11522 77588 11578 77644
rect 11626 77588 11682 77644
rect 18222 77588 18278 77644
rect 18326 77588 18382 77644
rect 18430 77588 18486 77644
rect 25026 77588 25082 77644
rect 25130 77588 25186 77644
rect 25234 77588 25290 77644
rect 21420 77308 21476 77364
rect 17836 77196 17892 77252
rect 22204 77084 22260 77140
rect 22652 77084 22708 77140
rect 8016 76804 8072 76860
rect 8120 76804 8176 76860
rect 8224 76804 8280 76860
rect 14820 76804 14876 76860
rect 14924 76804 14980 76860
rect 15028 76804 15084 76860
rect 21624 76804 21680 76860
rect 21728 76804 21784 76860
rect 21832 76804 21888 76860
rect 28428 76804 28484 76860
rect 28532 76804 28588 76860
rect 28636 76804 28692 76860
rect 14140 76412 14196 76468
rect 23884 76188 23940 76244
rect 26684 76188 26740 76244
rect 4614 76020 4670 76076
rect 4718 76020 4774 76076
rect 4822 76020 4878 76076
rect 11418 76020 11474 76076
rect 11522 76020 11578 76076
rect 11626 76020 11682 76076
rect 18222 76020 18278 76076
rect 18326 76020 18382 76076
rect 18430 76020 18486 76076
rect 25026 76020 25082 76076
rect 25130 76020 25186 76076
rect 25234 76020 25290 76076
rect 15260 75964 15316 76020
rect 13692 75404 13748 75460
rect 8016 75236 8072 75292
rect 8120 75236 8176 75292
rect 8224 75236 8280 75292
rect 14820 75236 14876 75292
rect 14924 75236 14980 75292
rect 15028 75236 15084 75292
rect 21624 75236 21680 75292
rect 21728 75236 21784 75292
rect 21832 75236 21888 75292
rect 26796 75180 26852 75236
rect 28428 75236 28484 75292
rect 28532 75236 28588 75292
rect 28636 75236 28692 75292
rect 11228 75068 11284 75124
rect 20860 75068 20916 75124
rect 24556 74956 24612 75012
rect 14364 74732 14420 74788
rect 19964 74732 20020 74788
rect 23212 74732 23268 74788
rect 23436 74732 23492 74788
rect 14028 74620 14084 74676
rect 4614 74452 4670 74508
rect 4718 74452 4774 74508
rect 4822 74452 4878 74508
rect 11418 74452 11474 74508
rect 11522 74452 11578 74508
rect 11626 74452 11682 74508
rect 18222 74452 18278 74508
rect 18326 74452 18382 74508
rect 18430 74452 18486 74508
rect 25026 74452 25082 74508
rect 25130 74452 25186 74508
rect 25234 74452 25290 74508
rect 23548 74396 23604 74452
rect 26572 74284 26628 74340
rect 26796 74284 26852 74340
rect 11228 74172 11284 74228
rect 12572 74060 12628 74116
rect 13804 73948 13860 74004
rect 23884 73836 23940 73892
rect 24556 73836 24612 73892
rect 8016 73668 8072 73724
rect 8120 73668 8176 73724
rect 8224 73668 8280 73724
rect 14820 73668 14876 73724
rect 14924 73668 14980 73724
rect 15028 73668 15084 73724
rect 21624 73668 21680 73724
rect 21728 73668 21784 73724
rect 21832 73668 21888 73724
rect 28428 73668 28484 73724
rect 28532 73668 28588 73724
rect 28636 73668 28692 73724
rect 19964 73612 20020 73668
rect 23548 73612 23604 73668
rect 18060 73388 18116 73444
rect 13916 73276 13972 73332
rect 15260 73164 15316 73220
rect 15820 73164 15876 73220
rect 4614 72884 4670 72940
rect 4718 72884 4774 72940
rect 4822 72884 4878 72940
rect 11418 72884 11474 72940
rect 11522 72884 11578 72940
rect 11626 72884 11682 72940
rect 18222 72884 18278 72940
rect 18326 72884 18382 72940
rect 18430 72884 18486 72940
rect 25026 72884 25082 72940
rect 25130 72884 25186 72940
rect 25234 72884 25290 72940
rect 16492 72828 16548 72884
rect 12796 72716 12852 72772
rect 23436 72716 23492 72772
rect 14476 72604 14532 72660
rect 21196 72492 21252 72548
rect 23212 72492 23268 72548
rect 22540 72380 22596 72436
rect 9100 72268 9156 72324
rect 15372 72268 15428 72324
rect 15596 72268 15652 72324
rect 12012 72156 12068 72212
rect 8016 72100 8072 72156
rect 8120 72100 8176 72156
rect 8224 72100 8280 72156
rect 14820 72100 14876 72156
rect 14924 72100 14980 72156
rect 15028 72100 15084 72156
rect 21624 72100 21680 72156
rect 21728 72100 21784 72156
rect 21832 72100 21888 72156
rect 28428 72100 28484 72156
rect 28532 72100 28588 72156
rect 28636 72100 28692 72156
rect 12012 71820 12068 71876
rect 15484 71820 15540 71876
rect 16492 71596 16548 71652
rect 14252 71484 14308 71540
rect 21420 71484 21476 71540
rect 22540 71484 22596 71540
rect 23324 71484 23380 71540
rect 4614 71316 4670 71372
rect 4718 71316 4774 71372
rect 4822 71316 4878 71372
rect 11418 71316 11474 71372
rect 11522 71316 11578 71372
rect 11626 71316 11682 71372
rect 18222 71316 18278 71372
rect 18326 71316 18382 71372
rect 18430 71316 18486 71372
rect 25026 71316 25082 71372
rect 25130 71316 25186 71372
rect 25234 71316 25290 71372
rect 23212 71260 23268 71316
rect 13916 71148 13972 71204
rect 14140 71148 14196 71204
rect 13692 70924 13748 70980
rect 15260 70924 15316 70980
rect 15484 70924 15540 70980
rect 16044 70924 16100 70980
rect 23324 70924 23380 70980
rect 13804 70812 13860 70868
rect 14140 70812 14196 70868
rect 15372 70812 15428 70868
rect 23436 70812 23492 70868
rect 14252 70700 14308 70756
rect 13244 70588 13300 70644
rect 14364 70588 14420 70644
rect 8016 70532 8072 70588
rect 8120 70532 8176 70588
rect 8224 70532 8280 70588
rect 15260 70588 15316 70644
rect 16044 70588 16100 70644
rect 20860 70588 20916 70644
rect 21980 70588 22036 70644
rect 14820 70532 14876 70588
rect 14924 70532 14980 70588
rect 15028 70532 15084 70588
rect 21624 70532 21680 70588
rect 21728 70532 21784 70588
rect 21832 70532 21888 70588
rect 28428 70532 28484 70588
rect 28532 70532 28588 70588
rect 28636 70532 28692 70588
rect 19740 70364 19796 70420
rect 23324 70028 23380 70084
rect 15484 69916 15540 69972
rect 9436 69804 9492 69860
rect 4614 69748 4670 69804
rect 4718 69748 4774 69804
rect 4822 69748 4878 69804
rect 11418 69748 11474 69804
rect 11522 69748 11578 69804
rect 11626 69748 11682 69804
rect 18222 69748 18278 69804
rect 18326 69748 18382 69804
rect 18430 69748 18486 69804
rect 25026 69748 25082 69804
rect 25130 69748 25186 69804
rect 25234 69748 25290 69804
rect 14140 69468 14196 69524
rect 13244 69356 13300 69412
rect 16940 69356 16996 69412
rect 9436 69132 9492 69188
rect 11228 69132 11284 69188
rect 14028 69132 14084 69188
rect 3836 69020 3892 69076
rect 8016 68964 8072 69020
rect 8120 68964 8176 69020
rect 8224 68964 8280 69020
rect 14820 68964 14876 69020
rect 14924 68964 14980 69020
rect 15028 68964 15084 69020
rect 21624 68964 21680 69020
rect 21728 68964 21784 69020
rect 21832 68964 21888 69020
rect 28428 68964 28484 69020
rect 28532 68964 28588 69020
rect 28636 68964 28692 69020
rect 15260 68908 15316 68964
rect 17164 68908 17220 68964
rect 18620 68796 18676 68852
rect 2492 68572 2548 68628
rect 14252 68572 14308 68628
rect 14588 68460 14644 68516
rect 3948 68348 4004 68404
rect 4396 68348 4452 68404
rect 4614 68180 4670 68236
rect 4718 68180 4774 68236
rect 4822 68180 4878 68236
rect 11418 68180 11474 68236
rect 11522 68180 11578 68236
rect 11626 68180 11682 68236
rect 18222 68180 18278 68236
rect 18326 68180 18382 68236
rect 18430 68180 18486 68236
rect 25026 68180 25082 68236
rect 25130 68180 25186 68236
rect 25234 68180 25290 68236
rect 20188 68124 20244 68180
rect 21420 68124 21476 68180
rect 22876 68012 22932 68068
rect 9660 67788 9716 67844
rect 10892 67676 10948 67732
rect 13916 67564 13972 67620
rect 19404 67564 19460 67620
rect 23324 67564 23380 67620
rect 8016 67396 8072 67452
rect 8120 67396 8176 67452
rect 8224 67396 8280 67452
rect 14820 67396 14876 67452
rect 14924 67396 14980 67452
rect 15028 67396 15084 67452
rect 21624 67396 21680 67452
rect 21728 67396 21784 67452
rect 21832 67396 21888 67452
rect 28428 67396 28484 67452
rect 28532 67396 28588 67452
rect 28636 67396 28692 67452
rect 13468 67116 13524 67172
rect 10780 67004 10836 67060
rect 17612 67004 17668 67060
rect 12796 66780 12852 66836
rect 4614 66612 4670 66668
rect 4718 66612 4774 66668
rect 4822 66612 4878 66668
rect 11418 66612 11474 66668
rect 11522 66612 11578 66668
rect 11626 66612 11682 66668
rect 18222 66612 18278 66668
rect 18326 66612 18382 66668
rect 18430 66612 18486 66668
rect 25026 66612 25082 66668
rect 25130 66612 25186 66668
rect 25234 66612 25290 66668
rect 13580 66444 13636 66500
rect 18956 65996 19012 66052
rect 8016 65828 8072 65884
rect 8120 65828 8176 65884
rect 8224 65828 8280 65884
rect 14820 65828 14876 65884
rect 14924 65828 14980 65884
rect 15028 65828 15084 65884
rect 21624 65828 21680 65884
rect 21728 65828 21784 65884
rect 21832 65828 21888 65884
rect 28428 65828 28484 65884
rect 28532 65828 28588 65884
rect 28636 65828 28692 65884
rect 14364 65772 14420 65828
rect 22428 65772 22484 65828
rect 22764 65660 22820 65716
rect 4172 65548 4228 65604
rect 13468 65548 13524 65604
rect 17948 65548 18004 65604
rect 19180 65548 19236 65604
rect 2492 65436 2548 65492
rect 23324 65100 23380 65156
rect 4614 65044 4670 65100
rect 4718 65044 4774 65100
rect 4822 65044 4878 65100
rect 11418 65044 11474 65100
rect 11522 65044 11578 65100
rect 11626 65044 11682 65100
rect 18222 65044 18278 65100
rect 18326 65044 18382 65100
rect 18430 65044 18486 65100
rect 25026 65044 25082 65100
rect 25130 65044 25186 65100
rect 25234 65044 25290 65100
rect 4172 64652 4228 64708
rect 17276 64652 17332 64708
rect 13468 64428 13524 64484
rect 13356 64316 13412 64372
rect 8016 64260 8072 64316
rect 8120 64260 8176 64316
rect 8224 64260 8280 64316
rect 14820 64260 14876 64316
rect 14924 64260 14980 64316
rect 15028 64260 15084 64316
rect 21624 64260 21680 64316
rect 21728 64260 21784 64316
rect 21832 64260 21888 64316
rect 28428 64260 28484 64316
rect 28532 64260 28588 64316
rect 28636 64260 28692 64316
rect 26684 64092 26740 64148
rect 9660 63644 9716 63700
rect 13580 63644 13636 63700
rect 15260 63644 15316 63700
rect 26684 63532 26740 63588
rect 4614 63476 4670 63532
rect 4718 63476 4774 63532
rect 4822 63476 4878 63532
rect 11418 63476 11474 63532
rect 11522 63476 11578 63532
rect 11626 63476 11682 63532
rect 18222 63476 18278 63532
rect 18326 63476 18382 63532
rect 18430 63476 18486 63532
rect 25026 63476 25082 63532
rect 25130 63476 25186 63532
rect 25234 63476 25290 63532
rect 22876 63420 22932 63476
rect 15260 63308 15316 63364
rect 17612 63196 17668 63252
rect 16268 63084 16324 63140
rect 17164 63084 17220 63140
rect 19068 63084 19124 63140
rect 3948 62860 4004 62916
rect 16268 62860 16324 62916
rect 8016 62692 8072 62748
rect 8120 62692 8176 62748
rect 8224 62692 8280 62748
rect 14820 62692 14876 62748
rect 14924 62692 14980 62748
rect 15028 62692 15084 62748
rect 21624 62692 21680 62748
rect 21728 62692 21784 62748
rect 21832 62692 21888 62748
rect 28428 62692 28484 62748
rect 28532 62692 28588 62748
rect 28636 62692 28692 62748
rect 11228 62636 11284 62692
rect 19740 62636 19796 62692
rect 14252 62524 14308 62580
rect 14476 62188 14532 62244
rect 17500 62188 17556 62244
rect 15372 62076 15428 62132
rect 4614 61908 4670 61964
rect 4718 61908 4774 61964
rect 4822 61908 4878 61964
rect 11418 61908 11474 61964
rect 11522 61908 11578 61964
rect 11626 61908 11682 61964
rect 14476 61852 14532 61908
rect 15932 61852 15988 61908
rect 18222 61908 18278 61964
rect 18326 61908 18382 61964
rect 18430 61908 18486 61964
rect 25026 61908 25082 61964
rect 25130 61908 25186 61964
rect 25234 61908 25290 61964
rect 15596 61740 15652 61796
rect 16940 61740 16996 61796
rect 4396 61628 4452 61684
rect 15372 61516 15428 61572
rect 15596 61516 15652 61572
rect 21420 61516 21476 61572
rect 13356 61404 13412 61460
rect 12796 61292 12852 61348
rect 8016 61124 8072 61180
rect 8120 61124 8176 61180
rect 8224 61124 8280 61180
rect 14820 61124 14876 61180
rect 14924 61124 14980 61180
rect 15028 61124 15084 61180
rect 21624 61124 21680 61180
rect 21728 61124 21784 61180
rect 21832 61124 21888 61180
rect 28428 61124 28484 61180
rect 28532 61124 28588 61180
rect 28636 61124 28692 61180
rect 16156 61068 16212 61124
rect 14476 60956 14532 61012
rect 11228 60844 11284 60900
rect 19404 60732 19460 60788
rect 20188 60732 20244 60788
rect 17164 60620 17220 60676
rect 3836 60508 3892 60564
rect 14252 60508 14308 60564
rect 15260 60508 15316 60564
rect 18620 60508 18676 60564
rect 17948 60396 18004 60452
rect 22428 60396 22484 60452
rect 4614 60340 4670 60396
rect 4718 60340 4774 60396
rect 4822 60340 4878 60396
rect 11418 60340 11474 60396
rect 11522 60340 11578 60396
rect 11626 60340 11682 60396
rect 18222 60340 18278 60396
rect 18326 60340 18382 60396
rect 18430 60340 18486 60396
rect 25026 60340 25082 60396
rect 25130 60340 25186 60396
rect 25234 60340 25290 60396
rect 22764 60284 22820 60340
rect 17276 60172 17332 60228
rect 14364 59948 14420 60004
rect 11788 59724 11844 59780
rect 14140 59724 14196 59780
rect 16156 59724 16212 59780
rect 19068 59612 19124 59668
rect 8016 59556 8072 59612
rect 8120 59556 8176 59612
rect 8224 59556 8280 59612
rect 14820 59556 14876 59612
rect 14924 59556 14980 59612
rect 15028 59556 15084 59612
rect 21624 59556 21680 59612
rect 21728 59556 21784 59612
rect 21832 59556 21888 59612
rect 28428 59556 28484 59612
rect 28532 59556 28588 59612
rect 28636 59556 28692 59612
rect 17500 59276 17556 59332
rect 14028 59164 14084 59220
rect 15932 59052 15988 59108
rect 10780 58828 10836 58884
rect 15260 58828 15316 58884
rect 22092 58828 22148 58884
rect 4614 58772 4670 58828
rect 4718 58772 4774 58828
rect 4822 58772 4878 58828
rect 11418 58772 11474 58828
rect 11522 58772 11578 58828
rect 11626 58772 11682 58828
rect 18222 58772 18278 58828
rect 18326 58772 18382 58828
rect 18430 58772 18486 58828
rect 25026 58772 25082 58828
rect 25130 58772 25186 58828
rect 25234 58772 25290 58828
rect 4172 58716 4228 58772
rect 15932 58716 15988 58772
rect 16380 58604 16436 58660
rect 13356 58492 13412 58548
rect 22316 58492 22372 58548
rect 16380 58380 16436 58436
rect 8876 58268 8932 58324
rect 9548 58268 9604 58324
rect 10556 58268 10612 58324
rect 2716 58156 2772 58212
rect 8016 57988 8072 58044
rect 8120 57988 8176 58044
rect 8224 57988 8280 58044
rect 14820 57988 14876 58044
rect 14924 57988 14980 58044
rect 15028 57988 15084 58044
rect 21624 57988 21680 58044
rect 21728 57988 21784 58044
rect 21832 57988 21888 58044
rect 28428 57988 28484 58044
rect 28532 57988 28588 58044
rect 28636 57988 28692 58044
rect 5852 57932 5908 57988
rect 12460 57932 12516 57988
rect 15260 57932 15316 57988
rect 23436 57932 23492 57988
rect 10108 57820 10164 57876
rect 13692 57820 13748 57876
rect 6300 57708 6356 57764
rect 3724 57260 3780 57316
rect 4614 57204 4670 57260
rect 4718 57204 4774 57260
rect 4822 57204 4878 57260
rect 13692 57260 13748 57316
rect 24108 57260 24164 57316
rect 11418 57204 11474 57260
rect 11522 57204 11578 57260
rect 11626 57204 11682 57260
rect 10780 57148 10836 57204
rect 14140 57148 14196 57204
rect 18222 57204 18278 57260
rect 18326 57204 18382 57260
rect 18430 57204 18486 57260
rect 25026 57204 25082 57260
rect 25130 57204 25186 57260
rect 25234 57204 25290 57260
rect 22204 57148 22260 57204
rect 24332 57148 24388 57204
rect 5404 56924 5460 56980
rect 25564 56924 25620 56980
rect 17052 56812 17108 56868
rect 3612 56700 3668 56756
rect 5292 56700 5348 56756
rect 5516 56700 5572 56756
rect 5852 56700 5908 56756
rect 16492 56700 16548 56756
rect 19516 56700 19572 56756
rect 4284 56476 4340 56532
rect 6636 56476 6692 56532
rect 8016 56420 8072 56476
rect 8120 56420 8176 56476
rect 8224 56420 8280 56476
rect 14820 56420 14876 56476
rect 14924 56420 14980 56476
rect 15028 56420 15084 56476
rect 21624 56420 21680 56476
rect 21728 56420 21784 56476
rect 21832 56420 21888 56476
rect 28428 56420 28484 56476
rect 28532 56420 28588 56476
rect 28636 56420 28692 56476
rect 16156 56364 16212 56420
rect 11116 56252 11172 56308
rect 22540 56252 22596 56308
rect 3836 56140 3892 56196
rect 10332 56140 10388 56196
rect 19068 56140 19124 56196
rect 26124 56140 26180 56196
rect 26348 56028 26404 56084
rect 17948 55916 18004 55972
rect 4614 55636 4670 55692
rect 4718 55636 4774 55692
rect 4822 55636 4878 55692
rect 4172 55580 4228 55636
rect 11788 55692 11844 55748
rect 11418 55636 11474 55692
rect 11522 55636 11578 55692
rect 11626 55636 11682 55692
rect 18222 55636 18278 55692
rect 18326 55636 18382 55692
rect 18430 55636 18486 55692
rect 25026 55636 25082 55692
rect 25130 55636 25186 55692
rect 25234 55636 25290 55692
rect 15484 55468 15540 55524
rect 21308 55468 21364 55524
rect 12460 55132 12516 55188
rect 17164 55132 17220 55188
rect 24108 55132 24164 55188
rect 10668 55020 10724 55076
rect 8016 54852 8072 54908
rect 8120 54852 8176 54908
rect 8224 54852 8280 54908
rect 14820 54852 14876 54908
rect 14924 54852 14980 54908
rect 15028 54852 15084 54908
rect 21624 54852 21680 54908
rect 21728 54852 21784 54908
rect 21832 54852 21888 54908
rect 28428 54852 28484 54908
rect 28532 54852 28588 54908
rect 28636 54852 28692 54908
rect 23212 54796 23268 54852
rect 24108 54796 24164 54852
rect 25788 54684 25844 54740
rect 2604 54572 2660 54628
rect 8540 54460 8596 54516
rect 6412 54348 6468 54404
rect 26684 54348 26740 54404
rect 10444 54236 10500 54292
rect 12908 54236 12964 54292
rect 19964 54236 20020 54292
rect 10332 54124 10388 54180
rect 23436 54124 23492 54180
rect 4614 54068 4670 54124
rect 4718 54068 4774 54124
rect 4822 54068 4878 54124
rect 11418 54068 11474 54124
rect 11522 54068 11578 54124
rect 11626 54068 11682 54124
rect 18222 54068 18278 54124
rect 18326 54068 18382 54124
rect 18430 54068 18486 54124
rect 25026 54068 25082 54124
rect 25130 54068 25186 54124
rect 25234 54068 25290 54124
rect 6412 54012 6468 54068
rect 6636 53788 6692 53844
rect 12908 53788 12964 53844
rect 19068 53676 19124 53732
rect 20300 53676 20356 53732
rect 4172 53564 4228 53620
rect 6300 53564 6356 53620
rect 8428 53564 8484 53620
rect 19852 53564 19908 53620
rect 26124 53564 26180 53620
rect 11004 53452 11060 53508
rect 16380 53452 16436 53508
rect 12012 53340 12068 53396
rect 8016 53284 8072 53340
rect 8120 53284 8176 53340
rect 8224 53284 8280 53340
rect 26684 53340 26740 53396
rect 14820 53284 14876 53340
rect 14924 53284 14980 53340
rect 15028 53284 15084 53340
rect 21624 53284 21680 53340
rect 21728 53284 21784 53340
rect 21832 53284 21888 53340
rect 28428 53284 28484 53340
rect 28532 53284 28588 53340
rect 28636 53284 28692 53340
rect 22540 53228 22596 53284
rect 8876 53116 8932 53172
rect 9548 53116 9604 53172
rect 21308 53116 21364 53172
rect 4396 53004 4452 53060
rect 5740 53004 5796 53060
rect 10108 53004 10164 53060
rect 11116 53004 11172 53060
rect 22428 53004 22484 53060
rect 10332 52892 10388 52948
rect 13692 52892 13748 52948
rect 18620 52892 18676 52948
rect 20188 52892 20244 52948
rect 2716 52668 2772 52724
rect 4614 52500 4670 52556
rect 4718 52500 4774 52556
rect 4822 52500 4878 52556
rect 17052 52556 17108 52612
rect 11418 52500 11474 52556
rect 11522 52500 11578 52556
rect 11626 52500 11682 52556
rect 18222 52500 18278 52556
rect 18326 52500 18382 52556
rect 18430 52500 18486 52556
rect 25026 52500 25082 52556
rect 25130 52500 25186 52556
rect 25234 52500 25290 52556
rect 5740 52444 5796 52500
rect 7420 52332 7476 52388
rect 13356 52332 13412 52388
rect 18844 52332 18900 52388
rect 2828 52220 2884 52276
rect 14140 52220 14196 52276
rect 17500 52220 17556 52276
rect 3500 52108 3556 52164
rect 11004 52108 11060 52164
rect 12908 52108 12964 52164
rect 7532 51996 7588 52052
rect 10108 51996 10164 52052
rect 15932 51996 15988 52052
rect 19292 51996 19348 52052
rect 22092 51996 22148 52052
rect 8016 51716 8072 51772
rect 8120 51716 8176 51772
rect 8224 51716 8280 51772
rect 14820 51716 14876 51772
rect 14924 51716 14980 51772
rect 15028 51716 15084 51772
rect 21624 51716 21680 51772
rect 21728 51716 21784 51772
rect 21832 51716 21888 51772
rect 28428 51716 28484 51772
rect 28532 51716 28588 51772
rect 28636 51716 28692 51772
rect 19292 51660 19348 51716
rect 5964 51548 6020 51604
rect 10780 51436 10836 51492
rect 18732 51436 18788 51492
rect 5852 51324 5908 51380
rect 6188 51212 6244 51268
rect 23212 51212 23268 51268
rect 3836 51100 3892 51156
rect 10780 51100 10836 51156
rect 22204 51100 22260 51156
rect 5292 50988 5348 51044
rect 4614 50932 4670 50988
rect 4718 50932 4774 50988
rect 4822 50932 4878 50988
rect 11418 50932 11474 50988
rect 11522 50932 11578 50988
rect 11626 50932 11682 50988
rect 18222 50932 18278 50988
rect 18326 50932 18382 50988
rect 18430 50932 18486 50988
rect 25026 50932 25082 50988
rect 25130 50932 25186 50988
rect 25234 50932 25290 50988
rect 5404 50876 5460 50932
rect 17948 50764 18004 50820
rect 19068 50652 19124 50708
rect 7420 50540 7476 50596
rect 22316 50540 22372 50596
rect 25788 50540 25844 50596
rect 14476 50428 14532 50484
rect 17724 50428 17780 50484
rect 20076 50428 20132 50484
rect 13916 50316 13972 50372
rect 19292 50316 19348 50372
rect 8428 50204 8484 50260
rect 8016 50148 8072 50204
rect 8120 50148 8176 50204
rect 8224 50148 8280 50204
rect 14820 50148 14876 50204
rect 14924 50148 14980 50204
rect 15028 50148 15084 50204
rect 21624 50148 21680 50204
rect 21728 50148 21784 50204
rect 21832 50148 21888 50204
rect 28428 50148 28484 50204
rect 28532 50148 28588 50204
rect 28636 50148 28692 50204
rect 6412 49980 6468 50036
rect 17500 49980 17556 50036
rect 12460 49868 12516 49924
rect 14364 49868 14420 49924
rect 2604 49756 2660 49812
rect 2828 49756 2884 49812
rect 21308 49756 21364 49812
rect 11004 49644 11060 49700
rect 18620 49644 18676 49700
rect 9772 49532 9828 49588
rect 4614 49364 4670 49420
rect 4718 49364 4774 49420
rect 4822 49364 4878 49420
rect 11418 49364 11474 49420
rect 11522 49364 11578 49420
rect 11626 49364 11682 49420
rect 18222 49364 18278 49420
rect 18326 49364 18382 49420
rect 18430 49364 18486 49420
rect 25026 49364 25082 49420
rect 25130 49364 25186 49420
rect 25234 49364 25290 49420
rect 10780 49308 10836 49364
rect 14364 49196 14420 49252
rect 3836 48972 3892 49028
rect 4172 48972 4228 49028
rect 11788 48972 11844 49028
rect 26348 48972 26404 49028
rect 14476 48860 14532 48916
rect 3612 48748 3668 48804
rect 6188 48748 6244 48804
rect 10444 48636 10500 48692
rect 14364 48636 14420 48692
rect 8016 48580 8072 48636
rect 8120 48580 8176 48636
rect 8224 48580 8280 48636
rect 4284 48524 4340 48580
rect 22428 48636 22484 48692
rect 24332 48636 24388 48692
rect 14820 48580 14876 48636
rect 14924 48580 14980 48636
rect 15028 48580 15084 48636
rect 21624 48580 21680 48636
rect 21728 48580 21784 48636
rect 21832 48580 21888 48636
rect 28428 48580 28484 48636
rect 28532 48580 28588 48636
rect 28636 48580 28692 48636
rect 17500 48524 17556 48580
rect 3724 48412 3780 48468
rect 7532 48412 7588 48468
rect 10444 48412 10500 48468
rect 11228 48412 11284 48468
rect 8540 48300 8596 48356
rect 17948 48300 18004 48356
rect 21308 48188 21364 48244
rect 10780 48076 10836 48132
rect 26124 48076 26180 48132
rect 4614 47796 4670 47852
rect 4718 47796 4774 47852
rect 4822 47796 4878 47852
rect 11418 47796 11474 47852
rect 11522 47796 11578 47852
rect 11626 47796 11682 47852
rect 10220 47740 10276 47796
rect 18222 47796 18278 47852
rect 18326 47796 18382 47852
rect 18430 47796 18486 47852
rect 25026 47796 25082 47852
rect 25130 47796 25186 47852
rect 25234 47796 25290 47852
rect 5516 47628 5572 47684
rect 9772 47628 9828 47684
rect 10556 47628 10612 47684
rect 12460 47628 12516 47684
rect 10780 47516 10836 47572
rect 13916 47516 13972 47572
rect 23436 47516 23492 47572
rect 3836 47404 3892 47460
rect 12012 47404 12068 47460
rect 17500 47404 17556 47460
rect 15932 47292 15988 47348
rect 10444 47180 10500 47236
rect 14364 47180 14420 47236
rect 17948 47180 18004 47236
rect 19964 47180 20020 47236
rect 10220 47068 10276 47124
rect 17164 47068 17220 47124
rect 17500 47068 17556 47124
rect 8016 47012 8072 47068
rect 8120 47012 8176 47068
rect 8224 47012 8280 47068
rect 9996 47012 10052 47068
rect 14820 47012 14876 47068
rect 14924 47012 14980 47068
rect 15028 47012 15084 47068
rect 11004 46956 11060 47012
rect 21624 47012 21680 47068
rect 21728 47012 21784 47068
rect 21832 47012 21888 47068
rect 28428 47012 28484 47068
rect 28532 47012 28588 47068
rect 28636 47012 28692 47068
rect 20748 46844 20804 46900
rect 22988 46844 23044 46900
rect 4060 46732 4116 46788
rect 5180 46732 5236 46788
rect 10332 46732 10388 46788
rect 13244 46732 13300 46788
rect 20076 46732 20132 46788
rect 4172 46620 4228 46676
rect 3164 46508 3220 46564
rect 5852 46508 5908 46564
rect 11228 46508 11284 46564
rect 23548 46508 23604 46564
rect 4614 46228 4670 46284
rect 4718 46228 4774 46284
rect 4822 46228 4878 46284
rect 11418 46228 11474 46284
rect 11522 46228 11578 46284
rect 11626 46228 11682 46284
rect 18222 46228 18278 46284
rect 18326 46228 18382 46284
rect 18430 46228 18486 46284
rect 25026 46228 25082 46284
rect 25130 46228 25186 46284
rect 25234 46228 25290 46284
rect 7868 46172 7924 46228
rect 22764 46172 22820 46228
rect 7084 46060 7140 46116
rect 17052 45948 17108 46004
rect 15260 45836 15316 45892
rect 2380 45724 2436 45780
rect 11004 45724 11060 45780
rect 14476 45612 14532 45668
rect 24780 45612 24836 45668
rect 6188 45500 6244 45556
rect 9660 45500 9716 45556
rect 11228 45500 11284 45556
rect 8016 45444 8072 45500
rect 8120 45444 8176 45500
rect 8224 45444 8280 45500
rect 14820 45444 14876 45500
rect 14924 45444 14980 45500
rect 15028 45444 15084 45500
rect 21624 45444 21680 45500
rect 21728 45444 21784 45500
rect 21832 45444 21888 45500
rect 28428 45444 28484 45500
rect 28532 45444 28588 45500
rect 28636 45444 28692 45500
rect 6748 45388 6804 45444
rect 6972 45388 7028 45444
rect 7644 45388 7700 45444
rect 20748 45276 20804 45332
rect 11788 44940 11844 44996
rect 3724 44716 3780 44772
rect 11004 44716 11060 44772
rect 13804 44716 13860 44772
rect 4614 44660 4670 44716
rect 4718 44660 4774 44716
rect 4822 44660 4878 44716
rect 11418 44660 11474 44716
rect 11522 44660 11578 44716
rect 11626 44660 11682 44716
rect 18222 44660 18278 44716
rect 18326 44660 18382 44716
rect 18430 44660 18486 44716
rect 25026 44660 25082 44716
rect 25130 44660 25186 44716
rect 25234 44660 25290 44716
rect 3836 44604 3892 44660
rect 12124 44604 12180 44660
rect 3612 44492 3668 44548
rect 10444 44492 10500 44548
rect 13580 44492 13636 44548
rect 7196 44380 7252 44436
rect 13916 44380 13972 44436
rect 14588 44380 14644 44436
rect 17500 44380 17556 44436
rect 5852 44268 5908 44324
rect 10892 44268 10948 44324
rect 17612 44268 17668 44324
rect 23772 44268 23828 44324
rect 5964 44156 6020 44212
rect 11004 44156 11060 44212
rect 19292 44156 19348 44212
rect 6748 43932 6804 43988
rect 8016 43876 8072 43932
rect 8120 43876 8176 43932
rect 8224 43876 8280 43932
rect 14820 43876 14876 43932
rect 14924 43876 14980 43932
rect 15028 43876 15084 43932
rect 21624 43876 21680 43932
rect 21728 43876 21784 43932
rect 21832 43876 21888 43932
rect 28428 43876 28484 43932
rect 28532 43876 28588 43932
rect 28636 43876 28692 43932
rect 10556 43820 10612 43876
rect 11228 43820 11284 43876
rect 23436 43820 23492 43876
rect 3164 43708 3220 43764
rect 20748 43708 20804 43764
rect 25452 43708 25508 43764
rect 16156 43596 16212 43652
rect 21308 43596 21364 43652
rect 5740 43484 5796 43540
rect 10892 43484 10948 43540
rect 13804 43484 13860 43540
rect 14588 43484 14644 43540
rect 15260 43484 15316 43540
rect 5964 43372 6020 43428
rect 9660 43372 9716 43428
rect 18620 43372 18676 43428
rect 16716 43260 16772 43316
rect 26572 43260 26628 43316
rect 20972 43148 21028 43204
rect 4614 43092 4670 43148
rect 4718 43092 4774 43148
rect 4822 43092 4878 43148
rect 11418 43092 11474 43148
rect 11522 43092 11578 43148
rect 11626 43092 11682 43148
rect 18222 43092 18278 43148
rect 18326 43092 18382 43148
rect 18430 43092 18486 43148
rect 25026 43092 25082 43148
rect 25130 43092 25186 43148
rect 25234 43092 25290 43148
rect 10332 43036 10388 43092
rect 12124 42924 12180 42980
rect 16716 42700 16772 42756
rect 23436 42700 23492 42756
rect 11116 42588 11172 42644
rect 9884 42364 9940 42420
rect 10556 42364 10612 42420
rect 12460 42364 12516 42420
rect 13916 42364 13972 42420
rect 8016 42308 8072 42364
rect 8120 42308 8176 42364
rect 8224 42308 8280 42364
rect 14820 42308 14876 42364
rect 14924 42308 14980 42364
rect 15028 42308 15084 42364
rect 21624 42308 21680 42364
rect 21728 42308 21784 42364
rect 21832 42308 21888 42364
rect 28428 42308 28484 42364
rect 28532 42308 28588 42364
rect 28636 42308 28692 42364
rect 12236 42140 12292 42196
rect 20860 42140 20916 42196
rect 24108 42140 24164 42196
rect 24668 42140 24724 42196
rect 11004 42028 11060 42084
rect 18620 42028 18676 42084
rect 19404 42028 19460 42084
rect 24332 42028 24388 42084
rect 7868 41916 7924 41972
rect 18060 41916 18116 41972
rect 21084 41916 21140 41972
rect 24780 41916 24836 41972
rect 9884 41804 9940 41860
rect 10332 41804 10388 41860
rect 25452 41804 25508 41860
rect 16716 41692 16772 41748
rect 24668 41580 24724 41636
rect 4614 41524 4670 41580
rect 4718 41524 4774 41580
rect 4822 41524 4878 41580
rect 11418 41524 11474 41580
rect 11522 41524 11578 41580
rect 11626 41524 11682 41580
rect 18222 41524 18278 41580
rect 18326 41524 18382 41580
rect 18430 41524 18486 41580
rect 25026 41524 25082 41580
rect 25130 41524 25186 41580
rect 25234 41524 25290 41580
rect 17724 41468 17780 41524
rect 15260 41356 15316 41412
rect 19292 41356 19348 41412
rect 23772 41132 23828 41188
rect 13244 41020 13300 41076
rect 18620 41020 18676 41076
rect 17948 40908 18004 40964
rect 23548 40908 23604 40964
rect 4172 40796 4228 40852
rect 7868 40796 7924 40852
rect 11228 40796 11284 40852
rect 11788 40796 11844 40852
rect 19404 40796 19460 40852
rect 25452 40796 25508 40852
rect 8016 40740 8072 40796
rect 8120 40740 8176 40796
rect 8224 40740 8280 40796
rect 14820 40740 14876 40796
rect 14924 40740 14980 40796
rect 15028 40740 15084 40796
rect 21624 40740 21680 40796
rect 21728 40740 21784 40796
rect 21832 40740 21888 40796
rect 28428 40740 28484 40796
rect 28532 40740 28588 40796
rect 28636 40740 28692 40796
rect 21084 40684 21140 40740
rect 9660 40572 9716 40628
rect 15260 40572 15316 40628
rect 24108 40460 24164 40516
rect 20300 40348 20356 40404
rect 7084 40236 7140 40292
rect 23436 40236 23492 40292
rect 4172 40124 4228 40180
rect 16828 40124 16884 40180
rect 4614 39956 4670 40012
rect 4718 39956 4774 40012
rect 4822 39956 4878 40012
rect 11418 39956 11474 40012
rect 11522 39956 11578 40012
rect 11626 39956 11682 40012
rect 18222 39956 18278 40012
rect 18326 39956 18382 40012
rect 18430 39956 18486 40012
rect 25026 39956 25082 40012
rect 25130 39956 25186 40012
rect 25234 39956 25290 40012
rect 11116 39788 11172 39844
rect 11788 39788 11844 39844
rect 13580 39676 13636 39732
rect 13692 39564 13748 39620
rect 15260 39452 15316 39508
rect 6076 39340 6132 39396
rect 21308 39340 21364 39396
rect 11788 39228 11844 39284
rect 17052 39228 17108 39284
rect 20300 39228 20356 39284
rect 8016 39172 8072 39228
rect 8120 39172 8176 39228
rect 8224 39172 8280 39228
rect 14820 39172 14876 39228
rect 14924 39172 14980 39228
rect 15028 39172 15084 39228
rect 21624 39172 21680 39228
rect 21728 39172 21784 39228
rect 21832 39172 21888 39228
rect 28428 39172 28484 39228
rect 28532 39172 28588 39228
rect 28636 39172 28692 39228
rect 10892 39116 10948 39172
rect 20860 39116 20916 39172
rect 22092 39116 22148 39172
rect 16828 39004 16884 39060
rect 3724 38892 3780 38948
rect 7644 38780 7700 38836
rect 16828 38780 16884 38836
rect 20076 38780 20132 38836
rect 11228 38668 11284 38724
rect 17948 38556 18004 38612
rect 21420 38556 21476 38612
rect 5740 38444 5796 38500
rect 21196 38444 21252 38500
rect 22092 38444 22148 38500
rect 4614 38388 4670 38444
rect 4718 38388 4774 38444
rect 4822 38388 4878 38444
rect 11418 38388 11474 38444
rect 11522 38388 11578 38444
rect 11626 38388 11682 38444
rect 18222 38388 18278 38444
rect 18326 38388 18382 38444
rect 18430 38388 18486 38444
rect 25026 38388 25082 38444
rect 25130 38388 25186 38444
rect 25234 38388 25290 38444
rect 12796 38332 12852 38388
rect 2380 38220 2436 38276
rect 11116 38108 11172 38164
rect 19292 38108 19348 38164
rect 4172 37996 4228 38052
rect 11228 37996 11284 38052
rect 21084 37884 21140 37940
rect 24108 37884 24164 37940
rect 21308 37772 21364 37828
rect 23660 37772 23716 37828
rect 7196 37660 7252 37716
rect 8016 37604 8072 37660
rect 8120 37604 8176 37660
rect 8224 37604 8280 37660
rect 14820 37604 14876 37660
rect 14924 37604 14980 37660
rect 15028 37604 15084 37660
rect 21624 37604 21680 37660
rect 21728 37604 21784 37660
rect 21832 37604 21888 37660
rect 28428 37604 28484 37660
rect 28532 37604 28588 37660
rect 28636 37604 28692 37660
rect 12236 37548 12292 37604
rect 20972 37548 21028 37604
rect 24332 37548 24388 37604
rect 5180 37436 5236 37492
rect 13580 37436 13636 37492
rect 15484 37436 15540 37492
rect 19292 37436 19348 37492
rect 25452 37436 25508 37492
rect 18956 37324 19012 37380
rect 26796 37324 26852 37380
rect 4614 36820 4670 36876
rect 4718 36820 4774 36876
rect 4822 36820 4878 36876
rect 24780 36988 24836 37044
rect 10444 36876 10500 36932
rect 11004 36876 11060 36932
rect 11418 36820 11474 36876
rect 11522 36820 11578 36876
rect 11626 36820 11682 36876
rect 18222 36820 18278 36876
rect 18326 36820 18382 36876
rect 18430 36820 18486 36876
rect 25026 36820 25082 36876
rect 25130 36820 25186 36876
rect 25234 36820 25290 36876
rect 9884 36764 9940 36820
rect 12796 36764 12852 36820
rect 18620 36764 18676 36820
rect 6972 36652 7028 36708
rect 11788 36652 11844 36708
rect 14364 36652 14420 36708
rect 18620 36540 18676 36596
rect 24780 36540 24836 36596
rect 13692 36428 13748 36484
rect 18956 36428 19012 36484
rect 13804 36316 13860 36372
rect 26796 36316 26852 36372
rect 11228 36204 11284 36260
rect 3836 36092 3892 36148
rect 6188 36092 6244 36148
rect 8016 36036 8072 36092
rect 8120 36036 8176 36092
rect 8224 36036 8280 36092
rect 17500 36092 17556 36148
rect 14820 36036 14876 36092
rect 14924 36036 14980 36092
rect 15028 36036 15084 36092
rect 21624 36036 21680 36092
rect 21728 36036 21784 36092
rect 21832 36036 21888 36092
rect 28428 36036 28484 36092
rect 28532 36036 28588 36092
rect 28636 36036 28692 36092
rect 4060 35980 4116 36036
rect 7868 35644 7924 35700
rect 12460 35644 12516 35700
rect 22764 35532 22820 35588
rect 11116 35420 11172 35476
rect 11788 35420 11844 35476
rect 14476 35420 14532 35476
rect 17724 35420 17780 35476
rect 18956 35420 19012 35476
rect 25452 35420 25508 35476
rect 14364 35308 14420 35364
rect 20860 35308 20916 35364
rect 22988 35308 23044 35364
rect 4614 35252 4670 35308
rect 4718 35252 4774 35308
rect 4822 35252 4878 35308
rect 11418 35252 11474 35308
rect 11522 35252 11578 35308
rect 11626 35252 11682 35308
rect 18222 35252 18278 35308
rect 18326 35252 18382 35308
rect 18430 35252 18486 35308
rect 25026 35252 25082 35308
rect 25130 35252 25186 35308
rect 25234 35252 25290 35308
rect 11004 35196 11060 35252
rect 24668 35196 24724 35252
rect 15820 35084 15876 35140
rect 16380 35084 16436 35140
rect 19180 35084 19236 35140
rect 13692 34972 13748 35028
rect 19740 34972 19796 35028
rect 20300 34972 20356 35028
rect 10444 34860 10500 34916
rect 22092 34860 22148 34916
rect 24668 34748 24724 34804
rect 3612 34636 3668 34692
rect 19964 34524 20020 34580
rect 22204 34524 22260 34580
rect 8016 34468 8072 34524
rect 8120 34468 8176 34524
rect 8224 34468 8280 34524
rect 14820 34468 14876 34524
rect 14924 34468 14980 34524
rect 15028 34468 15084 34524
rect 21624 34468 21680 34524
rect 21728 34468 21784 34524
rect 21832 34468 21888 34524
rect 28428 34468 28484 34524
rect 28532 34468 28588 34524
rect 28636 34468 28692 34524
rect 25452 34412 25508 34468
rect 11228 34300 11284 34356
rect 19628 33740 19684 33796
rect 4614 33684 4670 33740
rect 4718 33684 4774 33740
rect 4822 33684 4878 33740
rect 11418 33684 11474 33740
rect 11522 33684 11578 33740
rect 11626 33684 11682 33740
rect 18222 33684 18278 33740
rect 18326 33684 18382 33740
rect 18430 33684 18486 33740
rect 25026 33684 25082 33740
rect 25130 33684 25186 33740
rect 25234 33684 25290 33740
rect 8540 33628 8596 33684
rect 23324 33628 23380 33684
rect 23660 33628 23716 33684
rect 10556 33516 10612 33572
rect 24444 33404 24500 33460
rect 5180 33292 5236 33348
rect 10556 33292 10612 33348
rect 20748 33292 20804 33348
rect 16044 33068 16100 33124
rect 19964 33068 20020 33124
rect 8016 32900 8072 32956
rect 8120 32900 8176 32956
rect 8224 32900 8280 32956
rect 14820 32900 14876 32956
rect 14924 32900 14980 32956
rect 15028 32900 15084 32956
rect 21624 32900 21680 32956
rect 21728 32900 21784 32956
rect 21832 32900 21888 32956
rect 28428 32900 28484 32956
rect 28532 32900 28588 32956
rect 28636 32900 28692 32956
rect 10892 32844 10948 32900
rect 9212 32732 9268 32788
rect 11004 32732 11060 32788
rect 11228 32732 11284 32788
rect 16604 32732 16660 32788
rect 17500 32732 17556 32788
rect 17724 32732 17780 32788
rect 19404 32732 19460 32788
rect 25564 32620 25620 32676
rect 17500 32396 17556 32452
rect 20076 32396 20132 32452
rect 4614 32116 4670 32172
rect 4718 32116 4774 32172
rect 4822 32116 4878 32172
rect 24780 32172 24836 32228
rect 11418 32116 11474 32172
rect 11522 32116 11578 32172
rect 11626 32116 11682 32172
rect 18222 32116 18278 32172
rect 18326 32116 18382 32172
rect 18430 32116 18486 32172
rect 25026 32116 25082 32172
rect 25130 32116 25186 32172
rect 25234 32116 25290 32172
rect 20524 32060 20580 32116
rect 11228 31836 11284 31892
rect 11004 31724 11060 31780
rect 20300 31948 20356 32004
rect 23548 31836 23604 31892
rect 20748 31724 20804 31780
rect 21196 31612 21252 31668
rect 25788 31612 25844 31668
rect 20860 31500 20916 31556
rect 19740 31388 19796 31444
rect 8016 31332 8072 31388
rect 8120 31332 8176 31388
rect 8224 31332 8280 31388
rect 14820 31332 14876 31388
rect 14924 31332 14980 31388
rect 15028 31332 15084 31388
rect 21624 31332 21680 31388
rect 21728 31332 21784 31388
rect 21832 31332 21888 31388
rect 28428 31332 28484 31388
rect 28532 31332 28588 31388
rect 28636 31332 28692 31388
rect 7644 31276 7700 31332
rect 16492 31164 16548 31220
rect 21980 31164 22036 31220
rect 19740 31052 19796 31108
rect 26124 31052 26180 31108
rect 25788 30828 25844 30884
rect 23548 30716 23604 30772
rect 4614 30548 4670 30604
rect 4718 30548 4774 30604
rect 4822 30548 4878 30604
rect 11418 30548 11474 30604
rect 11522 30548 11578 30604
rect 11626 30548 11682 30604
rect 18222 30548 18278 30604
rect 18326 30548 18382 30604
rect 18430 30548 18486 30604
rect 25026 30548 25082 30604
rect 25130 30548 25186 30604
rect 25234 30548 25290 30604
rect 21420 30380 21476 30436
rect 20300 30044 20356 30100
rect 8016 29764 8072 29820
rect 8120 29764 8176 29820
rect 8224 29764 8280 29820
rect 14820 29764 14876 29820
rect 14924 29764 14980 29820
rect 15028 29764 15084 29820
rect 21624 29764 21680 29820
rect 21728 29764 21784 29820
rect 21832 29764 21888 29820
rect 28428 29764 28484 29820
rect 28532 29764 28588 29820
rect 28636 29764 28692 29820
rect 24780 29260 24836 29316
rect 8540 29036 8596 29092
rect 4614 28980 4670 29036
rect 4718 28980 4774 29036
rect 4822 28980 4878 29036
rect 11418 28980 11474 29036
rect 11522 28980 11578 29036
rect 11626 28980 11682 29036
rect 18222 28980 18278 29036
rect 18326 28980 18382 29036
rect 18430 28980 18486 29036
rect 25026 28980 25082 29036
rect 25130 28980 25186 29036
rect 25234 28980 25290 29036
rect 5180 28812 5236 28868
rect 25564 28812 25620 28868
rect 10556 28700 10612 28756
rect 11116 28700 11172 28756
rect 5068 28476 5124 28532
rect 13692 28476 13748 28532
rect 20524 28476 20580 28532
rect 24780 28476 24836 28532
rect 25788 28364 25844 28420
rect 25564 28252 25620 28308
rect 26684 28252 26740 28308
rect 8016 28196 8072 28252
rect 8120 28196 8176 28252
rect 8224 28196 8280 28252
rect 14820 28196 14876 28252
rect 14924 28196 14980 28252
rect 15028 28196 15084 28252
rect 21624 28196 21680 28252
rect 21728 28196 21784 28252
rect 21832 28196 21888 28252
rect 28428 28196 28484 28252
rect 28532 28196 28588 28252
rect 28636 28196 28692 28252
rect 23548 28140 23604 28196
rect 22092 28028 22148 28084
rect 13692 27804 13748 27860
rect 26684 27804 26740 27860
rect 17724 27468 17780 27524
rect 21196 27468 21252 27524
rect 4614 27412 4670 27468
rect 4718 27412 4774 27468
rect 4822 27412 4878 27468
rect 11418 27412 11474 27468
rect 11522 27412 11578 27468
rect 11626 27412 11682 27468
rect 18222 27412 18278 27468
rect 18326 27412 18382 27468
rect 18430 27412 18486 27468
rect 25026 27412 25082 27468
rect 25130 27412 25186 27468
rect 25234 27412 25290 27468
rect 10556 27356 10612 27412
rect 19964 27356 20020 27412
rect 20524 27356 20580 27412
rect 26124 27356 26180 27412
rect 7644 27244 7700 27300
rect 20748 27244 20804 27300
rect 9772 27132 9828 27188
rect 19292 27020 19348 27076
rect 20412 26796 20468 26852
rect 19180 26684 19236 26740
rect 23324 26684 23380 26740
rect 8016 26628 8072 26684
rect 8120 26628 8176 26684
rect 8224 26628 8280 26684
rect 14820 26628 14876 26684
rect 14924 26628 14980 26684
rect 15028 26628 15084 26684
rect 18620 26348 18676 26404
rect 19964 26348 20020 26404
rect 21624 26628 21680 26684
rect 21728 26628 21784 26684
rect 21832 26628 21888 26684
rect 28428 26628 28484 26684
rect 28532 26628 28588 26684
rect 28636 26628 28692 26684
rect 22204 26460 22260 26516
rect 14588 26124 14644 26180
rect 12684 26012 12740 26068
rect 19404 26012 19460 26068
rect 10892 25900 10948 25956
rect 23548 25900 23604 25956
rect 4614 25844 4670 25900
rect 4718 25844 4774 25900
rect 4822 25844 4878 25900
rect 11418 25844 11474 25900
rect 11522 25844 11578 25900
rect 11626 25844 11682 25900
rect 18222 25844 18278 25900
rect 18326 25844 18382 25900
rect 18430 25844 18486 25900
rect 19180 25788 19236 25844
rect 25026 25844 25082 25900
rect 25130 25844 25186 25900
rect 25234 25844 25290 25900
rect 14588 25452 14644 25508
rect 18620 25340 18676 25396
rect 19516 25116 19572 25172
rect 24444 25116 24500 25172
rect 8016 25060 8072 25116
rect 8120 25060 8176 25116
rect 8224 25060 8280 25116
rect 14820 25060 14876 25116
rect 14924 25060 14980 25116
rect 15028 25060 15084 25116
rect 21624 25060 21680 25116
rect 21728 25060 21784 25116
rect 21832 25060 21888 25116
rect 28428 25060 28484 25116
rect 28532 25060 28588 25116
rect 28636 25060 28692 25116
rect 11788 24892 11844 24948
rect 19068 24892 19124 24948
rect 20860 24892 20916 24948
rect 21196 24892 21252 24948
rect 25452 24892 25508 24948
rect 19628 24780 19684 24836
rect 20748 24668 20804 24724
rect 9772 24332 9828 24388
rect 19628 24332 19684 24388
rect 4614 24276 4670 24332
rect 4718 24276 4774 24332
rect 4822 24276 4878 24332
rect 11418 24276 11474 24332
rect 11522 24276 11578 24332
rect 11626 24276 11682 24332
rect 18222 24276 18278 24332
rect 18326 24276 18382 24332
rect 18430 24276 18486 24332
rect 25026 24276 25082 24332
rect 25130 24276 25186 24332
rect 25234 24276 25290 24332
rect 19740 24220 19796 24276
rect 26684 24220 26740 24276
rect 10444 23996 10500 24052
rect 19852 23996 19908 24052
rect 16604 23772 16660 23828
rect 9212 23660 9268 23716
rect 12684 23548 12740 23604
rect 22204 23548 22260 23604
rect 8016 23492 8072 23548
rect 8120 23492 8176 23548
rect 8224 23492 8280 23548
rect 14820 23492 14876 23548
rect 14924 23492 14980 23548
rect 15028 23492 15084 23548
rect 21624 23492 21680 23548
rect 21728 23492 21784 23548
rect 21832 23492 21888 23548
rect 28428 23492 28484 23548
rect 28532 23492 28588 23548
rect 28636 23492 28692 23548
rect 23772 23436 23828 23492
rect 11788 23324 11844 23380
rect 26684 23324 26740 23380
rect 22652 23212 22708 23268
rect 15484 22876 15540 22932
rect 17388 22764 17444 22820
rect 4614 22708 4670 22764
rect 4718 22708 4774 22764
rect 4822 22708 4878 22764
rect 11418 22708 11474 22764
rect 11522 22708 11578 22764
rect 11626 22708 11682 22764
rect 18222 22708 18278 22764
rect 18326 22708 18382 22764
rect 18430 22708 18486 22764
rect 25026 22708 25082 22764
rect 25130 22708 25186 22764
rect 25234 22708 25290 22764
rect 16380 22652 16436 22708
rect 19292 22540 19348 22596
rect 23772 22316 23828 22372
rect 17724 22092 17780 22148
rect 8016 21924 8072 21980
rect 8120 21924 8176 21980
rect 8224 21924 8280 21980
rect 14820 21924 14876 21980
rect 14924 21924 14980 21980
rect 15028 21924 15084 21980
rect 21624 21924 21680 21980
rect 21728 21924 21784 21980
rect 21832 21924 21888 21980
rect 28428 21924 28484 21980
rect 28532 21924 28588 21980
rect 28636 21924 28692 21980
rect 17724 21308 17780 21364
rect 16940 21196 16996 21252
rect 4614 21140 4670 21196
rect 4718 21140 4774 21196
rect 4822 21140 4878 21196
rect 11418 21140 11474 21196
rect 11522 21140 11578 21196
rect 11626 21140 11682 21196
rect 18222 21140 18278 21196
rect 18326 21140 18382 21196
rect 18430 21140 18486 21196
rect 25026 21140 25082 21196
rect 25130 21140 25186 21196
rect 25234 21140 25290 21196
rect 7084 20636 7140 20692
rect 8016 20356 8072 20412
rect 8120 20356 8176 20412
rect 8224 20356 8280 20412
rect 14820 20356 14876 20412
rect 14924 20356 14980 20412
rect 15028 20356 15084 20412
rect 21624 20356 21680 20412
rect 21728 20356 21784 20412
rect 21832 20356 21888 20412
rect 28428 20356 28484 20412
rect 28532 20356 28588 20412
rect 28636 20356 28692 20412
rect 4614 19572 4670 19628
rect 4718 19572 4774 19628
rect 4822 19572 4878 19628
rect 11418 19572 11474 19628
rect 11522 19572 11578 19628
rect 11626 19572 11682 19628
rect 18222 19572 18278 19628
rect 18326 19572 18382 19628
rect 18430 19572 18486 19628
rect 25026 19572 25082 19628
rect 25130 19572 25186 19628
rect 25234 19572 25290 19628
rect 15372 19292 15428 19348
rect 16268 19068 16324 19124
rect 8016 18788 8072 18844
rect 8120 18788 8176 18844
rect 8224 18788 8280 18844
rect 14820 18788 14876 18844
rect 14924 18788 14980 18844
rect 15028 18788 15084 18844
rect 21624 18788 21680 18844
rect 21728 18788 21784 18844
rect 21832 18788 21888 18844
rect 28428 18788 28484 18844
rect 28532 18788 28588 18844
rect 28636 18788 28692 18844
rect 4396 18396 4452 18452
rect 4614 18004 4670 18060
rect 4718 18004 4774 18060
rect 4822 18004 4878 18060
rect 11418 18004 11474 18060
rect 11522 18004 11578 18060
rect 11626 18004 11682 18060
rect 18222 18004 18278 18060
rect 18326 18004 18382 18060
rect 18430 18004 18486 18060
rect 25026 18004 25082 18060
rect 25130 18004 25186 18060
rect 25234 18004 25290 18060
rect 15484 17724 15540 17780
rect 8016 17220 8072 17276
rect 8120 17220 8176 17276
rect 8224 17220 8280 17276
rect 14820 17220 14876 17276
rect 14924 17220 14980 17276
rect 15028 17220 15084 17276
rect 21624 17220 21680 17276
rect 21728 17220 21784 17276
rect 21832 17220 21888 17276
rect 28428 17220 28484 17276
rect 28532 17220 28588 17276
rect 28636 17220 28692 17276
rect 16268 17164 16324 17220
rect 16268 16940 16324 16996
rect 5852 16716 5908 16772
rect 4614 16436 4670 16492
rect 4718 16436 4774 16492
rect 4822 16436 4878 16492
rect 11418 16436 11474 16492
rect 11522 16436 11578 16492
rect 11626 16436 11682 16492
rect 18222 16436 18278 16492
rect 18326 16436 18382 16492
rect 18430 16436 18486 16492
rect 25026 16436 25082 16492
rect 25130 16436 25186 16492
rect 25234 16436 25290 16492
rect 8016 15652 8072 15708
rect 8120 15652 8176 15708
rect 8224 15652 8280 15708
rect 14820 15652 14876 15708
rect 14924 15652 14980 15708
rect 15028 15652 15084 15708
rect 21624 15652 21680 15708
rect 21728 15652 21784 15708
rect 21832 15652 21888 15708
rect 28428 15652 28484 15708
rect 28532 15652 28588 15708
rect 28636 15652 28692 15708
rect 10668 15372 10724 15428
rect 14588 15148 14644 15204
rect 16940 14924 16996 14980
rect 4614 14868 4670 14924
rect 4718 14868 4774 14924
rect 4822 14868 4878 14924
rect 11418 14868 11474 14924
rect 11522 14868 11578 14924
rect 11626 14868 11682 14924
rect 18222 14868 18278 14924
rect 18326 14868 18382 14924
rect 18430 14868 18486 14924
rect 25026 14868 25082 14924
rect 25130 14868 25186 14924
rect 25234 14868 25290 14924
rect 9884 14700 9940 14756
rect 5852 14252 5908 14308
rect 8016 14084 8072 14140
rect 8120 14084 8176 14140
rect 8224 14084 8280 14140
rect 14820 14084 14876 14140
rect 14924 14084 14980 14140
rect 15028 14084 15084 14140
rect 21624 14084 21680 14140
rect 21728 14084 21784 14140
rect 21832 14084 21888 14140
rect 28428 14084 28484 14140
rect 28532 14084 28588 14140
rect 28636 14084 28692 14140
rect 3500 13916 3556 13972
rect 9884 13356 9940 13412
rect 4614 13300 4670 13356
rect 4718 13300 4774 13356
rect 4822 13300 4878 13356
rect 11418 13300 11474 13356
rect 11522 13300 11578 13356
rect 11626 13300 11682 13356
rect 18222 13300 18278 13356
rect 18326 13300 18382 13356
rect 18430 13300 18486 13356
rect 25026 13300 25082 13356
rect 25130 13300 25186 13356
rect 25234 13300 25290 13356
rect 7084 13132 7140 13188
rect 8016 12516 8072 12572
rect 8120 12516 8176 12572
rect 8224 12516 8280 12572
rect 14820 12516 14876 12572
rect 14924 12516 14980 12572
rect 15028 12516 15084 12572
rect 21624 12516 21680 12572
rect 21728 12516 21784 12572
rect 21832 12516 21888 12572
rect 28428 12516 28484 12572
rect 28532 12516 28588 12572
rect 28636 12516 28692 12572
rect 16380 12348 16436 12404
rect 18620 12348 18676 12404
rect 18956 12348 19012 12404
rect 17388 12124 17444 12180
rect 18620 11788 18676 11844
rect 4614 11732 4670 11788
rect 4718 11732 4774 11788
rect 4822 11732 4878 11788
rect 11418 11732 11474 11788
rect 11522 11732 11578 11788
rect 11626 11732 11682 11788
rect 18222 11732 18278 11788
rect 18326 11732 18382 11788
rect 18430 11732 18486 11788
rect 25026 11732 25082 11788
rect 25130 11732 25186 11788
rect 25234 11732 25290 11788
rect 20412 11676 20468 11732
rect 20972 11564 21028 11620
rect 5852 11340 5908 11396
rect 5852 11116 5908 11172
rect 8016 10948 8072 11004
rect 8120 10948 8176 11004
rect 8224 10948 8280 11004
rect 14820 10948 14876 11004
rect 14924 10948 14980 11004
rect 15028 10948 15084 11004
rect 21624 10948 21680 11004
rect 21728 10948 21784 11004
rect 21832 10948 21888 11004
rect 28428 10948 28484 11004
rect 28532 10948 28588 11004
rect 28636 10948 28692 11004
rect 18732 10780 18788 10836
rect 20300 10780 20356 10836
rect 16268 10556 16324 10612
rect 4614 10164 4670 10220
rect 4718 10164 4774 10220
rect 4822 10164 4878 10220
rect 11418 10164 11474 10220
rect 11522 10164 11578 10220
rect 11626 10164 11682 10220
rect 18222 10164 18278 10220
rect 18326 10164 18382 10220
rect 18430 10164 18486 10220
rect 25026 10164 25082 10220
rect 25130 10164 25186 10220
rect 25234 10164 25290 10220
rect 16268 10108 16324 10164
rect 8016 9380 8072 9436
rect 8120 9380 8176 9436
rect 8224 9380 8280 9436
rect 14820 9380 14876 9436
rect 14924 9380 14980 9436
rect 15028 9380 15084 9436
rect 21624 9380 21680 9436
rect 21728 9380 21784 9436
rect 21832 9380 21888 9436
rect 28428 9380 28484 9436
rect 28532 9380 28588 9436
rect 28636 9380 28692 9436
rect 16268 9100 16324 9156
rect 20972 8876 21028 8932
rect 4614 8596 4670 8652
rect 4718 8596 4774 8652
rect 4822 8596 4878 8652
rect 11418 8596 11474 8652
rect 11522 8596 11578 8652
rect 11626 8596 11682 8652
rect 18222 8596 18278 8652
rect 18326 8596 18382 8652
rect 18430 8596 18486 8652
rect 25026 8596 25082 8652
rect 25130 8596 25186 8652
rect 25234 8596 25290 8652
rect 3388 8204 3444 8260
rect 20636 7980 20692 8036
rect 8016 7812 8072 7868
rect 8120 7812 8176 7868
rect 8224 7812 8280 7868
rect 14820 7812 14876 7868
rect 14924 7812 14980 7868
rect 15028 7812 15084 7868
rect 21624 7812 21680 7868
rect 21728 7812 21784 7868
rect 21832 7812 21888 7868
rect 28428 7812 28484 7868
rect 28532 7812 28588 7868
rect 28636 7812 28692 7868
rect 4614 7028 4670 7084
rect 4718 7028 4774 7084
rect 4822 7028 4878 7084
rect 11418 7028 11474 7084
rect 11522 7028 11578 7084
rect 11626 7028 11682 7084
rect 18222 7028 18278 7084
rect 18326 7028 18382 7084
rect 18430 7028 18486 7084
rect 25026 7028 25082 7084
rect 25130 7028 25186 7084
rect 25234 7028 25290 7084
rect 15708 6636 15764 6692
rect 8016 6244 8072 6300
rect 8120 6244 8176 6300
rect 8224 6244 8280 6300
rect 14820 6244 14876 6300
rect 14924 6244 14980 6300
rect 15028 6244 15084 6300
rect 21624 6244 21680 6300
rect 21728 6244 21784 6300
rect 21832 6244 21888 6300
rect 28428 6244 28484 6300
rect 28532 6244 28588 6300
rect 28636 6244 28692 6300
rect 4614 5460 4670 5516
rect 4718 5460 4774 5516
rect 4822 5460 4878 5516
rect 11418 5460 11474 5516
rect 11522 5460 11578 5516
rect 11626 5460 11682 5516
rect 18222 5460 18278 5516
rect 18326 5460 18382 5516
rect 18430 5460 18486 5516
rect 25026 5460 25082 5516
rect 25130 5460 25186 5516
rect 25234 5460 25290 5516
rect 8016 4676 8072 4732
rect 8120 4676 8176 4732
rect 8224 4676 8280 4732
rect 14820 4676 14876 4732
rect 14924 4676 14980 4732
rect 15028 4676 15084 4732
rect 21624 4676 21680 4732
rect 21728 4676 21784 4732
rect 21832 4676 21888 4732
rect 28428 4676 28484 4732
rect 28532 4676 28588 4732
rect 28636 4676 28692 4732
rect 18060 4060 18116 4116
rect 4614 3892 4670 3948
rect 4718 3892 4774 3948
rect 4822 3892 4878 3948
rect 11418 3892 11474 3948
rect 11522 3892 11578 3948
rect 11626 3892 11682 3948
rect 18222 3892 18278 3948
rect 18326 3892 18382 3948
rect 18430 3892 18486 3948
rect 25026 3892 25082 3948
rect 25130 3892 25186 3948
rect 25234 3892 25290 3948
rect 23212 3500 23268 3556
rect 19852 3388 19908 3444
rect 8016 3108 8072 3164
rect 8120 3108 8176 3164
rect 8224 3108 8280 3164
rect 14820 3108 14876 3164
rect 14924 3108 14980 3164
rect 15028 3108 15084 3164
rect 21624 3108 21680 3164
rect 21728 3108 21784 3164
rect 21832 3108 21888 3164
rect 28428 3108 28484 3164
rect 28532 3108 28588 3164
rect 28636 3108 28692 3164
rect 19852 2716 19908 2772
rect 4614 2324 4670 2380
rect 4718 2324 4774 2380
rect 4822 2324 4878 2380
rect 11418 2324 11474 2380
rect 11522 2324 11578 2380
rect 11626 2324 11682 2380
rect 18222 2324 18278 2380
rect 18326 2324 18382 2380
rect 18430 2324 18486 2380
rect 25026 2324 25082 2380
rect 25130 2324 25186 2380
rect 25234 2324 25290 2380
rect 18060 2156 18116 2212
rect 8016 1540 8072 1596
rect 8120 1540 8176 1596
rect 8224 1540 8280 1596
rect 14820 1540 14876 1596
rect 14924 1540 14980 1596
rect 15028 1540 15084 1596
rect 21624 1540 21680 1596
rect 21728 1540 21784 1596
rect 21832 1540 21888 1596
rect 28428 1540 28484 1596
rect 28532 1540 28588 1596
rect 28636 1540 28692 1596
<< metal4 >>
rect 4586 118412 4906 118444
rect 4586 118356 4614 118412
rect 4670 118356 4718 118412
rect 4774 118356 4822 118412
rect 4878 118356 4906 118412
rect 4586 116844 4906 118356
rect 4586 116788 4614 116844
rect 4670 116788 4718 116844
rect 4774 116788 4822 116844
rect 4878 116788 4906 116844
rect 4586 115276 4906 116788
rect 4586 115220 4614 115276
rect 4670 115220 4718 115276
rect 4774 115220 4822 115276
rect 4878 115220 4906 115276
rect 4586 113708 4906 115220
rect 4586 113652 4614 113708
rect 4670 113652 4718 113708
rect 4774 113652 4822 113708
rect 4878 113652 4906 113708
rect 4586 112140 4906 113652
rect 4586 112084 4614 112140
rect 4670 112084 4718 112140
rect 4774 112084 4822 112140
rect 4878 112084 4906 112140
rect 4586 110572 4906 112084
rect 4586 110516 4614 110572
rect 4670 110516 4718 110572
rect 4774 110516 4822 110572
rect 4878 110516 4906 110572
rect 4586 109004 4906 110516
rect 4586 108948 4614 109004
rect 4670 108948 4718 109004
rect 4774 108948 4822 109004
rect 4878 108948 4906 109004
rect 4586 107436 4906 108948
rect 4586 107380 4614 107436
rect 4670 107380 4718 107436
rect 4774 107380 4822 107436
rect 4878 107380 4906 107436
rect 4586 105868 4906 107380
rect 4586 105812 4614 105868
rect 4670 105812 4718 105868
rect 4774 105812 4822 105868
rect 4878 105812 4906 105868
rect 4586 104300 4906 105812
rect 4586 104244 4614 104300
rect 4670 104244 4718 104300
rect 4774 104244 4822 104300
rect 4878 104244 4906 104300
rect 4586 102732 4906 104244
rect 4586 102676 4614 102732
rect 4670 102676 4718 102732
rect 4774 102676 4822 102732
rect 4878 102676 4906 102732
rect 4586 101164 4906 102676
rect 7988 117628 8308 118444
rect 7988 117572 8016 117628
rect 8072 117572 8120 117628
rect 8176 117572 8224 117628
rect 8280 117572 8308 117628
rect 7988 116060 8308 117572
rect 7988 116004 8016 116060
rect 8072 116004 8120 116060
rect 8176 116004 8224 116060
rect 8280 116004 8308 116060
rect 7988 114492 8308 116004
rect 7988 114436 8016 114492
rect 8072 114436 8120 114492
rect 8176 114436 8224 114492
rect 8280 114436 8308 114492
rect 7988 112924 8308 114436
rect 7988 112868 8016 112924
rect 8072 112868 8120 112924
rect 8176 112868 8224 112924
rect 8280 112868 8308 112924
rect 7988 111356 8308 112868
rect 7988 111300 8016 111356
rect 8072 111300 8120 111356
rect 8176 111300 8224 111356
rect 8280 111300 8308 111356
rect 7988 109788 8308 111300
rect 7988 109732 8016 109788
rect 8072 109732 8120 109788
rect 8176 109732 8224 109788
rect 8280 109732 8308 109788
rect 7988 108220 8308 109732
rect 7988 108164 8016 108220
rect 8072 108164 8120 108220
rect 8176 108164 8224 108220
rect 8280 108164 8308 108220
rect 7988 106652 8308 108164
rect 7988 106596 8016 106652
rect 8072 106596 8120 106652
rect 8176 106596 8224 106652
rect 8280 106596 8308 106652
rect 7988 105084 8308 106596
rect 7988 105028 8016 105084
rect 8072 105028 8120 105084
rect 8176 105028 8224 105084
rect 8280 105028 8308 105084
rect 7988 103516 8308 105028
rect 11390 118412 11710 118444
rect 11390 118356 11418 118412
rect 11474 118356 11522 118412
rect 11578 118356 11626 118412
rect 11682 118356 11710 118412
rect 11390 116844 11710 118356
rect 11390 116788 11418 116844
rect 11474 116788 11522 116844
rect 11578 116788 11626 116844
rect 11682 116788 11710 116844
rect 11390 115276 11710 116788
rect 11390 115220 11418 115276
rect 11474 115220 11522 115276
rect 11578 115220 11626 115276
rect 11682 115220 11710 115276
rect 11390 113708 11710 115220
rect 11390 113652 11418 113708
rect 11474 113652 11522 113708
rect 11578 113652 11626 113708
rect 11682 113652 11710 113708
rect 11390 112140 11710 113652
rect 11390 112084 11418 112140
rect 11474 112084 11522 112140
rect 11578 112084 11626 112140
rect 11682 112084 11710 112140
rect 11390 110572 11710 112084
rect 11390 110516 11418 110572
rect 11474 110516 11522 110572
rect 11578 110516 11626 110572
rect 11682 110516 11710 110572
rect 11390 109004 11710 110516
rect 11390 108948 11418 109004
rect 11474 108948 11522 109004
rect 11578 108948 11626 109004
rect 11682 108948 11710 109004
rect 11390 107436 11710 108948
rect 11390 107380 11418 107436
rect 11474 107380 11522 107436
rect 11578 107380 11626 107436
rect 11682 107380 11710 107436
rect 11390 105868 11710 107380
rect 11390 105812 11418 105868
rect 11474 105812 11522 105868
rect 11578 105812 11626 105868
rect 11682 105812 11710 105868
rect 8540 104356 8596 104366
rect 8540 103796 8596 104300
rect 11390 104300 11710 105812
rect 11390 104244 11418 104300
rect 11474 104244 11522 104300
rect 11578 104244 11626 104300
rect 11682 104244 11710 104300
rect 8540 103730 8596 103740
rect 9436 103796 9492 103806
rect 7988 103460 8016 103516
rect 8072 103460 8120 103516
rect 8176 103460 8224 103516
rect 8280 103460 8308 103516
rect 4586 101108 4614 101164
rect 4670 101108 4718 101164
rect 4774 101108 4822 101164
rect 4878 101108 4906 101164
rect 4586 99596 4906 101108
rect 4586 99540 4614 99596
rect 4670 99540 4718 99596
rect 4774 99540 4822 99596
rect 4878 99540 4906 99596
rect 4586 98028 4906 99540
rect 4586 97972 4614 98028
rect 4670 97972 4718 98028
rect 4774 97972 4822 98028
rect 4878 97972 4906 98028
rect 4586 96460 4906 97972
rect 4586 96404 4614 96460
rect 4670 96404 4718 96460
rect 4774 96404 4822 96460
rect 4878 96404 4906 96460
rect 4586 94892 4906 96404
rect 4586 94836 4614 94892
rect 4670 94836 4718 94892
rect 4774 94836 4822 94892
rect 4878 94836 4906 94892
rect 4586 93324 4906 94836
rect 6524 102564 6580 102574
rect 6524 94612 6580 102508
rect 6524 94546 6580 94556
rect 7988 101948 8308 103460
rect 9436 102228 9492 103740
rect 9436 102162 9492 102172
rect 9660 102788 9716 102798
rect 7988 101892 8016 101948
rect 8072 101892 8120 101948
rect 8176 101892 8224 101948
rect 8280 101892 8308 101948
rect 7988 100380 8308 101892
rect 7988 100324 8016 100380
rect 8072 100324 8120 100380
rect 8176 100324 8224 100380
rect 8280 100324 8308 100380
rect 7988 98812 8308 100324
rect 7988 98756 8016 98812
rect 8072 98756 8120 98812
rect 8176 98756 8224 98812
rect 8280 98756 8308 98812
rect 7988 97244 8308 98756
rect 7988 97188 8016 97244
rect 8072 97188 8120 97244
rect 8176 97188 8224 97244
rect 8280 97188 8308 97244
rect 7988 95676 8308 97188
rect 9660 97076 9716 102732
rect 9660 97010 9716 97020
rect 11390 102732 11710 104244
rect 11390 102676 11418 102732
rect 11474 102676 11522 102732
rect 11578 102676 11626 102732
rect 11682 102676 11710 102732
rect 11390 101164 11710 102676
rect 11390 101108 11418 101164
rect 11474 101108 11522 101164
rect 11578 101108 11626 101164
rect 11682 101108 11710 101164
rect 11390 99596 11710 101108
rect 11390 99540 11418 99596
rect 11474 99540 11522 99596
rect 11578 99540 11626 99596
rect 11682 99540 11710 99596
rect 11390 98028 11710 99540
rect 11390 97972 11418 98028
rect 11474 97972 11522 98028
rect 11578 97972 11626 98028
rect 11682 97972 11710 98028
rect 11390 96460 11710 97972
rect 14792 117628 15112 118444
rect 14792 117572 14820 117628
rect 14876 117572 14924 117628
rect 14980 117572 15028 117628
rect 15084 117572 15112 117628
rect 14792 116060 15112 117572
rect 14792 116004 14820 116060
rect 14876 116004 14924 116060
rect 14980 116004 15028 116060
rect 15084 116004 15112 116060
rect 14792 114492 15112 116004
rect 14792 114436 14820 114492
rect 14876 114436 14924 114492
rect 14980 114436 15028 114492
rect 15084 114436 15112 114492
rect 14792 112924 15112 114436
rect 14792 112868 14820 112924
rect 14876 112868 14924 112924
rect 14980 112868 15028 112924
rect 15084 112868 15112 112924
rect 14792 111356 15112 112868
rect 14792 111300 14820 111356
rect 14876 111300 14924 111356
rect 14980 111300 15028 111356
rect 15084 111300 15112 111356
rect 14792 109788 15112 111300
rect 14792 109732 14820 109788
rect 14876 109732 14924 109788
rect 14980 109732 15028 109788
rect 15084 109732 15112 109788
rect 14792 108220 15112 109732
rect 14792 108164 14820 108220
rect 14876 108164 14924 108220
rect 14980 108164 15028 108220
rect 15084 108164 15112 108220
rect 14792 106652 15112 108164
rect 14792 106596 14820 106652
rect 14876 106596 14924 106652
rect 14980 106596 15028 106652
rect 15084 106596 15112 106652
rect 14792 105084 15112 106596
rect 14792 105028 14820 105084
rect 14876 105028 14924 105084
rect 14980 105028 15028 105084
rect 15084 105028 15112 105084
rect 14792 103516 15112 105028
rect 14792 103460 14820 103516
rect 14876 103460 14924 103516
rect 14980 103460 15028 103516
rect 15084 103460 15112 103516
rect 14792 101948 15112 103460
rect 14792 101892 14820 101948
rect 14876 101892 14924 101948
rect 14980 101892 15028 101948
rect 15084 101892 15112 101948
rect 14792 100380 15112 101892
rect 14792 100324 14820 100380
rect 14876 100324 14924 100380
rect 14980 100324 15028 100380
rect 15084 100324 15112 100380
rect 14792 98812 15112 100324
rect 14792 98756 14820 98812
rect 14876 98756 14924 98812
rect 14980 98756 15028 98812
rect 15084 98756 15112 98812
rect 18194 118412 18514 118444
rect 18194 118356 18222 118412
rect 18278 118356 18326 118412
rect 18382 118356 18430 118412
rect 18486 118356 18514 118412
rect 18194 116844 18514 118356
rect 18194 116788 18222 116844
rect 18278 116788 18326 116844
rect 18382 116788 18430 116844
rect 18486 116788 18514 116844
rect 18194 115276 18514 116788
rect 18194 115220 18222 115276
rect 18278 115220 18326 115276
rect 18382 115220 18430 115276
rect 18486 115220 18514 115276
rect 18194 113708 18514 115220
rect 18194 113652 18222 113708
rect 18278 113652 18326 113708
rect 18382 113652 18430 113708
rect 18486 113652 18514 113708
rect 18194 112140 18514 113652
rect 18194 112084 18222 112140
rect 18278 112084 18326 112140
rect 18382 112084 18430 112140
rect 18486 112084 18514 112140
rect 18194 110572 18514 112084
rect 18194 110516 18222 110572
rect 18278 110516 18326 110572
rect 18382 110516 18430 110572
rect 18486 110516 18514 110572
rect 18194 109004 18514 110516
rect 18194 108948 18222 109004
rect 18278 108948 18326 109004
rect 18382 108948 18430 109004
rect 18486 108948 18514 109004
rect 18194 107436 18514 108948
rect 18194 107380 18222 107436
rect 18278 107380 18326 107436
rect 18382 107380 18430 107436
rect 18486 107380 18514 107436
rect 18194 105868 18514 107380
rect 18194 105812 18222 105868
rect 18278 105812 18326 105868
rect 18382 105812 18430 105868
rect 18486 105812 18514 105868
rect 18194 104300 18514 105812
rect 18194 104244 18222 104300
rect 18278 104244 18326 104300
rect 18382 104244 18430 104300
rect 18486 104244 18514 104300
rect 18194 102732 18514 104244
rect 18194 102676 18222 102732
rect 18278 102676 18326 102732
rect 18382 102676 18430 102732
rect 18486 102676 18514 102732
rect 18194 101164 18514 102676
rect 18194 101108 18222 101164
rect 18278 101108 18326 101164
rect 18382 101108 18430 101164
rect 18486 101108 18514 101164
rect 18194 99596 18514 101108
rect 18194 99540 18222 99596
rect 18278 99540 18326 99596
rect 18382 99540 18430 99596
rect 18486 99540 18514 99596
rect 14252 97300 14308 97310
rect 14028 97188 14084 97198
rect 7988 95620 8016 95676
rect 8072 95620 8120 95676
rect 8176 95620 8224 95676
rect 8280 95620 8308 95676
rect 4586 93268 4614 93324
rect 4670 93268 4718 93324
rect 4774 93268 4822 93324
rect 4878 93268 4906 93324
rect 4586 91756 4906 93268
rect 4586 91700 4614 91756
rect 4670 91700 4718 91756
rect 4774 91700 4822 91756
rect 4878 91700 4906 91756
rect 4586 90188 4906 91700
rect 4586 90132 4614 90188
rect 4670 90132 4718 90188
rect 4774 90132 4822 90188
rect 4878 90132 4906 90188
rect 4586 88620 4906 90132
rect 4586 88564 4614 88620
rect 4670 88564 4718 88620
rect 4774 88564 4822 88620
rect 4878 88564 4906 88620
rect 3388 88004 3444 88014
rect 2492 68628 2548 68638
rect 2492 65492 2548 68572
rect 2492 65426 2548 65436
rect 2716 58212 2772 58222
rect 2604 54628 2660 54638
rect 2604 49812 2660 54572
rect 2716 52724 2772 58156
rect 2716 52658 2772 52668
rect 2604 49746 2660 49756
rect 2828 52276 2884 52286
rect 2828 49812 2884 52220
rect 2828 49746 2884 49756
rect 3164 46564 3220 46574
rect 2380 45780 2436 45790
rect 2380 38276 2436 45724
rect 3164 43764 3220 46508
rect 3164 43698 3220 43708
rect 2380 38210 2436 38220
rect 3388 8260 3444 87948
rect 4586 87052 4906 88564
rect 4586 86996 4614 87052
rect 4670 86996 4718 87052
rect 4774 86996 4822 87052
rect 4878 86996 4906 87052
rect 4586 85484 4906 86996
rect 4586 85428 4614 85484
rect 4670 85428 4718 85484
rect 4774 85428 4822 85484
rect 4878 85428 4906 85484
rect 4586 83916 4906 85428
rect 4586 83860 4614 83916
rect 4670 83860 4718 83916
rect 4774 83860 4822 83916
rect 4878 83860 4906 83916
rect 4586 82348 4906 83860
rect 4586 82292 4614 82348
rect 4670 82292 4718 82348
rect 4774 82292 4822 82348
rect 4878 82292 4906 82348
rect 4586 80780 4906 82292
rect 4586 80724 4614 80780
rect 4670 80724 4718 80780
rect 4774 80724 4822 80780
rect 4878 80724 4906 80780
rect 4586 79212 4906 80724
rect 7988 94108 8308 95620
rect 7988 94052 8016 94108
rect 8072 94052 8120 94108
rect 8176 94052 8224 94108
rect 8280 94052 8308 94108
rect 7988 92540 8308 94052
rect 7988 92484 8016 92540
rect 8072 92484 8120 92540
rect 8176 92484 8224 92540
rect 8280 92484 8308 92540
rect 7988 90972 8308 92484
rect 7988 90916 8016 90972
rect 8072 90916 8120 90972
rect 8176 90916 8224 90972
rect 8280 90916 8308 90972
rect 7988 89404 8308 90916
rect 10892 96404 10948 96414
rect 10892 95844 10948 96348
rect 10892 90692 10948 95788
rect 10892 90626 10948 90636
rect 11390 96404 11418 96460
rect 11474 96404 11522 96460
rect 11578 96404 11626 96460
rect 11682 96404 11710 96460
rect 11390 94892 11710 96404
rect 13916 96964 13972 96974
rect 13916 95172 13972 96908
rect 14028 96404 14084 97132
rect 14252 96964 14308 97244
rect 14792 97244 15112 98756
rect 17948 98756 18004 98766
rect 14252 96898 14308 96908
rect 14364 97188 14420 97198
rect 14028 96338 14084 96348
rect 14364 95844 14420 97132
rect 14792 97188 14820 97244
rect 14876 97188 14924 97244
rect 14980 97188 15028 97244
rect 15084 97188 15112 97244
rect 14364 95778 14420 95788
rect 14588 96180 14644 96190
rect 14588 95284 14644 96124
rect 14588 95218 14644 95228
rect 14792 95676 15112 97188
rect 14792 95620 14820 95676
rect 14876 95620 14924 95676
rect 14980 95620 15028 95676
rect 15084 95620 15112 95676
rect 13916 95106 13972 95116
rect 11390 94836 11418 94892
rect 11474 94836 11522 94892
rect 11578 94836 11626 94892
rect 11682 94836 11710 94892
rect 11390 93324 11710 94836
rect 11390 93268 11418 93324
rect 11474 93268 11522 93324
rect 11578 93268 11626 93324
rect 11682 93268 11710 93324
rect 11390 91756 11710 93268
rect 11390 91700 11418 91756
rect 11474 91700 11522 91756
rect 11578 91700 11626 91756
rect 11682 91700 11710 91756
rect 7988 89348 8016 89404
rect 8072 89348 8120 89404
rect 8176 89348 8224 89404
rect 8280 89348 8308 89404
rect 7988 87836 8308 89348
rect 7988 87780 8016 87836
rect 8072 87780 8120 87836
rect 8176 87780 8224 87836
rect 8280 87780 8308 87836
rect 7988 86268 8308 87780
rect 7988 86212 8016 86268
rect 8072 86212 8120 86268
rect 8176 86212 8224 86268
rect 8280 86212 8308 86268
rect 7988 84700 8308 86212
rect 7988 84644 8016 84700
rect 8072 84644 8120 84700
rect 8176 84644 8224 84700
rect 8280 84644 8308 84700
rect 7988 83132 8308 84644
rect 7988 83076 8016 83132
rect 8072 83076 8120 83132
rect 8176 83076 8224 83132
rect 8280 83076 8308 83132
rect 7988 81564 8308 83076
rect 7988 81508 8016 81564
rect 8072 81508 8120 81564
rect 8176 81508 8224 81564
rect 8280 81508 8308 81564
rect 4586 79156 4614 79212
rect 4670 79156 4718 79212
rect 4774 79156 4822 79212
rect 4878 79156 4906 79212
rect 4586 77644 4906 79156
rect 4586 77588 4614 77644
rect 4670 77588 4718 77644
rect 4774 77588 4822 77644
rect 4878 77588 4906 77644
rect 4586 76076 4906 77588
rect 4586 76020 4614 76076
rect 4670 76020 4718 76076
rect 4774 76020 4822 76076
rect 4878 76020 4906 76076
rect 4586 74508 4906 76020
rect 4586 74452 4614 74508
rect 4670 74452 4718 74508
rect 4774 74452 4822 74508
rect 4878 74452 4906 74508
rect 4586 72940 4906 74452
rect 4586 72884 4614 72940
rect 4670 72884 4718 72940
rect 4774 72884 4822 72940
rect 4878 72884 4906 72940
rect 4586 71372 4906 72884
rect 4586 71316 4614 71372
rect 4670 71316 4718 71372
rect 4774 71316 4822 71372
rect 4878 71316 4906 71372
rect 4586 69804 4906 71316
rect 4586 69748 4614 69804
rect 4670 69748 4718 69804
rect 4774 69748 4822 69804
rect 4878 69748 4906 69804
rect 3836 69076 3892 69086
rect 3836 60564 3892 69020
rect 3948 68404 4004 68414
rect 3948 62916 4004 68348
rect 4396 68404 4452 68414
rect 4172 65604 4228 65614
rect 4172 64708 4228 65548
rect 4172 64642 4228 64652
rect 3948 62850 4004 62860
rect 4396 61684 4452 68348
rect 4396 61618 4452 61628
rect 4586 68236 4906 69748
rect 4586 68180 4614 68236
rect 4670 68180 4718 68236
rect 4774 68180 4822 68236
rect 4878 68180 4906 68236
rect 4586 66668 4906 68180
rect 4586 66612 4614 66668
rect 4670 66612 4718 66668
rect 4774 66612 4822 66668
rect 4878 66612 4906 66668
rect 4586 65100 4906 66612
rect 4586 65044 4614 65100
rect 4670 65044 4718 65100
rect 4774 65044 4822 65100
rect 4878 65044 4906 65100
rect 4586 63532 4906 65044
rect 4586 63476 4614 63532
rect 4670 63476 4718 63532
rect 4774 63476 4822 63532
rect 4878 63476 4906 63532
rect 4586 61964 4906 63476
rect 4586 61908 4614 61964
rect 4670 61908 4718 61964
rect 4774 61908 4822 61964
rect 4878 61908 4906 61964
rect 3836 60498 3892 60508
rect 4586 60396 4906 61908
rect 4586 60340 4614 60396
rect 4670 60340 4718 60396
rect 4774 60340 4822 60396
rect 4878 60340 4906 60396
rect 4586 58828 4906 60340
rect 4172 58772 4228 58782
rect 3724 57316 3780 57326
rect 3612 56756 3668 56766
rect 3500 52164 3556 52174
rect 3500 13972 3556 52108
rect 3612 48804 3668 56700
rect 3612 48738 3668 48748
rect 3724 48468 3780 57260
rect 3724 48402 3780 48412
rect 3836 56196 3892 56206
rect 3836 51156 3892 56140
rect 4172 55636 4228 58716
rect 4586 58772 4614 58828
rect 4670 58772 4718 58828
rect 4774 58772 4822 58828
rect 4878 58772 4906 58828
rect 4586 57260 4906 58772
rect 4586 57204 4614 57260
rect 4670 57204 4718 57260
rect 4774 57204 4822 57260
rect 4878 57204 4906 57260
rect 4172 55570 4228 55580
rect 4284 56532 4340 56542
rect 3836 49028 3892 51100
rect 3836 47460 3892 48972
rect 4172 53620 4228 53630
rect 4172 49028 4228 53564
rect 4172 48962 4228 48972
rect 4284 48580 4340 56476
rect 4586 55692 4906 57204
rect 4586 55636 4614 55692
rect 4670 55636 4718 55692
rect 4774 55636 4822 55692
rect 4878 55636 4906 55692
rect 4586 54124 4906 55636
rect 4586 54068 4614 54124
rect 4670 54068 4718 54124
rect 4774 54068 4822 54124
rect 4878 54068 4906 54124
rect 4284 48514 4340 48524
rect 4396 53060 4452 53070
rect 3836 47394 3892 47404
rect 4060 46788 4116 46798
rect 3724 44772 3780 44782
rect 3612 44548 3668 44558
rect 3612 34692 3668 44492
rect 3724 38948 3780 44716
rect 3724 38882 3780 38892
rect 3836 44660 3892 44670
rect 3836 36148 3892 44604
rect 3836 36082 3892 36092
rect 4060 36036 4116 46732
rect 4172 46676 4228 46686
rect 4172 40852 4228 46620
rect 4172 40180 4228 40796
rect 4172 38052 4228 40124
rect 4172 37986 4228 37996
rect 4060 35970 4116 35980
rect 3612 34626 3668 34636
rect 4396 18452 4452 53004
rect 4396 18386 4452 18396
rect 4586 52556 4906 54068
rect 4586 52500 4614 52556
rect 4670 52500 4718 52556
rect 4774 52500 4822 52556
rect 4878 52500 4906 52556
rect 4586 50988 4906 52500
rect 4586 50932 4614 50988
rect 4670 50932 4718 50988
rect 4774 50932 4822 50988
rect 4878 50932 4906 50988
rect 4586 49420 4906 50932
rect 4586 49364 4614 49420
rect 4670 49364 4718 49420
rect 4774 49364 4822 49420
rect 4878 49364 4906 49420
rect 4586 47852 4906 49364
rect 4586 47796 4614 47852
rect 4670 47796 4718 47852
rect 4774 47796 4822 47852
rect 4878 47796 4906 47852
rect 4586 46284 4906 47796
rect 4586 46228 4614 46284
rect 4670 46228 4718 46284
rect 4774 46228 4822 46284
rect 4878 46228 4906 46284
rect 4586 44716 4906 46228
rect 4586 44660 4614 44716
rect 4670 44660 4718 44716
rect 4774 44660 4822 44716
rect 4878 44660 4906 44716
rect 4586 43148 4906 44660
rect 4586 43092 4614 43148
rect 4670 43092 4718 43148
rect 4774 43092 4822 43148
rect 4878 43092 4906 43148
rect 4586 41580 4906 43092
rect 4586 41524 4614 41580
rect 4670 41524 4718 41580
rect 4774 41524 4822 41580
rect 4878 41524 4906 41580
rect 4586 40012 4906 41524
rect 4586 39956 4614 40012
rect 4670 39956 4718 40012
rect 4774 39956 4822 40012
rect 4878 39956 4906 40012
rect 4586 38444 4906 39956
rect 4586 38388 4614 38444
rect 4670 38388 4718 38444
rect 4774 38388 4822 38444
rect 4878 38388 4906 38444
rect 4586 36876 4906 38388
rect 4586 36820 4614 36876
rect 4670 36820 4718 36876
rect 4774 36820 4822 36876
rect 4878 36820 4906 36876
rect 4586 35308 4906 36820
rect 4586 35252 4614 35308
rect 4670 35252 4718 35308
rect 4774 35252 4822 35308
rect 4878 35252 4906 35308
rect 4586 33740 4906 35252
rect 4586 33684 4614 33740
rect 4670 33684 4718 33740
rect 4774 33684 4822 33740
rect 4878 33684 4906 33740
rect 4586 32172 4906 33684
rect 4586 32116 4614 32172
rect 4670 32116 4718 32172
rect 4774 32116 4822 32172
rect 4878 32116 4906 32172
rect 4586 30604 4906 32116
rect 4586 30548 4614 30604
rect 4670 30548 4718 30604
rect 4774 30548 4822 30604
rect 4878 30548 4906 30604
rect 4586 29036 4906 30548
rect 4586 28980 4614 29036
rect 4670 28980 4718 29036
rect 4774 28980 4822 29036
rect 4878 28980 4906 29036
rect 4586 27468 4906 28980
rect 5068 80052 5124 80062
rect 5068 28532 5124 79996
rect 7988 79996 8308 81508
rect 7988 79940 8016 79996
rect 8072 79940 8120 79996
rect 8176 79940 8224 79996
rect 8280 79940 8308 79996
rect 7988 78428 8308 79940
rect 7988 78372 8016 78428
rect 8072 78372 8120 78428
rect 8176 78372 8224 78428
rect 8280 78372 8308 78428
rect 7988 76860 8308 78372
rect 11390 90188 11710 91700
rect 11390 90132 11418 90188
rect 11474 90132 11522 90188
rect 11578 90132 11626 90188
rect 11682 90132 11710 90188
rect 11390 88620 11710 90132
rect 11390 88564 11418 88620
rect 11474 88564 11522 88620
rect 11578 88564 11626 88620
rect 11682 88564 11710 88620
rect 11390 87052 11710 88564
rect 11390 86996 11418 87052
rect 11474 86996 11522 87052
rect 11578 86996 11626 87052
rect 11682 86996 11710 87052
rect 11390 85484 11710 86996
rect 11390 85428 11418 85484
rect 11474 85428 11522 85484
rect 11578 85428 11626 85484
rect 11682 85428 11710 85484
rect 11390 83916 11710 85428
rect 11390 83860 11418 83916
rect 11474 83860 11522 83916
rect 11578 83860 11626 83916
rect 11682 83860 11710 83916
rect 11390 82348 11710 83860
rect 11390 82292 11418 82348
rect 11474 82292 11522 82348
rect 11578 82292 11626 82348
rect 11682 82292 11710 82348
rect 11390 80780 11710 82292
rect 14792 94108 15112 95620
rect 14792 94052 14820 94108
rect 14876 94052 14924 94108
rect 14980 94052 15028 94108
rect 15084 94052 15112 94108
rect 14792 92540 15112 94052
rect 15260 97748 15316 97758
rect 15260 94052 15316 97692
rect 17948 96852 18004 98700
rect 18060 98532 18116 98542
rect 18060 97636 18116 98476
rect 18060 97570 18116 97580
rect 18194 98028 18514 99540
rect 18194 97972 18222 98028
rect 18278 97972 18326 98028
rect 18382 97972 18430 98028
rect 18486 97972 18514 98028
rect 17948 96786 18004 96796
rect 18194 96460 18514 97972
rect 18194 96404 18222 96460
rect 18278 96404 18326 96460
rect 18382 96404 18430 96460
rect 18486 96404 18514 96460
rect 18194 94892 18514 96404
rect 21596 117628 21916 118444
rect 21596 117572 21624 117628
rect 21680 117572 21728 117628
rect 21784 117572 21832 117628
rect 21888 117572 21916 117628
rect 21596 116060 21916 117572
rect 21596 116004 21624 116060
rect 21680 116004 21728 116060
rect 21784 116004 21832 116060
rect 21888 116004 21916 116060
rect 21596 114492 21916 116004
rect 21596 114436 21624 114492
rect 21680 114436 21728 114492
rect 21784 114436 21832 114492
rect 21888 114436 21916 114492
rect 21596 112924 21916 114436
rect 21596 112868 21624 112924
rect 21680 112868 21728 112924
rect 21784 112868 21832 112924
rect 21888 112868 21916 112924
rect 21596 111356 21916 112868
rect 21596 111300 21624 111356
rect 21680 111300 21728 111356
rect 21784 111300 21832 111356
rect 21888 111300 21916 111356
rect 21596 109788 21916 111300
rect 21596 109732 21624 109788
rect 21680 109732 21728 109788
rect 21784 109732 21832 109788
rect 21888 109732 21916 109788
rect 21596 108220 21916 109732
rect 21596 108164 21624 108220
rect 21680 108164 21728 108220
rect 21784 108164 21832 108220
rect 21888 108164 21916 108220
rect 21596 106652 21916 108164
rect 21596 106596 21624 106652
rect 21680 106596 21728 106652
rect 21784 106596 21832 106652
rect 21888 106596 21916 106652
rect 21596 105084 21916 106596
rect 24998 118412 25318 118444
rect 24998 118356 25026 118412
rect 25082 118356 25130 118412
rect 25186 118356 25234 118412
rect 25290 118356 25318 118412
rect 24998 116844 25318 118356
rect 24998 116788 25026 116844
rect 25082 116788 25130 116844
rect 25186 116788 25234 116844
rect 25290 116788 25318 116844
rect 24998 115276 25318 116788
rect 24998 115220 25026 115276
rect 25082 115220 25130 115276
rect 25186 115220 25234 115276
rect 25290 115220 25318 115276
rect 24998 113708 25318 115220
rect 24998 113652 25026 113708
rect 25082 113652 25130 113708
rect 25186 113652 25234 113708
rect 25290 113652 25318 113708
rect 24998 112140 25318 113652
rect 24998 112084 25026 112140
rect 25082 112084 25130 112140
rect 25186 112084 25234 112140
rect 25290 112084 25318 112140
rect 24998 110572 25318 112084
rect 24998 110516 25026 110572
rect 25082 110516 25130 110572
rect 25186 110516 25234 110572
rect 25290 110516 25318 110572
rect 24998 109004 25318 110516
rect 24998 108948 25026 109004
rect 25082 108948 25130 109004
rect 25186 108948 25234 109004
rect 25290 108948 25318 109004
rect 24998 107436 25318 108948
rect 24998 107380 25026 107436
rect 25082 107380 25130 107436
rect 25186 107380 25234 107436
rect 25290 107380 25318 107436
rect 24998 105868 25318 107380
rect 24998 105812 25026 105868
rect 25082 105812 25130 105868
rect 25186 105812 25234 105868
rect 25290 105812 25318 105868
rect 21596 105028 21624 105084
rect 21680 105028 21728 105084
rect 21784 105028 21832 105084
rect 21888 105028 21916 105084
rect 21596 103516 21916 105028
rect 21596 103460 21624 103516
rect 21680 103460 21728 103516
rect 21784 103460 21832 103516
rect 21888 103460 21916 103516
rect 21596 101948 21916 103460
rect 21596 101892 21624 101948
rect 21680 101892 21728 101948
rect 21784 101892 21832 101948
rect 21888 101892 21916 101948
rect 21596 100380 21916 101892
rect 21596 100324 21624 100380
rect 21680 100324 21728 100380
rect 21784 100324 21832 100380
rect 21888 100324 21916 100380
rect 21596 98812 21916 100324
rect 21596 98756 21624 98812
rect 21680 98756 21728 98812
rect 21784 98756 21832 98812
rect 21888 98756 21916 98812
rect 21596 97244 21916 98756
rect 24444 105700 24500 105710
rect 24444 97412 24500 105644
rect 24444 97346 24500 97356
rect 24998 104300 25318 105812
rect 24998 104244 25026 104300
rect 25082 104244 25130 104300
rect 25186 104244 25234 104300
rect 25290 104244 25318 104300
rect 24998 102732 25318 104244
rect 24998 102676 25026 102732
rect 25082 102676 25130 102732
rect 25186 102676 25234 102732
rect 25290 102676 25318 102732
rect 24998 101164 25318 102676
rect 24998 101108 25026 101164
rect 25082 101108 25130 101164
rect 25186 101108 25234 101164
rect 25290 101108 25318 101164
rect 24998 99596 25318 101108
rect 24998 99540 25026 99596
rect 25082 99540 25130 99596
rect 25186 99540 25234 99596
rect 25290 99540 25318 99596
rect 24998 98028 25318 99540
rect 24998 97972 25026 98028
rect 25082 97972 25130 98028
rect 25186 97972 25234 98028
rect 25290 97972 25318 98028
rect 21596 97188 21624 97244
rect 21680 97188 21728 97244
rect 21784 97188 21832 97244
rect 21888 97188 21916 97244
rect 21596 95676 21916 97188
rect 21596 95620 21624 95676
rect 21680 95620 21728 95676
rect 21784 95620 21832 95676
rect 21888 95620 21916 95676
rect 18194 94836 18222 94892
rect 18278 94836 18326 94892
rect 18382 94836 18430 94892
rect 18486 94836 18514 94892
rect 15260 93986 15316 93996
rect 15372 94276 15428 94286
rect 15372 93898 15428 94220
rect 15260 93842 15428 93898
rect 15596 93940 15652 93950
rect 15260 93828 15316 93842
rect 15260 93762 15316 93772
rect 14792 92484 14820 92540
rect 14876 92484 14924 92540
rect 14980 92484 15028 92540
rect 15084 92484 15112 92540
rect 14792 90972 15112 92484
rect 15596 93268 15652 93884
rect 14792 90916 14820 90972
rect 14876 90916 14924 90972
rect 14980 90916 15028 90972
rect 15084 90916 15112 90972
rect 14792 89404 15112 90916
rect 14792 89348 14820 89404
rect 14876 89348 14924 89404
rect 14980 89348 15028 89404
rect 15084 89348 15112 89404
rect 14792 87836 15112 89348
rect 15372 91476 15428 91486
rect 15372 89236 15428 91420
rect 15372 89170 15428 89180
rect 14792 87780 14820 87836
rect 14876 87780 14924 87836
rect 14980 87780 15028 87836
rect 15084 87780 15112 87836
rect 14792 86268 15112 87780
rect 14792 86212 14820 86268
rect 14876 86212 14924 86268
rect 14980 86212 15028 86268
rect 15084 86212 15112 86268
rect 15484 88116 15540 88126
rect 15484 86324 15540 88060
rect 15596 87668 15652 93212
rect 18194 93324 18514 94836
rect 19068 95172 19124 95182
rect 19068 94500 19124 95116
rect 19068 94434 19124 94444
rect 19740 94724 19796 94734
rect 18194 93268 18222 93324
rect 18278 93268 18326 93324
rect 18382 93268 18430 93324
rect 18486 93268 18514 93324
rect 17836 92372 17892 92382
rect 15596 87602 15652 87612
rect 15708 89124 15764 89134
rect 15484 86258 15540 86268
rect 14792 84700 15112 86212
rect 15708 85988 15764 89068
rect 17836 88004 17892 92316
rect 17836 87938 17892 87948
rect 18194 91756 18514 93268
rect 18194 91700 18222 91756
rect 18278 91700 18326 91756
rect 18382 91700 18430 91756
rect 18486 91700 18514 91756
rect 18194 90188 18514 91700
rect 18194 90132 18222 90188
rect 18278 90132 18326 90188
rect 18382 90132 18430 90188
rect 18486 90132 18514 90188
rect 18194 88620 18514 90132
rect 19740 88788 19796 94668
rect 21596 94108 21916 95620
rect 21596 94052 21624 94108
rect 21680 94052 21728 94108
rect 21784 94052 21832 94108
rect 21888 94052 21916 94108
rect 20524 93716 20580 93726
rect 19740 88722 19796 88732
rect 20188 92708 20244 92718
rect 18194 88564 18222 88620
rect 18278 88564 18326 88620
rect 18382 88564 18430 88620
rect 18486 88564 18514 88620
rect 15708 85922 15764 85932
rect 18194 87052 18514 88564
rect 18194 86996 18222 87052
rect 18278 86996 18326 87052
rect 18382 86996 18430 87052
rect 18486 86996 18514 87052
rect 14792 84644 14820 84700
rect 14876 84644 14924 84700
rect 14980 84644 15028 84700
rect 15084 84644 15112 84700
rect 14792 83132 15112 84644
rect 14792 83076 14820 83132
rect 14876 83076 14924 83132
rect 14980 83076 15028 83132
rect 15084 83076 15112 83132
rect 14792 81564 15112 83076
rect 18194 85484 18514 86996
rect 18194 85428 18222 85484
rect 18278 85428 18326 85484
rect 18382 85428 18430 85484
rect 18486 85428 18514 85484
rect 18194 83916 18514 85428
rect 18194 83860 18222 83916
rect 18278 83860 18326 83916
rect 18382 83860 18430 83916
rect 18486 83860 18514 83916
rect 20188 83972 20244 92652
rect 20188 83906 20244 83916
rect 14792 81508 14820 81564
rect 14876 81508 14924 81564
rect 14980 81508 15028 81564
rect 15084 81508 15112 81564
rect 11390 80724 11418 80780
rect 11474 80724 11522 80780
rect 11578 80724 11626 80780
rect 11682 80724 11710 80780
rect 11390 79212 11710 80724
rect 11390 79156 11418 79212
rect 11474 79156 11522 79212
rect 11578 79156 11626 79212
rect 11682 79156 11710 79212
rect 7988 76804 8016 76860
rect 8072 76804 8120 76860
rect 8176 76804 8224 76860
rect 8280 76804 8308 76860
rect 7988 75292 8308 76804
rect 7988 75236 8016 75292
rect 8072 75236 8120 75292
rect 8176 75236 8224 75292
rect 8280 75236 8308 75292
rect 7988 73724 8308 75236
rect 7988 73668 8016 73724
rect 8072 73668 8120 73724
rect 8176 73668 8224 73724
rect 8280 73668 8308 73724
rect 7988 72156 8308 73668
rect 9100 77700 9156 77710
rect 9100 72324 9156 77644
rect 11390 77644 11710 79156
rect 12796 80948 12852 80958
rect 11390 77588 11418 77644
rect 11474 77588 11522 77644
rect 11578 77588 11626 77644
rect 11682 77588 11710 77644
rect 11390 76076 11710 77588
rect 11390 76020 11418 76076
rect 11474 76020 11522 76076
rect 11578 76020 11626 76076
rect 11682 76020 11710 76076
rect 11228 75124 11284 75134
rect 11228 74228 11284 75068
rect 11228 74162 11284 74172
rect 11390 74508 11710 76020
rect 11390 74452 11418 74508
rect 11474 74452 11522 74508
rect 11578 74452 11626 74508
rect 11682 74452 11710 74508
rect 9100 72258 9156 72268
rect 11390 72940 11710 74452
rect 12572 78820 12628 78830
rect 12572 74116 12628 78764
rect 12572 74050 12628 74060
rect 11390 72884 11418 72940
rect 11474 72884 11522 72940
rect 11578 72884 11626 72940
rect 11682 72884 11710 72940
rect 7988 72100 8016 72156
rect 8072 72100 8120 72156
rect 8176 72100 8224 72156
rect 8280 72100 8308 72156
rect 7988 70588 8308 72100
rect 7988 70532 8016 70588
rect 8072 70532 8120 70588
rect 8176 70532 8224 70588
rect 8280 70532 8308 70588
rect 7988 69020 8308 70532
rect 11390 71372 11710 72884
rect 12796 72772 12852 80892
rect 14028 80612 14084 80622
rect 12796 72706 12852 72716
rect 13692 75460 13748 75470
rect 12012 72212 12068 72222
rect 12012 71876 12068 72156
rect 12012 71810 12068 71820
rect 11390 71316 11418 71372
rect 11474 71316 11522 71372
rect 11578 71316 11626 71372
rect 11682 71316 11710 71372
rect 9436 69860 9492 69870
rect 9436 69188 9492 69804
rect 11390 69804 11710 71316
rect 13692 70980 13748 75404
rect 14028 74676 14084 80556
rect 14792 79996 15112 81508
rect 14792 79940 14820 79996
rect 14876 79940 14924 79996
rect 14980 79940 15028 79996
rect 15084 79940 15112 79996
rect 14588 79716 14644 79726
rect 14252 79156 14308 79166
rect 13692 70914 13748 70924
rect 13804 74004 13860 74014
rect 13804 70868 13860 73948
rect 13916 73332 13972 73342
rect 13916 71204 13972 73276
rect 13916 71138 13972 71148
rect 13804 70802 13860 70812
rect 11390 69748 11418 69804
rect 11474 69748 11522 69804
rect 11578 69748 11626 69804
rect 11682 69748 11710 69804
rect 9436 69122 9492 69132
rect 11228 69188 11284 69198
rect 7988 68964 8016 69020
rect 8072 68964 8120 69020
rect 8176 68964 8224 69020
rect 8280 68964 8308 69020
rect 7988 67452 8308 68964
rect 7988 67396 8016 67452
rect 8072 67396 8120 67452
rect 8176 67396 8224 67452
rect 8280 67396 8308 67452
rect 7988 65884 8308 67396
rect 7988 65828 8016 65884
rect 8072 65828 8120 65884
rect 8176 65828 8224 65884
rect 8280 65828 8308 65884
rect 7988 64316 8308 65828
rect 7988 64260 8016 64316
rect 8072 64260 8120 64316
rect 8176 64260 8224 64316
rect 8280 64260 8308 64316
rect 7988 62748 8308 64260
rect 9660 67844 9716 67854
rect 9660 63700 9716 67788
rect 10892 67732 10948 67742
rect 9660 63634 9716 63644
rect 10780 67060 10836 67070
rect 7988 62692 8016 62748
rect 8072 62692 8120 62748
rect 8176 62692 8224 62748
rect 8280 62692 8308 62748
rect 7988 61180 8308 62692
rect 7988 61124 8016 61180
rect 8072 61124 8120 61180
rect 8176 61124 8224 61180
rect 8280 61124 8308 61180
rect 7988 59612 8308 61124
rect 7988 59556 8016 59612
rect 8072 59556 8120 59612
rect 8176 59556 8224 59612
rect 8280 59556 8308 59612
rect 7988 58044 8308 59556
rect 10780 58884 10836 67004
rect 10780 58818 10836 58828
rect 5852 57988 5908 57998
rect 5404 56980 5460 56990
rect 5292 56756 5348 56766
rect 5292 51044 5348 56700
rect 5292 50978 5348 50988
rect 5404 50932 5460 56924
rect 5404 50866 5460 50876
rect 5516 56756 5572 56766
rect 5516 47684 5572 56700
rect 5852 56756 5908 57932
rect 7988 57988 8016 58044
rect 8072 57988 8120 58044
rect 8176 57988 8224 58044
rect 8280 57988 8308 58044
rect 5740 53060 5796 53070
rect 5740 52500 5796 53004
rect 5740 52434 5796 52444
rect 5852 51380 5908 56700
rect 6300 57764 6356 57774
rect 6300 53620 6356 57708
rect 6636 56532 6692 56542
rect 6300 53554 6356 53564
rect 6412 54404 6468 54414
rect 6412 54068 6468 54348
rect 5852 51314 5908 51324
rect 5964 51604 6020 51614
rect 5516 47618 5572 47628
rect 5964 47068 6020 51548
rect 6188 51268 6244 51278
rect 6188 48804 6244 51212
rect 6412 50036 6468 54012
rect 6636 53844 6692 56476
rect 6636 53778 6692 53788
rect 7988 56476 8308 57988
rect 7988 56420 8016 56476
rect 8072 56420 8120 56476
rect 8176 56420 8224 56476
rect 8280 56420 8308 56476
rect 7988 54908 8308 56420
rect 7988 54852 8016 54908
rect 8072 54852 8120 54908
rect 8176 54852 8224 54908
rect 8280 54852 8308 54908
rect 7988 53340 8308 54852
rect 8876 58324 8932 58334
rect 8540 54516 8596 54526
rect 7988 53284 8016 53340
rect 8072 53284 8120 53340
rect 8176 53284 8224 53340
rect 8280 53284 8308 53340
rect 7420 52388 7476 52398
rect 7420 50596 7476 52332
rect 7420 50530 7476 50540
rect 7532 52052 7588 52062
rect 6412 49970 6468 49980
rect 6188 48738 6244 48748
rect 7532 48468 7588 51996
rect 7532 48402 7588 48412
rect 7988 51772 8308 53284
rect 7988 51716 8016 51772
rect 8072 51716 8120 51772
rect 8176 51716 8224 51772
rect 8280 51716 8308 51772
rect 7988 50204 8308 51716
rect 7988 50148 8016 50204
rect 8072 50148 8120 50204
rect 8176 50148 8224 50204
rect 8280 50148 8308 50204
rect 8428 53620 8484 53630
rect 8428 50260 8484 53564
rect 8428 50194 8484 50204
rect 7988 48636 8308 50148
rect 7988 48580 8016 48636
rect 8072 48580 8120 48636
rect 8176 48580 8224 48636
rect 8280 48580 8308 48636
rect 7988 47068 8308 48580
rect 8540 48356 8596 54460
rect 8876 53172 8932 58268
rect 8876 53106 8932 53116
rect 9548 58324 9604 58334
rect 9548 53172 9604 58268
rect 10556 58324 10612 58334
rect 9548 53106 9604 53116
rect 10108 57876 10164 57886
rect 10108 53060 10164 57820
rect 10332 56196 10388 56206
rect 10332 54180 10388 56140
rect 10332 54114 10388 54124
rect 10444 54292 10500 54302
rect 10108 52052 10164 53004
rect 10108 51986 10164 51996
rect 10332 52948 10388 52958
rect 8540 48290 8596 48300
rect 9772 49588 9828 49598
rect 5964 47012 6132 47068
rect 5180 46788 5236 46798
rect 5180 37492 5236 46732
rect 5852 46564 5908 46574
rect 5852 44324 5908 46508
rect 5852 44258 5908 44268
rect 5964 44212 6020 44222
rect 5740 43540 5796 43550
rect 5740 38500 5796 43484
rect 5964 43428 6020 44156
rect 5964 43362 6020 43372
rect 6076 39396 6132 47012
rect 7988 47012 8016 47068
rect 8072 47012 8120 47068
rect 8176 47012 8224 47068
rect 8280 47012 8308 47068
rect 9772 47684 9828 49532
rect 9772 47068 9828 47628
rect 10220 47796 10276 47806
rect 10220 47124 10276 47740
rect 9996 47068 10052 47078
rect 9772 47012 9996 47068
rect 10220 47058 10276 47068
rect 7868 46228 7924 46238
rect 7084 46116 7140 46126
rect 6076 39330 6132 39340
rect 6188 45556 6244 45566
rect 5740 38434 5796 38444
rect 5180 37426 5236 37436
rect 6188 36148 6244 45500
rect 6748 45444 6804 45454
rect 6748 43988 6804 45388
rect 6748 43922 6804 43932
rect 6972 45444 7028 45454
rect 6972 36708 7028 45388
rect 7084 40292 7140 46060
rect 7644 45444 7700 45454
rect 7084 40226 7140 40236
rect 7196 44436 7252 44446
rect 7196 37716 7252 44380
rect 7644 38836 7700 45388
rect 7868 41972 7924 46172
rect 7868 41906 7924 41916
rect 7988 45500 8308 47012
rect 9996 47002 10052 47012
rect 10332 46788 10388 52892
rect 10444 48692 10500 54236
rect 10444 48626 10500 48636
rect 10444 48468 10500 48478
rect 10444 47236 10500 48412
rect 10556 47684 10612 58268
rect 10780 57204 10836 57214
rect 10556 47618 10612 47628
rect 10668 55076 10724 55086
rect 10444 47170 10500 47180
rect 10332 46722 10388 46732
rect 7988 45444 8016 45500
rect 8072 45444 8120 45500
rect 8176 45444 8224 45500
rect 8280 45444 8308 45500
rect 7988 43932 8308 45444
rect 7988 43876 8016 43932
rect 8072 43876 8120 43932
rect 8176 43876 8224 43932
rect 8280 43876 8308 43932
rect 7988 42364 8308 43876
rect 7988 42308 8016 42364
rect 8072 42308 8120 42364
rect 8176 42308 8224 42364
rect 8280 42308 8308 42364
rect 7644 38770 7700 38780
rect 7868 40852 7924 40862
rect 7196 37650 7252 37660
rect 6972 36642 7028 36652
rect 6188 36082 6244 36092
rect 7868 35700 7924 40796
rect 7868 35634 7924 35644
rect 7988 40796 8308 42308
rect 7988 40740 8016 40796
rect 8072 40740 8120 40796
rect 8176 40740 8224 40796
rect 8280 40740 8308 40796
rect 7988 39228 8308 40740
rect 9660 45556 9716 45566
rect 9660 43428 9716 45500
rect 9660 40628 9716 43372
rect 10444 44548 10500 44558
rect 10332 43092 10388 43102
rect 9660 40562 9716 40572
rect 9884 42420 9940 42430
rect 9884 41860 9940 42364
rect 7988 39172 8016 39228
rect 8072 39172 8120 39228
rect 8176 39172 8224 39228
rect 8280 39172 8308 39228
rect 7988 37660 8308 39172
rect 7988 37604 8016 37660
rect 8072 37604 8120 37660
rect 8176 37604 8224 37660
rect 8280 37604 8308 37660
rect 7988 36092 8308 37604
rect 9884 36820 9940 41804
rect 10332 41860 10388 43036
rect 10332 41794 10388 41804
rect 10444 36932 10500 44492
rect 10556 43876 10612 43886
rect 10556 42420 10612 43820
rect 10556 42354 10612 42364
rect 10444 36866 10500 36876
rect 9884 36754 9940 36764
rect 7988 36036 8016 36092
rect 8072 36036 8120 36092
rect 8176 36036 8224 36092
rect 8280 36036 8308 36092
rect 7988 34524 8308 36036
rect 7988 34468 8016 34524
rect 8072 34468 8120 34524
rect 8176 34468 8224 34524
rect 8280 34468 8308 34524
rect 5180 33348 5236 33358
rect 5180 28868 5236 33292
rect 7988 32956 8308 34468
rect 10444 34916 10500 34926
rect 7988 32900 8016 32956
rect 8072 32900 8120 32956
rect 8176 32900 8224 32956
rect 8280 32900 8308 32956
rect 7988 31388 8308 32900
rect 5180 28802 5236 28812
rect 7644 31332 7700 31342
rect 5068 28466 5124 28476
rect 4586 27412 4614 27468
rect 4670 27412 4718 27468
rect 4774 27412 4822 27468
rect 4878 27412 4906 27468
rect 4586 25900 4906 27412
rect 7644 27300 7700 31276
rect 7644 27234 7700 27244
rect 7988 31332 8016 31388
rect 8072 31332 8120 31388
rect 8176 31332 8224 31388
rect 8280 31332 8308 31388
rect 7988 29820 8308 31332
rect 7988 29764 8016 29820
rect 8072 29764 8120 29820
rect 8176 29764 8224 29820
rect 8280 29764 8308 29820
rect 7988 28252 8308 29764
rect 8540 33684 8596 33694
rect 8540 29092 8596 33628
rect 8540 29026 8596 29036
rect 9212 32788 9268 32798
rect 7988 28196 8016 28252
rect 8072 28196 8120 28252
rect 8176 28196 8224 28252
rect 8280 28196 8308 28252
rect 4586 25844 4614 25900
rect 4670 25844 4718 25900
rect 4774 25844 4822 25900
rect 4878 25844 4906 25900
rect 4586 24332 4906 25844
rect 4586 24276 4614 24332
rect 4670 24276 4718 24332
rect 4774 24276 4822 24332
rect 4878 24276 4906 24332
rect 4586 22764 4906 24276
rect 4586 22708 4614 22764
rect 4670 22708 4718 22764
rect 4774 22708 4822 22764
rect 4878 22708 4906 22764
rect 4586 21196 4906 22708
rect 4586 21140 4614 21196
rect 4670 21140 4718 21196
rect 4774 21140 4822 21196
rect 4878 21140 4906 21196
rect 4586 19628 4906 21140
rect 7988 26684 8308 28196
rect 7988 26628 8016 26684
rect 8072 26628 8120 26684
rect 8176 26628 8224 26684
rect 8280 26628 8308 26684
rect 7988 25116 8308 26628
rect 7988 25060 8016 25116
rect 8072 25060 8120 25116
rect 8176 25060 8224 25116
rect 8280 25060 8308 25116
rect 7988 23548 8308 25060
rect 9212 23716 9268 32732
rect 9772 27188 9828 27198
rect 9772 24388 9828 27132
rect 9772 24322 9828 24332
rect 10444 24052 10500 34860
rect 10556 33572 10612 33582
rect 10556 33348 10612 33516
rect 10556 33282 10612 33292
rect 10556 28756 10612 28766
rect 10556 27412 10612 28700
rect 10556 27346 10612 27356
rect 10444 23986 10500 23996
rect 9212 23650 9268 23660
rect 7988 23492 8016 23548
rect 8072 23492 8120 23548
rect 8176 23492 8224 23548
rect 8280 23492 8308 23548
rect 7988 21980 8308 23492
rect 7988 21924 8016 21980
rect 8072 21924 8120 21980
rect 8176 21924 8224 21980
rect 8280 21924 8308 21980
rect 4586 19572 4614 19628
rect 4670 19572 4718 19628
rect 4774 19572 4822 19628
rect 4878 19572 4906 19628
rect 3500 13906 3556 13916
rect 4586 18060 4906 19572
rect 4586 18004 4614 18060
rect 4670 18004 4718 18060
rect 4774 18004 4822 18060
rect 4878 18004 4906 18060
rect 4586 16492 4906 18004
rect 7084 20692 7140 20702
rect 4586 16436 4614 16492
rect 4670 16436 4718 16492
rect 4774 16436 4822 16492
rect 4878 16436 4906 16492
rect 4586 14924 4906 16436
rect 4586 14868 4614 14924
rect 4670 14868 4718 14924
rect 4774 14868 4822 14924
rect 4878 14868 4906 14924
rect 3388 8194 3444 8204
rect 4586 13356 4906 14868
rect 5852 16772 5908 16782
rect 5852 14308 5908 16716
rect 5852 14242 5908 14252
rect 4586 13300 4614 13356
rect 4670 13300 4718 13356
rect 4774 13300 4822 13356
rect 4878 13300 4906 13356
rect 4586 11788 4906 13300
rect 7084 13188 7140 20636
rect 7084 13122 7140 13132
rect 7988 20412 8308 21924
rect 7988 20356 8016 20412
rect 8072 20356 8120 20412
rect 8176 20356 8224 20412
rect 8280 20356 8308 20412
rect 7988 18844 8308 20356
rect 7988 18788 8016 18844
rect 8072 18788 8120 18844
rect 8176 18788 8224 18844
rect 8280 18788 8308 18844
rect 7988 17276 8308 18788
rect 7988 17220 8016 17276
rect 8072 17220 8120 17276
rect 8176 17220 8224 17276
rect 8280 17220 8308 17276
rect 7988 15708 8308 17220
rect 7988 15652 8016 15708
rect 8072 15652 8120 15708
rect 8176 15652 8224 15708
rect 8280 15652 8308 15708
rect 7988 14140 8308 15652
rect 10668 15428 10724 55020
rect 10780 51492 10836 57148
rect 10780 51426 10836 51436
rect 10780 51156 10836 51166
rect 10780 49364 10836 51100
rect 10780 49298 10836 49308
rect 10780 48132 10836 48142
rect 10780 47572 10836 48076
rect 10780 47506 10836 47516
rect 10892 44324 10948 67676
rect 11228 62692 11284 69132
rect 11228 60900 11284 62636
rect 11228 60834 11284 60844
rect 11390 68236 11710 69748
rect 13244 70644 13300 70654
rect 13244 69412 13300 70588
rect 13244 69346 13300 69356
rect 11390 68180 11418 68236
rect 11474 68180 11522 68236
rect 11578 68180 11626 68236
rect 11682 68180 11710 68236
rect 11390 66668 11710 68180
rect 14028 69188 14084 74620
rect 14140 76468 14196 76478
rect 14140 71398 14196 76412
rect 14252 71540 14308 79100
rect 14588 79044 14644 79660
rect 14476 78820 14532 78830
rect 14476 78484 14532 78764
rect 14476 78418 14532 78428
rect 14252 71474 14308 71484
rect 14364 74788 14420 74798
rect 14140 71342 14308 71398
rect 14140 71204 14196 71214
rect 14140 70868 14196 71148
rect 14140 70802 14196 70812
rect 14252 70756 14308 71342
rect 14252 70690 14308 70700
rect 14364 70644 14420 74732
rect 14364 70578 14420 70588
rect 14476 72660 14532 72670
rect 13916 67620 13972 67630
rect 13468 67172 13524 67182
rect 11390 66612 11418 66668
rect 11474 66612 11522 66668
rect 11578 66612 11626 66668
rect 11682 66612 11710 66668
rect 11390 65100 11710 66612
rect 11390 65044 11418 65100
rect 11474 65044 11522 65100
rect 11578 65044 11626 65100
rect 11682 65044 11710 65100
rect 11390 63532 11710 65044
rect 11390 63476 11418 63532
rect 11474 63476 11522 63532
rect 11578 63476 11626 63532
rect 11682 63476 11710 63532
rect 11390 61964 11710 63476
rect 11390 61908 11418 61964
rect 11474 61908 11522 61964
rect 11578 61908 11626 61964
rect 11682 61908 11710 61964
rect 11390 60396 11710 61908
rect 12796 66836 12852 66846
rect 12796 61348 12852 66780
rect 13468 65604 13524 67116
rect 13468 64484 13524 65548
rect 13468 64418 13524 64428
rect 13580 66500 13636 66510
rect 13356 64372 13412 64382
rect 13356 61460 13412 64316
rect 13580 63700 13636 66444
rect 13580 63634 13636 63644
rect 13356 61394 13412 61404
rect 12796 61282 12852 61292
rect 11390 60340 11418 60396
rect 11474 60340 11522 60396
rect 11578 60340 11626 60396
rect 11682 60340 11710 60396
rect 11390 58828 11710 60340
rect 11390 58772 11418 58828
rect 11474 58772 11522 58828
rect 11578 58772 11626 58828
rect 11682 58772 11710 58828
rect 11390 57260 11710 58772
rect 11390 57204 11418 57260
rect 11474 57204 11522 57260
rect 11578 57204 11626 57260
rect 11682 57204 11710 57260
rect 11116 56308 11172 56318
rect 11004 53508 11060 53518
rect 11004 52164 11060 53452
rect 11116 53060 11172 56252
rect 11116 52994 11172 53004
rect 11390 55692 11710 57204
rect 11390 55636 11418 55692
rect 11474 55636 11522 55692
rect 11578 55636 11626 55692
rect 11682 55636 11710 55692
rect 11788 59780 11844 59790
rect 11788 55748 11844 59724
rect 13356 58548 13412 58558
rect 11788 55682 11844 55692
rect 12460 57988 12516 57998
rect 11390 54124 11710 55636
rect 12460 55188 12516 57932
rect 12460 55122 12516 55132
rect 11390 54068 11418 54124
rect 11474 54068 11522 54124
rect 11578 54068 11626 54124
rect 11682 54068 11710 54124
rect 11004 50428 11060 52108
rect 11390 52556 11710 54068
rect 12908 54292 12964 54302
rect 12908 53844 12964 54236
rect 11390 52500 11418 52556
rect 11474 52500 11522 52556
rect 11578 52500 11626 52556
rect 11682 52500 11710 52556
rect 11390 50988 11710 52500
rect 11390 50932 11418 50988
rect 11474 50932 11522 50988
rect 11578 50932 11626 50988
rect 11682 50932 11710 50988
rect 11004 50372 11284 50428
rect 11004 49700 11060 49710
rect 11004 48358 11060 49644
rect 11228 48468 11284 50372
rect 11228 48402 11284 48412
rect 11390 49420 11710 50932
rect 11390 49364 11418 49420
rect 11474 49364 11522 49420
rect 11578 49364 11626 49420
rect 11682 49364 11710 49420
rect 11004 48302 11172 48358
rect 10892 44258 10948 44268
rect 11004 47012 11060 47022
rect 11004 45780 11060 46956
rect 11004 44772 11060 45724
rect 11004 44212 11060 44716
rect 11004 44146 11060 44156
rect 10892 43540 10948 43550
rect 10892 39172 10948 43484
rect 11116 42644 11172 48302
rect 11390 47852 11710 49364
rect 12012 53396 12068 53406
rect 11390 47796 11418 47852
rect 11474 47796 11522 47852
rect 11578 47796 11626 47852
rect 11682 47796 11710 47852
rect 11228 46564 11284 46574
rect 11228 45556 11284 46508
rect 11228 45490 11284 45500
rect 11390 46284 11710 47796
rect 11390 46228 11418 46284
rect 11474 46228 11522 46284
rect 11578 46228 11626 46284
rect 11682 46228 11710 46284
rect 11390 44716 11710 46228
rect 11788 49028 11844 49038
rect 11788 44996 11844 48972
rect 12012 47460 12068 53340
rect 12908 52164 12964 53788
rect 13356 52388 13412 58492
rect 13692 57876 13748 57886
rect 13692 57316 13748 57820
rect 13692 52948 13748 57260
rect 13692 52882 13748 52892
rect 13356 52322 13412 52332
rect 12908 52098 12964 52108
rect 13916 50372 13972 67564
rect 14028 59220 14084 69132
rect 14140 69524 14196 69534
rect 14140 59780 14196 69468
rect 14252 68628 14308 68638
rect 14252 62580 14308 68572
rect 14252 60564 14308 62524
rect 14252 60498 14308 60508
rect 14364 65828 14420 65838
rect 14364 60004 14420 65772
rect 14476 62244 14532 72604
rect 14588 68516 14644 78988
rect 14588 68450 14644 68460
rect 14792 78428 15112 79940
rect 14792 78372 14820 78428
rect 14876 78372 14924 78428
rect 14980 78372 15028 78428
rect 15084 78372 15112 78428
rect 14792 76860 15112 78372
rect 14792 76804 14820 76860
rect 14876 76804 14924 76860
rect 14980 76804 15028 76860
rect 15084 76804 15112 76860
rect 14792 75292 15112 76804
rect 15708 82740 15764 82750
rect 14792 75236 14820 75292
rect 14876 75236 14924 75292
rect 14980 75236 15028 75292
rect 15084 75236 15112 75292
rect 14792 73724 15112 75236
rect 14792 73668 14820 73724
rect 14876 73668 14924 73724
rect 14980 73668 15028 73724
rect 15084 73668 15112 73724
rect 14792 72156 15112 73668
rect 15260 76020 15316 76030
rect 15260 73220 15316 75964
rect 15260 73154 15316 73164
rect 14792 72100 14820 72156
rect 14876 72100 14924 72156
rect 14980 72100 15028 72156
rect 15084 72100 15112 72156
rect 14792 70588 15112 72100
rect 15372 72324 15428 72334
rect 14792 70532 14820 70588
rect 14876 70532 14924 70588
rect 14980 70532 15028 70588
rect 15084 70532 15112 70588
rect 15260 70980 15316 70990
rect 15260 70644 15316 70924
rect 15372 70868 15428 72268
rect 15596 72324 15652 72334
rect 15484 71876 15540 71886
rect 15484 70980 15540 71820
rect 15484 70914 15540 70924
rect 15372 70802 15428 70812
rect 15596 70588 15652 72268
rect 15260 70578 15316 70588
rect 14792 69020 15112 70532
rect 15484 70532 15652 70588
rect 15484 69972 15540 70532
rect 15484 69906 15540 69916
rect 14792 68964 14820 69020
rect 14876 68964 14924 69020
rect 14980 68964 15028 69020
rect 15084 68964 15112 69020
rect 14476 62178 14532 62188
rect 14792 67452 15112 68964
rect 14792 67396 14820 67452
rect 14876 67396 14924 67452
rect 14980 67396 15028 67452
rect 15084 67396 15112 67452
rect 14792 65884 15112 67396
rect 14792 65828 14820 65884
rect 14876 65828 14924 65884
rect 14980 65828 15028 65884
rect 15084 65828 15112 65884
rect 14792 64316 15112 65828
rect 14792 64260 14820 64316
rect 14876 64260 14924 64316
rect 14980 64260 15028 64316
rect 15084 64260 15112 64316
rect 14792 62748 15112 64260
rect 15260 68964 15316 68974
rect 15260 63700 15316 68908
rect 15260 63634 15316 63644
rect 14792 62692 14820 62748
rect 14876 62692 14924 62748
rect 14980 62692 15028 62748
rect 15084 62692 15112 62748
rect 14476 61908 14532 61918
rect 14476 61012 14532 61852
rect 14476 60946 14532 60956
rect 14792 61180 15112 62692
rect 14792 61124 14820 61180
rect 14876 61124 14924 61180
rect 14980 61124 15028 61180
rect 15084 61124 15112 61180
rect 14364 59938 14420 59948
rect 14140 59714 14196 59724
rect 14028 59154 14084 59164
rect 14792 59612 15112 61124
rect 15260 63364 15316 63374
rect 15260 60564 15316 63308
rect 15260 60498 15316 60508
rect 15372 62132 15428 62142
rect 15372 61572 15428 62076
rect 14792 59556 14820 59612
rect 14876 59556 14924 59612
rect 14980 59556 15028 59612
rect 15084 59556 15112 59612
rect 14792 58044 15112 59556
rect 14792 57988 14820 58044
rect 14876 57988 14924 58044
rect 14980 57988 15028 58044
rect 15084 57988 15112 58044
rect 14140 57204 14196 57214
rect 14140 52276 14196 57148
rect 14140 52210 14196 52220
rect 14792 56476 15112 57988
rect 15260 58884 15316 58894
rect 15260 57988 15316 58828
rect 15260 57922 15316 57932
rect 14792 56420 14820 56476
rect 14876 56420 14924 56476
rect 14980 56420 15028 56476
rect 15084 56420 15112 56476
rect 14792 54908 15112 56420
rect 14792 54852 14820 54908
rect 14876 54852 14924 54908
rect 14980 54852 15028 54908
rect 15084 54852 15112 54908
rect 14792 53340 15112 54852
rect 14792 53284 14820 53340
rect 14876 53284 14924 53340
rect 14980 53284 15028 53340
rect 15084 53284 15112 53340
rect 14792 51772 15112 53284
rect 14792 51716 14820 51772
rect 14876 51716 14924 51772
rect 14980 51716 15028 51772
rect 15084 51716 15112 51772
rect 13916 50306 13972 50316
rect 14476 50484 14532 50494
rect 12460 49924 12516 49934
rect 12460 47684 12516 49868
rect 12460 47618 12516 47628
rect 14364 49924 14420 49934
rect 14364 49252 14420 49868
rect 14364 48692 14420 49196
rect 14476 48916 14532 50428
rect 14476 48850 14532 48860
rect 14792 50204 15112 51716
rect 14792 50148 14820 50204
rect 14876 50148 14924 50204
rect 14980 50148 15028 50204
rect 15084 50148 15112 50204
rect 12012 47394 12068 47404
rect 13916 47572 13972 47582
rect 11788 44930 11844 44940
rect 13244 46788 13300 46798
rect 11390 44660 11418 44716
rect 11474 44660 11522 44716
rect 11578 44660 11626 44716
rect 11682 44660 11710 44716
rect 11116 42578 11172 42588
rect 11228 43876 11284 43886
rect 10892 39106 10948 39116
rect 11004 42084 11060 42094
rect 11004 36932 11060 42028
rect 11228 40852 11284 43820
rect 11116 39844 11172 39854
rect 11116 38164 11172 39788
rect 11116 38098 11172 38108
rect 11228 38724 11284 40796
rect 11004 36866 11060 36876
rect 11228 38052 11284 38668
rect 11228 36260 11284 37996
rect 11228 36194 11284 36204
rect 11390 43148 11710 44660
rect 11390 43092 11418 43148
rect 11474 43092 11522 43148
rect 11578 43092 11626 43148
rect 11682 43092 11710 43148
rect 11390 41580 11710 43092
rect 12124 44660 12180 44670
rect 12124 42980 12180 44604
rect 12124 42914 12180 42924
rect 12460 42420 12516 42430
rect 11390 41524 11418 41580
rect 11474 41524 11522 41580
rect 11578 41524 11626 41580
rect 11682 41524 11710 41580
rect 11390 40012 11710 41524
rect 12236 42196 12292 42206
rect 11390 39956 11418 40012
rect 11474 39956 11522 40012
rect 11578 39956 11626 40012
rect 11682 39956 11710 40012
rect 11390 38444 11710 39956
rect 11788 40852 11844 40862
rect 11788 39844 11844 40796
rect 11788 39778 11844 39788
rect 11390 38388 11418 38444
rect 11474 38388 11522 38444
rect 11578 38388 11626 38444
rect 11682 38388 11710 38444
rect 11390 36876 11710 38388
rect 11390 36820 11418 36876
rect 11474 36820 11522 36876
rect 11578 36820 11626 36876
rect 11682 36820 11710 36876
rect 11116 35476 11172 35486
rect 11004 35252 11060 35262
rect 10892 32900 10948 32910
rect 10892 25956 10948 32844
rect 11004 32788 11060 35196
rect 11004 31780 11060 32732
rect 11004 31714 11060 31724
rect 11116 28756 11172 35420
rect 11390 35308 11710 36820
rect 11788 39284 11844 39294
rect 11788 36708 11844 39228
rect 12236 37604 12292 42140
rect 12236 37538 12292 37548
rect 11788 35476 11844 36652
rect 12460 35700 12516 42364
rect 13244 41076 13300 46732
rect 13804 44772 13860 44782
rect 13244 41010 13300 41020
rect 13580 44548 13636 44558
rect 13580 39732 13636 44492
rect 12796 38388 12852 38398
rect 12796 36820 12852 38332
rect 13580 37492 13636 39676
rect 13804 43540 13860 44716
rect 13580 37426 13636 37436
rect 13692 39620 13748 39630
rect 12796 36754 12852 36764
rect 13692 36484 13748 39564
rect 13692 36418 13748 36428
rect 13804 36372 13860 43484
rect 13916 44436 13972 47516
rect 14364 47236 14420 48636
rect 14364 47170 14420 47180
rect 14792 48636 15112 50148
rect 14792 48580 14820 48636
rect 14876 48580 14924 48636
rect 14980 48580 15028 48636
rect 15084 48580 15112 48636
rect 14792 47068 15112 48580
rect 14792 47012 14820 47068
rect 14876 47012 14924 47068
rect 14980 47012 15028 47068
rect 15084 47012 15112 47068
rect 13916 42420 13972 44380
rect 13916 42354 13972 42364
rect 14476 45668 14532 45678
rect 13804 36306 13860 36316
rect 14364 36708 14420 36718
rect 12460 35634 12516 35644
rect 11788 35410 11844 35420
rect 11390 35252 11418 35308
rect 11474 35252 11522 35308
rect 11578 35252 11626 35308
rect 11682 35252 11710 35308
rect 14364 35364 14420 36652
rect 14476 35476 14532 45612
rect 14792 45500 15112 47012
rect 14792 45444 14820 45500
rect 14876 45444 14924 45500
rect 14980 45444 15028 45500
rect 15084 45444 15112 45500
rect 14588 44436 14644 44446
rect 14588 43540 14644 44380
rect 14588 43474 14644 43484
rect 14792 43932 15112 45444
rect 14792 43876 14820 43932
rect 14876 43876 14924 43932
rect 14980 43876 15028 43932
rect 15084 43876 15112 43932
rect 14476 35410 14532 35420
rect 14792 42364 15112 43876
rect 15260 45892 15316 45902
rect 15260 43540 15316 45836
rect 15260 43474 15316 43484
rect 14792 42308 14820 42364
rect 14876 42308 14924 42364
rect 14980 42308 15028 42364
rect 15084 42308 15112 42364
rect 14792 40796 15112 42308
rect 14792 40740 14820 40796
rect 14876 40740 14924 40796
rect 14980 40740 15028 40796
rect 15084 40740 15112 40796
rect 14792 39228 15112 40740
rect 15260 41412 15316 41422
rect 15260 40628 15316 41356
rect 15260 39508 15316 40572
rect 15260 39442 15316 39452
rect 14792 39172 14820 39228
rect 14876 39172 14924 39228
rect 14980 39172 15028 39228
rect 15084 39172 15112 39228
rect 14792 37660 15112 39172
rect 14792 37604 14820 37660
rect 14876 37604 14924 37660
rect 14980 37604 15028 37660
rect 15084 37604 15112 37660
rect 14792 36092 15112 37604
rect 14792 36036 14820 36092
rect 14876 36036 14924 36092
rect 14980 36036 15028 36092
rect 15084 36036 15112 36092
rect 14364 35298 14420 35308
rect 11228 34356 11284 34366
rect 11228 32788 11284 34300
rect 11228 31892 11284 32732
rect 11228 31826 11284 31836
rect 11390 33740 11710 35252
rect 11390 33684 11418 33740
rect 11474 33684 11522 33740
rect 11578 33684 11626 33740
rect 11682 33684 11710 33740
rect 11390 32172 11710 33684
rect 11390 32116 11418 32172
rect 11474 32116 11522 32172
rect 11578 32116 11626 32172
rect 11682 32116 11710 32172
rect 11116 28690 11172 28700
rect 11390 30604 11710 32116
rect 11390 30548 11418 30604
rect 11474 30548 11522 30604
rect 11578 30548 11626 30604
rect 11682 30548 11710 30604
rect 11390 29036 11710 30548
rect 11390 28980 11418 29036
rect 11474 28980 11522 29036
rect 11578 28980 11626 29036
rect 11682 28980 11710 29036
rect 10892 25890 10948 25900
rect 11390 27468 11710 28980
rect 13692 35028 13748 35038
rect 13692 28532 13748 34972
rect 13692 27860 13748 28476
rect 13692 27794 13748 27804
rect 14792 34524 15112 36036
rect 14792 34468 14820 34524
rect 14876 34468 14924 34524
rect 14980 34468 15028 34524
rect 15084 34468 15112 34524
rect 14792 32956 15112 34468
rect 14792 32900 14820 32956
rect 14876 32900 14924 32956
rect 14980 32900 15028 32956
rect 15084 32900 15112 32956
rect 14792 31388 15112 32900
rect 14792 31332 14820 31388
rect 14876 31332 14924 31388
rect 14980 31332 15028 31388
rect 15084 31332 15112 31388
rect 14792 29820 15112 31332
rect 14792 29764 14820 29820
rect 14876 29764 14924 29820
rect 14980 29764 15028 29820
rect 15084 29764 15112 29820
rect 14792 28252 15112 29764
rect 14792 28196 14820 28252
rect 14876 28196 14924 28252
rect 14980 28196 15028 28252
rect 15084 28196 15112 28252
rect 11390 27412 11418 27468
rect 11474 27412 11522 27468
rect 11578 27412 11626 27468
rect 11682 27412 11710 27468
rect 11390 25900 11710 27412
rect 14792 26684 15112 28196
rect 14792 26628 14820 26684
rect 14876 26628 14924 26684
rect 14980 26628 15028 26684
rect 15084 26628 15112 26684
rect 14588 26180 14644 26190
rect 10668 15362 10724 15372
rect 11390 25844 11418 25900
rect 11474 25844 11522 25900
rect 11578 25844 11626 25900
rect 11682 25844 11710 25900
rect 11390 24332 11710 25844
rect 12684 26068 12740 26078
rect 11390 24276 11418 24332
rect 11474 24276 11522 24332
rect 11578 24276 11626 24332
rect 11682 24276 11710 24332
rect 11390 22764 11710 24276
rect 11788 24948 11844 24958
rect 11788 23380 11844 24892
rect 12684 23604 12740 26012
rect 12684 23538 12740 23548
rect 14588 25508 14644 26124
rect 11788 23314 11844 23324
rect 11390 22708 11418 22764
rect 11474 22708 11522 22764
rect 11578 22708 11626 22764
rect 11682 22708 11710 22764
rect 11390 21196 11710 22708
rect 11390 21140 11418 21196
rect 11474 21140 11522 21196
rect 11578 21140 11626 21196
rect 11682 21140 11710 21196
rect 11390 19628 11710 21140
rect 11390 19572 11418 19628
rect 11474 19572 11522 19628
rect 11578 19572 11626 19628
rect 11682 19572 11710 19628
rect 11390 18060 11710 19572
rect 11390 18004 11418 18060
rect 11474 18004 11522 18060
rect 11578 18004 11626 18060
rect 11682 18004 11710 18060
rect 11390 16492 11710 18004
rect 11390 16436 11418 16492
rect 11474 16436 11522 16492
rect 11578 16436 11626 16492
rect 11682 16436 11710 16492
rect 11390 14924 11710 16436
rect 14588 15204 14644 25452
rect 14588 15138 14644 15148
rect 14792 25116 15112 26628
rect 14792 25060 14820 25116
rect 14876 25060 14924 25116
rect 14980 25060 15028 25116
rect 15084 25060 15112 25116
rect 14792 23548 15112 25060
rect 14792 23492 14820 23548
rect 14876 23492 14924 23548
rect 14980 23492 15028 23548
rect 15084 23492 15112 23548
rect 14792 21980 15112 23492
rect 14792 21924 14820 21980
rect 14876 21924 14924 21980
rect 14980 21924 15028 21980
rect 15084 21924 15112 21980
rect 14792 20412 15112 21924
rect 14792 20356 14820 20412
rect 14876 20356 14924 20412
rect 14980 20356 15028 20412
rect 15084 20356 15112 20412
rect 14792 18844 15112 20356
rect 15372 19348 15428 61516
rect 15596 61796 15652 61806
rect 15596 61572 15652 61740
rect 15596 61506 15652 61516
rect 15484 55524 15540 55534
rect 15484 37492 15540 55468
rect 15484 37426 15540 37436
rect 15372 19282 15428 19292
rect 15484 22932 15540 22942
rect 14792 18788 14820 18844
rect 14876 18788 14924 18844
rect 14980 18788 15028 18844
rect 15084 18788 15112 18844
rect 14792 17276 15112 18788
rect 15484 17780 15540 22876
rect 15484 17714 15540 17724
rect 14792 17220 14820 17276
rect 14876 17220 14924 17276
rect 14980 17220 15028 17276
rect 15084 17220 15112 17276
rect 14792 15708 15112 17220
rect 14792 15652 14820 15708
rect 14876 15652 14924 15708
rect 14980 15652 15028 15708
rect 15084 15652 15112 15708
rect 11390 14868 11418 14924
rect 11474 14868 11522 14924
rect 11578 14868 11626 14924
rect 11682 14868 11710 14924
rect 7988 14084 8016 14140
rect 8072 14084 8120 14140
rect 8176 14084 8224 14140
rect 8280 14084 8308 14140
rect 4586 11732 4614 11788
rect 4670 11732 4718 11788
rect 4774 11732 4822 11788
rect 4878 11732 4906 11788
rect 4586 10220 4906 11732
rect 7988 12572 8308 14084
rect 9884 14756 9940 14766
rect 9884 13412 9940 14700
rect 9884 13346 9940 13356
rect 11390 13356 11710 14868
rect 7988 12516 8016 12572
rect 8072 12516 8120 12572
rect 8176 12516 8224 12572
rect 8280 12516 8308 12572
rect 5852 11396 5908 11406
rect 5852 11172 5908 11340
rect 5852 11106 5908 11116
rect 4586 10164 4614 10220
rect 4670 10164 4718 10220
rect 4774 10164 4822 10220
rect 4878 10164 4906 10220
rect 4586 8652 4906 10164
rect 4586 8596 4614 8652
rect 4670 8596 4718 8652
rect 4774 8596 4822 8652
rect 4878 8596 4906 8652
rect 4586 7084 4906 8596
rect 4586 7028 4614 7084
rect 4670 7028 4718 7084
rect 4774 7028 4822 7084
rect 4878 7028 4906 7084
rect 4586 5516 4906 7028
rect 4586 5460 4614 5516
rect 4670 5460 4718 5516
rect 4774 5460 4822 5516
rect 4878 5460 4906 5516
rect 4586 3948 4906 5460
rect 4586 3892 4614 3948
rect 4670 3892 4718 3948
rect 4774 3892 4822 3948
rect 4878 3892 4906 3948
rect 4586 2380 4906 3892
rect 4586 2324 4614 2380
rect 4670 2324 4718 2380
rect 4774 2324 4822 2380
rect 4878 2324 4906 2380
rect 4586 1508 4906 2324
rect 7988 11004 8308 12516
rect 7988 10948 8016 11004
rect 8072 10948 8120 11004
rect 8176 10948 8224 11004
rect 8280 10948 8308 11004
rect 7988 9436 8308 10948
rect 7988 9380 8016 9436
rect 8072 9380 8120 9436
rect 8176 9380 8224 9436
rect 8280 9380 8308 9436
rect 7988 7868 8308 9380
rect 7988 7812 8016 7868
rect 8072 7812 8120 7868
rect 8176 7812 8224 7868
rect 8280 7812 8308 7868
rect 7988 6300 8308 7812
rect 7988 6244 8016 6300
rect 8072 6244 8120 6300
rect 8176 6244 8224 6300
rect 8280 6244 8308 6300
rect 7988 4732 8308 6244
rect 7988 4676 8016 4732
rect 8072 4676 8120 4732
rect 8176 4676 8224 4732
rect 8280 4676 8308 4732
rect 7988 3164 8308 4676
rect 7988 3108 8016 3164
rect 8072 3108 8120 3164
rect 8176 3108 8224 3164
rect 8280 3108 8308 3164
rect 7988 1596 8308 3108
rect 7988 1540 8016 1596
rect 8072 1540 8120 1596
rect 8176 1540 8224 1596
rect 8280 1540 8308 1596
rect 7988 1508 8308 1540
rect 11390 13300 11418 13356
rect 11474 13300 11522 13356
rect 11578 13300 11626 13356
rect 11682 13300 11710 13356
rect 11390 11788 11710 13300
rect 11390 11732 11418 11788
rect 11474 11732 11522 11788
rect 11578 11732 11626 11788
rect 11682 11732 11710 11788
rect 11390 10220 11710 11732
rect 11390 10164 11418 10220
rect 11474 10164 11522 10220
rect 11578 10164 11626 10220
rect 11682 10164 11710 10220
rect 11390 8652 11710 10164
rect 11390 8596 11418 8652
rect 11474 8596 11522 8652
rect 11578 8596 11626 8652
rect 11682 8596 11710 8652
rect 11390 7084 11710 8596
rect 11390 7028 11418 7084
rect 11474 7028 11522 7084
rect 11578 7028 11626 7084
rect 11682 7028 11710 7084
rect 11390 5516 11710 7028
rect 11390 5460 11418 5516
rect 11474 5460 11522 5516
rect 11578 5460 11626 5516
rect 11682 5460 11710 5516
rect 11390 3948 11710 5460
rect 11390 3892 11418 3948
rect 11474 3892 11522 3948
rect 11578 3892 11626 3948
rect 11682 3892 11710 3948
rect 11390 2380 11710 3892
rect 11390 2324 11418 2380
rect 11474 2324 11522 2380
rect 11578 2324 11626 2380
rect 11682 2324 11710 2380
rect 11390 1508 11710 2324
rect 14792 14140 15112 15652
rect 14792 14084 14820 14140
rect 14876 14084 14924 14140
rect 14980 14084 15028 14140
rect 15084 14084 15112 14140
rect 14792 12572 15112 14084
rect 14792 12516 14820 12572
rect 14876 12516 14924 12572
rect 14980 12516 15028 12572
rect 15084 12516 15112 12572
rect 14792 11004 15112 12516
rect 14792 10948 14820 11004
rect 14876 10948 14924 11004
rect 14980 10948 15028 11004
rect 15084 10948 15112 11004
rect 14792 9436 15112 10948
rect 14792 9380 14820 9436
rect 14876 9380 14924 9436
rect 14980 9380 15028 9436
rect 15084 9380 15112 9436
rect 14792 7868 15112 9380
rect 14792 7812 14820 7868
rect 14876 7812 14924 7868
rect 14980 7812 15028 7868
rect 15084 7812 15112 7868
rect 14792 6300 15112 7812
rect 15708 6692 15764 82684
rect 18194 82348 18514 83860
rect 18194 82292 18222 82348
rect 18278 82292 18326 82348
rect 18382 82292 18430 82348
rect 18486 82292 18514 82348
rect 18194 80780 18514 82292
rect 18194 80724 18222 80780
rect 18278 80724 18326 80780
rect 18382 80724 18430 80780
rect 18486 80724 18514 80780
rect 18194 79212 18514 80724
rect 18194 79156 18222 79212
rect 18278 79156 18326 79212
rect 18382 79156 18430 79212
rect 18486 79156 18514 79212
rect 16044 78596 16100 78606
rect 15820 73220 15876 73230
rect 15820 35140 15876 73164
rect 16044 70980 16100 78540
rect 18194 77644 18514 79156
rect 18194 77588 18222 77644
rect 18278 77588 18326 77644
rect 18382 77588 18430 77644
rect 18486 77588 18514 77644
rect 17836 77252 17892 77262
rect 16492 72884 16548 72894
rect 16492 71652 16548 72828
rect 16492 71586 16548 71596
rect 16044 70914 16100 70924
rect 16044 70644 16100 70654
rect 15932 61908 15988 61918
rect 15932 59108 15988 61852
rect 15932 59042 15988 59052
rect 15932 58772 15988 58782
rect 15932 52052 15988 58716
rect 15932 47348 15988 51996
rect 15932 47282 15988 47292
rect 15820 35074 15876 35084
rect 16044 33124 16100 70588
rect 16940 69412 16996 69422
rect 16268 63140 16324 63150
rect 16268 62916 16324 63084
rect 16268 62850 16324 62860
rect 16940 61796 16996 69356
rect 16940 61730 16996 61740
rect 17164 68964 17220 68974
rect 17164 63140 17220 68908
rect 17612 67060 17668 67070
rect 16156 61124 16212 61134
rect 16156 59780 16212 61068
rect 17164 60676 17220 63084
rect 17164 60610 17220 60620
rect 17276 64708 17332 64718
rect 17276 60228 17332 64652
rect 17612 63252 17668 67004
rect 17612 63186 17668 63196
rect 17276 60162 17332 60172
rect 17500 62244 17556 62254
rect 16156 59714 16212 59724
rect 17500 59332 17556 62188
rect 17500 59266 17556 59276
rect 17836 58828 17892 77196
rect 18194 76076 18514 77588
rect 18194 76020 18222 76076
rect 18278 76020 18326 76076
rect 18382 76020 18430 76076
rect 18486 76020 18514 76076
rect 18194 74508 18514 76020
rect 18194 74452 18222 74508
rect 18278 74452 18326 74508
rect 18382 74452 18430 74508
rect 18486 74452 18514 74508
rect 18060 73444 18116 73454
rect 17948 65604 18004 65614
rect 17948 60452 18004 65548
rect 17948 60386 18004 60396
rect 17164 58772 17892 58828
rect 16380 58660 16436 58670
rect 16380 58436 16436 58604
rect 16380 58370 16436 58380
rect 17052 56868 17108 56878
rect 16492 56756 16548 56766
rect 16156 56420 16212 56430
rect 16156 43652 16212 56364
rect 16156 43586 16212 43596
rect 16380 53508 16436 53518
rect 16380 35140 16436 53452
rect 16380 35074 16436 35084
rect 16044 33058 16100 33068
rect 16492 31220 16548 56700
rect 17052 52612 17108 56812
rect 17052 52546 17108 52556
rect 17164 55188 17220 58772
rect 17164 47124 17220 55132
rect 17948 55972 18004 55982
rect 17164 47058 17220 47068
rect 17500 52276 17556 52286
rect 17500 50036 17556 52220
rect 17948 50820 18004 55916
rect 17948 50754 18004 50764
rect 17724 50484 17780 50494
rect 17500 48580 17556 49980
rect 17500 47460 17556 48524
rect 17500 47124 17556 47404
rect 17500 47058 17556 47068
rect 17612 50372 17780 50428
rect 17052 46004 17108 46014
rect 16716 43316 16772 43326
rect 16716 42756 16772 43260
rect 16716 41748 16772 42700
rect 16716 41682 16772 41692
rect 16828 40180 16884 40190
rect 16828 39060 16884 40124
rect 17052 39284 17108 45948
rect 17052 39218 17108 39228
rect 17500 44436 17556 44446
rect 16828 38836 16884 39004
rect 16828 38770 16884 38780
rect 17500 36148 17556 44380
rect 17612 44324 17668 50372
rect 17948 48356 18004 48366
rect 17948 47236 18004 48300
rect 17948 47170 18004 47180
rect 17612 44258 17668 44268
rect 18060 41972 18116 73388
rect 18060 41906 18116 41916
rect 18194 72940 18514 74452
rect 19964 74788 20020 74798
rect 19964 73668 20020 74732
rect 19964 73602 20020 73612
rect 18194 72884 18222 72940
rect 18278 72884 18326 72940
rect 18382 72884 18430 72940
rect 18486 72884 18514 72940
rect 18194 71372 18514 72884
rect 18194 71316 18222 71372
rect 18278 71316 18326 71372
rect 18382 71316 18430 71372
rect 18486 71316 18514 71372
rect 18194 69804 18514 71316
rect 18194 69748 18222 69804
rect 18278 69748 18326 69804
rect 18382 69748 18430 69804
rect 18486 69748 18514 69804
rect 18194 68236 18514 69748
rect 19740 70420 19796 70430
rect 18194 68180 18222 68236
rect 18278 68180 18326 68236
rect 18382 68180 18430 68236
rect 18486 68180 18514 68236
rect 18194 66668 18514 68180
rect 18194 66612 18222 66668
rect 18278 66612 18326 66668
rect 18382 66612 18430 66668
rect 18486 66612 18514 66668
rect 18194 65100 18514 66612
rect 18194 65044 18222 65100
rect 18278 65044 18326 65100
rect 18382 65044 18430 65100
rect 18486 65044 18514 65100
rect 18194 63532 18514 65044
rect 18194 63476 18222 63532
rect 18278 63476 18326 63532
rect 18382 63476 18430 63532
rect 18486 63476 18514 63532
rect 18194 61964 18514 63476
rect 18194 61908 18222 61964
rect 18278 61908 18326 61964
rect 18382 61908 18430 61964
rect 18486 61908 18514 61964
rect 18194 60396 18514 61908
rect 18620 68852 18676 68862
rect 18620 60564 18676 68796
rect 19404 67620 19460 67630
rect 18620 60498 18676 60508
rect 18956 66052 19012 66062
rect 18194 60340 18222 60396
rect 18278 60340 18326 60396
rect 18382 60340 18430 60396
rect 18486 60340 18514 60396
rect 18194 58828 18514 60340
rect 18194 58772 18222 58828
rect 18278 58772 18326 58828
rect 18382 58772 18430 58828
rect 18486 58772 18514 58828
rect 18194 57260 18514 58772
rect 18194 57204 18222 57260
rect 18278 57204 18326 57260
rect 18382 57204 18430 57260
rect 18486 57204 18514 57260
rect 18194 55692 18514 57204
rect 18194 55636 18222 55692
rect 18278 55636 18326 55692
rect 18382 55636 18430 55692
rect 18486 55636 18514 55692
rect 18194 54124 18514 55636
rect 18194 54068 18222 54124
rect 18278 54068 18326 54124
rect 18382 54068 18430 54124
rect 18486 54068 18514 54124
rect 18194 52556 18514 54068
rect 18194 52500 18222 52556
rect 18278 52500 18326 52556
rect 18382 52500 18430 52556
rect 18486 52500 18514 52556
rect 18194 50988 18514 52500
rect 18194 50932 18222 50988
rect 18278 50932 18326 50988
rect 18382 50932 18430 50988
rect 18486 50932 18514 50988
rect 18194 49420 18514 50932
rect 18620 52948 18676 52958
rect 18620 49700 18676 52892
rect 18844 52388 18900 52398
rect 18620 49634 18676 49644
rect 18732 51492 18788 51502
rect 18194 49364 18222 49420
rect 18278 49364 18326 49420
rect 18382 49364 18430 49420
rect 18486 49364 18514 49420
rect 18194 47852 18514 49364
rect 18194 47796 18222 47852
rect 18278 47796 18326 47852
rect 18382 47796 18430 47852
rect 18486 47796 18514 47852
rect 18194 46284 18514 47796
rect 18194 46228 18222 46284
rect 18278 46228 18326 46284
rect 18382 46228 18430 46284
rect 18486 46228 18514 46284
rect 18194 44716 18514 46228
rect 18194 44660 18222 44716
rect 18278 44660 18326 44716
rect 18382 44660 18430 44716
rect 18486 44660 18514 44716
rect 18194 43148 18514 44660
rect 18194 43092 18222 43148
rect 18278 43092 18326 43148
rect 18382 43092 18430 43148
rect 18486 43092 18514 43148
rect 18194 41580 18514 43092
rect 18620 43428 18676 43438
rect 18620 42084 18676 43372
rect 18620 42018 18676 42028
rect 17500 36082 17556 36092
rect 17724 41524 17780 41534
rect 17724 35476 17780 41468
rect 18194 41524 18222 41580
rect 18278 41524 18326 41580
rect 18382 41524 18430 41580
rect 18486 41524 18514 41580
rect 17948 40964 18004 40974
rect 17948 38612 18004 40908
rect 17948 38546 18004 38556
rect 18194 40012 18514 41524
rect 18194 39956 18222 40012
rect 18278 39956 18326 40012
rect 18382 39956 18430 40012
rect 18486 39956 18514 40012
rect 17724 35410 17780 35420
rect 18194 38444 18514 39956
rect 18194 38388 18222 38444
rect 18278 38388 18326 38444
rect 18382 38388 18430 38444
rect 18486 38388 18514 38444
rect 18194 36876 18514 38388
rect 18194 36820 18222 36876
rect 18278 36820 18326 36876
rect 18382 36820 18430 36876
rect 18486 36820 18514 36876
rect 18194 35308 18514 36820
rect 18620 41076 18676 41086
rect 18620 36820 18676 41020
rect 18620 36596 18676 36764
rect 18620 36530 18676 36540
rect 18194 35252 18222 35308
rect 18278 35252 18326 35308
rect 18382 35252 18430 35308
rect 18486 35252 18514 35308
rect 18194 33740 18514 35252
rect 18194 33684 18222 33740
rect 18278 33684 18326 33740
rect 18382 33684 18430 33740
rect 18486 33684 18514 33740
rect 16492 31154 16548 31164
rect 16604 32788 16660 32798
rect 16604 23828 16660 32732
rect 17500 32788 17556 32798
rect 17500 32452 17556 32732
rect 17500 32386 17556 32396
rect 17724 32788 17780 32798
rect 17724 27524 17780 32732
rect 17724 27458 17780 27468
rect 18194 32172 18514 33684
rect 18194 32116 18222 32172
rect 18278 32116 18326 32172
rect 18382 32116 18430 32172
rect 18486 32116 18514 32172
rect 18194 30604 18514 32116
rect 18194 30548 18222 30604
rect 18278 30548 18326 30604
rect 18382 30548 18430 30604
rect 18486 30548 18514 30604
rect 18194 29036 18514 30548
rect 18194 28980 18222 29036
rect 18278 28980 18326 29036
rect 18382 28980 18430 29036
rect 18486 28980 18514 29036
rect 18194 27468 18514 28980
rect 16604 23762 16660 23772
rect 18194 27412 18222 27468
rect 18278 27412 18326 27468
rect 18382 27412 18430 27468
rect 18486 27412 18514 27468
rect 18194 25900 18514 27412
rect 18194 25844 18222 25900
rect 18278 25844 18326 25900
rect 18382 25844 18430 25900
rect 18486 25844 18514 25900
rect 18194 24332 18514 25844
rect 18620 26404 18676 26414
rect 18620 25396 18676 26348
rect 18620 25330 18676 25340
rect 18194 24276 18222 24332
rect 18278 24276 18326 24332
rect 18382 24276 18430 24332
rect 18486 24276 18514 24332
rect 17388 22820 17444 22830
rect 16380 22708 16436 22718
rect 16268 19124 16324 19134
rect 16268 17220 16324 19068
rect 16268 16996 16324 17164
rect 16268 16930 16324 16940
rect 16380 12404 16436 22652
rect 16940 21252 16996 21262
rect 16940 14980 16996 21196
rect 16940 14914 16996 14924
rect 16380 12338 16436 12348
rect 17388 12180 17444 22764
rect 18194 22764 18514 24276
rect 18194 22708 18222 22764
rect 18278 22708 18326 22764
rect 18382 22708 18430 22764
rect 18486 22708 18514 22764
rect 17724 22148 17780 22158
rect 17724 21364 17780 22092
rect 17724 21298 17780 21308
rect 17388 12114 17444 12124
rect 18194 21196 18514 22708
rect 18194 21140 18222 21196
rect 18278 21140 18326 21196
rect 18382 21140 18430 21196
rect 18486 21140 18514 21196
rect 18194 19628 18514 21140
rect 18194 19572 18222 19628
rect 18278 19572 18326 19628
rect 18382 19572 18430 19628
rect 18486 19572 18514 19628
rect 18194 18060 18514 19572
rect 18194 18004 18222 18060
rect 18278 18004 18326 18060
rect 18382 18004 18430 18060
rect 18486 18004 18514 18060
rect 18194 16492 18514 18004
rect 18194 16436 18222 16492
rect 18278 16436 18326 16492
rect 18382 16436 18430 16492
rect 18486 16436 18514 16492
rect 18194 14924 18514 16436
rect 18194 14868 18222 14924
rect 18278 14868 18326 14924
rect 18382 14868 18430 14924
rect 18486 14868 18514 14924
rect 18194 13356 18514 14868
rect 18194 13300 18222 13356
rect 18278 13300 18326 13356
rect 18382 13300 18430 13356
rect 18486 13300 18514 13356
rect 18194 11788 18514 13300
rect 18194 11732 18222 11788
rect 18278 11732 18326 11788
rect 18382 11732 18430 11788
rect 18486 11732 18514 11788
rect 18620 12404 18676 12414
rect 18620 11844 18676 12348
rect 18620 11778 18676 11788
rect 16268 10612 16324 10622
rect 16268 10164 16324 10556
rect 16268 9156 16324 10108
rect 16268 9090 16324 9100
rect 18194 10220 18514 11732
rect 18732 10836 18788 51436
rect 18844 26908 18900 52332
rect 18956 37380 19012 65996
rect 19180 65604 19236 65614
rect 19068 63140 19124 63150
rect 19068 59668 19124 63084
rect 19068 59602 19124 59612
rect 19068 56196 19124 56206
rect 19068 53732 19124 56140
rect 19068 53666 19124 53676
rect 18956 37314 19012 37324
rect 19068 50708 19124 50718
rect 18956 36484 19012 36494
rect 18956 35476 19012 36428
rect 18956 35410 19012 35420
rect 18844 26852 19012 26908
rect 18956 12404 19012 26852
rect 19068 24948 19124 50652
rect 19180 35140 19236 65548
rect 19404 60788 19460 67564
rect 19740 62692 19796 70364
rect 19740 62626 19796 62636
rect 20188 68180 20244 68190
rect 19404 60722 19460 60732
rect 20188 60788 20244 68124
rect 20188 60722 20244 60732
rect 19516 56756 19572 56766
rect 19292 52052 19348 52062
rect 19292 51716 19348 51996
rect 19292 50372 19348 51660
rect 19292 50306 19348 50316
rect 19292 44212 19348 44222
rect 19292 41412 19348 44156
rect 19292 38164 19348 41356
rect 19404 42084 19460 42094
rect 19404 40852 19460 42028
rect 19404 40786 19460 40796
rect 19292 37492 19348 38108
rect 19292 37426 19348 37436
rect 19180 35074 19236 35084
rect 19404 32788 19460 32798
rect 19292 27076 19348 27086
rect 19180 26740 19236 26750
rect 19180 25844 19236 26684
rect 19180 25778 19236 25788
rect 19068 24882 19124 24892
rect 19292 22596 19348 27020
rect 19404 26068 19460 32732
rect 19404 26002 19460 26012
rect 19516 25172 19572 56700
rect 19964 54292 20020 54302
rect 19852 53620 19908 53630
rect 19740 35028 19796 35038
rect 19516 25106 19572 25116
rect 19628 33796 19684 33806
rect 19628 24836 19684 33740
rect 19740 31444 19796 34972
rect 19740 31378 19796 31388
rect 19628 24388 19684 24780
rect 19628 24322 19684 24332
rect 19740 31108 19796 31118
rect 19740 24276 19796 31052
rect 19740 24210 19796 24220
rect 19852 24052 19908 53564
rect 19964 47236 20020 54236
rect 20300 53732 20356 53742
rect 20188 52948 20244 52958
rect 19964 47170 20020 47180
rect 20076 50484 20132 50494
rect 20076 46788 20132 50428
rect 20076 46722 20132 46732
rect 20076 38836 20132 38846
rect 19964 34580 20020 34590
rect 19964 33124 20020 34524
rect 19964 33058 20020 33068
rect 20076 32452 20132 38780
rect 20076 32386 20132 32396
rect 19964 27412 20020 27422
rect 19964 26404 20020 27356
rect 19964 26338 20020 26348
rect 19852 23986 19908 23996
rect 19292 22530 19348 22540
rect 20188 15148 20244 52892
rect 20300 50428 20356 53676
rect 20300 50372 20468 50428
rect 20300 40404 20356 40414
rect 20300 39284 20356 40348
rect 20300 35028 20356 39228
rect 20300 34962 20356 34972
rect 20300 32004 20356 32014
rect 20300 30100 20356 31948
rect 20300 30034 20356 30044
rect 20412 28378 20468 50372
rect 20524 38668 20580 93660
rect 20860 92820 20916 92830
rect 20748 84420 20804 84430
rect 20748 83748 20804 84364
rect 20748 83682 20804 83692
rect 20860 83076 20916 92764
rect 20860 83010 20916 83020
rect 21596 92540 21916 94052
rect 24998 96460 25318 97972
rect 24998 96404 25026 96460
rect 25082 96404 25130 96460
rect 25186 96404 25234 96460
rect 25290 96404 25318 96460
rect 24998 94892 25318 96404
rect 24998 94836 25026 94892
rect 25082 94836 25130 94892
rect 25186 94836 25234 94892
rect 25290 94836 25318 94892
rect 21596 92484 21624 92540
rect 21680 92484 21728 92540
rect 21784 92484 21832 92540
rect 21888 92484 21916 92540
rect 21596 90972 21916 92484
rect 23100 93604 23156 93614
rect 22988 91700 23044 91710
rect 21596 90916 21624 90972
rect 21680 90916 21728 90972
rect 21784 90916 21832 90972
rect 21888 90916 21916 90972
rect 21596 89404 21916 90916
rect 22876 91588 22932 91598
rect 22876 90020 22932 91532
rect 22876 89954 22932 89964
rect 21596 89348 21624 89404
rect 21680 89348 21728 89404
rect 21784 89348 21832 89404
rect 21888 89348 21916 89404
rect 21596 87836 21916 89348
rect 22988 89236 23044 91644
rect 22988 89170 23044 89180
rect 21596 87780 21624 87836
rect 21680 87780 21728 87836
rect 21784 87780 21832 87836
rect 21888 87780 21916 87836
rect 21596 86268 21916 87780
rect 21596 86212 21624 86268
rect 21680 86212 21728 86268
rect 21784 86212 21832 86268
rect 21888 86212 21916 86268
rect 21596 84700 21916 86212
rect 21596 84644 21624 84700
rect 21680 84644 21728 84700
rect 21784 84644 21832 84700
rect 21888 84644 21916 84700
rect 21596 83132 21916 84644
rect 21596 83076 21624 83132
rect 21680 83076 21728 83132
rect 21784 83076 21832 83132
rect 21888 83076 21916 83132
rect 21596 81564 21916 83076
rect 21596 81508 21624 81564
rect 21680 81508 21728 81564
rect 21784 81508 21832 81564
rect 21888 81508 21916 81564
rect 21196 80276 21252 80286
rect 20860 75124 20916 75134
rect 20860 70644 20916 75068
rect 21196 72548 21252 80220
rect 21596 79996 21916 81508
rect 21596 79940 21624 79996
rect 21680 79940 21728 79996
rect 21784 79940 21832 79996
rect 21888 79940 21916 79996
rect 21596 78428 21916 79940
rect 21596 78372 21624 78428
rect 21680 78372 21728 78428
rect 21784 78372 21832 78428
rect 21888 78372 21916 78428
rect 21196 72482 21252 72492
rect 21420 77364 21476 77374
rect 21420 71540 21476 77308
rect 21420 71474 21476 71484
rect 21596 76860 21916 78372
rect 22204 81060 22260 81070
rect 22204 77140 22260 81004
rect 22204 77074 22260 77084
rect 22652 77140 22708 77150
rect 21596 76804 21624 76860
rect 21680 76804 21728 76860
rect 21784 76804 21832 76860
rect 21888 76804 21916 76860
rect 21596 75292 21916 76804
rect 21596 75236 21624 75292
rect 21680 75236 21728 75292
rect 21784 75236 21832 75292
rect 21888 75236 21916 75292
rect 21596 73724 21916 75236
rect 21596 73668 21624 73724
rect 21680 73668 21728 73724
rect 21784 73668 21832 73724
rect 21888 73668 21916 73724
rect 21596 72156 21916 73668
rect 21596 72100 21624 72156
rect 21680 72100 21728 72156
rect 21784 72100 21832 72156
rect 21888 72100 21916 72156
rect 20860 70578 20916 70588
rect 21596 70588 21916 72100
rect 22540 72436 22596 72446
rect 22540 71540 22596 72380
rect 22540 71474 22596 71484
rect 21596 70532 21624 70588
rect 21680 70532 21728 70588
rect 21784 70532 21832 70588
rect 21888 70532 21916 70588
rect 21596 69020 21916 70532
rect 21596 68964 21624 69020
rect 21680 68964 21728 69020
rect 21784 68964 21832 69020
rect 21888 68964 21916 69020
rect 21420 68180 21476 68190
rect 21420 61572 21476 68124
rect 21420 61506 21476 61516
rect 21596 67452 21916 68964
rect 21596 67396 21624 67452
rect 21680 67396 21728 67452
rect 21784 67396 21832 67452
rect 21888 67396 21916 67452
rect 21596 65884 21916 67396
rect 21596 65828 21624 65884
rect 21680 65828 21728 65884
rect 21784 65828 21832 65884
rect 21888 65828 21916 65884
rect 21596 64316 21916 65828
rect 21596 64260 21624 64316
rect 21680 64260 21728 64316
rect 21784 64260 21832 64316
rect 21888 64260 21916 64316
rect 21596 62748 21916 64260
rect 21596 62692 21624 62748
rect 21680 62692 21728 62748
rect 21784 62692 21832 62748
rect 21888 62692 21916 62748
rect 21596 61180 21916 62692
rect 21596 61124 21624 61180
rect 21680 61124 21728 61180
rect 21784 61124 21832 61180
rect 21888 61124 21916 61180
rect 21596 59612 21916 61124
rect 21596 59556 21624 59612
rect 21680 59556 21728 59612
rect 21784 59556 21832 59612
rect 21888 59556 21916 59612
rect 21596 58044 21916 59556
rect 21596 57988 21624 58044
rect 21680 57988 21728 58044
rect 21784 57988 21832 58044
rect 21888 57988 21916 58044
rect 21596 56476 21916 57988
rect 21596 56420 21624 56476
rect 21680 56420 21728 56476
rect 21784 56420 21832 56476
rect 21888 56420 21916 56476
rect 21308 55524 21364 55534
rect 21308 53172 21364 55468
rect 21308 53106 21364 53116
rect 21596 54908 21916 56420
rect 21596 54852 21624 54908
rect 21680 54852 21728 54908
rect 21784 54852 21832 54908
rect 21888 54852 21916 54908
rect 21596 53340 21916 54852
rect 21596 53284 21624 53340
rect 21680 53284 21728 53340
rect 21784 53284 21832 53340
rect 21888 53284 21916 53340
rect 21596 51772 21916 53284
rect 21596 51716 21624 51772
rect 21680 51716 21728 51772
rect 21784 51716 21832 51772
rect 21888 51716 21916 51772
rect 21596 50204 21916 51716
rect 21596 50148 21624 50204
rect 21680 50148 21728 50204
rect 21784 50148 21832 50204
rect 21888 50148 21916 50204
rect 21308 49812 21364 49822
rect 21308 48244 21364 49756
rect 20748 46900 20804 46910
rect 20748 45332 20804 46844
rect 20748 43764 20804 45276
rect 20748 43698 20804 43708
rect 21308 43652 21364 48188
rect 21308 43586 21364 43596
rect 21596 48636 21916 50148
rect 21596 48580 21624 48636
rect 21680 48580 21728 48636
rect 21784 48580 21832 48636
rect 21888 48580 21916 48636
rect 21596 47068 21916 48580
rect 21596 47012 21624 47068
rect 21680 47012 21728 47068
rect 21784 47012 21832 47068
rect 21888 47012 21916 47068
rect 21596 45500 21916 47012
rect 21596 45444 21624 45500
rect 21680 45444 21728 45500
rect 21784 45444 21832 45500
rect 21888 45444 21916 45500
rect 21596 43932 21916 45444
rect 21596 43876 21624 43932
rect 21680 43876 21728 43932
rect 21784 43876 21832 43932
rect 21888 43876 21916 43932
rect 20972 43204 21028 43214
rect 20860 42196 20916 42206
rect 20860 39172 20916 42140
rect 20524 38612 20692 38668
rect 20524 32116 20580 32126
rect 20524 28532 20580 32060
rect 20524 28466 20580 28476
rect 20300 28322 20468 28378
rect 20300 20998 20356 28322
rect 20524 27412 20580 27422
rect 20524 26908 20580 27356
rect 20412 26852 20580 26908
rect 20412 26786 20468 26796
rect 20300 20942 20468 20998
rect 20188 15092 20356 15148
rect 18956 12338 19012 12348
rect 18732 10770 18788 10780
rect 20300 10836 20356 15092
rect 20412 11732 20468 20942
rect 20412 11666 20468 11676
rect 20300 10770 20356 10780
rect 18194 10164 18222 10220
rect 18278 10164 18326 10220
rect 18382 10164 18430 10220
rect 18486 10164 18514 10220
rect 15708 6626 15764 6636
rect 18194 8652 18514 10164
rect 18194 8596 18222 8652
rect 18278 8596 18326 8652
rect 18382 8596 18430 8652
rect 18486 8596 18514 8652
rect 18194 7084 18514 8596
rect 20636 8036 20692 38612
rect 20860 35364 20916 39116
rect 20972 37604 21028 43148
rect 21596 42364 21916 43876
rect 21596 42308 21624 42364
rect 21680 42308 21728 42364
rect 21784 42308 21832 42364
rect 21888 42308 21916 42364
rect 21084 41972 21140 41982
rect 21084 40740 21140 41916
rect 21084 37940 21140 40684
rect 21596 40796 21916 42308
rect 21596 40740 21624 40796
rect 21680 40740 21728 40796
rect 21784 40740 21832 40796
rect 21888 40740 21916 40796
rect 21308 39396 21364 39406
rect 21084 37874 21140 37884
rect 21196 38500 21252 38510
rect 20972 37538 21028 37548
rect 20860 35298 20916 35308
rect 20748 33348 20804 33358
rect 20748 31780 20804 33292
rect 20748 31714 20804 31724
rect 21196 31668 21252 38444
rect 21308 37828 21364 39340
rect 21596 39228 21916 40740
rect 21596 39172 21624 39228
rect 21680 39172 21728 39228
rect 21784 39172 21832 39228
rect 21888 39172 21916 39228
rect 21308 37762 21364 37772
rect 21420 38612 21476 38622
rect 21196 31602 21252 31612
rect 20860 31556 20916 31566
rect 20748 27300 20804 27310
rect 20748 24724 20804 27244
rect 20860 24948 20916 31500
rect 21420 30436 21476 38556
rect 21420 30370 21476 30380
rect 21596 37660 21916 39172
rect 21596 37604 21624 37660
rect 21680 37604 21728 37660
rect 21784 37604 21832 37660
rect 21888 37604 21916 37660
rect 21596 36092 21916 37604
rect 21596 36036 21624 36092
rect 21680 36036 21728 36092
rect 21784 36036 21832 36092
rect 21888 36036 21916 36092
rect 21596 34524 21916 36036
rect 21596 34468 21624 34524
rect 21680 34468 21728 34524
rect 21784 34468 21832 34524
rect 21888 34468 21916 34524
rect 21596 32956 21916 34468
rect 21596 32900 21624 32956
rect 21680 32900 21728 32956
rect 21784 32900 21832 32956
rect 21888 32900 21916 32956
rect 21596 31388 21916 32900
rect 21596 31332 21624 31388
rect 21680 31332 21728 31388
rect 21784 31332 21832 31388
rect 21888 31332 21916 31388
rect 21596 29820 21916 31332
rect 21980 70644 22036 70654
rect 21980 31220 22036 70588
rect 22428 65828 22484 65838
rect 22428 60452 22484 65772
rect 22428 60386 22484 60396
rect 22092 58884 22148 58894
rect 22092 52052 22148 58828
rect 22316 58548 22372 58558
rect 22092 51986 22148 51996
rect 22204 57204 22260 57214
rect 22204 51156 22260 57148
rect 22204 51090 22260 51100
rect 22316 50596 22372 58492
rect 22540 56308 22596 56318
rect 22540 53284 22596 56252
rect 22540 53218 22596 53228
rect 22316 50530 22372 50540
rect 22428 53060 22484 53070
rect 22428 48692 22484 53004
rect 22428 48626 22484 48636
rect 22092 39172 22148 39182
rect 22092 38500 22148 39116
rect 22092 38434 22148 38444
rect 21980 31154 22036 31164
rect 22092 34916 22148 34926
rect 21596 29764 21624 29820
rect 21680 29764 21728 29820
rect 21784 29764 21832 29820
rect 21888 29764 21916 29820
rect 21596 28252 21916 29764
rect 21596 28196 21624 28252
rect 21680 28196 21728 28252
rect 21784 28196 21832 28252
rect 21888 28196 21916 28252
rect 20860 24882 20916 24892
rect 21196 27524 21252 27534
rect 21196 24948 21252 27468
rect 21196 24882 21252 24892
rect 21596 26684 21916 28196
rect 22092 28084 22148 34860
rect 22092 28018 22148 28028
rect 22204 34580 22260 34590
rect 21596 26628 21624 26684
rect 21680 26628 21728 26684
rect 21784 26628 21832 26684
rect 21888 26628 21916 26684
rect 21596 25116 21916 26628
rect 21596 25060 21624 25116
rect 21680 25060 21728 25116
rect 21784 25060 21832 25116
rect 21888 25060 21916 25116
rect 20748 24658 20804 24668
rect 21596 23548 21916 25060
rect 21596 23492 21624 23548
rect 21680 23492 21728 23548
rect 21784 23492 21832 23548
rect 21888 23492 21916 23548
rect 22204 26516 22260 34524
rect 22204 23604 22260 26460
rect 22204 23538 22260 23548
rect 21596 21980 21916 23492
rect 22652 23268 22708 77084
rect 22876 68068 22932 68078
rect 22764 65716 22820 65726
rect 22764 60340 22820 65660
rect 22876 63476 22932 68012
rect 22876 63410 22932 63420
rect 22764 60274 22820 60284
rect 22988 46900 23044 46910
rect 22764 46228 22820 46238
rect 22764 35588 22820 46172
rect 22764 35522 22820 35532
rect 22988 35364 23044 46844
rect 23100 38668 23156 93548
rect 24998 93324 25318 94836
rect 24998 93268 25026 93324
rect 25082 93268 25130 93324
rect 25186 93268 25234 93324
rect 25290 93268 25318 93324
rect 24998 91756 25318 93268
rect 24998 91700 25026 91756
rect 25082 91700 25130 91756
rect 25186 91700 25234 91756
rect 25290 91700 25318 91756
rect 28400 117628 28720 118444
rect 28400 117572 28428 117628
rect 28484 117572 28532 117628
rect 28588 117572 28636 117628
rect 28692 117572 28720 117628
rect 28400 116060 28720 117572
rect 28400 116004 28428 116060
rect 28484 116004 28532 116060
rect 28588 116004 28636 116060
rect 28692 116004 28720 116060
rect 28400 114492 28720 116004
rect 28400 114436 28428 114492
rect 28484 114436 28532 114492
rect 28588 114436 28636 114492
rect 28692 114436 28720 114492
rect 28400 112924 28720 114436
rect 28400 112868 28428 112924
rect 28484 112868 28532 112924
rect 28588 112868 28636 112924
rect 28692 112868 28720 112924
rect 28400 111356 28720 112868
rect 28400 111300 28428 111356
rect 28484 111300 28532 111356
rect 28588 111300 28636 111356
rect 28692 111300 28720 111356
rect 28400 109788 28720 111300
rect 28400 109732 28428 109788
rect 28484 109732 28532 109788
rect 28588 109732 28636 109788
rect 28692 109732 28720 109788
rect 28400 108220 28720 109732
rect 28400 108164 28428 108220
rect 28484 108164 28532 108220
rect 28588 108164 28636 108220
rect 28692 108164 28720 108220
rect 28400 106652 28720 108164
rect 28400 106596 28428 106652
rect 28484 106596 28532 106652
rect 28588 106596 28636 106652
rect 28692 106596 28720 106652
rect 28400 105084 28720 106596
rect 28400 105028 28428 105084
rect 28484 105028 28532 105084
rect 28588 105028 28636 105084
rect 28692 105028 28720 105084
rect 28400 103516 28720 105028
rect 28400 103460 28428 103516
rect 28484 103460 28532 103516
rect 28588 103460 28636 103516
rect 28692 103460 28720 103516
rect 28400 101948 28720 103460
rect 28400 101892 28428 101948
rect 28484 101892 28532 101948
rect 28588 101892 28636 101948
rect 28692 101892 28720 101948
rect 28400 100380 28720 101892
rect 28400 100324 28428 100380
rect 28484 100324 28532 100380
rect 28588 100324 28636 100380
rect 28692 100324 28720 100380
rect 28400 98812 28720 100324
rect 28400 98756 28428 98812
rect 28484 98756 28532 98812
rect 28588 98756 28636 98812
rect 28692 98756 28720 98812
rect 28400 97244 28720 98756
rect 28400 97188 28428 97244
rect 28484 97188 28532 97244
rect 28588 97188 28636 97244
rect 28692 97188 28720 97244
rect 28400 95676 28720 97188
rect 28400 95620 28428 95676
rect 28484 95620 28532 95676
rect 28588 95620 28636 95676
rect 28692 95620 28720 95676
rect 28400 94108 28720 95620
rect 28400 94052 28428 94108
rect 28484 94052 28532 94108
rect 28588 94052 28636 94108
rect 28692 94052 28720 94108
rect 28400 92540 28720 94052
rect 28400 92484 28428 92540
rect 28484 92484 28532 92540
rect 28588 92484 28636 92540
rect 28692 92484 28720 92540
rect 24998 90188 25318 91700
rect 24998 90132 25026 90188
rect 25082 90132 25130 90188
rect 25186 90132 25234 90188
rect 25290 90132 25318 90188
rect 24998 88620 25318 90132
rect 24998 88564 25026 88620
rect 25082 88564 25130 88620
rect 25186 88564 25234 88620
rect 25290 88564 25318 88620
rect 24998 87052 25318 88564
rect 24998 86996 25026 87052
rect 25082 86996 25130 87052
rect 25186 86996 25234 87052
rect 25290 86996 25318 87052
rect 24998 85484 25318 86996
rect 24998 85428 25026 85484
rect 25082 85428 25130 85484
rect 25186 85428 25234 85484
rect 25290 85428 25318 85484
rect 24998 83916 25318 85428
rect 24998 83860 25026 83916
rect 25082 83860 25130 83916
rect 25186 83860 25234 83916
rect 25290 83860 25318 83916
rect 25564 91700 25620 91710
rect 25564 83972 25620 91644
rect 25564 83906 25620 83916
rect 28400 90972 28720 92484
rect 28400 90916 28428 90972
rect 28484 90916 28532 90972
rect 28588 90916 28636 90972
rect 28692 90916 28720 90972
rect 28400 89404 28720 90916
rect 28400 89348 28428 89404
rect 28484 89348 28532 89404
rect 28588 89348 28636 89404
rect 28692 89348 28720 89404
rect 28400 87836 28720 89348
rect 28400 87780 28428 87836
rect 28484 87780 28532 87836
rect 28588 87780 28636 87836
rect 28692 87780 28720 87836
rect 28400 86268 28720 87780
rect 28400 86212 28428 86268
rect 28484 86212 28532 86268
rect 28588 86212 28636 86268
rect 28692 86212 28720 86268
rect 28400 84700 28720 86212
rect 28400 84644 28428 84700
rect 28484 84644 28532 84700
rect 28588 84644 28636 84700
rect 28692 84644 28720 84700
rect 24998 82348 25318 83860
rect 28400 83132 28720 84644
rect 28400 83076 28428 83132
rect 28484 83076 28532 83132
rect 28588 83076 28636 83132
rect 28692 83076 28720 83132
rect 24998 82292 25026 82348
rect 25082 82292 25130 82348
rect 25186 82292 25234 82348
rect 25290 82292 25318 82348
rect 24998 80780 25318 82292
rect 24998 80724 25026 80780
rect 25082 80724 25130 80780
rect 25186 80724 25234 80780
rect 25290 80724 25318 80780
rect 28028 82852 28084 82862
rect 28028 80836 28084 82796
rect 28028 80770 28084 80780
rect 28400 81564 28720 83076
rect 28400 81508 28428 81564
rect 28484 81508 28532 81564
rect 28588 81508 28636 81564
rect 28692 81508 28720 81564
rect 24998 79212 25318 80724
rect 24998 79156 25026 79212
rect 25082 79156 25130 79212
rect 25186 79156 25234 79212
rect 25290 79156 25318 79212
rect 24998 77644 25318 79156
rect 24998 77588 25026 77644
rect 25082 77588 25130 77644
rect 25186 77588 25234 77644
rect 25290 77588 25318 77644
rect 23884 76244 23940 76254
rect 23212 74788 23268 74798
rect 23212 72548 23268 74732
rect 23212 71316 23268 72492
rect 23436 74788 23492 74798
rect 23436 72772 23492 74732
rect 23548 74452 23604 74462
rect 23548 73668 23604 74396
rect 23884 73892 23940 76188
rect 24998 76076 25318 77588
rect 26684 80164 26740 80174
rect 26684 76244 26740 80108
rect 26684 76178 26740 76188
rect 28400 79996 28720 81508
rect 28400 79940 28428 79996
rect 28484 79940 28532 79996
rect 28588 79940 28636 79996
rect 28692 79940 28720 79996
rect 28400 78428 28720 79940
rect 28400 78372 28428 78428
rect 28484 78372 28532 78428
rect 28588 78372 28636 78428
rect 28692 78372 28720 78428
rect 28400 76860 28720 78372
rect 28400 76804 28428 76860
rect 28484 76804 28532 76860
rect 28588 76804 28636 76860
rect 28692 76804 28720 76860
rect 24998 76020 25026 76076
rect 25082 76020 25130 76076
rect 25186 76020 25234 76076
rect 25290 76020 25318 76076
rect 23884 73826 23940 73836
rect 24556 75012 24612 75022
rect 24556 73892 24612 74956
rect 24556 73826 24612 73836
rect 24998 74508 25318 76020
rect 28400 75292 28720 76804
rect 24998 74452 25026 74508
rect 25082 74452 25130 74508
rect 25186 74452 25234 74508
rect 25290 74452 25318 74508
rect 23548 73602 23604 73612
rect 23212 71250 23268 71260
rect 23324 71540 23380 71550
rect 23324 70980 23380 71484
rect 23324 70914 23380 70924
rect 23436 70868 23492 72716
rect 23436 70802 23492 70812
rect 24998 72940 25318 74452
rect 26796 75236 26852 75246
rect 24998 72884 25026 72940
rect 25082 72884 25130 72940
rect 25186 72884 25234 72940
rect 25290 72884 25318 72940
rect 24998 71372 25318 72884
rect 24998 71316 25026 71372
rect 25082 71316 25130 71372
rect 25186 71316 25234 71372
rect 25290 71316 25318 71372
rect 23324 70084 23380 70094
rect 23324 67620 23380 70028
rect 23324 65156 23380 67564
rect 23324 65090 23380 65100
rect 24998 69804 25318 71316
rect 24998 69748 25026 69804
rect 25082 69748 25130 69804
rect 25186 69748 25234 69804
rect 25290 69748 25318 69804
rect 24998 68236 25318 69748
rect 24998 68180 25026 68236
rect 25082 68180 25130 68236
rect 25186 68180 25234 68236
rect 25290 68180 25318 68236
rect 24998 66668 25318 68180
rect 24998 66612 25026 66668
rect 25082 66612 25130 66668
rect 25186 66612 25234 66668
rect 25290 66612 25318 66668
rect 24998 65100 25318 66612
rect 24998 65044 25026 65100
rect 25082 65044 25130 65100
rect 25186 65044 25234 65100
rect 25290 65044 25318 65100
rect 24998 63532 25318 65044
rect 24998 63476 25026 63532
rect 25082 63476 25130 63532
rect 25186 63476 25234 63532
rect 25290 63476 25318 63532
rect 24998 61964 25318 63476
rect 24998 61908 25026 61964
rect 25082 61908 25130 61964
rect 25186 61908 25234 61964
rect 25290 61908 25318 61964
rect 24998 60396 25318 61908
rect 24998 60340 25026 60396
rect 25082 60340 25130 60396
rect 25186 60340 25234 60396
rect 25290 60340 25318 60396
rect 24998 58828 25318 60340
rect 24998 58772 25026 58828
rect 25082 58772 25130 58828
rect 25186 58772 25234 58828
rect 25290 58772 25318 58828
rect 23436 57988 23492 57998
rect 23212 54852 23268 54862
rect 23212 51268 23268 54796
rect 23436 54180 23492 57932
rect 24108 57316 24164 57326
rect 24108 55188 24164 57260
rect 24998 57260 25318 58772
rect 24108 54852 24164 55132
rect 24108 54786 24164 54796
rect 24332 57204 24388 57214
rect 23436 54114 23492 54124
rect 23212 51202 23268 51212
rect 24332 48692 24388 57148
rect 24332 48626 24388 48636
rect 24998 57204 25026 57260
rect 25082 57204 25130 57260
rect 25186 57204 25234 57260
rect 25290 57204 25318 57260
rect 24998 55692 25318 57204
rect 26572 74340 26628 74350
rect 24998 55636 25026 55692
rect 25082 55636 25130 55692
rect 25186 55636 25234 55692
rect 25290 55636 25318 55692
rect 24998 54124 25318 55636
rect 24998 54068 25026 54124
rect 25082 54068 25130 54124
rect 25186 54068 25234 54124
rect 25290 54068 25318 54124
rect 24998 52556 25318 54068
rect 24998 52500 25026 52556
rect 25082 52500 25130 52556
rect 25186 52500 25234 52556
rect 25290 52500 25318 52556
rect 24998 50988 25318 52500
rect 24998 50932 25026 50988
rect 25082 50932 25130 50988
rect 25186 50932 25234 50988
rect 25290 50932 25318 50988
rect 24998 49420 25318 50932
rect 25564 56980 25620 56990
rect 25564 50428 25620 56924
rect 26124 56196 26180 56206
rect 25788 54740 25844 54750
rect 25788 50596 25844 54684
rect 25788 50530 25844 50540
rect 26124 53620 26180 56140
rect 25564 50372 25844 50428
rect 24998 49364 25026 49420
rect 25082 49364 25130 49420
rect 25186 49364 25234 49420
rect 25290 49364 25318 49420
rect 24998 47852 25318 49364
rect 24998 47796 25026 47852
rect 25082 47796 25130 47852
rect 25186 47796 25234 47852
rect 25290 47796 25318 47852
rect 23436 47572 23492 47582
rect 23436 43876 23492 47516
rect 23436 43810 23492 43820
rect 23548 46564 23604 46574
rect 23436 42756 23492 42766
rect 23436 40292 23492 42700
rect 23548 40964 23604 46508
rect 24998 46284 25318 47796
rect 24998 46228 25026 46284
rect 25082 46228 25130 46284
rect 25186 46228 25234 46284
rect 25290 46228 25318 46284
rect 24780 45668 24836 45678
rect 23772 44324 23828 44334
rect 23772 41188 23828 44268
rect 23772 41122 23828 41132
rect 24108 42196 24164 42206
rect 23548 40898 23604 40908
rect 23436 40226 23492 40236
rect 24108 40516 24164 42140
rect 24668 42196 24724 42206
rect 23100 38612 23268 38668
rect 22988 35298 23044 35308
rect 22652 23202 22708 23212
rect 21596 21924 21624 21980
rect 21680 21924 21728 21980
rect 21784 21924 21832 21980
rect 21888 21924 21916 21980
rect 21596 20412 21916 21924
rect 21596 20356 21624 20412
rect 21680 20356 21728 20412
rect 21784 20356 21832 20412
rect 21888 20356 21916 20412
rect 21596 18844 21916 20356
rect 21596 18788 21624 18844
rect 21680 18788 21728 18844
rect 21784 18788 21832 18844
rect 21888 18788 21916 18844
rect 21596 17276 21916 18788
rect 21596 17220 21624 17276
rect 21680 17220 21728 17276
rect 21784 17220 21832 17276
rect 21888 17220 21916 17276
rect 21596 15708 21916 17220
rect 21596 15652 21624 15708
rect 21680 15652 21728 15708
rect 21784 15652 21832 15708
rect 21888 15652 21916 15708
rect 21596 14140 21916 15652
rect 21596 14084 21624 14140
rect 21680 14084 21728 14140
rect 21784 14084 21832 14140
rect 21888 14084 21916 14140
rect 21596 12572 21916 14084
rect 21596 12516 21624 12572
rect 21680 12516 21728 12572
rect 21784 12516 21832 12572
rect 21888 12516 21916 12572
rect 20972 11620 21028 11630
rect 20972 8932 21028 11564
rect 20972 8866 21028 8876
rect 21596 11004 21916 12516
rect 21596 10948 21624 11004
rect 21680 10948 21728 11004
rect 21784 10948 21832 11004
rect 21888 10948 21916 11004
rect 21596 9436 21916 10948
rect 21596 9380 21624 9436
rect 21680 9380 21728 9436
rect 21784 9380 21832 9436
rect 21888 9380 21916 9436
rect 20636 7970 20692 7980
rect 18194 7028 18222 7084
rect 18278 7028 18326 7084
rect 18382 7028 18430 7084
rect 18486 7028 18514 7084
rect 14792 6244 14820 6300
rect 14876 6244 14924 6300
rect 14980 6244 15028 6300
rect 15084 6244 15112 6300
rect 14792 4732 15112 6244
rect 14792 4676 14820 4732
rect 14876 4676 14924 4732
rect 14980 4676 15028 4732
rect 15084 4676 15112 4732
rect 14792 3164 15112 4676
rect 18194 5516 18514 7028
rect 18194 5460 18222 5516
rect 18278 5460 18326 5516
rect 18382 5460 18430 5516
rect 18486 5460 18514 5516
rect 14792 3108 14820 3164
rect 14876 3108 14924 3164
rect 14980 3108 15028 3164
rect 15084 3108 15112 3164
rect 14792 1596 15112 3108
rect 18060 4116 18116 4126
rect 18060 2212 18116 4060
rect 18060 2146 18116 2156
rect 18194 3948 18514 5460
rect 18194 3892 18222 3948
rect 18278 3892 18326 3948
rect 18382 3892 18430 3948
rect 18486 3892 18514 3948
rect 18194 2380 18514 3892
rect 21596 7868 21916 9380
rect 21596 7812 21624 7868
rect 21680 7812 21728 7868
rect 21784 7812 21832 7868
rect 21888 7812 21916 7868
rect 21596 6300 21916 7812
rect 21596 6244 21624 6300
rect 21680 6244 21728 6300
rect 21784 6244 21832 6300
rect 21888 6244 21916 6300
rect 21596 4732 21916 6244
rect 21596 4676 21624 4732
rect 21680 4676 21728 4732
rect 21784 4676 21832 4732
rect 21888 4676 21916 4732
rect 19852 3444 19908 3454
rect 19852 2772 19908 3388
rect 19852 2706 19908 2716
rect 21596 3164 21916 4676
rect 23212 3556 23268 38612
rect 24108 37940 24164 40460
rect 24108 37874 24164 37884
rect 24332 42084 24388 42094
rect 23660 37828 23716 37838
rect 23324 33684 23380 33694
rect 23324 26740 23380 33628
rect 23660 33684 23716 37772
rect 24332 37604 24388 42028
rect 24668 41636 24724 42140
rect 24780 41972 24836 45612
rect 24780 41906 24836 41916
rect 24998 44716 25318 46228
rect 24998 44660 25026 44716
rect 25082 44660 25130 44716
rect 25186 44660 25234 44716
rect 25290 44660 25318 44716
rect 24998 43148 25318 44660
rect 24998 43092 25026 43148
rect 25082 43092 25130 43148
rect 25186 43092 25234 43148
rect 25290 43092 25318 43148
rect 24668 41570 24724 41580
rect 24998 41580 25318 43092
rect 25452 43764 25508 43774
rect 25452 41860 25508 43708
rect 25452 41794 25508 41804
rect 24332 37538 24388 37548
rect 24998 41524 25026 41580
rect 25082 41524 25130 41580
rect 25186 41524 25234 41580
rect 25290 41524 25318 41580
rect 24998 40012 25318 41524
rect 24998 39956 25026 40012
rect 25082 39956 25130 40012
rect 25186 39956 25234 40012
rect 25290 39956 25318 40012
rect 24998 38444 25318 39956
rect 24998 38388 25026 38444
rect 25082 38388 25130 38444
rect 25186 38388 25234 38444
rect 25290 38388 25318 38444
rect 24780 37044 24836 37054
rect 24780 36596 24836 36988
rect 24780 36530 24836 36540
rect 24998 36876 25318 38388
rect 24998 36820 25026 36876
rect 25082 36820 25130 36876
rect 25186 36820 25234 36876
rect 25290 36820 25318 36876
rect 24998 35308 25318 36820
rect 25452 40852 25508 40862
rect 25452 37492 25508 40796
rect 25452 35476 25508 37436
rect 25452 35410 25508 35420
rect 24668 35252 24724 35262
rect 24668 34804 24724 35196
rect 24668 34738 24724 34748
rect 24998 35252 25026 35308
rect 25082 35252 25130 35308
rect 25186 35252 25234 35308
rect 25290 35252 25318 35308
rect 23660 33618 23716 33628
rect 24998 33740 25318 35252
rect 24998 33684 25026 33740
rect 25082 33684 25130 33740
rect 25186 33684 25234 33740
rect 25290 33684 25318 33740
rect 24444 33460 24500 33470
rect 23548 31892 23604 31902
rect 23548 30772 23604 31836
rect 23548 30706 23604 30716
rect 23324 26674 23380 26684
rect 23548 28196 23604 28206
rect 23548 25956 23604 28140
rect 23548 25890 23604 25900
rect 24444 25172 24500 33404
rect 24780 32228 24836 32238
rect 24780 29316 24836 32172
rect 24780 28532 24836 29260
rect 24780 28466 24836 28476
rect 24998 32172 25318 33684
rect 24998 32116 25026 32172
rect 25082 32116 25130 32172
rect 25186 32116 25234 32172
rect 25290 32116 25318 32172
rect 24998 30604 25318 32116
rect 24998 30548 25026 30604
rect 25082 30548 25130 30604
rect 25186 30548 25234 30604
rect 25290 30548 25318 30604
rect 24998 29036 25318 30548
rect 24998 28980 25026 29036
rect 25082 28980 25130 29036
rect 25186 28980 25234 29036
rect 25290 28980 25318 29036
rect 24444 25106 24500 25116
rect 24998 27468 25318 28980
rect 24998 27412 25026 27468
rect 25082 27412 25130 27468
rect 25186 27412 25234 27468
rect 25290 27412 25318 27468
rect 24998 25900 25318 27412
rect 24998 25844 25026 25900
rect 25082 25844 25130 25900
rect 25186 25844 25234 25900
rect 25290 25844 25318 25900
rect 24998 24332 25318 25844
rect 25452 34468 25508 34478
rect 25452 24948 25508 34412
rect 25564 32676 25620 32686
rect 25564 28868 25620 32620
rect 25788 31668 25844 50372
rect 26124 48132 26180 53564
rect 26348 56084 26404 56094
rect 26348 49028 26404 56028
rect 26348 48962 26404 48972
rect 26124 48066 26180 48076
rect 26572 43316 26628 74284
rect 26796 74340 26852 75180
rect 26796 74274 26852 74284
rect 28400 75236 28428 75292
rect 28484 75236 28532 75292
rect 28588 75236 28636 75292
rect 28692 75236 28720 75292
rect 28400 73724 28720 75236
rect 28400 73668 28428 73724
rect 28484 73668 28532 73724
rect 28588 73668 28636 73724
rect 28692 73668 28720 73724
rect 28400 72156 28720 73668
rect 28400 72100 28428 72156
rect 28484 72100 28532 72156
rect 28588 72100 28636 72156
rect 28692 72100 28720 72156
rect 28400 70588 28720 72100
rect 28400 70532 28428 70588
rect 28484 70532 28532 70588
rect 28588 70532 28636 70588
rect 28692 70532 28720 70588
rect 28400 69020 28720 70532
rect 28400 68964 28428 69020
rect 28484 68964 28532 69020
rect 28588 68964 28636 69020
rect 28692 68964 28720 69020
rect 28400 67452 28720 68964
rect 28400 67396 28428 67452
rect 28484 67396 28532 67452
rect 28588 67396 28636 67452
rect 28692 67396 28720 67452
rect 28400 65884 28720 67396
rect 28400 65828 28428 65884
rect 28484 65828 28532 65884
rect 28588 65828 28636 65884
rect 28692 65828 28720 65884
rect 28400 64316 28720 65828
rect 28400 64260 28428 64316
rect 28484 64260 28532 64316
rect 28588 64260 28636 64316
rect 28692 64260 28720 64316
rect 26684 64148 26740 64158
rect 26684 63588 26740 64092
rect 26684 63522 26740 63532
rect 28400 62748 28720 64260
rect 28400 62692 28428 62748
rect 28484 62692 28532 62748
rect 28588 62692 28636 62748
rect 28692 62692 28720 62748
rect 28400 61180 28720 62692
rect 28400 61124 28428 61180
rect 28484 61124 28532 61180
rect 28588 61124 28636 61180
rect 28692 61124 28720 61180
rect 28400 59612 28720 61124
rect 28400 59556 28428 59612
rect 28484 59556 28532 59612
rect 28588 59556 28636 59612
rect 28692 59556 28720 59612
rect 28400 58044 28720 59556
rect 28400 57988 28428 58044
rect 28484 57988 28532 58044
rect 28588 57988 28636 58044
rect 28692 57988 28720 58044
rect 28400 56476 28720 57988
rect 28400 56420 28428 56476
rect 28484 56420 28532 56476
rect 28588 56420 28636 56476
rect 28692 56420 28720 56476
rect 28400 54908 28720 56420
rect 28400 54852 28428 54908
rect 28484 54852 28532 54908
rect 28588 54852 28636 54908
rect 28692 54852 28720 54908
rect 26684 54404 26740 54414
rect 26684 53396 26740 54348
rect 26684 53330 26740 53340
rect 28400 53340 28720 54852
rect 26572 43250 26628 43260
rect 28400 53284 28428 53340
rect 28484 53284 28532 53340
rect 28588 53284 28636 53340
rect 28692 53284 28720 53340
rect 28400 51772 28720 53284
rect 28400 51716 28428 51772
rect 28484 51716 28532 51772
rect 28588 51716 28636 51772
rect 28692 51716 28720 51772
rect 28400 50204 28720 51716
rect 28400 50148 28428 50204
rect 28484 50148 28532 50204
rect 28588 50148 28636 50204
rect 28692 50148 28720 50204
rect 28400 48636 28720 50148
rect 28400 48580 28428 48636
rect 28484 48580 28532 48636
rect 28588 48580 28636 48636
rect 28692 48580 28720 48636
rect 28400 47068 28720 48580
rect 28400 47012 28428 47068
rect 28484 47012 28532 47068
rect 28588 47012 28636 47068
rect 28692 47012 28720 47068
rect 28400 45500 28720 47012
rect 28400 45444 28428 45500
rect 28484 45444 28532 45500
rect 28588 45444 28636 45500
rect 28692 45444 28720 45500
rect 28400 43932 28720 45444
rect 28400 43876 28428 43932
rect 28484 43876 28532 43932
rect 28588 43876 28636 43932
rect 28692 43876 28720 43932
rect 28400 42364 28720 43876
rect 28400 42308 28428 42364
rect 28484 42308 28532 42364
rect 28588 42308 28636 42364
rect 28692 42308 28720 42364
rect 28400 40796 28720 42308
rect 28400 40740 28428 40796
rect 28484 40740 28532 40796
rect 28588 40740 28636 40796
rect 28692 40740 28720 40796
rect 28400 39228 28720 40740
rect 28400 39172 28428 39228
rect 28484 39172 28532 39228
rect 28588 39172 28636 39228
rect 28692 39172 28720 39228
rect 28400 37660 28720 39172
rect 28400 37604 28428 37660
rect 28484 37604 28532 37660
rect 28588 37604 28636 37660
rect 28692 37604 28720 37660
rect 26796 37380 26852 37390
rect 26796 36372 26852 37324
rect 26796 36306 26852 36316
rect 25788 31602 25844 31612
rect 28400 36092 28720 37604
rect 28400 36036 28428 36092
rect 28484 36036 28532 36092
rect 28588 36036 28636 36092
rect 28692 36036 28720 36092
rect 28400 34524 28720 36036
rect 28400 34468 28428 34524
rect 28484 34468 28532 34524
rect 28588 34468 28636 34524
rect 28692 34468 28720 34524
rect 28400 32956 28720 34468
rect 28400 32900 28428 32956
rect 28484 32900 28532 32956
rect 28588 32900 28636 32956
rect 28692 32900 28720 32956
rect 28400 31388 28720 32900
rect 28400 31332 28428 31388
rect 28484 31332 28532 31388
rect 28588 31332 28636 31388
rect 28692 31332 28720 31388
rect 26124 31108 26180 31118
rect 25564 28308 25620 28812
rect 25788 30884 25844 30894
rect 25788 28420 25844 30828
rect 25788 28354 25844 28364
rect 25564 28242 25620 28252
rect 26124 27412 26180 31052
rect 28400 29820 28720 31332
rect 28400 29764 28428 29820
rect 28484 29764 28532 29820
rect 28588 29764 28636 29820
rect 28692 29764 28720 29820
rect 26684 28308 26740 28318
rect 26684 27860 26740 28252
rect 26684 27794 26740 27804
rect 28400 28252 28720 29764
rect 28400 28196 28428 28252
rect 28484 28196 28532 28252
rect 28588 28196 28636 28252
rect 28692 28196 28720 28252
rect 26124 27346 26180 27356
rect 25452 24882 25508 24892
rect 28400 26684 28720 28196
rect 28400 26628 28428 26684
rect 28484 26628 28532 26684
rect 28588 26628 28636 26684
rect 28692 26628 28720 26684
rect 28400 25116 28720 26628
rect 28400 25060 28428 25116
rect 28484 25060 28532 25116
rect 28588 25060 28636 25116
rect 28692 25060 28720 25116
rect 24998 24276 25026 24332
rect 25082 24276 25130 24332
rect 25186 24276 25234 24332
rect 25290 24276 25318 24332
rect 23772 23492 23828 23502
rect 23772 22372 23828 23436
rect 23772 22306 23828 22316
rect 24998 22764 25318 24276
rect 26684 24276 26740 24286
rect 26684 23380 26740 24220
rect 26684 23314 26740 23324
rect 28400 23548 28720 25060
rect 28400 23492 28428 23548
rect 28484 23492 28532 23548
rect 28588 23492 28636 23548
rect 28692 23492 28720 23548
rect 24998 22708 25026 22764
rect 25082 22708 25130 22764
rect 25186 22708 25234 22764
rect 25290 22708 25318 22764
rect 23212 3490 23268 3500
rect 24998 21196 25318 22708
rect 24998 21140 25026 21196
rect 25082 21140 25130 21196
rect 25186 21140 25234 21196
rect 25290 21140 25318 21196
rect 24998 19628 25318 21140
rect 24998 19572 25026 19628
rect 25082 19572 25130 19628
rect 25186 19572 25234 19628
rect 25290 19572 25318 19628
rect 24998 18060 25318 19572
rect 24998 18004 25026 18060
rect 25082 18004 25130 18060
rect 25186 18004 25234 18060
rect 25290 18004 25318 18060
rect 24998 16492 25318 18004
rect 24998 16436 25026 16492
rect 25082 16436 25130 16492
rect 25186 16436 25234 16492
rect 25290 16436 25318 16492
rect 24998 14924 25318 16436
rect 24998 14868 25026 14924
rect 25082 14868 25130 14924
rect 25186 14868 25234 14924
rect 25290 14868 25318 14924
rect 24998 13356 25318 14868
rect 24998 13300 25026 13356
rect 25082 13300 25130 13356
rect 25186 13300 25234 13356
rect 25290 13300 25318 13356
rect 24998 11788 25318 13300
rect 24998 11732 25026 11788
rect 25082 11732 25130 11788
rect 25186 11732 25234 11788
rect 25290 11732 25318 11788
rect 24998 10220 25318 11732
rect 24998 10164 25026 10220
rect 25082 10164 25130 10220
rect 25186 10164 25234 10220
rect 25290 10164 25318 10220
rect 24998 8652 25318 10164
rect 24998 8596 25026 8652
rect 25082 8596 25130 8652
rect 25186 8596 25234 8652
rect 25290 8596 25318 8652
rect 24998 7084 25318 8596
rect 24998 7028 25026 7084
rect 25082 7028 25130 7084
rect 25186 7028 25234 7084
rect 25290 7028 25318 7084
rect 24998 5516 25318 7028
rect 24998 5460 25026 5516
rect 25082 5460 25130 5516
rect 25186 5460 25234 5516
rect 25290 5460 25318 5516
rect 24998 3948 25318 5460
rect 24998 3892 25026 3948
rect 25082 3892 25130 3948
rect 25186 3892 25234 3948
rect 25290 3892 25318 3948
rect 21596 3108 21624 3164
rect 21680 3108 21728 3164
rect 21784 3108 21832 3164
rect 21888 3108 21916 3164
rect 18194 2324 18222 2380
rect 18278 2324 18326 2380
rect 18382 2324 18430 2380
rect 18486 2324 18514 2380
rect 14792 1540 14820 1596
rect 14876 1540 14924 1596
rect 14980 1540 15028 1596
rect 15084 1540 15112 1596
rect 14792 1508 15112 1540
rect 18194 1508 18514 2324
rect 21596 1596 21916 3108
rect 21596 1540 21624 1596
rect 21680 1540 21728 1596
rect 21784 1540 21832 1596
rect 21888 1540 21916 1596
rect 21596 1508 21916 1540
rect 24998 2380 25318 3892
rect 24998 2324 25026 2380
rect 25082 2324 25130 2380
rect 25186 2324 25234 2380
rect 25290 2324 25318 2380
rect 24998 1508 25318 2324
rect 28400 21980 28720 23492
rect 28400 21924 28428 21980
rect 28484 21924 28532 21980
rect 28588 21924 28636 21980
rect 28692 21924 28720 21980
rect 28400 20412 28720 21924
rect 28400 20356 28428 20412
rect 28484 20356 28532 20412
rect 28588 20356 28636 20412
rect 28692 20356 28720 20412
rect 28400 18844 28720 20356
rect 28400 18788 28428 18844
rect 28484 18788 28532 18844
rect 28588 18788 28636 18844
rect 28692 18788 28720 18844
rect 28400 17276 28720 18788
rect 28400 17220 28428 17276
rect 28484 17220 28532 17276
rect 28588 17220 28636 17276
rect 28692 17220 28720 17276
rect 28400 15708 28720 17220
rect 28400 15652 28428 15708
rect 28484 15652 28532 15708
rect 28588 15652 28636 15708
rect 28692 15652 28720 15708
rect 28400 14140 28720 15652
rect 28400 14084 28428 14140
rect 28484 14084 28532 14140
rect 28588 14084 28636 14140
rect 28692 14084 28720 14140
rect 28400 12572 28720 14084
rect 28400 12516 28428 12572
rect 28484 12516 28532 12572
rect 28588 12516 28636 12572
rect 28692 12516 28720 12572
rect 28400 11004 28720 12516
rect 28400 10948 28428 11004
rect 28484 10948 28532 11004
rect 28588 10948 28636 11004
rect 28692 10948 28720 11004
rect 28400 9436 28720 10948
rect 28400 9380 28428 9436
rect 28484 9380 28532 9436
rect 28588 9380 28636 9436
rect 28692 9380 28720 9436
rect 28400 7868 28720 9380
rect 28400 7812 28428 7868
rect 28484 7812 28532 7868
rect 28588 7812 28636 7868
rect 28692 7812 28720 7868
rect 28400 6300 28720 7812
rect 28400 6244 28428 6300
rect 28484 6244 28532 6300
rect 28588 6244 28636 6300
rect 28692 6244 28720 6300
rect 28400 4732 28720 6244
rect 28400 4676 28428 4732
rect 28484 4676 28532 4732
rect 28588 4676 28636 4732
rect 28692 4676 28720 4732
rect 28400 3164 28720 4676
rect 28400 3108 28428 3164
rect 28484 3108 28532 3164
rect 28588 3108 28636 3164
rect 28692 3108 28720 3164
rect 28400 1596 28720 3108
rect 28400 1540 28428 1596
rect 28484 1540 28532 1596
rect 28588 1540 28636 1596
rect 28692 1540 28720 1596
rect 28400 1508 28720 1540
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _0979_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0980_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0981_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4592 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _0982_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7504 0 1 101920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  _0983_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 1 101920
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0984_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7728 0 1 100352
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0985_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 -1 95648
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0986_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6832 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0987_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10864 0 -1 94080
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0988_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 95648
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0989_
timestamp 1698431365
transform 1 0 21392 0 1 98784
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0990_
timestamp 1698431365
transform 1 0 23744 0 -1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0991_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23744 0 1 97216
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0992_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23520 0 1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0993_
timestamp 1698431365
transform -1 0 7728 0 1 100352
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0994_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 1 95648
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0995_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21952 0 -1 97216
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0996_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10640 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0997_
timestamp 1698431365
transform 1 0 9408 0 -1 100352
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0998_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 95648
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0999_
timestamp 1698431365
transform 1 0 14224 0 -1 97216
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1000_
timestamp 1698431365
transform -1 0 12880 0 -1 97216
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1001_
timestamp 1698431365
transform -1 0 11424 0 -1 101920
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1002_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 100352
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1003_
timestamp 1698431365
transform -1 0 16688 0 -1 103488
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1004_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10192 0 -1 103488
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1005_
timestamp 1698431365
transform -1 0 9072 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1006_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8512 0 -1 105056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1007_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9520 0 1 84672
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  _1008_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14336 0 -1 84672
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1009_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16240 0 -1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1010_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _1011_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 87808
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  _1012_
timestamp 1698431365
transform 1 0 13440 0 1 86240
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  _1013_
timestamp 1698431365
transform 1 0 17472 0 -1 84672
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1014_
timestamp 1698431365
transform -1 0 21616 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _1015_
timestamp 1698431365
transform 1 0 12096 0 -1 81536
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1016_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16576 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1017_
timestamp 1698431365
transform 1 0 10192 0 1 89376
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_12  _1018_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 87808
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _1019_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1020_
timestamp 1698431365
transform -1 0 16800 0 1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1021_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  _1022_
timestamp 1698431365
transform 1 0 9408 0 -1 78400
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1023_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15456 0 1 51744
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1024_
timestamp 1698431365
transform -1 0 11424 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  _1025_
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1026_
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1027_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14560 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1028_
timestamp 1698431365
transform -1 0 13776 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1029_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3920 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1030_
timestamp 1698431365
transform 1 0 20832 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  _1031_
timestamp 1698431365
transform 1 0 11088 0 -1 79968
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1032_
timestamp 1698431365
transform -1 0 16688 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1033_
timestamp 1698431365
transform -1 0 14672 0 -1 68992
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1034_
timestamp 1698431365
transform -1 0 26992 0 1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1035_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1036_
timestamp 1698431365
transform 1 0 16016 0 1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1037_
timestamp 1698431365
transform 1 0 15232 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1038_
timestamp 1698431365
transform 1 0 14000 0 1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1039_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1040_
timestamp 1698431365
transform 1 0 12880 0 -1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1041_
timestamp 1698431365
transform -1 0 25088 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1042_
timestamp 1698431365
transform 1 0 20160 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1043_
timestamp 1698431365
transform -1 0 22064 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1044_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20160 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1045_
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1046_
timestamp 1698431365
transform 1 0 14560 0 1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1047_
timestamp 1698431365
transform -1 0 24192 0 -1 72128
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1048_
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1049_
timestamp 1698431365
transform 1 0 12880 0 -1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1050_
timestamp 1698431365
transform -1 0 24416 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1051_
timestamp 1698431365
transform 1 0 15232 0 1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1052_
timestamp 1698431365
transform -1 0 17024 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1053_
timestamp 1698431365
transform 1 0 10416 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1054_
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1055_
timestamp 1698431365
transform 1 0 11424 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1056_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14784 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1057_
timestamp 1698431365
transform -1 0 20832 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1058_
timestamp 1698431365
transform 1 0 16800 0 1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1059_
timestamp 1698431365
transform 1 0 21392 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1060_
timestamp 1698431365
transform -1 0 19824 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1061_
timestamp 1698431365
transform -1 0 20496 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1062_
timestamp 1698431365
transform 1 0 7616 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1063_
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1064_
timestamp 1698431365
transform -1 0 14336 0 1 68992
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1065_
timestamp 1698431365
transform 1 0 12432 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1066_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12096 0 -1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1067_
timestamp 1698431365
transform 1 0 13440 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1068_
timestamp 1698431365
transform -1 0 17024 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1069_
timestamp 1698431365
transform -1 0 18592 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1070_
timestamp 1698431365
transform 1 0 13440 0 1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1071_
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1072_
timestamp 1698431365
transform -1 0 13104 0 -1 61152
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1073_
timestamp 1698431365
transform 1 0 13104 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1074_
timestamp 1698431365
transform 1 0 15344 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1075_
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1076_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9296 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1077_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13216 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1078_
timestamp 1698431365
transform 1 0 15120 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1079_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10416 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1080_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12768 0 1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1081_
timestamp 1698431365
transform -1 0 14784 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1082_
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1083_
timestamp 1698431365
transform -1 0 12880 0 -1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1084_
timestamp 1698431365
transform -1 0 17024 0 -1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1085_
timestamp 1698431365
transform 1 0 9184 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1086_
timestamp 1698431365
transform 1 0 15680 0 1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1087_
timestamp 1698431365
transform -1 0 17024 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1088_
timestamp 1698431365
transform 1 0 11536 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1089_
timestamp 1698431365
transform 1 0 10192 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1090_
timestamp 1698431365
transform -1 0 18480 0 -1 72128
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1091_
timestamp 1698431365
transform 1 0 19152 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1092_
timestamp 1698431365
transform 1 0 21168 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1093_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 86240
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1094_
timestamp 1698431365
transform 1 0 13440 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1095_
timestamp 1698431365
transform 1 0 4928 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1096_
timestamp 1698431365
transform -1 0 26992 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1097_
timestamp 1698431365
transform -1 0 20272 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1098_
timestamp 1698431365
transform -1 0 23968 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1099_
timestamp 1698431365
transform 1 0 21056 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1100_
timestamp 1698431365
transform -1 0 23184 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1101_
timestamp 1698431365
transform 1 0 19600 0 1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1102_
timestamp 1698431365
transform 1 0 22848 0 1 72128
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1103_
timestamp 1698431365
transform 1 0 22512 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1104_
timestamp 1698431365
transform 1 0 9856 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1105_
timestamp 1698431365
transform 1 0 17472 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1106_
timestamp 1698431365
transform 1 0 18144 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1107_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1108_
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1109_
timestamp 1698431365
transform 1 0 12432 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1110_
timestamp 1698431365
transform 1 0 4816 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1111_
timestamp 1698431365
transform 1 0 10416 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1112_
timestamp 1698431365
transform 1 0 12320 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1113_
timestamp 1698431365
transform -1 0 15120 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1114_
timestamp 1698431365
transform 1 0 12992 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1115_
timestamp 1698431365
transform 1 0 8176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1116_
timestamp 1698431365
transform 1 0 8176 0 1 72128
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1117_
timestamp 1698431365
transform -1 0 9184 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1118_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1119_
timestamp 1698431365
transform -1 0 10528 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1120_
timestamp 1698431365
transform 1 0 7952 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1121_
timestamp 1698431365
transform 1 0 10192 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1122_
timestamp 1698431365
transform 1 0 11872 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1123_
timestamp 1698431365
transform 1 0 10528 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1124_
timestamp 1698431365
transform -1 0 18480 0 -1 73696
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1125_
timestamp 1698431365
transform -1 0 19936 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1126_
timestamp 1698431365
transform 1 0 18816 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1127_
timestamp 1698431365
transform 1 0 17472 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1128_
timestamp 1698431365
transform -1 0 23408 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1129_
timestamp 1698431365
transform 1 0 3920 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1130_
timestamp 1698431365
transform -1 0 28000 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1131_
timestamp 1698431365
transform -1 0 19040 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1132_
timestamp 1698431365
transform -1 0 19936 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1133_
timestamp 1698431365
transform 1 0 17808 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1134_
timestamp 1698431365
transform -1 0 19488 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1135_
timestamp 1698431365
transform 1 0 18256 0 -1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1136_
timestamp 1698431365
transform 1 0 22624 0 1 67424
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1137_
timestamp 1698431365
transform -1 0 23744 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1138_
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1139_
timestamp 1698431365
transform -1 0 20720 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1140_
timestamp 1698431365
transform 1 0 19488 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1141_
timestamp 1698431365
transform -1 0 20384 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1142_
timestamp 1698431365
transform 1 0 16016 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1143_
timestamp 1698431365
transform 1 0 9520 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1144_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11088 0 -1 79968
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1145_
timestamp 1698431365
transform -1 0 24640 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1146_
timestamp 1698431365
transform -1 0 25872 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1147_
timestamp 1698431365
transform 1 0 15344 0 -1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1148_
timestamp 1698431365
transform 1 0 8064 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1149_
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1150_
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1151_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 70560
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1152_
timestamp 1698431365
transform 1 0 11088 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1153_
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1154_
timestamp 1698431365
transform 1 0 9408 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1155_
timestamp 1698431365
transform 1 0 9968 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1156_
timestamp 1698431365
transform 1 0 9856 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1157_
timestamp 1698431365
transform -1 0 19936 0 -1 67424
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1158_
timestamp 1698431365
transform 1 0 19152 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1159_
timestamp 1698431365
transform 1 0 21168 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1160_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23072 0 -1 79968
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1161_
timestamp 1698431365
transform -1 0 18368 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1162_
timestamp 1698431365
transform 1 0 4032 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1163_
timestamp 1698431365
transform -1 0 22400 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1164_
timestamp 1698431365
transform 1 0 14336 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1165_
timestamp 1698431365
transform 1 0 12320 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1166_
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1167_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1168_
timestamp 1698431365
transform -1 0 20832 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1169_
timestamp 1698431365
transform 1 0 22736 0 -1 65856
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1170_
timestamp 1698431365
transform -1 0 19600 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1171_
timestamp 1698431365
transform -1 0 17024 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1172_
timestamp 1698431365
transform -1 0 19264 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1173_
timestamp 1698431365
transform 1 0 19264 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1174_
timestamp 1698431365
transform -1 0 19264 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1175_
timestamp 1698431365
transform 1 0 15120 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1176_
timestamp 1698431365
transform -1 0 7056 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1177_
timestamp 1698431365
transform -1 0 13104 0 1 78400
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1178_
timestamp 1698431365
transform 1 0 14112 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1179_
timestamp 1698431365
transform -1 0 27216 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1180_
timestamp 1698431365
transform 1 0 14784 0 1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1181_
timestamp 1698431365
transform 1 0 8176 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1182_
timestamp 1698431365
transform 1 0 8176 0 -1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1183_
timestamp 1698431365
transform -1 0 9632 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1184_
timestamp 1698431365
transform 1 0 15120 0 1 68992
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1185_
timestamp 1698431365
transform 1 0 10080 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1186_
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1187_
timestamp 1698431365
transform 1 0 10304 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1188_
timestamp 1698431365
transform 1 0 10304 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1189_
timestamp 1698431365
transform 1 0 9856 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1190_
timestamp 1698431365
transform -1 0 18480 0 -1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1191_
timestamp 1698431365
transform -1 0 19152 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1192_
timestamp 1698431365
transform 1 0 21168 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1193_
timestamp 1698431365
transform 1 0 19600 0 -1 81536
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1194_
timestamp 1698431365
transform 1 0 19152 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1195_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18592 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1196_
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1197_
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1198_
timestamp 1698431365
transform -1 0 18928 0 1 56448
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1199_
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1200_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1201_
timestamp 1698431365
transform -1 0 23072 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1202_
timestamp 1698431365
transform 1 0 7728 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1203_
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1204_
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1205_
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1206_
timestamp 1698431365
transform -1 0 21840 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1207_
timestamp 1698431365
transform -1 0 11648 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1208_
timestamp 1698431365
transform -1 0 21168 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1209_
timestamp 1698431365
transform 1 0 20272 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1210_
timestamp 1698431365
transform 1 0 19488 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1211_
timestamp 1698431365
transform -1 0 20720 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1212_
timestamp 1698431365
transform -1 0 22624 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1213_
timestamp 1698431365
transform -1 0 23856 0 -1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1214_
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1215_
timestamp 1698431365
transform 1 0 9632 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1216_
timestamp 1698431365
transform 1 0 14448 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1217_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13776 0 1 61152
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1218_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14000 0 -1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1219_
timestamp 1698431365
transform -1 0 14672 0 1 59584
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1220_
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1221_
timestamp 1698431365
transform 1 0 15904 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1222_
timestamp 1698431365
transform -1 0 19040 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1223_
timestamp 1698431365
transform -1 0 14672 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1224_
timestamp 1698431365
transform 1 0 13328 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1225_
timestamp 1698431365
transform 1 0 14560 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1226_
timestamp 1698431365
transform -1 0 15568 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1227_
timestamp 1698431365
transform 1 0 16240 0 1 58016
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1228_
timestamp 1698431365
transform -1 0 24864 0 1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1229_
timestamp 1698431365
transform 1 0 11984 0 1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1230_
timestamp 1698431365
transform 1 0 14224 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1231_
timestamp 1698431365
transform 1 0 14672 0 1 59584
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1232_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22960 0 -1 72128
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1233_
timestamp 1698431365
transform 1 0 17696 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1234_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20720 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1235_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1236_
timestamp 1698431365
transform 1 0 12432 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1237_
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1238_
timestamp 1698431365
transform -1 0 9408 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1239_
timestamp 1698431365
transform -1 0 19040 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1240_
timestamp 1698431365
transform 1 0 13440 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1241_
timestamp 1698431365
transform -1 0 12432 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1242_
timestamp 1698431365
transform -1 0 24080 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1243_
timestamp 1698431365
transform 1 0 15568 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1244_
timestamp 1698431365
transform -1 0 17696 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1245_
timestamp 1698431365
transform -1 0 12880 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1246_
timestamp 1698431365
transform -1 0 16912 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1247_
timestamp 1698431365
transform 1 0 15792 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1248_
timestamp 1698431365
transform -1 0 19712 0 1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1249_
timestamp 1698431365
transform -1 0 11424 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1250_
timestamp 1698431365
transform 1 0 9632 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1251_
timestamp 1698431365
transform 1 0 15904 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1252_
timestamp 1698431365
transform -1 0 15344 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1253_
timestamp 1698431365
transform -1 0 15904 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1254_
timestamp 1698431365
transform 1 0 15456 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1255_
timestamp 1698431365
transform -1 0 17024 0 -1 59584
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1256_
timestamp 1698431365
transform -1 0 13104 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1257_
timestamp 1698431365
transform 1 0 11312 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1258_
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1259_
timestamp 1698431365
transform 1 0 14560 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1260_
timestamp 1698431365
transform -1 0 23408 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1261_
timestamp 1698431365
transform 1 0 14112 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1262_
timestamp 1698431365
transform 1 0 15232 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1263_
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1264_
timestamp 1698431365
transform -1 0 18144 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1265_
timestamp 1698431365
transform 1 0 17696 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1266_
timestamp 1698431365
transform 1 0 19152 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1267_
timestamp 1698431365
transform 1 0 12208 0 -1 83104
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1268_
timestamp 1698431365
transform -1 0 16016 0 1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1269_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18480 0 1 84672
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1270_
timestamp 1698431365
transform -1 0 14224 0 1 92512
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1271_
timestamp 1698431365
transform -1 0 12656 0 -1 94080
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1272_
timestamp 1698431365
transform 1 0 15456 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1273_
timestamp 1698431365
transform -1 0 13888 0 1 90944
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1274_
timestamp 1698431365
transform 1 0 13104 0 -1 90944
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1275_
timestamp 1698431365
transform -1 0 13104 0 1 90944
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1276_
timestamp 1698431365
transform -1 0 15904 0 1 90944
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1277_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20160 0 -1 94080
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1278_
timestamp 1698431365
transform -1 0 19376 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1279_
timestamp 1698431365
transform 1 0 15456 0 -1 89376
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1280_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 1 89376
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1281_
timestamp 1698431365
transform 1 0 15792 0 -1 86240
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1282_
timestamp 1698431365
transform -1 0 18816 0 1 87808
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1283_
timestamp 1698431365
transform 1 0 15456 0 1 86240
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1284_
timestamp 1698431365
transform 1 0 18704 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1285_
timestamp 1698431365
transform -1 0 18704 0 1 90944
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1286_
timestamp 1698431365
transform -1 0 20272 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1287_
timestamp 1698431365
transform -1 0 17360 0 1 90944
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1288_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17808 0 1 94080
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1289_
timestamp 1698431365
transform 1 0 15792 0 1 92512
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1290_
timestamp 1698431365
transform -1 0 18816 0 1 92512
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1291_
timestamp 1698431365
transform -1 0 14224 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1292_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13552 0 1 94080
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1293_
timestamp 1698431365
transform 1 0 13440 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1294_
timestamp 1698431365
transform -1 0 12320 0 1 92512
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1295_
timestamp 1698431365
transform 1 0 10976 0 -1 95648
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1296_
timestamp 1698431365
transform 1 0 19936 0 1 86240
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1297_
timestamp 1698431365
transform 1 0 19600 0 -1 84672
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1298_
timestamp 1698431365
transform 1 0 20608 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1299_
timestamp 1698431365
transform -1 0 20608 0 -1 90944
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1300_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19936 0 -1 97216
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1301_
timestamp 1698431365
transform 1 0 15232 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1302_
timestamp 1698431365
transform -1 0 14448 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1303_
timestamp 1698431365
transform -1 0 14224 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1304_
timestamp 1698431365
transform -1 0 13104 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1305_
timestamp 1698431365
transform -1 0 11200 0 -1 97216
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1306_
timestamp 1698431365
transform -1 0 13552 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1307_
timestamp 1698431365
transform -1 0 13104 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1308_
timestamp 1698431365
transform 1 0 15568 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1309_
timestamp 1698431365
transform 1 0 14336 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1310_
timestamp 1698431365
transform 1 0 11872 0 1 95648
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1311_
timestamp 1698431365
transform -1 0 10976 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1312_
timestamp 1698431365
transform -1 0 8288 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1313_
timestamp 1698431365
transform 1 0 25200 0 -1 117600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1314_
timestamp 1698431365
transform -1 0 18704 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1315_
timestamp 1698431365
transform 1 0 16688 0 1 79968
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1316_
timestamp 1698431365
transform 1 0 19488 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1317_
timestamp 1698431365
transform -1 0 19376 0 -1 89376
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1318_
timestamp 1698431365
transform 1 0 18704 0 1 97216
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1319_
timestamp 1698431365
transform -1 0 19040 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1320_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14224 0 1 92512
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1321_
timestamp 1698431365
transform -1 0 18368 0 -1 97216
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1322_
timestamp 1698431365
transform -1 0 15456 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1323_
timestamp 1698431365
transform -1 0 9184 0 -1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1324_
timestamp 1698431365
transform -1 0 9184 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1325_
timestamp 1698431365
transform 1 0 11984 0 1 101920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1326_
timestamp 1698431365
transform 1 0 9520 0 1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1327_
timestamp 1698431365
transform 1 0 23184 0 -1 103488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform 1 0 19488 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1329_
timestamp 1698431365
transform 1 0 18368 0 -1 79968
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1330_
timestamp 1698431365
transform 1 0 21168 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1331_
timestamp 1698431365
transform 1 0 21168 0 1 92512
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1332_
timestamp 1698431365
transform 1 0 19936 0 -1 98784
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1333_
timestamp 1698431365
transform -1 0 19264 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1334_
timestamp 1698431365
transform -1 0 18480 0 -1 98784
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1335_
timestamp 1698431365
transform -1 0 15456 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1336_
timestamp 1698431365
transform -1 0 9968 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1337_
timestamp 1698431365
transform -1 0 20496 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1338_
timestamp 1698431365
transform -1 0 13104 0 1 103488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1339_
timestamp 1698431365
transform -1 0 22960 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1340_
timestamp 1698431365
transform 1 0 21840 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1341_
timestamp 1698431365
transform -1 0 24528 0 -1 103488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_
timestamp 1698431365
transform -1 0 19600 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1343_
timestamp 1698431365
transform -1 0 20720 0 1 79968
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1344_
timestamp 1698431365
transform 1 0 20160 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1345_
timestamp 1698431365
transform -1 0 20608 0 1 92512
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1346_
timestamp 1698431365
transform 1 0 19264 0 1 95648
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1347_
timestamp 1698431365
transform 1 0 16128 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1348_
timestamp 1698431365
transform -1 0 18144 0 1 97216
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1349_
timestamp 1698431365
transform -1 0 15344 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1350_
timestamp 1698431365
transform 1 0 18480 0 -1 98784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1351_
timestamp 1698431365
transform 1 0 17248 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1352_
timestamp 1698431365
transform 1 0 16128 0 -1 106624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1353_
timestamp 1698431365
transform 1 0 20608 0 -1 108192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1354_
timestamp 1698431365
transform 1 0 20272 0 1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1355_
timestamp 1698431365
transform -1 0 20272 0 1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1356_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19936 0 1 86240
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1357_
timestamp 1698431365
transform -1 0 16912 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1358_
timestamp 1698431365
transform 1 0 17360 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1359_
timestamp 1698431365
transform 1 0 16912 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1360_
timestamp 1698431365
transform 1 0 14784 0 1 94080
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1361_
timestamp 1698431365
transform 1 0 15008 0 -1 94080
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1362_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15568 0 -1 94080
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1363_
timestamp 1698431365
transform -1 0 14224 0 1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1364_
timestamp 1698431365
transform -1 0 9184 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1365_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 -1 103488
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1366_
timestamp 1698431365
transform 1 0 17472 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1367_
timestamp 1698431365
transform 1 0 17248 0 1 84672
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1368_
timestamp 1698431365
transform 1 0 18368 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1369_
timestamp 1698431365
transform -1 0 18144 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1370_
timestamp 1698431365
transform 1 0 18928 0 1 98784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1371_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 1 97216
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1372_
timestamp 1698431365
transform -1 0 11536 0 1 103488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1373_
timestamp 1698431365
transform -1 0 13104 0 1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1374_
timestamp 1698431365
transform -1 0 16240 0 -1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1375_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17920 0 1 89376
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1376_
timestamp 1698431365
transform 1 0 14112 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1377_
timestamp 1698431365
transform 1 0 13328 0 1 101920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1378_
timestamp 1698431365
transform -1 0 14560 0 1 103488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1379_
timestamp 1698431365
transform 1 0 11984 0 -1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1380_
timestamp 1698431365
transform 1 0 14560 0 1 103488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1381_
timestamp 1698431365
transform -1 0 8288 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  _1382_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1383_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25760 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1384_
timestamp 1698431365
transform 1 0 15008 0 1 3136
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1385_
timestamp 1698431365
transform -1 0 19712 0 -1 3136
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1386_
timestamp 1698431365
transform 1 0 18144 0 1 1568
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1387_
timestamp 1698431365
transform 1 0 23296 0 -1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1388_
timestamp 1698431365
transform -1 0 24192 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1389_
timestamp 1698431365
transform 1 0 10192 0 -1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1390_
timestamp 1698431365
transform 1 0 12320 0 -1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1391_
timestamp 1698431365
transform 1 0 11312 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1392_
timestamp 1698431365
transform 1 0 5488 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1393_
timestamp 1698431365
transform -1 0 7168 0 -1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1394_
timestamp 1698431365
transform 1 0 7504 0 1 3136
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1395_
timestamp 1698431365
transform -1 0 13104 0 1 3136
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1396_
timestamp 1698431365
transform 1 0 25088 0 -1 3136
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1397_
timestamp 1698431365
transform 1 0 17248 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1398_
timestamp 1698431365
transform -1 0 21728 0 1 1568
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1399_
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1400_
timestamp 1698431365
transform 1 0 21616 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1401_
timestamp 1698431365
transform 1 0 21952 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1402_
timestamp 1698431365
transform 1 0 23296 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1403_
timestamp 1698431365
transform -1 0 27328 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1404_
timestamp 1698431365
transform -1 0 28336 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1405_
timestamp 1698431365
transform 1 0 2688 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1406_
timestamp 1698431365
transform 1 0 21504 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1407_
timestamp 1698431365
transform 1 0 21952 0 -1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1408_
timestamp 1698431365
transform 1 0 19376 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1409_
timestamp 1698431365
transform 1 0 18704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  _1410_
timestamp 1698431365
transform 1 0 3248 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1411_
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1412_
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1413_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4144 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1414_
timestamp 1698431365
transform 1 0 21504 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1415_
timestamp 1698431365
transform 1 0 21056 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  _1416_
timestamp 1698431365
transform 1 0 7952 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1417_
timestamp 1698431365
transform 1 0 16688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1418_
timestamp 1698431365
transform 1 0 15792 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1419_
timestamp 1698431365
transform 1 0 3472 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1420_
timestamp 1698431365
transform 1 0 12208 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1421_
timestamp 1698431365
transform 1 0 11648 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1422_
timestamp 1698431365
transform 1 0 4032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1423_
timestamp 1698431365
transform 1 0 21952 0 -1 68992
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1424_
timestamp 1698431365
transform 1 0 25424 0 1 72128
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1425_
timestamp 1698431365
transform 1 0 11088 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1426_
timestamp 1698431365
transform 1 0 9968 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1427_
timestamp 1698431365
transform 1 0 3808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1428_
timestamp 1698431365
transform 1 0 24416 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1429_
timestamp 1698431365
transform 1 0 23296 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1430_
timestamp 1698431365
transform 1 0 4368 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1431_
timestamp 1698431365
transform 1 0 11312 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1432_
timestamp 1698431365
transform 1 0 10304 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1433_
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1434_
timestamp 1698431365
transform -1 0 28336 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1435_
timestamp 1698431365
transform 1 0 23296 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1436_
timestamp 1698431365
transform 1 0 22400 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1437_
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1438_
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1439_
timestamp 1698431365
transform 1 0 8176 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1440_
timestamp 1698431365
transform 1 0 4592 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1441_
timestamp 1698431365
transform 1 0 9520 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1442_
timestamp 1698431365
transform 1 0 8736 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1443_
timestamp 1698431365
transform -1 0 3248 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1444_
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1445_
timestamp 1698431365
transform 1 0 8176 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1446_
timestamp 1698431365
transform 1 0 6608 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1447_
timestamp 1698431365
transform -1 0 9184 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1448_
timestamp 1698431365
transform 1 0 8288 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1449_
timestamp 1698431365
transform 1 0 3472 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1450_
timestamp 1698431365
transform 1 0 19040 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1451_
timestamp 1698431365
transform 1 0 15456 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1452_
timestamp 1698431365
transform 1 0 3920 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1453_
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1454_
timestamp 1698431365
transform 1 0 11872 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1455_
timestamp 1698431365
transform 1 0 3584 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1456_
timestamp 1698431365
transform 1 0 11984 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1457_
timestamp 1698431365
transform 1 0 10976 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1458_
timestamp 1698431365
transform 1 0 5600 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1459_
timestamp 1698431365
transform 1 0 19264 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1460_
timestamp 1698431365
transform 1 0 18144 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1461_
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1462_
timestamp 1698431365
transform 1 0 14000 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1463_
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1464_
timestamp 1698431365
transform 1 0 2352 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1465_
timestamp 1698431365
transform 1 0 18816 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1466_
timestamp 1698431365
transform 1 0 17808 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1467_
timestamp 1698431365
transform 1 0 2352 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1468_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1469_
timestamp 1698431365
transform 1 0 14784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1470_
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1471_
timestamp 1698431365
transform 1 0 21728 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1472_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1473_
timestamp 1698431365
transform 1 0 3024 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1474_
timestamp 1698431365
transform 1 0 20160 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1475_
timestamp 1698431365
transform 1 0 19824 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1476_
timestamp 1698431365
transform 1 0 3808 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1477_
timestamp 1698431365
transform 1 0 26656 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1478_
timestamp 1698431365
transform 1 0 25760 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1479_
timestamp 1698431365
transform 1 0 2912 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1480_
timestamp 1698431365
transform 1 0 26432 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1481_
timestamp 1698431365
transform 1 0 25760 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1482_
timestamp 1698431365
transform 1 0 2576 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1483_
timestamp 1698431365
transform 1 0 26544 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1484_
timestamp 1698431365
transform 1 0 25984 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1485_
timestamp 1698431365
transform 1 0 3024 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1486_
timestamp 1698431365
transform 1 0 25424 0 1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1487_
timestamp 1698431365
transform 1 0 22064 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1488_
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1489_
timestamp 1698431365
transform 1 0 3472 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1490_
timestamp 1698431365
transform 1 0 26992 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1491_
timestamp 1698431365
transform 1 0 26096 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1492_
timestamp 1698431365
transform 1 0 3360 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1493_
timestamp 1698431365
transform 1 0 23632 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1494_
timestamp 1698431365
transform 1 0 22736 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1495_
timestamp 1698431365
transform 1 0 17920 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1496_
timestamp 1698431365
transform 1 0 26992 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1497_
timestamp 1698431365
transform 1 0 25088 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1498_
timestamp 1698431365
transform 1 0 2912 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1499_
timestamp 1698431365
transform 1 0 26544 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1500_
timestamp 1698431365
transform 1 0 25648 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1501_
timestamp 1698431365
transform 1 0 21952 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1502_
timestamp 1698431365
transform 1 0 26096 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1503_
timestamp 1698431365
transform 1 0 25424 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1504_
timestamp 1698431365
transform 1 0 20048 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1505_
timestamp 1698431365
transform -1 0 24416 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1506_
timestamp 1698431365
transform 1 0 22624 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1507_
timestamp 1698431365
transform 1 0 23744 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1508_
timestamp 1698431365
transform 1 0 22848 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1509_
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1510_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1511_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1512_
timestamp 1698431365
transform 1 0 8288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1513_
timestamp 1698431365
transform 1 0 7392 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1514_
timestamp 1698431365
transform 1 0 6272 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1515_
timestamp 1698431365
transform 1 0 7504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1516_
timestamp 1698431365
transform 1 0 6272 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1517_
timestamp 1698431365
transform 1 0 9520 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1518_
timestamp 1698431365
transform -1 0 10304 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1519_
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1520_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1521_
timestamp 1698431365
transform 1 0 7616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1522_
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1523_
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1524_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1525_
timestamp 1698431365
transform 1 0 21840 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1526_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1527_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1528_
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1529_
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1530_
timestamp 1698431365
transform 1 0 18592 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1531_
timestamp 1698431365
transform 1 0 17920 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1532_
timestamp 1698431365
transform 1 0 13216 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1533_
timestamp 1698431365
transform -1 0 14224 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1534_
timestamp 1698431365
transform 1 0 12208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1535_
timestamp 1698431365
transform 1 0 10416 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1536_
timestamp 1698431365
transform 1 0 9856 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1537_
timestamp 1698431365
transform 1 0 7616 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1538_
timestamp 1698431365
transform -1 0 26768 0 1 67424
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1539_
timestamp 1698431365
transform 1 0 7280 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1540_
timestamp 1698431365
transform 1 0 5936 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1541_
timestamp 1698431365
transform 1 0 7168 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1542_
timestamp 1698431365
transform 1 0 5824 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1543_
timestamp 1698431365
transform 1 0 7728 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1544_
timestamp 1698431365
transform 1 0 5712 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1545_
timestamp 1698431365
transform 1 0 12096 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1546_
timestamp 1698431365
transform 1 0 11088 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1547_
timestamp 1698431365
transform 1 0 6272 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1548_
timestamp 1698431365
transform 1 0 5712 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1549_
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1550_
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1551_
timestamp 1698431365
transform -1 0 12992 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1552_
timestamp 1698431365
transform -1 0 14224 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1553_
timestamp 1698431365
transform 1 0 8064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1554_
timestamp 1698431365
transform 1 0 7056 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1555_
timestamp 1698431365
transform 1 0 7616 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1556_
timestamp 1698431365
transform 1 0 6608 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1557_
timestamp 1698431365
transform 1 0 23296 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1558_
timestamp 1698431365
transform 1 0 22848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1559_
timestamp 1698431365
transform 1 0 23968 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1560_
timestamp 1698431365
transform 1 0 23632 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1561_
timestamp 1698431365
transform 1 0 23856 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1562_
timestamp 1698431365
transform 1 0 23520 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1563_
timestamp 1698431365
transform -1 0 18144 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1564_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1565_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1566_
timestamp 1698431365
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1567_
timestamp 1698431365
transform -1 0 26768 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1568_
timestamp 1698431365
transform 1 0 24976 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1569_
timestamp 1698431365
transform 1 0 23968 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1570_
timestamp 1698431365
transform -1 0 24976 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1571_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1572_
timestamp 1698431365
transform 1 0 23856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1573_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1574_
timestamp 1698431365
transform 1 0 23856 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1575_
timestamp 1698431365
transform -1 0 23520 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1576_
timestamp 1698431365
transform 1 0 21952 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1577_
timestamp 1698431365
transform 1 0 4704 0 1 100352
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1578_
timestamp 1698431365
transform -1 0 6608 0 1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1579_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5936 0 -1 87808
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1580_
timestamp 1698431365
transform -1 0 4928 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1581_
timestamp 1698431365
transform -1 0 4032 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1582_
timestamp 1698431365
transform -1 0 6384 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1583_
timestamp 1698431365
transform 1 0 6608 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1584_
timestamp 1698431365
transform 1 0 6720 0 -1 95648
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1585_
timestamp 1698431365
transform -1 0 6496 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1586_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6944 0 1 90944
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1587_
timestamp 1698431365
transform -1 0 3584 0 -1 92512
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1588_
timestamp 1698431365
transform -1 0 7504 0 1 90944
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1589_
timestamp 1698431365
transform 1 0 5936 0 -1 90944
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1590_
timestamp 1698431365
transform 1 0 7280 0 -1 90944
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1591_
timestamp 1698431365
transform 1 0 7840 0 -1 95648
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1592_
timestamp 1698431365
transform 1 0 9408 0 -1 95648
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1593_
timestamp 1698431365
transform 1 0 19040 0 1 100352
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1594_
timestamp 1698431365
transform -1 0 20384 0 1 98784
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1595_
timestamp 1698431365
transform 1 0 23296 0 -1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1596_
timestamp 1698431365
transform -1 0 23744 0 -1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1698431365
transform 1 0 24192 0 -1 101920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1598_
timestamp 1698431365
transform 1 0 25088 0 -1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1599_
timestamp 1698431365
transform -1 0 26544 0 1 97216
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1600_
timestamp 1698431365
transform -1 0 24192 0 -1 98784
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1601_
timestamp 1698431365
transform -1 0 24752 0 -1 98784
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1602_
timestamp 1698431365
transform 1 0 23744 0 1 97216
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1603_
timestamp 1698431365
transform 1 0 26544 0 1 97216
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1604_
timestamp 1698431365
transform 1 0 23072 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1605_
timestamp 1698431365
transform 1 0 25088 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1606_
timestamp 1698431365
transform -1 0 24752 0 -1 95648
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1607_
timestamp 1698431365
transform 1 0 25200 0 -1 95648
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1608_
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1609_
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1610_
timestamp 1698431365
transform -1 0 22736 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1611_
timestamp 1698431365
transform -1 0 26208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1612_
timestamp 1698431365
transform 1 0 11200 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1613_
timestamp 1698431365
transform -1 0 23968 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1614_
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1615_
timestamp 1698431365
transform -1 0 26208 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1616_
timestamp 1698431365
transform 1 0 22176 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1617_
timestamp 1698431365
transform -1 0 23072 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1618_
timestamp 1698431365
transform -1 0 24416 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1619_
timestamp 1698431365
transform 1 0 25424 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1620_
timestamp 1698431365
transform 1 0 20272 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1621_
timestamp 1698431365
transform 1 0 2352 0 1 84672
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1622_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19488 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1623_
timestamp 1698431365
transform 1 0 14112 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1624_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1625_
timestamp 1698431365
transform -1 0 24640 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1626_
timestamp 1698431365
transform 1 0 22288 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1627_
timestamp 1698431365
transform -1 0 19040 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1628_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1629_
timestamp 1698431365
transform -1 0 20608 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1630_
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1631_
timestamp 1698431365
transform 1 0 18032 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1632_
timestamp 1698431365
transform 1 0 15904 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1633_
timestamp 1698431365
transform -1 0 23184 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1634_
timestamp 1698431365
transform 1 0 22064 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1635_
timestamp 1698431365
transform 1 0 14672 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1636_
timestamp 1698431365
transform 1 0 13552 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1637_
timestamp 1698431365
transform 1 0 25424 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1638_
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1639_
timestamp 1698431365
transform -1 0 7952 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1640_
timestamp 1698431365
transform 1 0 10080 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1641_
timestamp 1698431365
transform 1 0 9296 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1642_
timestamp 1698431365
transform -1 0 8848 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1643_
timestamp 1698431365
transform -1 0 7504 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1644_
timestamp 1698431365
transform -1 0 12208 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1645_
timestamp 1698431365
transform 1 0 10416 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1646_
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1647_
timestamp 1698431365
transform 1 0 22400 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1648_
timestamp 1698431365
transform 1 0 7952 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1649_
timestamp 1698431365
transform -1 0 15456 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1650_
timestamp 1698431365
transform 1 0 13888 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1651_
timestamp 1698431365
transform -1 0 12992 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1652_
timestamp 1698431365
transform 1 0 11200 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1653_
timestamp 1698431365
transform 1 0 12096 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1654_
timestamp 1698431365
transform 1 0 10976 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1655_
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1656_
timestamp 1698431365
transform 1 0 8064 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1657_
timestamp 1698431365
transform -1 0 10192 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1658_
timestamp 1698431365
transform 1 0 7616 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1659_
timestamp 1698431365
transform 1 0 18368 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1660_
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1661_
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1662_
timestamp 1698431365
transform -1 0 15120 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1663_
timestamp 1698431365
transform -1 0 22736 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1664_
timestamp 1698431365
transform 1 0 20944 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1665_
timestamp 1698431365
transform 1 0 16352 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1666_
timestamp 1698431365
transform 1 0 15568 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1667_
timestamp 1698431365
transform -1 0 26880 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1668_
timestamp 1698431365
transform 1 0 25760 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1669_
timestamp 1698431365
transform -1 0 27888 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1670_
timestamp 1698431365
transform 1 0 26096 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1671_
timestamp 1698431365
transform 1 0 25424 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1672_
timestamp 1698431365
transform -1 0 27104 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1673_
timestamp 1698431365
transform 1 0 14672 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1674_
timestamp 1698431365
transform 1 0 13888 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1675_
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1676_
timestamp 1698431365
transform -1 0 26992 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1677_
timestamp 1698431365
transform -1 0 27664 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1678_
timestamp 1698431365
transform 1 0 25648 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1679_
timestamp 1698431365
transform -1 0 27552 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1680_
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1681_
timestamp 1698431365
transform 1 0 26432 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1682_
timestamp 1698431365
transform -1 0 27552 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1683_
timestamp 1698431365
transform -1 0 27552 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1684_
timestamp 1698431365
transform 1 0 25760 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1685_
timestamp 1698431365
transform 1 0 22064 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1686_
timestamp 1698431365
transform 1 0 21280 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1687_
timestamp 1698431365
transform -1 0 8400 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1688_
timestamp 1698431365
transform -1 0 23744 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1689_
timestamp 1698431365
transform -1 0 20272 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1690_
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1691_
timestamp 1698431365
transform 1 0 2352 0 -1 81536
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1692_
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1693_
timestamp 1698431365
transform 1 0 3024 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1694_
timestamp 1698431365
transform 1 0 6160 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1695_
timestamp 1698431365
transform -1 0 5264 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1696_
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1697_
timestamp 1698431365
transform -1 0 3248 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1698_
timestamp 1698431365
transform 1 0 4592 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1699_
timestamp 1698431365
transform 1 0 4144 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1700_
timestamp 1698431365
transform -1 0 5712 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1701_
timestamp 1698431365
transform -1 0 7952 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1702_
timestamp 1698431365
transform 1 0 6160 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1703_
timestamp 1698431365
transform 1 0 5936 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform -1 0 3584 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1705_
timestamp 1698431365
transform 1 0 2352 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1706_
timestamp 1698431365
transform -1 0 3248 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1707_
timestamp 1698431365
transform -1 0 3696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1708_
timestamp 1698431365
transform 1 0 2576 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1709_
timestamp 1698431365
transform -1 0 3472 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1710_
timestamp 1698431365
transform -1 0 3696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1711_
timestamp 1698431365
transform -1 0 3248 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1712_
timestamp 1698431365
transform -1 0 3472 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1713_
timestamp 1698431365
transform -1 0 4032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1714_
timestamp 1698431365
transform -1 0 3584 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1715_
timestamp 1698431365
transform -1 0 3696 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1716_
timestamp 1698431365
transform -1 0 3808 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1717_
timestamp 1698431365
transform -1 0 3584 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1718_
timestamp 1698431365
transform 1 0 2352 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1719_
timestamp 1698431365
transform -1 0 3360 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1720_
timestamp 1698431365
transform -1 0 6608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1721_
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1722_
timestamp 1698431365
transform -1 0 6608 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1723_
timestamp 1698431365
transform -1 0 3584 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1724_
timestamp 1698431365
transform 1 0 2352 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1725_
timestamp 1698431365
transform -1 0 3248 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1726_
timestamp 1698431365
transform -1 0 3696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1727_
timestamp 1698431365
transform -1 0 3920 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1728_
timestamp 1698431365
transform -1 0 3248 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1729_
timestamp 1698431365
transform -1 0 6160 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1730_
timestamp 1698431365
transform 1 0 4592 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1731_
timestamp 1698431365
transform -1 0 6608 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1732_
timestamp 1698431365
transform -1 0 4704 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1733_
timestamp 1698431365
transform -1 0 3248 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1734_
timestamp 1698431365
transform -1 0 3472 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1735_
timestamp 1698431365
transform -1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1736_
timestamp 1698431365
transform -1 0 4032 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1737_
timestamp 1698431365
transform -1 0 3360 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1738_
timestamp 1698431365
transform -1 0 3696 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1739_
timestamp 1698431365
transform 1 0 2352 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1740_
timestamp 1698431365
transform -1 0 3360 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1741_
timestamp 1698431365
transform -1 0 6720 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1742_
timestamp 1698431365
transform 1 0 4704 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1743_
timestamp 1698431365
transform -1 0 6160 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1744_
timestamp 1698431365
transform -1 0 6496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1745_
timestamp 1698431365
transform 1 0 4816 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1746_
timestamp 1698431365
transform -1 0 6608 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1747_
timestamp 1698431365
transform -1 0 3472 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1748_
timestamp 1698431365
transform -1 0 2912 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1749_
timestamp 1698431365
transform -1 0 3136 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1750_
timestamp 1698431365
transform -1 0 3696 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1751_
timestamp 1698431365
transform -1 0 2912 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1752_
timestamp 1698431365
transform -1 0 3248 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1753_
timestamp 1698431365
transform -1 0 3808 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1754_
timestamp 1698431365
transform -1 0 4256 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1755_
timestamp 1698431365
transform 1 0 2912 0 1 79968
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1756_
timestamp 1698431365
transform -1 0 3584 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1757_
timestamp 1698431365
transform -1 0 3472 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1758_
timestamp 1698431365
transform -1 0 3920 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1759_
timestamp 1698431365
transform -1 0 3248 0 -1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1760_
timestamp 1698431365
transform -1 0 3808 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1761_
timestamp 1698431365
transform -1 0 3248 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1762_
timestamp 1698431365
transform -1 0 3472 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1763_
timestamp 1698431365
transform -1 0 3696 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1764_
timestamp 1698431365
transform 1 0 2240 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1765_
timestamp 1698431365
transform -1 0 3248 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1766_
timestamp 1698431365
transform -1 0 3696 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1767_
timestamp 1698431365
transform 1 0 1904 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1768_
timestamp 1698431365
transform -1 0 3248 0 -1 68992
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1769_
timestamp 1698431365
transform -1 0 3696 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1770_
timestamp 1698431365
transform 1 0 2240 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1771_
timestamp 1698431365
transform 1 0 2128 0 -1 72128
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1772_
timestamp 1698431365
transform -1 0 5264 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1773_
timestamp 1698431365
transform 1 0 2464 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1774_
timestamp 1698431365
transform -1 0 3360 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1775_
timestamp 1698431365
transform -1 0 3808 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1776_
timestamp 1698431365
transform 1 0 2352 0 1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1777_
timestamp 1698431365
transform -1 0 3360 0 -1 78400
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1778_
timestamp 1698431365
transform 1 0 5600 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1779_
timestamp 1698431365
transform -1 0 6608 0 1 78400
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1780_
timestamp 1698431365
transform -1 0 3920 0 -1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1781_
timestamp 1698431365
transform 1 0 2128 0 -1 83104
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1782_
timestamp 1698431365
transform -1 0 7840 0 -1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1783_
timestamp 1698431365
transform 1 0 6832 0 -1 81536
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1784_
timestamp 1698431365
transform 1 0 5488 0 1 81536
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1785_
timestamp 1698431365
transform -1 0 6608 0 1 83104
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1786_
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1787_
timestamp 1698431365
transform -1 0 25312 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1788_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1789_
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1790_
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1791_
timestamp 1698431365
transform 1 0 22176 0 1 68992
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1792_
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1793_
timestamp 1698431365
transform 1 0 11760 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1794_
timestamp 1698431365
transform 1 0 21056 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1795_
timestamp 1698431365
transform 1 0 19600 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1796_
timestamp 1698431365
transform 1 0 17808 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1797_
timestamp 1698431365
transform 1 0 16688 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1798_
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1799_
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1800_
timestamp 1698431365
transform 1 0 14336 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1801_
timestamp 1698431365
transform 1 0 13440 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1802_
timestamp 1698431365
transform 1 0 13664 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1803_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1804_
timestamp 1698431365
transform 1 0 15008 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1805_
timestamp 1698431365
transform 1 0 14112 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1806_
timestamp 1698431365
transform 1 0 24528 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1807_
timestamp 1698431365
transform 1 0 22064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1808_
timestamp 1698431365
transform -1 0 22736 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1809_
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1810_
timestamp 1698431365
transform 1 0 17248 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1811_
timestamp 1698431365
transform 1 0 13440 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1812_
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1813_
timestamp 1698431365
transform 1 0 11536 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1814_
timestamp 1698431365
transform 1 0 10416 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1815_
timestamp 1698431365
transform 1 0 11424 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1816_
timestamp 1698431365
transform 1 0 9968 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1817_
timestamp 1698431365
transform 1 0 15456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1818_
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1819_
timestamp 1698431365
transform 1 0 11312 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1820_
timestamp 1698431365
transform 1 0 10192 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1821_
timestamp 1698431365
transform 1 0 11200 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1822_
timestamp 1698431365
transform 1 0 10080 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1823_
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1824_
timestamp 1698431365
transform -1 0 18144 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1825_
timestamp 1698431365
transform 1 0 14336 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1826_
timestamp 1698431365
transform 1 0 13328 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1827_
timestamp 1698431365
transform 1 0 11088 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1828_
timestamp 1698431365
transform 1 0 9968 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1829_
timestamp 1698431365
transform 1 0 11536 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1830_
timestamp 1698431365
transform 1 0 10416 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1831_
timestamp 1698431365
transform 1 0 19152 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1832_
timestamp 1698431365
transform 1 0 18256 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1833_
timestamp 1698431365
transform 1 0 14784 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1834_
timestamp 1698431365
transform 1 0 13888 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1835_
timestamp 1698431365
transform 1 0 26768 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1836_
timestamp 1698431365
transform 1 0 25872 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1837_
timestamp 1698431365
transform 1 0 26320 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1838_
timestamp 1698431365
transform 1 0 25872 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1839_
timestamp 1698431365
transform 1 0 26880 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1840_
timestamp 1698431365
transform 1 0 25648 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1841_
timestamp 1698431365
transform 1 0 16016 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1842_
timestamp 1698431365
transform 1 0 15120 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1843_
timestamp 1698431365
transform 1 0 26208 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1844_
timestamp 1698431365
transform 1 0 25872 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1845_
timestamp 1698431365
transform 1 0 26768 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1846_
timestamp 1698431365
transform 1 0 24192 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1847_
timestamp 1698431365
transform -1 0 24864 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1848_
timestamp 1698431365
transform -1 0 28000 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1849_
timestamp 1698431365
transform 1 0 26768 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1850_
timestamp 1698431365
transform 1 0 26208 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1851_
timestamp 1698431365
transform -1 0 25984 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1852_
timestamp 1698431365
transform -1 0 26880 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1853_
timestamp 1698431365
transform -1 0 23968 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 22176 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1855_
timestamp 1698431365
transform -1 0 20832 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1856_
timestamp 1698431365
transform -1 0 20384 0 1 1568
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1857_
timestamp 1698431365
transform -1 0 20944 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1858_
timestamp 1698431365
transform -1 0 20944 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1859_
timestamp 1698431365
transform -1 0 3024 0 1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1860_
timestamp 1698431365
transform -1 0 21616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1861_
timestamp 1698431365
transform 1 0 19712 0 -1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1862_
timestamp 1698431365
transform -1 0 22288 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1863_
timestamp 1698431365
transform 1 0 19152 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1864_
timestamp 1698431365
transform -1 0 16912 0 -1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1865_
timestamp 1698431365
transform 1 0 15456 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1866_
timestamp 1698431365
transform 1 0 20272 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1867_
timestamp 1698431365
transform -1 0 24080 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1868_
timestamp 1698431365
transform 1 0 21168 0 -1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1869_
timestamp 1698431365
transform 1 0 20272 0 1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1870_
timestamp 1698431365
transform 1 0 19488 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform 1 0 10864 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1872_
timestamp 1698431365
transform 1 0 8064 0 -1 78400
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1873_
timestamp 1698431365
transform 1 0 22400 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1874_
timestamp 1698431365
transform 1 0 21840 0 1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1875_
timestamp 1698431365
transform -1 0 19040 0 -1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1876_
timestamp 1698431365
transform 1 0 17248 0 -1 78400
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1877_
timestamp 1698431365
transform 1 0 18480 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1878_
timestamp 1698431365
transform 1 0 17584 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1879_
timestamp 1698431365
transform -1 0 17024 0 -1 81536
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1880_
timestamp 1698431365
transform 1 0 13552 0 1 78400
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1881_
timestamp 1698431365
transform -1 0 24864 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1882_
timestamp 1698431365
transform 1 0 21728 0 1 72128
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1883_
timestamp 1698431365
transform 1 0 22064 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1884_
timestamp 1698431365
transform 1 0 20944 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1885_
timestamp 1698431365
transform -1 0 24080 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1886_
timestamp 1698431365
transform 1 0 21392 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1887_
timestamp 1698431365
transform 1 0 3472 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1888_
timestamp 1698431365
transform -1 0 22288 0 1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1889_
timestamp 1698431365
transform 1 0 21504 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1890_
timestamp 1698431365
transform 1 0 19824 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1891_
timestamp 1698431365
transform 1 0 12432 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1892_
timestamp 1698431365
transform 1 0 11200 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1893_
timestamp 1698431365
transform 1 0 3696 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1894_
timestamp 1698431365
transform 1 0 2688 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1895_
timestamp 1698431365
transform 1 0 8176 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1896_
timestamp 1698431365
transform 1 0 7056 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1897_
timestamp 1698431365
transform 1 0 4592 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1898_
timestamp 1698431365
transform -1 0 6608 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1899_
timestamp 1698431365
transform 1 0 7952 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1900_
timestamp 1698431365
transform 1 0 6832 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1901_
timestamp 1698431365
transform 1 0 6608 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1902_
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1903_
timestamp 1698431365
transform 1 0 7392 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1904_
timestamp 1698431365
transform 1 0 6384 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1905_
timestamp 1698431365
transform 1 0 6160 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1906_
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1907_
timestamp 1698431365
transform 1 0 3696 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1908_
timestamp 1698431365
transform 1 0 2688 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1909_
timestamp 1698431365
transform 1 0 3808 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1910_
timestamp 1698431365
transform 1 0 2800 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1911_
timestamp 1698431365
transform 1 0 6832 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1912_
timestamp 1698431365
transform 1 0 5936 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1913_
timestamp 1698431365
transform -1 0 20384 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1914_
timestamp 1698431365
transform -1 0 20944 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1915_
timestamp 1698431365
transform 1 0 6608 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1916_
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1917_
timestamp 1698431365
transform -1 0 19376 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1918_
timestamp 1698431365
transform 1 0 18256 0 1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1919_
timestamp 1698431365
transform 1 0 6608 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1920_
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1921_
timestamp 1698431365
transform 1 0 6720 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1922_
timestamp 1698431365
transform 1 0 5600 0 1 72128
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1923_
timestamp 1698431365
transform 1 0 6608 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1924_
timestamp 1698431365
transform 1 0 5488 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1925_
timestamp 1698431365
transform 1 0 7504 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1926_
timestamp 1698431365
transform 1 0 6384 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1927_
timestamp 1698431365
transform -1 0 20832 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1928_
timestamp 1698431365
transform 1 0 19040 0 -1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1929_
timestamp 1698431365
transform -1 0 20608 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1930_
timestamp 1698431365
transform 1 0 18816 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1931_
timestamp 1698431365
transform -1 0 25760 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1932_
timestamp 1698431365
transform 1 0 23184 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1933_
timestamp 1698431365
transform -1 0 24640 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1934_
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1935_
timestamp 1698431365
transform -1 0 24864 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1936_
timestamp 1698431365
transform -1 0 26768 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1937_
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1938_
timestamp 1698431365
transform -1 0 22176 0 -1 94080
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1939_
timestamp 1698431365
transform -1 0 4144 0 1 94080
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1940_
timestamp 1698431365
transform -1 0 3360 0 -1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1698431365
transform 1 0 2016 0 -1 97216
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1942_
timestamp 1698431365
transform 1 0 10976 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1943_
timestamp 1698431365
transform -1 0 3472 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1944_
timestamp 1698431365
transform -1 0 3584 0 -1 98784
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1945_
timestamp 1698431365
transform -1 0 11088 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1946_
timestamp 1698431365
transform -1 0 3696 0 -1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1947_
timestamp 1698431365
transform 1 0 3248 0 1 101920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1948_
timestamp 1698431365
transform 1 0 21168 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1949_
timestamp 1698431365
transform -1 0 4032 0 1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1950_
timestamp 1698431365
transform -1 0 4592 0 -1 103488
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1951_
timestamp 1698431365
transform 1 0 17136 0 1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1952_
timestamp 1698431365
transform -1 0 4032 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1953_
timestamp 1698431365
transform -1 0 8512 0 -1 105056
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1954_
timestamp 1698431365
transform -1 0 7392 0 -1 103488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1955_
timestamp 1698431365
transform -1 0 4480 0 -1 105056
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1956_
timestamp 1698431365
transform -1 0 3584 0 -1 106624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1957_
timestamp 1698431365
transform -1 0 7280 0 -1 105056
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1958_
timestamp 1698431365
transform -1 0 6608 0 -1 106624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform -1 0 15120 0 1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1960_
timestamp 1698431365
transform 1 0 13664 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1961_
timestamp 1698431365
transform -1 0 13104 0 1 84672
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1962_
timestamp 1698431365
transform 1 0 11872 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1963_
timestamp 1698431365
transform -1 0 13104 0 1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1964_
timestamp 1698431365
transform 1 0 10976 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1965_
timestamp 1698431365
transform 1 0 5936 0 1 98784
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1966_
timestamp 1698431365
transform -1 0 5712 0 -1 98784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1967_
timestamp 1698431365
transform 1 0 7616 0 1 92512
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1968_
timestamp 1698431365
transform 1 0 9408 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1969_
timestamp 1698431365
transform 1 0 7952 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1970_
timestamp 1698431365
transform 1 0 11312 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1971_
timestamp 1698431365
transform 1 0 10416 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1972_
timestamp 1698431365
transform 1 0 8848 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1973_
timestamp 1698431365
transform 1 0 7840 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1974_
timestamp 1698431365
transform 1 0 9520 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1975_
timestamp 1698431365
transform 1 0 8288 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1976_
timestamp 1698431365
transform 1 0 10640 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1977_
timestamp 1698431365
transform 1 0 8512 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1978_
timestamp 1698431365
transform 1 0 9968 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1979_
timestamp 1698431365
transform 1 0 8288 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1980_
timestamp 1698431365
transform 1 0 9408 0 -1 98784
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1981_
timestamp 1698431365
transform -1 0 7504 0 1 98784
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1982_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1983_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1984_
timestamp 1698431365
transform -1 0 24416 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1985_
timestamp 1698431365
transform 1 0 14896 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1986_
timestamp 1698431365
transform 1 0 9856 0 1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1987_
timestamp 1698431365
transform 1 0 8848 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1988_
timestamp 1698431365
transform 1 0 22624 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1989_
timestamp 1698431365
transform 1 0 9184 0 1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1990_
timestamp 1698431365
transform -1 0 24752 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1991_
timestamp 1698431365
transform 1 0 6608 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1992_
timestamp 1698431365
transform 1 0 7280 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1993_
timestamp 1698431365
transform 1 0 6496 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1994_
timestamp 1698431365
transform 1 0 7168 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1995_
timestamp 1698431365
transform 1 0 14896 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1996_
timestamp 1698431365
transform 1 0 11200 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1997_
timestamp 1698431365
transform 1 0 10192 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1998_
timestamp 1698431365
transform 1 0 17584 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1999_
timestamp 1698431365
transform 1 0 12096 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2000_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2001_
timestamp 1698431365
transform 1 0 13776 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2002_
timestamp 1698431365
transform -1 0 23968 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2003_
timestamp 1698431365
transform -1 0 21504 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2004_
timestamp 1698431365
transform 1 0 25088 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2005_
timestamp 1698431365
transform 1 0 25088 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2006_
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2007_
timestamp 1698431365
transform 1 0 19264 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2008_
timestamp 1698431365
transform -1 0 28336 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2009_
timestamp 1698431365
transform 1 0 21728 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2010_
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2011_
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2012_
timestamp 1698431365
transform 1 0 24752 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2013_
timestamp 1698431365
transform -1 0 24864 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2014_
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2015_
timestamp 1698431365
transform 1 0 5040 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2016_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2017_
timestamp 1698431365
transform -1 0 10976 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2018_
timestamp 1698431365
transform 1 0 4256 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2019_
timestamp 1698431365
transform 1 0 4368 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2020_
timestamp 1698431365
transform -1 0 26208 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2021_
timestamp 1698431365
transform 1 0 20048 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2022_
timestamp 1698431365
transform 1 0 22624 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2023_
timestamp 1698431365
transform 1 0 16800 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2024_
timestamp 1698431365
transform 1 0 11760 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2025_
timestamp 1698431365
transform 1 0 9632 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2026_
timestamp 1698431365
transform 1 0 6608 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2027_
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2028_
timestamp 1698431365
transform 1 0 4592 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2029_
timestamp 1698431365
transform 1 0 4480 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2030_
timestamp 1698431365
transform 1 0 9968 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2031_
timestamp 1698431365
transform 1 0 4368 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2032_
timestamp 1698431365
transform 1 0 9408 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2033_
timestamp 1698431365
transform -1 0 13104 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2034_
timestamp 1698431365
transform 1 0 6048 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2035_
timestamp 1698431365
transform 1 0 5376 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2036_
timestamp 1698431365
transform 1 0 21616 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2037_
timestamp 1698431365
transform -1 0 26096 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2038_
timestamp 1698431365
transform -1 0 27664 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2039_
timestamp 1698431365
transform 1 0 15344 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2040_
timestamp 1698431365
transform -1 0 28000 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2041_
timestamp 1698431365
transform -1 0 28336 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2042_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2043_
timestamp 1698431365
transform 1 0 23184 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2044_
timestamp 1698431365
transform 1 0 23296 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2045_
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2046_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 -1 100352
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2047_
timestamp 1698431365
transform 1 0 5712 0 -1 101920
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2048_
timestamp 1698431365
transform 1 0 2800 0 -1 86240
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2049_
timestamp 1698431365
transform -1 0 7280 0 -1 97216
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2050_
timestamp 1698431365
transform 1 0 4592 0 -1 94080
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2051_
timestamp 1698431365
transform 1 0 1568 0 1 90944
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2052_
timestamp 1698431365
transform -1 0 8960 0 1 89376
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2053_
timestamp 1698431365
transform -1 0 10752 0 1 94080
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2054_
timestamp 1698431365
transform 1 0 18592 0 -1 103488
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2055_
timestamp 1698431365
transform -1 0 24416 0 1 100352
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2056_
timestamp 1698431365
transform -1 0 27664 0 1 100352
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2057_
timestamp 1698431365
transform -1 0 28336 0 -1 98784
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2058_
timestamp 1698431365
transform -1 0 28336 0 -1 97216
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2059_
timestamp 1698431365
transform 1 0 24864 0 1 94080
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2060_
timestamp 1698431365
transform 1 0 18816 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2061_
timestamp 1698431365
transform 1 0 12096 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2062_
timestamp 1698431365
transform 1 0 22400 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2063_
timestamp 1698431365
transform 1 0 15792 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2064_
timestamp 1698431365
transform 1 0 18256 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2065_
timestamp 1698431365
transform 1 0 15568 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2066_
timestamp 1698431365
transform -1 0 24752 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2067_
timestamp 1698431365
transform 1 0 12656 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2068_
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2069_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2070_
timestamp 1698431365
transform 1 0 4928 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2071_
timestamp 1698431365
transform 1 0 8848 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2072_
timestamp 1698431365
transform 1 0 6944 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2073_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2074_
timestamp 1698431365
transform 1 0 10416 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2075_
timestamp 1698431365
transform 1 0 9856 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2076_
timestamp 1698431365
transform 1 0 7504 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2077_
timestamp 1698431365
transform 1 0 6272 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2078_
timestamp 1698431365
transform 1 0 16688 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2079_
timestamp 1698431365
transform 1 0 13216 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2080_
timestamp 1698431365
transform -1 0 24416 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2081_
timestamp 1698431365
transform 1 0 14672 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2082_
timestamp 1698431365
transform -1 0 28336 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2083_
timestamp 1698431365
transform -1 0 28336 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2084_
timestamp 1698431365
transform -1 0 28336 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2085_
timestamp 1698431365
transform 1 0 12768 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2086_
timestamp 1698431365
transform -1 0 28336 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2087_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2088_
timestamp 1698431365
transform -1 0 28336 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2089_
timestamp 1698431365
transform -1 0 28336 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2090_
timestamp 1698431365
transform -1 0 28336 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2091_
timestamp 1698431365
transform 1 0 20384 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2092_
timestamp 1698431365
transform 1 0 5936 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2093_
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2094_
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2095_
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2096_
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2097_
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2098_
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2099_
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2100_
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2101_
timestamp 1698431365
transform 1 0 4256 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2102_
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2103_
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2104_
timestamp 1698431365
transform 1 0 3920 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2105_
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2106_
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2107_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2108_
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2109_
timestamp 1698431365
transform 1 0 4144 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2110_
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2111_
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2112_
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2113_
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2114_
timestamp 1698431365
transform 1 0 1568 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2115_
timestamp 1698431365
transform 1 0 1568 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2116_
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2117_
timestamp 1698431365
transform 1 0 1568 0 1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2118_
timestamp 1698431365
transform 1 0 1568 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2119_
timestamp 1698431365
transform 1 0 1568 0 1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2120_
timestamp 1698431365
transform 1 0 4368 0 -1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2121_
timestamp 1698431365
transform 1 0 1568 0 1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2122_
timestamp 1698431365
transform 1 0 6272 0 1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2123_
timestamp 1698431365
transform 1 0 3920 0 -1 83104
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2124_
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2125_
timestamp 1698431365
transform 1 0 9856 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2126_
timestamp 1698431365
transform 1 0 17696 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2127_
timestamp 1698431365
transform 1 0 15904 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2128_
timestamp 1698431365
transform 1 0 13776 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2129_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2130_
timestamp 1698431365
transform 1 0 11872 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2131_
timestamp 1698431365
transform 1 0 13440 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2132_
timestamp 1698431365
transform -1 0 24416 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2133_
timestamp 1698431365
transform 1 0 16128 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2134_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2135_
timestamp 1698431365
transform 1 0 9520 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2136_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2137_
timestamp 1698431365
transform 1 0 13328 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2138_
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2139_
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2140_
timestamp 1698431365
transform -1 0 19152 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2141_
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2142_
timestamp 1698431365
transform 1 0 8736 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2143_
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2144_
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2145_
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2146_
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2147_
timestamp 1698431365
transform 1 0 25088 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2148_
timestamp 1698431365
transform 1 0 25088 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2149_
timestamp 1698431365
transform 1 0 13776 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2150_
timestamp 1698431365
transform -1 0 28336 0 1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2151_
timestamp 1698431365
transform 1 0 25088 0 -1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2152_
timestamp 1698431365
transform -1 0 28336 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2153_
timestamp 1698431365
transform -1 0 28336 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2154_
timestamp 1698431365
transform -1 0 28336 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2155_
timestamp 1698431365
transform 1 0 21168 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2156_
timestamp 1698431365
transform -1 0 4816 0 -1 89376
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2157_
timestamp 1698431365
transform 1 0 14672 0 1 81536
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2158_
timestamp 1698431365
transform 1 0 18704 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2159_
timestamp 1698431365
transform 1 0 8176 0 1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2160_
timestamp 1698431365
transform 1 0 21616 0 -1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2161_
timestamp 1698431365
transform 1 0 14672 0 1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2162_
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2163_
timestamp 1698431365
transform 1 0 13440 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2164_
timestamp 1698431365
transform 1 0 21280 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2165_
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2166_
timestamp 1698431365
transform 1 0 19936 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2167_
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2168_
timestamp 1698431365
transform 1 0 10304 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2169_
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2170_
timestamp 1698431365
transform 1 0 5936 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2171_
timestamp 1698431365
transform 1 0 2688 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2172_
timestamp 1698431365
transform 1 0 6048 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2173_
timestamp 1698431365
transform 1 0 3920 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2174_
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2175_
timestamp 1698431365
transform 1 0 4368 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2176_
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2177_
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2178_
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2179_
timestamp 1698431365
transform -1 0 20496 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2180_
timestamp 1698431365
transform 1 0 4144 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2181_
timestamp 1698431365
transform -1 0 20720 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2182_
timestamp 1698431365
transform 1 0 4144 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2183_
timestamp 1698431365
transform 1 0 4816 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2184_
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2185_
timestamp 1698431365
transform 1 0 5488 0 1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2186_
timestamp 1698431365
transform -1 0 20944 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2187_
timestamp 1698431365
transform -1 0 21280 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2188_
timestamp 1698431365
transform 1 0 21616 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2189_
timestamp 1698431365
transform 1 0 19936 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2190_
timestamp 1698431365
transform -1 0 4816 0 1 92512
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2191_
timestamp 1698431365
transform -1 0 4816 0 1 95648
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2192_
timestamp 1698431365
transform -1 0 4816 0 1 98784
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2193_
timestamp 1698431365
transform -1 0 4816 0 -1 101920
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2194_
timestamp 1698431365
transform -1 0 4816 0 1 103488
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2195_
timestamp 1698431365
transform -1 0 8960 0 1 103488
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2196_
timestamp 1698431365
transform -1 0 4816 0 1 105056
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2197_
timestamp 1698431365
transform -1 0 8736 0 1 105056
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2198_
timestamp 1698431365
transform 1 0 13552 0 1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2199_
timestamp 1698431365
transform 1 0 10864 0 -1 84672
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2200_
timestamp 1698431365
transform 1 0 9296 0 1 83104
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2201_
timestamp 1698431365
transform 1 0 6272 0 1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2202_
timestamp 1698431365
transform 1 0 9856 0 1 87808
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2203_
timestamp 1698431365
transform 1 0 5936 0 -1 87808
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2204_
timestamp 1698431365
transform 1 0 7728 0 1 90944
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2205_
timestamp 1698431365
transform 1 0 9184 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2206_
timestamp 1698431365
transform 1 0 8288 0 1 92512
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2207_
timestamp 1698431365
transform 1 0 5712 0 -1 98784
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__I open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27776 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__I
timestamp 1698431365
transform 1 0 16800 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__A1
timestamp 1698431365
transform -1 0 2912 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__A2
timestamp 1698431365
transform -1 0 3360 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__A3
timestamp 1698431365
transform -1 0 2464 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A1
timestamp 1698431365
transform 1 0 4480 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__A1
timestamp 1698431365
transform -1 0 4592 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__A2
timestamp 1698431365
transform -1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__A1
timestamp 1698431365
transform -1 0 23632 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A1
timestamp 1698431365
transform 1 0 26208 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__I
timestamp 1698431365
transform -1 0 5936 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__A1
timestamp 1698431365
transform 1 0 7616 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__A1
timestamp 1698431365
transform 1 0 21392 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1000__A1
timestamp 1698431365
transform 1 0 5040 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__A1
timestamp 1698431365
transform -1 0 5264 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__A1
timestamp 1698431365
transform -1 0 5712 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A1
timestamp 1698431365
transform 1 0 7280 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1004__A3
timestamp 1698431365
transform 1 0 5600 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1008__I
timestamp 1698431365
transform 1 0 10192 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__A1
timestamp 1698431365
transform 1 0 18816 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__I
timestamp 1698431365
transform 1 0 16800 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A1
timestamp 1698431365
transform -1 0 8288 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A2
timestamp 1698431365
transform 1 0 19600 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A3
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__A1
timestamp 1698431365
transform 1 0 11312 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__A2
timestamp 1698431365
transform -1 0 7840 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__I
timestamp 1698431365
transform 1 0 16464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1022__I
timestamp 1698431365
transform 1 0 7840 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A1
timestamp 1698431365
transform 1 0 10640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A2
timestamp 1698431365
transform 1 0 11088 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A3
timestamp 1698431365
transform 1 0 24752 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A4
timestamp 1698431365
transform -1 0 10976 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__A1
timestamp 1698431365
transform -1 0 7392 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__A2
timestamp 1698431365
transform -1 0 6832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__I
timestamp 1698431365
transform 1 0 24528 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A1
timestamp 1698431365
transform 1 0 12880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A2
timestamp 1698431365
transform 1 0 14560 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A3
timestamp 1698431365
transform 1 0 19824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A4
timestamp 1698431365
transform 1 0 20272 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__A1
timestamp 1698431365
transform 1 0 11200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__A2
timestamp 1698431365
transform -1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1029__B1
timestamp 1698431365
transform -1 0 3472 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1029__B2
timestamp 1698431365
transform 1 0 3696 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__A1
timestamp 1698431365
transform 1 0 24640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__A2
timestamp 1698431365
transform 1 0 23632 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__I
timestamp 1698431365
transform 1 0 11872 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__A1
timestamp 1698431365
transform 1 0 12432 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__A2
timestamp 1698431365
transform 1 0 11984 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__A3
timestamp 1698431365
transform 1 0 18368 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__A4
timestamp 1698431365
transform 1 0 17472 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__A1
timestamp 1698431365
transform 1 0 14896 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__B1
timestamp 1698431365
transform 1 0 27104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A1
timestamp 1698431365
transform 1 0 12208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A2
timestamp 1698431365
transform 1 0 9968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A1
timestamp 1698431365
transform -1 0 11984 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A2
timestamp 1698431365
transform -1 0 11536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A3
timestamp 1698431365
transform 1 0 10752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__A1
timestamp 1698431365
transform 1 0 14000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__A2
timestamp 1698431365
transform 1 0 11536 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A2
timestamp 1698431365
transform -1 0 19600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__B1
timestamp 1698431365
transform -1 0 19152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A1
timestamp 1698431365
transform 1 0 8624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A2
timestamp 1698431365
transform 1 0 8176 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A3
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A4
timestamp 1698431365
transform 1 0 17920 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A1
timestamp 1698431365
transform 1 0 26656 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A3
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A1
timestamp 1698431365
transform 1 0 20160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A3
timestamp 1698431365
transform 1 0 21728 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A3
timestamp 1698431365
transform 1 0 23856 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__A1
timestamp 1698431365
transform 1 0 17472 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A1
timestamp 1698431365
transform 1 0 20048 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A2
timestamp 1698431365
transform 1 0 22848 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A3
timestamp 1698431365
transform 1 0 19712 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__A2
timestamp 1698431365
transform 1 0 25312 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__B1
timestamp 1698431365
transform 1 0 24528 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A2
timestamp 1698431365
transform 1 0 22736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A3
timestamp 1698431365
transform 1 0 13776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A2
timestamp 1698431365
transform -1 0 24192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__B1
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A1
timestamp 1698431365
transform 1 0 13888 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A2
timestamp 1698431365
transform 1 0 12880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A3
timestamp 1698431365
transform 1 0 12432 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A1
timestamp 1698431365
transform 1 0 19376 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__B1
timestamp 1698431365
transform 1 0 9968 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__A2
timestamp 1698431365
transform 1 0 22288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__A3
timestamp 1698431365
transform 1 0 11984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698431365
transform -1 0 10640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A2
timestamp 1698431365
transform -1 0 5936 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1056__A1
timestamp 1698431365
transform -1 0 13328 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1056__A2
timestamp 1698431365
transform -1 0 11088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1056__A3
timestamp 1698431365
transform 1 0 10304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A1
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A2
timestamp 1698431365
transform 1 0 21504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__B1
timestamp 1698431365
transform -1 0 20496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__A2
timestamp 1698431365
transform 1 0 10864 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__A3
timestamp 1698431365
transform -1 0 16016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698431365
transform -1 0 23296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A2
timestamp 1698431365
transform -1 0 21392 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__A2
timestamp 1698431365
transform 1 0 21952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__B1
timestamp 1698431365
transform 1 0 22400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1061__A1
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A1
timestamp 1698431365
transform 1 0 12880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A2
timestamp 1698431365
transform 1 0 13552 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A1
timestamp 1698431365
transform 1 0 15344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A2
timestamp 1698431365
transform 1 0 14448 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A3
timestamp 1698431365
transform 1 0 11760 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A4
timestamp 1698431365
transform 1 0 14784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__A1
timestamp 1698431365
transform 1 0 11872 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1068__A1
timestamp 1698431365
transform 1 0 20720 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1068__A2
timestamp 1698431365
transform 1 0 17808 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1068__A3
timestamp 1698431365
transform 1 0 17360 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1068__A4
timestamp 1698431365
transform 1 0 16800 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A1
timestamp 1698431365
transform 1 0 12432 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A3
timestamp 1698431365
transform 1 0 12880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1072__A1
timestamp 1698431365
transform 1 0 12432 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1072__A2
timestamp 1698431365
transform 1 0 12880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698431365
transform 1 0 19264 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A2
timestamp 1698431365
transform 1 0 17136 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A3
timestamp 1698431365
transform 1 0 17472 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A1
timestamp 1698431365
transform 1 0 16352 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A2
timestamp 1698431365
transform 1 0 20272 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A3
timestamp 1698431365
transform 1 0 14000 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A1
timestamp 1698431365
transform 1 0 11312 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A2
timestamp 1698431365
transform 1 0 10416 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A4
timestamp 1698431365
transform 1 0 10864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A2
timestamp 1698431365
transform -1 0 15120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A3
timestamp 1698431365
transform -1 0 12880 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__A2
timestamp 1698431365
transform 1 0 11536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__B
timestamp 1698431365
transform -1 0 12208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A1
timestamp 1698431365
transform -1 0 12432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__A1
timestamp 1698431365
transform 1 0 11536 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__A2
timestamp 1698431365
transform -1 0 7952 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__A3
timestamp 1698431365
transform -1 0 7504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A1
timestamp 1698431365
transform 1 0 12432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A2
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__B1
timestamp 1698431365
transform -1 0 10192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__A1
timestamp 1698431365
transform 1 0 9072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__A3
timestamp 1698431365
transform -1 0 11312 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__A1
timestamp 1698431365
transform 1 0 16800 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__A2
timestamp 1698431365
transform 1 0 17920 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__A3
timestamp 1698431365
transform 1 0 7056 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A2
timestamp 1698431365
transform -1 0 9968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__B1
timestamp 1698431365
transform 1 0 10192 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__A2
timestamp 1698431365
transform -1 0 23184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__A3
timestamp 1698431365
transform -1 0 14672 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A1
timestamp 1698431365
transform 1 0 22064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A2
timestamp 1698431365
transform 1 0 13552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__B1
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A2
timestamp 1698431365
transform 1 0 20608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A4
timestamp 1698431365
transform -1 0 16464 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A2
timestamp 1698431365
transform 1 0 20160 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__B1
timestamp 1698431365
transform 1 0 24752 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A1
timestamp 1698431365
transform 1 0 23632 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A1
timestamp 1698431365
transform 1 0 22848 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A2
timestamp 1698431365
transform -1 0 21840 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__B1
timestamp 1698431365
transform -1 0 6160 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__B2
timestamp 1698431365
transform -1 0 2240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__B1
timestamp 1698431365
transform 1 0 27552 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__A2
timestamp 1698431365
transform 1 0 19264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__B1
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A1
timestamp 1698431365
transform 1 0 27216 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A3
timestamp 1698431365
transform 1 0 25760 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A1
timestamp 1698431365
transform 1 0 23968 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A3
timestamp 1698431365
transform 1 0 21616 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A3
timestamp 1698431365
transform 1 0 24304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A2
timestamp 1698431365
transform -1 0 23072 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__B1
timestamp 1698431365
transform -1 0 22624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A2
timestamp 1698431365
transform -1 0 23744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__B1
timestamp 1698431365
transform 1 0 22064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__B1
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__A2
timestamp 1698431365
transform 1 0 19264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__B1
timestamp 1698431365
transform -1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A2
timestamp 1698431365
transform 1 0 20384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__B1
timestamp 1698431365
transform 1 0 19376 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A1
timestamp 1698431365
transform 1 0 18592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__A1
timestamp 1698431365
transform 1 0 13440 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__A2
timestamp 1698431365
transform 1 0 12992 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__A3
timestamp 1698431365
transform 1 0 19040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__A1
timestamp 1698431365
transform 1 0 10640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__A1
timestamp 1698431365
transform 1 0 13552 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__A3
timestamp 1698431365
transform -1 0 14672 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A1
timestamp 1698431365
transform 1 0 10080 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A2
timestamp 1698431365
transform 1 0 8960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A4
timestamp 1698431365
transform 1 0 9632 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A2
timestamp 1698431365
transform 1 0 10752 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__B
timestamp 1698431365
transform -1 0 9632 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A2
timestamp 1698431365
transform 1 0 7728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__B1
timestamp 1698431365
transform 1 0 8512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A2
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__B1
timestamp 1698431365
transform 1 0 11424 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__A2
timestamp 1698431365
transform 1 0 11648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__B1
timestamp 1698431365
transform 1 0 12432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__A2
timestamp 1698431365
transform 1 0 20720 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__A4
timestamp 1698431365
transform -1 0 16016 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A2
timestamp 1698431365
transform -1 0 19600 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__B1
timestamp 1698431365
transform 1 0 20720 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__A1
timestamp 1698431365
transform 1 0 18816 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698431365
transform -1 0 18144 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A2
timestamp 1698431365
transform 1 0 19264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A1
timestamp 1698431365
transform -1 0 2352 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__B1
timestamp 1698431365
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__B2
timestamp 1698431365
transform 1 0 4144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1130__B1
timestamp 1698431365
transform 1 0 27664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__A2
timestamp 1698431365
transform -1 0 20048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__B1
timestamp 1698431365
transform -1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1132__A1
timestamp 1698431365
transform -1 0 20160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1132__A3
timestamp 1698431365
transform 1 0 19488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__A1
timestamp 1698431365
transform 1 0 17920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__A2
timestamp 1698431365
transform -1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__A3
timestamp 1698431365
transform 1 0 17920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__A3
timestamp 1698431365
transform 1 0 23408 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__A4
timestamp 1698431365
transform 1 0 24304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__A2
timestamp 1698431365
transform 1 0 21728 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__B1
timestamp 1698431365
transform 1 0 21728 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A2
timestamp 1698431365
transform 1 0 23856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__B1
timestamp 1698431365
transform 1 0 23408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__B1
timestamp 1698431365
transform -1 0 8176 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__A2
timestamp 1698431365
transform 1 0 21392 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__B1
timestamp 1698431365
transform 1 0 19488 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__A2
timestamp 1698431365
transform -1 0 18704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__B1
timestamp 1698431365
transform 1 0 20720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__A2
timestamp 1698431365
transform -1 0 19152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__A1
timestamp 1698431365
transform 1 0 11088 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__A1
timestamp 1698431365
transform 1 0 15120 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__A3
timestamp 1698431365
transform 1 0 16688 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A1
timestamp 1698431365
transform 1 0 10416 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A2
timestamp 1698431365
transform 1 0 9968 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A4
timestamp 1698431365
transform 1 0 10864 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__A2
timestamp 1698431365
transform 1 0 12208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__B
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__A1
timestamp 1698431365
transform 1 0 9632 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__A2
timestamp 1698431365
transform 1 0 8960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__B1
timestamp 1698431365
transform 1 0 10080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__A2
timestamp 1698431365
transform 1 0 10416 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__B1
timestamp 1698431365
transform 1 0 11424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__A2
timestamp 1698431365
transform 1 0 11648 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__B1
timestamp 1698431365
transform 1 0 11200 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__A2
timestamp 1698431365
transform 1 0 19936 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__A4
timestamp 1698431365
transform 1 0 19376 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__A2
timestamp 1698431365
transform 1 0 18928 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__A1
timestamp 1698431365
transform 1 0 24192 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A1
timestamp 1698431365
transform 1 0 23296 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A2
timestamp 1698431365
transform 1 0 23744 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__A1
timestamp 1698431365
transform 1 0 5264 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__B1
timestamp 1698431365
transform 1 0 4368 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__B2
timestamp 1698431365
transform -1 0 5040 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__B1
timestamp 1698431365
transform 1 0 24640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__A2
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__B1
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A1
timestamp 1698431365
transform -1 0 13328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A3
timestamp 1698431365
transform 1 0 13328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A1
timestamp 1698431365
transform -1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A2
timestamp 1698431365
transform 1 0 11872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A3
timestamp 1698431365
transform -1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1168__A3
timestamp 1698431365
transform 1 0 23744 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1168__A4
timestamp 1698431365
transform 1 0 23296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1169__A2
timestamp 1698431365
transform 1 0 21840 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1169__B1
timestamp 1698431365
transform 1 0 22288 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A2
timestamp 1698431365
transform 1 0 21280 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__B1
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__B2
timestamp 1698431365
transform 1 0 21728 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__B1
timestamp 1698431365
transform -1 0 14000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__A2
timestamp 1698431365
transform 1 0 20944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__B1
timestamp 1698431365
transform 1 0 18032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__A2
timestamp 1698431365
transform 1 0 19824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__B1
timestamp 1698431365
transform 1 0 20832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__A1
timestamp 1698431365
transform 1 0 14000 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1180__A1
timestamp 1698431365
transform 1 0 15120 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1180__A3
timestamp 1698431365
transform 1 0 18816 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A1
timestamp 1698431365
transform 1 0 9072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A2
timestamp 1698431365
transform 1 0 7952 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A4
timestamp 1698431365
transform 1 0 9520 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__A2
timestamp 1698431365
transform 1 0 10752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__B
timestamp 1698431365
transform 1 0 10304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1186__A1
timestamp 1698431365
transform -1 0 7728 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1186__A2
timestamp 1698431365
transform -1 0 6832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1186__B1
timestamp 1698431365
transform -1 0 7280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__A1
timestamp 1698431365
transform 1 0 11760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__A2
timestamp 1698431365
transform 1 0 9856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__B1
timestamp 1698431365
transform 1 0 12208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__A2
timestamp 1698431365
transform 1 0 11312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__B1
timestamp 1698431365
transform 1 0 11200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__A2
timestamp 1698431365
transform 1 0 18704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__A4
timestamp 1698431365
transform -1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__A2
timestamp 1698431365
transform 1 0 16352 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__A1
timestamp 1698431365
transform 1 0 25760 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A1
timestamp 1698431365
transform -1 0 23408 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A2
timestamp 1698431365
transform 1 0 24976 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__A2
timestamp 1698431365
transform 1 0 18816 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1196__A2
timestamp 1698431365
transform 1 0 20160 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1197__A1
timestamp 1698431365
transform 1 0 22624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1197__A3
timestamp 1698431365
transform -1 0 23184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1198__A1
timestamp 1698431365
transform 1 0 11984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1198__A2
timestamp 1698431365
transform 1 0 13888 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1198__A3
timestamp 1698431365
transform 1 0 14336 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1198__A4
timestamp 1698431365
transform 1 0 13552 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A1
timestamp 1698431365
transform 1 0 16128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A2
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A3
timestamp 1698431365
transform -1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__A2
timestamp 1698431365
transform 1 0 19040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__B1
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__A1
timestamp 1698431365
transform 1 0 7504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__A2
timestamp 1698431365
transform -1 0 9632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__B1
timestamp 1698431365
transform -1 0 9184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__B2
timestamp 1698431365
transform -1 0 7280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1204__A1
timestamp 1698431365
transform 1 0 19488 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1204__A2
timestamp 1698431365
transform 1 0 17472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1204__A3
timestamp 1698431365
transform -1 0 20160 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1204__A4
timestamp 1698431365
transform 1 0 11760 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__A1
timestamp 1698431365
transform 1 0 21392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__A3
timestamp 1698431365
transform 1 0 21392 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__A1
timestamp 1698431365
transform 1 0 22736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__A3
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A2
timestamp 1698431365
transform 1 0 12320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__B1
timestamp 1698431365
transform -1 0 11872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__A1
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__A3
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__A1
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__A2
timestamp 1698431365
transform 1 0 18368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__A3
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__A2
timestamp 1698431365
transform 1 0 21168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__B1
timestamp 1698431365
transform 1 0 19488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1215__A2
timestamp 1698431365
transform 1 0 10080 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A2
timestamp 1698431365
transform 1 0 16464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__B1
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__C
timestamp 1698431365
transform 1 0 15792 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1218__A1
timestamp 1698431365
transform -1 0 15232 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__A1
timestamp 1698431365
transform 1 0 13776 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__A3
timestamp 1698431365
transform 1 0 14896 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__A2
timestamp 1698431365
transform 1 0 13888 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__A1
timestamp 1698431365
transform 1 0 15344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__A2
timestamp 1698431365
transform 1 0 16240 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__A4
timestamp 1698431365
transform 1 0 17696 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A1
timestamp 1698431365
transform -1 0 16240 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__A2
timestamp 1698431365
transform 1 0 14896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1224__A1
timestamp 1698431365
transform 1 0 12432 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1224__A2
timestamp 1698431365
transform -1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1224__A3
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__A2
timestamp 1698431365
transform 1 0 15568 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A1
timestamp 1698431365
transform -1 0 11872 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__A1
timestamp 1698431365
transform 1 0 14560 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__A2
timestamp 1698431365
transform 1 0 14000 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__A3
timestamp 1698431365
transform 1 0 14448 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__B1
timestamp 1698431365
transform 1 0 24304 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1229__B1
timestamp 1698431365
transform 1 0 13552 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__A2
timestamp 1698431365
transform 1 0 18704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__B1
timestamp 1698431365
transform 1 0 24976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__C
timestamp 1698431365
transform 1 0 19824 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1233__A2
timestamp 1698431365
transform -1 0 20944 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__B1
timestamp 1698431365
transform -1 0 11312 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1237__A2
timestamp 1698431365
transform 1 0 23408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__A1
timestamp 1698431365
transform -1 0 4928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__A2
timestamp 1698431365
transform 1 0 6160 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__B1
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__B2
timestamp 1698431365
transform -1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__B1
timestamp 1698431365
transform 1 0 16800 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1241__A2
timestamp 1698431365
transform 1 0 10192 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1241__B1
timestamp 1698431365
transform -1 0 9968 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__A2
timestamp 1698431365
transform 1 0 24080 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__A2
timestamp 1698431365
transform 1 0 14672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__A1
timestamp 1698431365
transform 1 0 18816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__A3
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1245__A1
timestamp 1698431365
transform 1 0 7616 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1245__A2
timestamp 1698431365
transform -1 0 11424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1245__A3
timestamp 1698431365
transform 1 0 8064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__A1
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__A3
timestamp 1698431365
transform -1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1247__A3
timestamp 1698431365
transform -1 0 15792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__A3
timestamp 1698431365
transform 1 0 21392 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1249__A1
timestamp 1698431365
transform 1 0 8848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1249__A2
timestamp 1698431365
transform -1 0 9520 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1250__B1
timestamp 1698431365
transform -1 0 8176 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1251__A2
timestamp 1698431365
transform 1 0 17584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1251__B1
timestamp 1698431365
transform 1 0 17136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__A2
timestamp 1698431365
transform -1 0 14336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__B1
timestamp 1698431365
transform -1 0 15792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1253__A2
timestamp 1698431365
transform 1 0 16016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1253__B1
timestamp 1698431365
transform -1 0 13664 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A1
timestamp 1698431365
transform 1 0 14560 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__B
timestamp 1698431365
transform 1 0 15568 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__C
timestamp 1698431365
transform 1 0 13552 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1256__A1
timestamp 1698431365
transform -1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1256__A2
timestamp 1698431365
transform 1 0 8512 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1257__A1
timestamp 1698431365
transform 1 0 10752 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A1
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A2
timestamp 1698431365
transform 1 0 12096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A3
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1259__A2
timestamp 1698431365
transform 1 0 16240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1259__B1
timestamp 1698431365
transform -1 0 16016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__A2
timestamp 1698431365
transform 1 0 24192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__B1
timestamp 1698431365
transform 1 0 22848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A3
timestamp 1698431365
transform 1 0 15568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A2
timestamp 1698431365
transform 1 0 18928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A4
timestamp 1698431365
transform 1 0 20608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__A2
timestamp 1698431365
transform -1 0 17248 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__A1
timestamp 1698431365
transform -1 0 17248 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1285__A1
timestamp 1698431365
transform 1 0 18480 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__B
timestamp 1698431365
transform 1 0 20608 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__A1
timestamp 1698431365
transform 1 0 15568 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__A2
timestamp 1698431365
transform 1 0 13888 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__A1
timestamp 1698431365
transform 1 0 7056 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__A2
timestamp 1698431365
transform -1 0 16912 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A1
timestamp 1698431365
transform -1 0 21392 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A2
timestamp 1698431365
transform 1 0 20720 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__A1
timestamp 1698431365
transform -1 0 19600 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1299__A1
timestamp 1698431365
transform 1 0 19376 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1301__B
timestamp 1698431365
transform 1 0 16688 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1303__A1
timestamp 1698431365
transform 1 0 19264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1303__A2
timestamp 1698431365
transform 1 0 18368 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__A2
timestamp 1698431365
transform 1 0 13104 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__B
timestamp 1698431365
transform 1 0 18368 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1310__A1
timestamp 1698431365
transform 1 0 6048 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1313__I
timestamp 1698431365
transform 1 0 24640 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1314__A1
timestamp 1698431365
transform 1 0 18928 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1314__A2
timestamp 1698431365
transform 1 0 16800 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__A1
timestamp 1698431365
transform 1 0 19376 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A1
timestamp 1698431365
transform 1 0 19600 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1319__A1
timestamp 1698431365
transform 1 0 19600 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__A1
timestamp 1698431365
transform 1 0 20272 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__A2
timestamp 1698431365
transform -1 0 20048 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1323__A2
timestamp 1698431365
transform -1 0 4368 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1323__B
timestamp 1698431365
transform -1 0 5264 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1325__A3
timestamp 1698431365
transform 1 0 6832 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__A1
timestamp 1698431365
transform 1 0 23296 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__A2
timestamp 1698431365
transform 1 0 19712 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1329__A1
timestamp 1698431365
transform 1 0 24192 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__A1
timestamp 1698431365
transform 1 0 21280 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1333__A1
timestamp 1698431365
transform -1 0 19824 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1335__A1
timestamp 1698431365
transform -1 0 12096 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1335__A2
timestamp 1698431365
transform 1 0 17920 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1336__A2
timestamp 1698431365
transform 1 0 6048 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1336__B
timestamp 1698431365
transform 1 0 5936 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1339__A1
timestamp 1698431365
transform 1 0 24752 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__A1
timestamp 1698431365
transform 1 0 24640 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__A2
timestamp 1698431365
transform -1 0 15680 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__A1
timestamp 1698431365
transform 1 0 18480 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A1
timestamp 1698431365
transform 1 0 19376 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1347__A1
timestamp 1698431365
transform -1 0 19712 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A1
timestamp 1698431365
transform -1 0 17696 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A2
timestamp 1698431365
transform 1 0 16576 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__A1
timestamp 1698431365
transform 1 0 20608 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__A2
timestamp 1698431365
transform 1 0 22288 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__B
timestamp 1698431365
transform 1 0 21840 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__A1
timestamp 1698431365
transform 1 0 18928 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__A1
timestamp 1698431365
transform 1 0 13664 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A1
timestamp 1698431365
transform 1 0 9408 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A1
timestamp 1698431365
transform -1 0 5376 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A2
timestamp 1698431365
transform 1 0 8512 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__B
timestamp 1698431365
transform 1 0 6048 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1367__A1
timestamp 1698431365
transform -1 0 17920 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A1
timestamp 1698431365
transform 1 0 20496 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A1
timestamp 1698431365
transform 1 0 20720 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__C
timestamp 1698431365
transform 1 0 21840 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A2
timestamp 1698431365
transform 1 0 5040 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__C
timestamp 1698431365
transform 1 0 8512 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__A1
timestamp 1698431365
transform -1 0 9184 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__A2
timestamp 1698431365
transform -1 0 9184 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A1
timestamp 1698431365
transform 1 0 13216 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__A2
timestamp 1698431365
transform 1 0 17472 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A1
timestamp 1698431365
transform -1 0 17696 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__C
timestamp 1698431365
transform 1 0 9856 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__A1
timestamp 1698431365
transform 1 0 13104 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__A2
timestamp 1698431365
transform 1 0 8960 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__A2
timestamp 1698431365
transform -1 0 13104 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__A1
timestamp 1698431365
transform 1 0 7616 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__I
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__I
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__I
timestamp 1698431365
transform 1 0 21280 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__A2
timestamp 1698431365
transform 1 0 20272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__B
timestamp 1698431365
transform 1 0 20720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698431365
transform 1 0 18480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A2
timestamp 1698431365
transform 1 0 19824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__A2
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__B
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A1
timestamp 1698431365
transform 1 0 10080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A2
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__A2
timestamp 1698431365
transform 1 0 22624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__B
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A1
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A2
timestamp 1698431365
transform -1 0 21840 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__A2
timestamp 1698431365
transform 1 0 17584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__B
timestamp 1698431365
transform 1 0 18032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A1
timestamp 1698431365
transform 1 0 15344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A2
timestamp 1698431365
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__A2
timestamp 1698431365
transform 1 0 12320 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__B
timestamp 1698431365
transform 1 0 13104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__A1
timestamp 1698431365
transform 1 0 8512 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__A2
timestamp 1698431365
transform 1 0 9744 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1424__I
timestamp 1698431365
transform 1 0 25312 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__A2
timestamp 1698431365
transform -1 0 11088 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__B
timestamp 1698431365
transform 1 0 12096 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1426__A1
timestamp 1698431365
transform 1 0 8624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1426__A2
timestamp 1698431365
transform -1 0 9408 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1428__A2
timestamp 1698431365
transform -1 0 24192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1428__B
timestamp 1698431365
transform -1 0 25760 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A1
timestamp 1698431365
transform -1 0 23296 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A2
timestamp 1698431365
transform 1 0 26096 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A2
timestamp 1698431365
transform 1 0 12880 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__B
timestamp 1698431365
transform 1 0 12432 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__A1
timestamp 1698431365
transform 1 0 10416 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__A2
timestamp 1698431365
transform 1 0 11200 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1434__I
timestamp 1698431365
transform 1 0 25760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__A2
timestamp 1698431365
transform 1 0 24416 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__B
timestamp 1698431365
transform 1 0 24416 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1436__A1
timestamp 1698431365
transform 1 0 22736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1436__A2
timestamp 1698431365
transform 1 0 23296 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A2
timestamp 1698431365
transform 1 0 9184 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__B
timestamp 1698431365
transform 1 0 8512 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A1
timestamp 1698431365
transform 1 0 7952 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A2
timestamp 1698431365
transform 1 0 8400 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A2
timestamp 1698431365
transform 1 0 9520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__B
timestamp 1698431365
transform 1 0 6160 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1442__A1
timestamp 1698431365
transform 1 0 6160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1442__A2
timestamp 1698431365
transform 1 0 6608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__A2
timestamp 1698431365
transform 1 0 7056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__B
timestamp 1698431365
transform 1 0 7504 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__A1
timestamp 1698431365
transform 1 0 7952 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__A2
timestamp 1698431365
transform -1 0 5936 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1447__A2
timestamp 1698431365
transform -1 0 5264 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1447__B
timestamp 1698431365
transform -1 0 5712 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1448__A1
timestamp 1698431365
transform -1 0 6608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1448__A2
timestamp 1698431365
transform 1 0 6832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1450__A2
timestamp 1698431365
transform 1 0 21392 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1450__B
timestamp 1698431365
transform 1 0 22288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__A1
timestamp 1698431365
transform 1 0 16016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__A2
timestamp 1698431365
transform 1 0 20608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1453__A2
timestamp 1698431365
transform 1 0 11984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1453__B
timestamp 1698431365
transform 1 0 10080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A1
timestamp 1698431365
transform 1 0 11648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A2
timestamp 1698431365
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A2
timestamp 1698431365
transform 1 0 9408 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__B
timestamp 1698431365
transform 1 0 9856 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A1
timestamp 1698431365
transform 1 0 9632 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A2
timestamp 1698431365
transform 1 0 9632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__A2
timestamp 1698431365
transform 1 0 20160 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__B
timestamp 1698431365
transform 1 0 20384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__A1
timestamp 1698431365
transform -1 0 17920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__A2
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A2
timestamp 1698431365
transform 1 0 11536 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__B
timestamp 1698431365
transform 1 0 15120 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__A1
timestamp 1698431365
transform -1 0 13328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__A2
timestamp 1698431365
transform 1 0 14000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__A2
timestamp 1698431365
transform 1 0 20608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__B
timestamp 1698431365
transform 1 0 22736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__A1
timestamp 1698431365
transform 1 0 17584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__A2
timestamp 1698431365
transform 1 0 18928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__A2
timestamp 1698431365
transform 1 0 18368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__B
timestamp 1698431365
transform 1 0 19936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A1
timestamp 1698431365
transform 1 0 14112 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A2
timestamp 1698431365
transform 1 0 14560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1471__A2
timestamp 1698431365
transform -1 0 23408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1471__B
timestamp 1698431365
transform -1 0 21840 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__A1
timestamp 1698431365
transform -1 0 21616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__A2
timestamp 1698431365
transform 1 0 22064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1474__A2
timestamp 1698431365
transform 1 0 22064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1474__B
timestamp 1698431365
transform 1 0 25088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A1
timestamp 1698431365
transform 1 0 22512 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A2
timestamp 1698431365
transform 1 0 21056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A2
timestamp 1698431365
transform 1 0 26432 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__B
timestamp 1698431365
transform 1 0 27776 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__A1
timestamp 1698431365
transform 1 0 25536 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__A2
timestamp 1698431365
transform 1 0 26880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1480__A2
timestamp 1698431365
transform 1 0 26208 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1480__B
timestamp 1698431365
transform 1 0 27552 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__A1
timestamp 1698431365
transform 1 0 26880 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__A2
timestamp 1698431365
transform 1 0 27328 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__A2
timestamp 1698431365
transform 1 0 26320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__B
timestamp 1698431365
transform 1 0 27440 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A1
timestamp 1698431365
transform 1 0 25760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A2
timestamp 1698431365
transform 1 0 27328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__I
timestamp 1698431365
transform -1 0 25536 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__A2
timestamp 1698431365
transform 1 0 25312 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__B
timestamp 1698431365
transform 1 0 25760 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A1
timestamp 1698431365
transform 1 0 23184 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A2
timestamp 1698431365
transform 1 0 24528 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A2
timestamp 1698431365
transform 1 0 26992 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__B
timestamp 1698431365
transform 1 0 27888 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1491__A1
timestamp 1698431365
transform 1 0 26096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1491__A2
timestamp 1698431365
transform 1 0 27440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__A2
timestamp 1698431365
transform 1 0 25312 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__B
timestamp 1698431365
transform 1 0 24864 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A1
timestamp 1698431365
transform 1 0 22512 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A2
timestamp 1698431365
transform 1 0 23744 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__A2
timestamp 1698431365
transform 1 0 27552 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__B
timestamp 1698431365
transform 1 0 27888 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A1
timestamp 1698431365
transform 1 0 26208 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A2
timestamp 1698431365
transform 1 0 28112 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1499__A2
timestamp 1698431365
transform 1 0 26992 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1499__B
timestamp 1698431365
transform 1 0 28000 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A1
timestamp 1698431365
transform 1 0 28000 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A2
timestamp 1698431365
transform 1 0 27440 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__I
timestamp 1698431365
transform 1 0 27104 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__A2
timestamp 1698431365
transform 1 0 26208 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__B
timestamp 1698431365
transform 1 0 27552 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A1
timestamp 1698431365
transform 1 0 27104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A2
timestamp 1698431365
transform 1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__I
timestamp 1698431365
transform 1 0 23744 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__A2
timestamp 1698431365
transform 1 0 28112 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__B
timestamp 1698431365
transform 1 0 27664 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__A1
timestamp 1698431365
transform 1 0 25088 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__A2
timestamp 1698431365
transform 1 0 26656 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__I
timestamp 1698431365
transform 1 0 26992 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1510__I
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A1
timestamp 1698431365
transform -1 0 10976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A2
timestamp 1698431365
transform 1 0 10528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__B
timestamp 1698431365
transform 1 0 9296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__A1
timestamp 1698431365
transform -1 0 8288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__A2
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A2
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__B
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A1
timestamp 1698431365
transform 1 0 6048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A2
timestamp 1698431365
transform 1 0 7168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__A1
timestamp 1698431365
transform -1 0 9072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__A2
timestamp 1698431365
transform 1 0 9632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__B
timestamp 1698431365
transform 1 0 9408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A1
timestamp 1698431365
transform 1 0 5600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A2
timestamp 1698431365
transform 1 0 6048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__A1
timestamp 1698431365
transform 1 0 11760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__A2
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__B
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1518__A1
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1518__A2
timestamp 1698431365
transform -1 0 12096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__A1
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__A2
timestamp 1698431365
transform -1 0 7728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__B
timestamp 1698431365
transform -1 0 7280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A1
timestamp 1698431365
transform 1 0 4144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1698431365
transform 1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A1
timestamp 1698431365
transform 1 0 6048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A2
timestamp 1698431365
transform 1 0 6496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__B
timestamp 1698431365
transform 1 0 8512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A1
timestamp 1698431365
transform 1 0 4592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A2
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__A2
timestamp 1698431365
transform 1 0 27104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__B
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A1
timestamp 1698431365
transform -1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A2
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__A2
timestamp 1698431365
transform 1 0 23520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__B
timestamp 1698431365
transform 1 0 22400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A1
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A2
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__I
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__A2
timestamp 1698431365
transform -1 0 26320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__B
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A1
timestamp 1698431365
transform 1 0 21168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A2
timestamp 1698431365
transform -1 0 24192 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A1
timestamp 1698431365
transform 1 0 20608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A2
timestamp 1698431365
transform 1 0 20160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__B
timestamp 1698431365
transform 1 0 19712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A1
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A2
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A2
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__B
timestamp 1698431365
transform 1 0 13664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1533__A1
timestamp 1698431365
transform 1 0 12208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1533__A2
timestamp 1698431365
transform 1 0 14896 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__A2
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__B
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__A1
timestamp 1698431365
transform 1 0 8064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__A2
timestamp 1698431365
transform 1 0 11312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1536__A2
timestamp 1698431365
transform 1 0 10976 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1536__B
timestamp 1698431365
transform 1 0 10528 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__A1
timestamp 1698431365
transform 1 0 7392 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__A2
timestamp 1698431365
transform 1 0 8736 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__I
timestamp 1698431365
transform 1 0 27888 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__A2
timestamp 1698431365
transform 1 0 8848 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__B
timestamp 1698431365
transform 1 0 8400 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__A1
timestamp 1698431365
transform 1 0 5712 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__A2
timestamp 1698431365
transform 1 0 7056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__A2
timestamp 1698431365
transform 1 0 8736 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__B
timestamp 1698431365
transform 1 0 8288 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__A1
timestamp 1698431365
transform -1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__A2
timestamp 1698431365
transform -1 0 7168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__A2
timestamp 1698431365
transform 1 0 9632 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__B
timestamp 1698431365
transform 1 0 8848 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1544__A1
timestamp 1698431365
transform -1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1544__A2
timestamp 1698431365
transform 1 0 6832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__A2
timestamp 1698431365
transform 1 0 12992 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__B
timestamp 1698431365
transform 1 0 14000 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A1
timestamp 1698431365
transform 1 0 11424 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A2
timestamp 1698431365
transform 1 0 12432 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__A2
timestamp 1698431365
transform 1 0 6608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__B
timestamp 1698431365
transform -1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A1
timestamp 1698431365
transform -1 0 3696 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A2
timestamp 1698431365
transform -1 0 4816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__A2
timestamp 1698431365
transform 1 0 12768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__B
timestamp 1698431365
transform 1 0 12320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__A1
timestamp 1698431365
transform -1 0 10304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__A2
timestamp 1698431365
transform 1 0 11200 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A2
timestamp 1698431365
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__B
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A1
timestamp 1698431365
transform 1 0 13552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A2
timestamp 1698431365
transform 1 0 14112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__A2
timestamp 1698431365
transform 1 0 9296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__B
timestamp 1698431365
transform 1 0 9632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1554__A1
timestamp 1698431365
transform 1 0 6384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1554__A2
timestamp 1698431365
transform 1 0 6832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A2
timestamp 1698431365
transform -1 0 6160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__B
timestamp 1698431365
transform 1 0 6384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A1
timestamp 1698431365
transform 1 0 5712 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A2
timestamp 1698431365
transform -1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A2
timestamp 1698431365
transform 1 0 24192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__B
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__A1
timestamp 1698431365
transform 1 0 24640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__A2
timestamp 1698431365
transform 1 0 22512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A2
timestamp 1698431365
transform 1 0 27328 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__B
timestamp 1698431365
transform 1 0 25088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__A1
timestamp 1698431365
transform -1 0 23968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__A2
timestamp 1698431365
transform 1 0 24640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A2
timestamp 1698431365
transform 1 0 24752 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__B
timestamp 1698431365
transform 1 0 25200 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A1
timestamp 1698431365
transform 1 0 23408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A2
timestamp 1698431365
transform 1 0 26544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__A2
timestamp 1698431365
transform 1 0 19264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__B
timestamp 1698431365
transform 1 0 18816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__A1
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__A2
timestamp 1698431365
transform 1 0 18480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__A2
timestamp 1698431365
transform 1 0 24528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__B
timestamp 1698431365
transform -1 0 24640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A1
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A2
timestamp 1698431365
transform 1 0 27888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__A2
timestamp 1698431365
transform 1 0 27216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__B
timestamp 1698431365
transform 1 0 26208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A1
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A2
timestamp 1698431365
transform 1 0 27328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__A2
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__B
timestamp 1698431365
transform 1 0 24864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__A1
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__A2
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A2
timestamp 1698431365
transform 1 0 24192 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__B
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1572__A1
timestamp 1698431365
transform 1 0 23632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1572__A2
timestamp 1698431365
transform 1 0 25312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__A2
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__B
timestamp 1698431365
transform 1 0 24640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A1
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A2
timestamp 1698431365
transform 1 0 25088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__A2
timestamp 1698431365
transform 1 0 23520 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__B
timestamp 1698431365
transform 1 0 23968 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1698431365
transform 1 0 22736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1698431365
transform 1 0 22848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A2
timestamp 1698431365
transform -1 0 4368 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__A1
timestamp 1698431365
transform -1 0 3136 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__B
timestamp 1698431365
transform -1 0 4816 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A1
timestamp 1698431365
transform 1 0 6160 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A2
timestamp 1698431365
transform 1 0 6608 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A1
timestamp 1698431365
transform -1 0 4592 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A1
timestamp 1698431365
transform -1 0 3920 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A2
timestamp 1698431365
transform 1 0 4368 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__B
timestamp 1698431365
transform 1 0 4144 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__B
timestamp 1698431365
transform 1 0 4592 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__A1
timestamp 1698431365
transform -1 0 3808 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1585__B
timestamp 1698431365
transform 1 0 4928 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__A1
timestamp 1698431365
transform -1 0 4592 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__A1
timestamp 1698431365
transform -1 0 2576 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A1
timestamp 1698431365
transform -1 0 6944 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__A1
timestamp 1698431365
transform 1 0 7168 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__A1
timestamp 1698431365
transform 1 0 5712 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1591__A1
timestamp 1698431365
transform 1 0 4032 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A1
timestamp 1698431365
transform 1 0 5376 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__A1
timestamp 1698431365
transform 1 0 22736 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__B
timestamp 1698431365
transform 1 0 26656 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__B
timestamp 1698431365
transform 1 0 25312 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__A1
timestamp 1698431365
transform 1 0 26208 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A1
timestamp 1698431365
transform 1 0 27328 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1698431365
transform -1 0 24192 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__A1
timestamp 1698431365
transform 1 0 25984 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__I
timestamp 1698431365
transform 1 0 26992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__I
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A2
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__I
timestamp 1698431365
transform 1 0 5712 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A1
timestamp 1698431365
transform 1 0 19040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A2
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__C
timestamp 1698431365
transform 1 0 18592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__A2
timestamp 1698431365
transform 1 0 15008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A1
timestamp 1698431365
transform 1 0 12432 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A2
timestamp 1698431365
transform 1 0 15456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__C
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A1
timestamp 1698431365
transform 1 0 28000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A2
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A1
timestamp 1698431365
transform 1 0 21840 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A2
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__C
timestamp 1698431365
transform 1 0 22288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A2
timestamp 1698431365
transform 1 0 19264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A1
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A2
timestamp 1698431365
transform 1 0 19712 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__C
timestamp 1698431365
transform 1 0 16352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__A2
timestamp 1698431365
transform 1 0 22624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A1
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A2
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__C
timestamp 1698431365
transform 1 0 17920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A2
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A1
timestamp 1698431365
transform 1 0 15344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__C
timestamp 1698431365
transform 1 0 15680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A2
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A1
timestamp 1698431365
transform 1 0 21840 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A2
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__C
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__A2
timestamp 1698431365
transform 1 0 16016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A1
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A2
timestamp 1698431365
transform 1 0 15680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__C
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1637__I
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1638__A2
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A1
timestamp 1698431365
transform 1 0 6608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A2
timestamp 1698431365
transform 1 0 7952 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__C
timestamp 1698431365
transform 1 0 6160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__A2
timestamp 1698431365
transform 1 0 10976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A1
timestamp 1698431365
transform 1 0 8624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A2
timestamp 1698431365
transform 1 0 10416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__C
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A2
timestamp 1698431365
transform 1 0 8848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A1
timestamp 1698431365
transform 1 0 6160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A2
timestamp 1698431365
transform 1 0 7728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__C
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A1
timestamp 1698431365
transform 1 0 13328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A2
timestamp 1698431365
transform 1 0 11872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A2
timestamp 1698431365
transform 1 0 11424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__C
timestamp 1698431365
transform 1 0 9968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A2
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__I
timestamp 1698431365
transform 1 0 18144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A1
timestamp 1698431365
transform 1 0 7728 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A2
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__C
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A2
timestamp 1698431365
transform 1 0 16128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A1
timestamp 1698431365
transform 1 0 12544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A2
timestamp 1698431365
transform 1 0 15680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__C
timestamp 1698431365
transform 1 0 15232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__A2
timestamp 1698431365
transform 1 0 12544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A1
timestamp 1698431365
transform 1 0 10976 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A2
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__C
timestamp 1698431365
transform 1 0 12096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A2
timestamp 1698431365
transform 1 0 13552 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A1
timestamp 1698431365
transform -1 0 11424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A2
timestamp 1698431365
transform 1 0 12768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__C
timestamp 1698431365
transform 1 0 12320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A2
timestamp 1698431365
transform 1 0 10080 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A1
timestamp 1698431365
transform -1 0 7840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A2
timestamp 1698431365
transform 1 0 8064 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__C
timestamp 1698431365
transform 1 0 8512 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__A2
timestamp 1698431365
transform -1 0 7616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A1
timestamp 1698431365
transform 1 0 6832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A2
timestamp 1698431365
transform 1 0 7840 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__C
timestamp 1698431365
transform 1 0 8960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A2
timestamp 1698431365
transform 1 0 19264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A1
timestamp 1698431365
transform -1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A2
timestamp 1698431365
transform 1 0 18592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__C
timestamp 1698431365
transform 1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A2
timestamp 1698431365
transform 1 0 13888 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A1
timestamp 1698431365
transform -1 0 14000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A2
timestamp 1698431365
transform 1 0 15792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__C
timestamp 1698431365
transform 1 0 15344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A2
timestamp 1698431365
transform 1 0 24080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A2
timestamp 1698431365
transform 1 0 23632 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__C
timestamp 1698431365
transform 1 0 22960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A2
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform -1 0 16128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1698431365
transform 1 0 16688 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__C
timestamp 1698431365
transform 1 0 16912 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__A2
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A1
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A2
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__C
timestamp 1698431365
transform 1 0 24416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A2
timestamp 1698431365
transform 1 0 27888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1698431365
transform -1 0 26320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A2
timestamp 1698431365
transform 1 0 27776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__C
timestamp 1698431365
transform 1 0 25648 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__A2
timestamp 1698431365
transform 1 0 28112 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A1
timestamp 1698431365
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A2
timestamp 1698431365
transform 1 0 27104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__C
timestamp 1698431365
transform 1 0 26208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__A2
timestamp 1698431365
transform 1 0 15568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A1
timestamp 1698431365
transform -1 0 12656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A2
timestamp 1698431365
transform -1 0 13888 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__C
timestamp 1698431365
transform 1 0 14112 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A2
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__A1
timestamp 1698431365
transform -1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__A2
timestamp 1698431365
transform 1 0 27552 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__C
timestamp 1698431365
transform 1 0 26432 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A2
timestamp 1698431365
transform -1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1698431365
transform 1 0 27552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A2
timestamp 1698431365
transform -1 0 27664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__C
timestamp 1698431365
transform -1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A2
timestamp 1698431365
transform 1 0 27664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A1
timestamp 1698431365
transform -1 0 25088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A2
timestamp 1698431365
transform 1 0 23968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__C
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A2
timestamp 1698431365
transform 1 0 27104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A1
timestamp 1698431365
transform -1 0 25760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A2
timestamp 1698431365
transform 1 0 27552 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__C
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A2
timestamp 1698431365
transform 1 0 27440 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1698431365
transform -1 0 25760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A2
timestamp 1698431365
transform 1 0 27776 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__C
timestamp 1698431365
transform 1 0 18032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A2
timestamp 1698431365
transform 1 0 22736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A1
timestamp 1698431365
transform -1 0 22512 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A2
timestamp 1698431365
transform 1 0 23296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__C
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__I
timestamp 1698431365
transform 1 0 8624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__I
timestamp 1698431365
transform 1 0 3808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__I
timestamp 1698431365
transform 1 0 5040 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__A2
timestamp 1698431365
transform -1 0 6160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__I
timestamp 1698431365
transform 1 0 4368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A2
timestamp 1698431365
transform 1 0 6608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__C
timestamp 1698431365
transform -1 0 5936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__I
timestamp 1698431365
transform -1 0 2128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A2
timestamp 1698431365
transform -1 0 2128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A2
timestamp 1698431365
transform -1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__C
timestamp 1698431365
transform 1 0 5488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__I
timestamp 1698431365
transform -1 0 5264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A2
timestamp 1698431365
transform 1 0 4032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A2
timestamp 1698431365
transform 1 0 2800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__C
timestamp 1698431365
transform 1 0 3360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__I
timestamp 1698431365
transform -1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A2
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A2
timestamp 1698431365
transform -1 0 5936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__C
timestamp 1698431365
transform 1 0 6160 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__I
timestamp 1698431365
transform -1 0 2352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__A2
timestamp 1698431365
transform 1 0 3024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A2
timestamp 1698431365
transform 1 0 3920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__C
timestamp 1698431365
transform 1 0 3472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__I
timestamp 1698431365
transform 1 0 3696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A2
timestamp 1698431365
transform 1 0 3248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A2
timestamp 1698431365
transform 1 0 4144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__C
timestamp 1698431365
transform 1 0 3696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__I
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A2
timestamp 1698431365
transform 1 0 2352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__A2
timestamp 1698431365
transform 1 0 5376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__C
timestamp 1698431365
transform 1 0 4928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__I
timestamp 1698431365
transform 1 0 5488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__A2
timestamp 1698431365
transform 1 0 3920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__A2
timestamp 1698431365
transform 1 0 4368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__C
timestamp 1698431365
transform 1 0 3920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__I
timestamp 1698431365
transform 1 0 4032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__I
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__A2
timestamp 1698431365
transform -1 0 2352 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A2
timestamp 1698431365
transform 1 0 2688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__C
timestamp 1698431365
transform 1 0 2016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__I
timestamp 1698431365
transform 1 0 6608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A2
timestamp 1698431365
transform 1 0 5040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A2
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__C
timestamp 1698431365
transform 1 0 4592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A2
timestamp 1698431365
transform 1 0 2576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A2
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__C
timestamp 1698431365
transform -1 0 2128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A2
timestamp 1698431365
transform 1 0 3024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__A2
timestamp 1698431365
transform 1 0 3920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__C
timestamp 1698431365
transform 1 0 3472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__A2
timestamp 1698431365
transform 1 0 3696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A2
timestamp 1698431365
transform 1 0 4368 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__C
timestamp 1698431365
transform 1 0 3920 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A2
timestamp 1698431365
transform -1 0 2128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A2
timestamp 1698431365
transform 1 0 2352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__C
timestamp 1698431365
transform 1 0 4368 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A2
timestamp 1698431365
transform 1 0 3808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A2
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__C
timestamp 1698431365
transform 1 0 2016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__A2
timestamp 1698431365
transform 1 0 3920 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A2
timestamp 1698431365
transform 1 0 4368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__C
timestamp 1698431365
transform 1 0 3920 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A2
timestamp 1698431365
transform 1 0 4256 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A2
timestamp 1698431365
transform 1 0 4816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__C
timestamp 1698431365
transform 1 0 4368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__A2
timestamp 1698431365
transform 1 0 3584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__A2
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__C
timestamp 1698431365
transform 1 0 5040 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A2
timestamp 1698431365
transform 1 0 2912 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__A2
timestamp 1698431365
transform 1 0 3808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__C
timestamp 1698431365
transform 1 0 3360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A2
timestamp 1698431365
transform 1 0 2016 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__A2
timestamp 1698431365
transform 1 0 3472 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__C
timestamp 1698431365
transform 1 0 3696 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__I
timestamp 1698431365
transform 1 0 4032 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__A2
timestamp 1698431365
transform 1 0 2240 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__I
timestamp 1698431365
transform -1 0 2912 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A2
timestamp 1698431365
transform 1 0 3696 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__C
timestamp 1698431365
transform -1 0 4704 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A2
timestamp 1698431365
transform -1 0 2128 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__A2
timestamp 1698431365
transform 1 0 2800 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__C
timestamp 1698431365
transform 1 0 4144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A2
timestamp 1698431365
transform 1 0 4592 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A2
timestamp 1698431365
transform 1 0 4144 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__C
timestamp 1698431365
transform 1 0 3696 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__A2
timestamp 1698431365
transform 1 0 3808 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A2
timestamp 1698431365
transform 1 0 4368 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__C
timestamp 1698431365
transform 1 0 3920 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__I
timestamp 1698431365
transform 1 0 3920 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A2
timestamp 1698431365
transform 1 0 2576 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__A2
timestamp 1698431365
transform 1 0 3248 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__C
timestamp 1698431365
transform 1 0 4368 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__I
timestamp 1698431365
transform 1 0 3920 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A2
timestamp 1698431365
transform 1 0 2912 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A2
timestamp 1698431365
transform 1 0 3920 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__C
timestamp 1698431365
transform 1 0 3472 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__I
timestamp 1698431365
transform -1 0 4816 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__A2
timestamp 1698431365
transform 1 0 2240 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__A2
timestamp 1698431365
transform 1 0 4032 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__C
timestamp 1698431365
transform 1 0 3584 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__I
timestamp 1698431365
transform 1 0 4032 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A2
timestamp 1698431365
transform 1 0 2128 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__A2
timestamp 1698431365
transform 1 0 6384 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__C
timestamp 1698431365
transform 1 0 4032 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A2
timestamp 1698431365
transform 1 0 6496 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A2
timestamp 1698431365
transform 1 0 5040 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__C
timestamp 1698431365
transform 1 0 6832 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A2
timestamp 1698431365
transform -1 0 3920 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__A2
timestamp 1698431365
transform 1 0 2800 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__C
timestamp 1698431365
transform 1 0 3248 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__A1
timestamp 1698431365
transform 1 0 7728 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__A2
timestamp 1698431365
transform 1 0 8064 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__A2
timestamp 1698431365
transform 1 0 6608 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__C
timestamp 1698431365
transform 1 0 6160 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__A1
timestamp 1698431365
transform 1 0 5040 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__A2
timestamp 1698431365
transform 1 0 5712 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A2
timestamp 1698431365
transform -1 0 5488 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__C
timestamp 1698431365
transform 1 0 4144 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__I
timestamp 1698431365
transform 1 0 25984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__I
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A2
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__B
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A1
timestamp 1698431365
transform 1 0 20160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A2
timestamp 1698431365
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A2
timestamp 1698431365
transform -1 0 12656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__B
timestamp 1698431365
transform 1 0 12880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A1
timestamp 1698431365
transform 1 0 8960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A2
timestamp 1698431365
transform 1 0 11088 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A2
timestamp 1698431365
transform 1 0 21952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__B
timestamp 1698431365
transform 1 0 23184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A1
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A2
timestamp 1698431365
transform 1 0 20944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__A2
timestamp 1698431365
transform -1 0 18928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__B
timestamp 1698431365
transform -1 0 19376 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A1
timestamp 1698431365
transform -1 0 17024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A2
timestamp 1698431365
transform -1 0 17920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__A2
timestamp 1698431365
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__B
timestamp 1698431365
transform -1 0 17472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A1
timestamp 1698431365
transform -1 0 13440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A2
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__A2
timestamp 1698431365
transform 1 0 15232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__B
timestamp 1698431365
transform 1 0 15456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A1
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A2
timestamp 1698431365
transform 1 0 14336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A2
timestamp 1698431365
transform 1 0 14560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__B
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A1
timestamp 1698431365
transform 1 0 12432 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A2
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A2
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__B
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A1
timestamp 1698431365
transform -1 0 14672 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A2
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__I
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__A2
timestamp 1698431365
transform 1 0 24080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__B
timestamp 1698431365
transform 1 0 23632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__A1
timestamp 1698431365
transform -1 0 21840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__A2
timestamp 1698431365
transform 1 0 22960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__A2
timestamp 1698431365
transform 1 0 20160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__B
timestamp 1698431365
transform 1 0 19712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__A1
timestamp 1698431365
transform 1 0 17024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__A2
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__A2
timestamp 1698431365
transform -1 0 14784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__B
timestamp 1698431365
transform 1 0 12768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__A1
timestamp 1698431365
transform -1 0 12544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__A2
timestamp 1698431365
transform 1 0 14112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A2
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__B
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__A1
timestamp 1698431365
transform -1 0 9968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__A2
timestamp 1698431365
transform 1 0 10192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A2
timestamp 1698431365
transform 1 0 12880 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__B
timestamp 1698431365
transform 1 0 11200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__A1
timestamp 1698431365
transform 1 0 9744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__A2
timestamp 1698431365
transform 1 0 10864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__A2
timestamp 1698431365
transform 1 0 17472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__B
timestamp 1698431365
transform 1 0 17024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1698431365
transform 1 0 14224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A2
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A2
timestamp 1698431365
transform 1 0 14000 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__B
timestamp 1698431365
transform 1 0 12208 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__A1
timestamp 1698431365
transform -1 0 9744 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__A2
timestamp 1698431365
transform 1 0 9968 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__A2
timestamp 1698431365
transform 1 0 12432 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__B
timestamp 1698431365
transform 1 0 10976 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A1
timestamp 1698431365
transform 1 0 9856 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A2
timestamp 1698431365
transform 1 0 11200 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A2
timestamp 1698431365
transform 1 0 19824 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__B
timestamp 1698431365
transform 1 0 19376 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__A1
timestamp 1698431365
transform 1 0 18368 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__A2
timestamp 1698431365
transform -1 0 18592 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__A2
timestamp 1698431365
transform 1 0 15456 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__B
timestamp 1698431365
transform 1 0 15904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__A1
timestamp 1698431365
transform 1 0 13104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__A2
timestamp 1698431365
transform 1 0 14224 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A2
timestamp 1698431365
transform 1 0 10864 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__B
timestamp 1698431365
transform 1 0 10416 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A1
timestamp 1698431365
transform 1 0 8960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A2
timestamp 1698431365
transform 1 0 9744 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A2
timestamp 1698431365
transform -1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__B
timestamp 1698431365
transform -1 0 8736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A1
timestamp 1698431365
transform -1 0 7728 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A2
timestamp 1698431365
transform -1 0 8288 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__A2
timestamp 1698431365
transform 1 0 21168 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__B
timestamp 1698431365
transform 1 0 20720 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A1
timestamp 1698431365
transform -1 0 20496 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A2
timestamp 1698431365
transform 1 0 20720 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A2
timestamp 1698431365
transform 1 0 16800 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__B
timestamp 1698431365
transform 1 0 15904 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A1
timestamp 1698431365
transform 1 0 12768 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A2
timestamp 1698431365
transform 1 0 13216 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__A2
timestamp 1698431365
transform 1 0 26880 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__B
timestamp 1698431365
transform 1 0 26432 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A1
timestamp 1698431365
transform -1 0 26208 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A2
timestamp 1698431365
transform 1 0 27328 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A2
timestamp 1698431365
transform 1 0 27776 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__B
timestamp 1698431365
transform 1 0 27328 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A1
timestamp 1698431365
transform -1 0 25872 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A2
timestamp 1698431365
transform 1 0 27552 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A2
timestamp 1698431365
transform 1 0 27440 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__B
timestamp 1698431365
transform 1 0 28000 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A1
timestamp 1698431365
transform 1 0 27328 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A2
timestamp 1698431365
transform 1 0 27776 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A2
timestamp 1698431365
transform 1 0 16912 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__B
timestamp 1698431365
transform 1 0 17360 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A1
timestamp 1698431365
transform 1 0 14448 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A2
timestamp 1698431365
transform 1 0 14896 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A2
timestamp 1698431365
transform 1 0 28000 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__B
timestamp 1698431365
transform 1 0 26656 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__A1
timestamp 1698431365
transform 1 0 27552 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__A2
timestamp 1698431365
transform 1 0 28000 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__A2
timestamp 1698431365
transform -1 0 28112 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__B
timestamp 1698431365
transform 1 0 26768 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A1
timestamp 1698431365
transform -1 0 25536 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A2
timestamp 1698431365
transform 1 0 28000 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__A2
timestamp 1698431365
transform 1 0 25760 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__B
timestamp 1698431365
transform 1 0 25312 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A1
timestamp 1698431365
transform 1 0 27888 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A2
timestamp 1698431365
transform 1 0 26656 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__A2
timestamp 1698431365
transform 1 0 27440 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__B
timestamp 1698431365
transform 1 0 25648 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__A1
timestamp 1698431365
transform 1 0 25984 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__A2
timestamp 1698431365
transform 1 0 27104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A2
timestamp 1698431365
transform 1 0 25312 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__B
timestamp 1698431365
transform 1 0 24640 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A1
timestamp 1698431365
transform 1 0 26992 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A2
timestamp 1698431365
transform 1 0 26880 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A2
timestamp 1698431365
transform 1 0 24192 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__B
timestamp 1698431365
transform 1 0 24640 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A1
timestamp 1698431365
transform 1 0 23296 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A2
timestamp 1698431365
transform 1 0 25088 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A2
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__I
timestamp 1698431365
transform -1 0 3472 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A1
timestamp 1698431365
transform 1 0 20944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A2
timestamp 1698431365
transform 1 0 15904 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__A1
timestamp 1698431365
transform -1 0 14560 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__A2
timestamp 1698431365
transform 1 0 16352 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__I
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__I
timestamp 1698431365
transform 1 0 21392 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A2
timestamp 1698431365
transform 1 0 22176 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A1
timestamp 1698431365
transform 1 0 19936 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A2
timestamp 1698431365
transform 1 0 21392 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__C
timestamp 1698431365
transform 1 0 22288 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A2
timestamp 1698431365
transform 1 0 8960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A1
timestamp 1698431365
transform 1 0 6944 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A2
timestamp 1698431365
transform 1 0 7392 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__C
timestamp 1698431365
transform 1 0 7840 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__A2
timestamp 1698431365
transform 1 0 25088 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A1
timestamp 1698431365
transform 1 0 23632 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A2
timestamp 1698431365
transform 1 0 24640 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__C
timestamp 1698431365
transform 1 0 23520 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A2
timestamp 1698431365
transform 1 0 22064 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A1
timestamp 1698431365
transform 1 0 19264 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A2
timestamp 1698431365
transform 1 0 20608 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__C
timestamp 1698431365
transform 1 0 19712 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A2
timestamp 1698431365
transform 1 0 19152 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__A1
timestamp 1698431365
transform 1 0 17248 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__A2
timestamp 1698431365
transform 1 0 21840 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__C
timestamp 1698431365
transform 1 0 17472 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__A2
timestamp 1698431365
transform -1 0 17696 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__A1
timestamp 1698431365
transform -1 0 13104 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__A2
timestamp 1698431365
transform -1 0 13104 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__C
timestamp 1698431365
transform 1 0 13552 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__A2
timestamp 1698431365
transform 1 0 24192 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A1
timestamp 1698431365
transform 1 0 24080 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A2
timestamp 1698431365
transform 1 0 23296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__C
timestamp 1698431365
transform 1 0 22960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__A2
timestamp 1698431365
transform 1 0 24640 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__A1
timestamp 1698431365
transform -1 0 21392 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__A2
timestamp 1698431365
transform 1 0 21952 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__C
timestamp 1698431365
transform 1 0 20720 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__I
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__A2
timestamp 1698431365
transform 1 0 22288 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__I
timestamp 1698431365
transform 1 0 5040 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A1
timestamp 1698431365
transform 1 0 21392 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A2
timestamp 1698431365
transform 1 0 22512 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__C
timestamp 1698431365
transform 1 0 20720 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__A2
timestamp 1698431365
transform 1 0 22848 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__A1
timestamp 1698431365
transform -1 0 20048 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__A2
timestamp 1698431365
transform 1 0 20944 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__C
timestamp 1698431365
transform 1 0 19600 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A2
timestamp 1698431365
transform 1 0 10976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A1
timestamp 1698431365
transform 1 0 10640 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A2
timestamp 1698431365
transform 1 0 10528 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__C
timestamp 1698431365
transform 1 0 9632 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__A2
timestamp 1698431365
transform -1 0 3696 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A1
timestamp 1698431365
transform -1 0 2240 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A2
timestamp 1698431365
transform -1 0 2688 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__C
timestamp 1698431365
transform 1 0 3360 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A2
timestamp 1698431365
transform 1 0 9632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__A1
timestamp 1698431365
transform 1 0 6832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__A2
timestamp 1698431365
transform 1 0 6832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__C
timestamp 1698431365
transform 1 0 4368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__A2
timestamp 1698431365
transform 1 0 3920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__A1
timestamp 1698431365
transform -1 0 3696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__A2
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__C
timestamp 1698431365
transform -1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__A2
timestamp 1698431365
transform 1 0 8848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A1
timestamp 1698431365
transform -1 0 6384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A2
timestamp 1698431365
transform 1 0 6608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__C
timestamp 1698431365
transform 1 0 5712 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A2
timestamp 1698431365
transform 1 0 7280 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A1
timestamp 1698431365
transform -1 0 3136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A2
timestamp 1698431365
transform 1 0 3360 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__C
timestamp 1698431365
transform -1 0 2240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__A2
timestamp 1698431365
transform 1 0 8288 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A1
timestamp 1698431365
transform 1 0 6160 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A2
timestamp 1698431365
transform 1 0 7728 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__C
timestamp 1698431365
transform 1 0 5712 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__A2
timestamp 1698431365
transform 1 0 7056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__A1
timestamp 1698431365
transform 1 0 5936 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__A2
timestamp 1698431365
transform 1 0 7504 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__C
timestamp 1698431365
transform 1 0 5040 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__A2
timestamp 1698431365
transform 1 0 3584 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__A1
timestamp 1698431365
transform 1 0 4704 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__A2
timestamp 1698431365
transform -1 0 2688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__C
timestamp 1698431365
transform 1 0 4256 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A2
timestamp 1698431365
transform 1 0 4480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A1
timestamp 1698431365
transform -1 0 2128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A2
timestamp 1698431365
transform 1 0 2688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__C
timestamp 1698431365
transform 1 0 3136 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__A2
timestamp 1698431365
transform 1 0 6608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A1
timestamp 1698431365
transform -1 0 3920 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A2
timestamp 1698431365
transform 1 0 5712 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__C
timestamp 1698431365
transform 1 0 3248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A2
timestamp 1698431365
transform 1 0 21616 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1698431365
transform 1 0 22400 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A2
timestamp 1698431365
transform 1 0 22736 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__C
timestamp 1698431365
transform 1 0 21952 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__A2
timestamp 1698431365
transform 1 0 7504 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A1
timestamp 1698431365
transform 1 0 5040 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A2
timestamp 1698431365
transform 1 0 6608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__C
timestamp 1698431365
transform 1 0 4592 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A2
timestamp 1698431365
transform 1 0 19376 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__A1
timestamp 1698431365
transform 1 0 20048 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__A2
timestamp 1698431365
transform 1 0 20496 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__C
timestamp 1698431365
transform 1 0 19600 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__A2
timestamp 1698431365
transform 1 0 7504 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A1
timestamp 1698431365
transform -1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A2
timestamp 1698431365
transform 1 0 7952 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__C
timestamp 1698431365
transform 1 0 4592 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A2
timestamp 1698431365
transform 1 0 8064 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__A1
timestamp 1698431365
transform 1 0 5040 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__A2
timestamp 1698431365
transform 1 0 6720 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__C
timestamp 1698431365
transform 1 0 4592 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A2
timestamp 1698431365
transform 1 0 7504 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A1
timestamp 1698431365
transform 1 0 5264 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A2
timestamp 1698431365
transform 1 0 7168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__C
timestamp 1698431365
transform 1 0 4816 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__A2
timestamp 1698431365
transform -1 0 6384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A1
timestamp 1698431365
transform 1 0 5264 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A2
timestamp 1698431365
transform 1 0 5712 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__C
timestamp 1698431365
transform -1 0 6160 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__A2
timestamp 1698431365
transform -1 0 22064 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A1
timestamp 1698431365
transform 1 0 20160 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A2
timestamp 1698431365
transform 1 0 20608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__C
timestamp 1698431365
transform 1 0 19712 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__A2
timestamp 1698431365
transform 1 0 21840 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A1
timestamp 1698431365
transform 1 0 20608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A2
timestamp 1698431365
transform 1 0 21952 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__C
timestamp 1698431365
transform 1 0 21504 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A2
timestamp 1698431365
transform 1 0 28112 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A1
timestamp 1698431365
transform 1 0 24640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A2
timestamp 1698431365
transform -1 0 23744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__C
timestamp 1698431365
transform 1 0 27104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__A2
timestamp 1698431365
transform 1 0 26544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__A1
timestamp 1698431365
transform 1 0 25648 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__A2
timestamp 1698431365
transform 1 0 25312 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__C
timestamp 1698431365
transform 1 0 25200 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__A1
timestamp 1698431365
transform 1 0 22400 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__A2
timestamp 1698431365
transform 1 0 23072 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1939__A2
timestamp 1698431365
transform 1 0 2464 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1939__B1
timestamp 1698431365
transform -1 0 3136 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__A1
timestamp 1698431365
transform 1 0 2464 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__A2
timestamp 1698431365
transform -1 0 2016 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__B
timestamp 1698431365
transform 1 0 5712 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__B
timestamp 1698431365
transform 1 0 2800 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A2
timestamp 1698431365
transform 1 0 2352 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__B
timestamp 1698431365
transform 1 0 6496 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__B
timestamp 1698431365
transform 1 0 2128 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A2
timestamp 1698431365
transform 1 0 2576 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__B
timestamp 1698431365
transform 1 0 23184 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A2
timestamp 1698431365
transform -1 0 2688 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__B
timestamp 1698431365
transform -1 0 2240 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__A2
timestamp 1698431365
transform 1 0 2912 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__B
timestamp 1698431365
transform -1 0 18256 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A2
timestamp 1698431365
transform -1 0 2688 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__B
timestamp 1698431365
transform -1 0 2240 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__A2
timestamp 1698431365
transform 1 0 5152 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__B1
timestamp 1698431365
transform 1 0 8064 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1954__A1
timestamp 1698431365
transform 1 0 4704 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__A2
timestamp 1698431365
transform 1 0 2800 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__B1
timestamp 1698431365
transform 1 0 4704 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__A1
timestamp 1698431365
transform 1 0 3808 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__A2
timestamp 1698431365
transform -1 0 5264 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__B1
timestamp 1698431365
transform 1 0 7504 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1958__A1
timestamp 1698431365
transform 1 0 5712 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A2
timestamp 1698431365
transform 1 0 15232 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A1
timestamp 1698431365
transform -1 0 9184 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A2
timestamp 1698431365
transform -1 0 16352 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__A2
timestamp 1698431365
transform 1 0 8960 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__A1
timestamp 1698431365
transform -1 0 7616 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__A2
timestamp 1698431365
transform -1 0 8512 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1963__A2
timestamp 1698431365
transform 1 0 10752 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A1
timestamp 1698431365
transform 1 0 10192 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A2
timestamp 1698431365
transform 1 0 10304 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__A2
timestamp 1698431365
transform 1 0 2800 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__A3
timestamp 1698431365
transform -1 0 4144 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__A1
timestamp 1698431365
transform 1 0 7280 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__B
timestamp 1698431365
transform -1 0 7168 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A1
timestamp 1698431365
transform -1 0 7056 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A1
timestamp 1698431365
transform -1 0 12768 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__B
timestamp 1698431365
transform 1 0 11424 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A1
timestamp 1698431365
transform -1 0 8736 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A1
timestamp 1698431365
transform -1 0 7840 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__B
timestamp 1698431365
transform 1 0 9520 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A1
timestamp 1698431365
transform 1 0 7168 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A1
timestamp 1698431365
transform 1 0 8064 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__B
timestamp 1698431365
transform 1 0 9744 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A1
timestamp 1698431365
transform -1 0 7840 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A1
timestamp 1698431365
transform 1 0 7728 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__B
timestamp 1698431365
transform 1 0 7840 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__A1
timestamp 1698431365
transform 1 0 6496 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__B
timestamp 1698431365
transform -1 0 7616 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__A1
timestamp 1698431365
transform -1 0 4144 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__A1
timestamp 1698431365
transform -1 0 6608 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__CLK
timestamp 1698431365
transform 1 0 23072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__CLK
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__CLK
timestamp 1698431365
transform 1 0 26096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__CLK
timestamp 1698431365
transform 1 0 18368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__CLK
timestamp 1698431365
transform 1 0 9632 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__CLK
timestamp 1698431365
transform 1 0 11648 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__CLK
timestamp 1698431365
transform 1 0 26208 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__CLK
timestamp 1698431365
transform 1 0 7952 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__CLK
timestamp 1698431365
transform 1 0 8512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__CLK
timestamp 1698431365
transform -1 0 6272 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__CLK
timestamp 1698431365
transform 1 0 18144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__CLK
timestamp 1698431365
transform 1 0 14448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1999__CLK
timestamp 1698431365
transform 1 0 16352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__CLK
timestamp 1698431365
transform 1 0 17024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__CLK
timestamp 1698431365
transform 1 0 24864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__CLK
timestamp 1698431365
transform 1 0 21840 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__CLK
timestamp 1698431365
transform 1 0 28112 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__CLK
timestamp 1698431365
transform 1 0 24304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__CLK
timestamp 1698431365
transform 1 0 28112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__CLK
timestamp 1698431365
transform 1 0 25984 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__CLK
timestamp 1698431365
transform 1 0 27664 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__CLK
timestamp 1698431365
transform 1 0 28000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__CLK
timestamp 1698431365
transform 1 0 8960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__CLK
timestamp 1698431365
transform 1 0 11200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__CLK
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__CLK
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__CLK
timestamp 1698431365
transform 1 0 26544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__CLK
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__CLK
timestamp 1698431365
transform 1 0 26544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__CLK
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__CLK
timestamp 1698431365
transform 1 0 15680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__CLK
timestamp 1698431365
transform 1 0 11536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__CLK
timestamp 1698431365
transform 1 0 9856 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2027__CLK
timestamp 1698431365
transform 1 0 8960 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__CLK
timestamp 1698431365
transform 1 0 7840 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__CLK
timestamp 1698431365
transform 1 0 7728 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__CLK
timestamp 1698431365
transform 1 0 13552 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__CLK
timestamp 1698431365
transform 1 0 6160 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__CLK
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2033__CLK
timestamp 1698431365
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2034__CLK
timestamp 1698431365
transform 1 0 5824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__CLK
timestamp 1698431365
transform 1 0 5152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__CLK
timestamp 1698431365
transform -1 0 27216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__CLK
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__CLK
timestamp 1698431365
transform 1 0 27664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__CLK
timestamp 1698431365
transform -1 0 19936 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__CLK
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__CLK
timestamp 1698431365
transform 1 0 28112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__CLK
timestamp 1698431365
transform 1 0 27328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__CLK
timestamp 1698431365
transform 1 0 27104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__CLK
timestamp 1698431365
transform 1 0 26768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__CLK
timestamp 1698431365
transform -1 0 23968 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__CLK
timestamp 1698431365
transform 1 0 4480 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__CLK
timestamp 1698431365
transform 1 0 5040 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__CLK
timestamp 1698431365
transform 1 0 6048 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__CLK
timestamp 1698431365
transform 1 0 5040 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__CLK
timestamp 1698431365
transform 1 0 4592 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2051__CLK
timestamp 1698431365
transform 1 0 4816 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__CLK
timestamp 1698431365
transform 1 0 8064 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__CLK
timestamp 1698431365
transform 1 0 5040 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2054__CLK
timestamp 1698431365
transform -1 0 24192 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2060__CLK
timestamp 1698431365
transform -1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__CLK
timestamp 1698431365
transform 1 0 14896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__CLK
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__CLK
timestamp 1698431365
transform 1 0 19712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__CLK
timestamp 1698431365
transform 1 0 22176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__CLK
timestamp 1698431365
transform 1 0 18928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2066__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2067__CLK
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2068__CLK
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2069__CLK
timestamp 1698431365
transform 1 0 12880 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__CLK
timestamp 1698431365
transform 1 0 8176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__CLK
timestamp 1698431365
transform 1 0 8624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__CLK
timestamp 1698431365
transform 1 0 10416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__CLK
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__CLK
timestamp 1698431365
transform 1 0 11984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__CLK
timestamp 1698431365
transform 1 0 13552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__CLK
timestamp 1698431365
transform -1 0 10976 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__CLK
timestamp 1698431365
transform 1 0 9520 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__CLK
timestamp 1698431365
transform 1 0 19824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__CLK
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__CLK
timestamp 1698431365
transform 1 0 25648 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2081__CLK
timestamp 1698431365
transform 1 0 19824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__CLK
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__CLK
timestamp 1698431365
transform 1 0 16240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__CLK
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__CLK
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__CLK
timestamp 1698431365
transform -1 0 18368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__CLK
timestamp 1698431365
transform 1 0 28112 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__CLK
timestamp 1698431365
transform 1 0 24192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2092__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__CLK
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__CLK
timestamp 1698431365
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__CLK
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__CLK
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2101__CLK
timestamp 1698431365
transform 1 0 7728 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__CLK
timestamp 1698431365
transform 1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__CLK
timestamp 1698431365
transform 1 0 7392 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2105__CLK
timestamp 1698431365
transform 1 0 4816 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2106__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2107__CLK
timestamp 1698431365
transform 1 0 5488 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__CLK
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2109__CLK
timestamp 1698431365
transform 1 0 7168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2111__CLK
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__CLK
timestamp 1698431365
transform 1 0 5040 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__CLK
timestamp 1698431365
transform 1 0 5040 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__CLK
timestamp 1698431365
transform 1 0 5040 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__CLK
timestamp 1698431365
transform 1 0 4144 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__CLK
timestamp 1698431365
transform 1 0 4816 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2120__CLK
timestamp 1698431365
transform 1 0 8288 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__CLK
timestamp 1698431365
transform 1 0 4592 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__CLK
timestamp 1698431365
transform -1 0 7168 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__CLK
timestamp 1698431365
transform 1 0 7280 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__CLK
timestamp 1698431365
transform 1 0 19264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__CLK
timestamp 1698431365
transform 1 0 11536 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__CLK
timestamp 1698431365
transform -1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__CLK
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__CLK
timestamp 1698431365
transform 1 0 13552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__CLK
timestamp 1698431365
transform 1 0 15008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__CLK
timestamp 1698431365
transform 1 0 14112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__CLK
timestamp 1698431365
transform 1 0 13216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__CLK
timestamp 1698431365
transform 1 0 23520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2133__CLK
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2134__CLK
timestamp 1698431365
transform 1 0 18144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2135__CLK
timestamp 1698431365
transform 1 0 12768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__CLK
timestamp 1698431365
transform 1 0 16576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__CLK
timestamp 1698431365
transform 1 0 12656 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__CLK
timestamp 1698431365
transform 1 0 20272 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2141__CLK
timestamp 1698431365
transform 1 0 16800 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__CLK
timestamp 1698431365
transform 1 0 11984 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__CLK
timestamp 1698431365
transform 1 0 10192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2144__CLK
timestamp 1698431365
transform 1 0 21392 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__CLK
timestamp 1698431365
transform 1 0 16800 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2146__CLK
timestamp 1698431365
transform 1 0 28112 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2148__CLK
timestamp 1698431365
transform 1 0 28112 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__CLK
timestamp 1698431365
transform 1 0 13552 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__CLK
timestamp 1698431365
transform 1 0 24192 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2152__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__CLK
timestamp 1698431365
transform 1 0 28112 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__CLK
timestamp 1698431365
transform 1 0 28112 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__CLK
timestamp 1698431365
transform 1 0 13888 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__CLK
timestamp 1698431365
transform 1 0 22624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2159__CLK
timestamp 1698431365
transform -1 0 9184 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__CLK
timestamp 1698431365
transform 1 0 28000 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2161__CLK
timestamp 1698431365
transform 1 0 14448 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2162__CLK
timestamp 1698431365
transform 1 0 23744 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__CLK
timestamp 1698431365
transform 1 0 11536 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2164__CLK
timestamp 1698431365
transform 1 0 27440 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2165__CLK
timestamp 1698431365
transform 1 0 24416 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__CLK
timestamp 1698431365
transform 1 0 23968 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__CLK
timestamp 1698431365
transform 1 0 24416 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2168__CLK
timestamp 1698431365
transform 1 0 13552 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__CLK
timestamp 1698431365
transform 1 0 5040 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__CLK
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__CLK
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__CLK
timestamp 1698431365
transform 1 0 5824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__CLK
timestamp 1698431365
transform 1 0 5824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__CLK
timestamp 1698431365
transform 1 0 8960 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2175__CLK
timestamp 1698431365
transform -1 0 7280 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__CLK
timestamp 1698431365
transform 1 0 2464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__CLK
timestamp 1698431365
transform 1 0 4032 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2178__CLK
timestamp 1698431365
transform 1 0 3808 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2180__CLK
timestamp 1698431365
transform 1 0 7952 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__CLK
timestamp 1698431365
transform 1 0 22400 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__CLK
timestamp 1698431365
transform 1 0 7616 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__CLK
timestamp 1698431365
transform 1 0 8288 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__CLK
timestamp 1698431365
transform 1 0 5712 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__CLK
timestamp 1698431365
transform 1 0 5264 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__CLK
timestamp 1698431365
transform 1 0 21392 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__CLK
timestamp 1698431365
transform 1 0 22288 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__CLK
timestamp 1698431365
transform 1 0 28112 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__CLK
timestamp 1698431365
transform 1 0 27664 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__CLK
timestamp 1698431365
transform 1 0 2800 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__CLK
timestamp 1698431365
transform 1 0 3248 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2192__CLK
timestamp 1698431365
transform 1 0 2576 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__CLK
timestamp 1698431365
transform 1 0 3024 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__CLK
timestamp 1698431365
transform 1 0 3248 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__CLK
timestamp 1698431365
transform 1 0 5600 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__CLK
timestamp 1698431365
transform -1 0 5376 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2197__CLK
timestamp 1698431365
transform -1 0 7392 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2198__CLK
timestamp 1698431365
transform 1 0 9744 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2199__CLK
timestamp 1698431365
transform 1 0 10640 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__CLK
timestamp 1698431365
transform 1 0 9856 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__CLK
timestamp 1698431365
transform 1 0 6048 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__CLK
timestamp 1698431365
transform 1 0 9968 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__CLK
timestamp 1698431365
transform 1 0 5712 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2204__CLK
timestamp 1698431365
transform 1 0 11088 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2205__CLK
timestamp 1698431365
transform 1 0 10192 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2206__CLK
timestamp 1698431365
transform 1 0 6944 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 10640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_clk_I
timestamp 1698431365
transform -1 0 19600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_clk_I
timestamp 1698431365
transform 1 0 21056 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_clk_I
timestamp 1698431365
transform 1 0 10752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_clk_I
timestamp 1698431365
transform 1 0 6048 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_clk_I
timestamp 1698431365
transform 1 0 12656 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_clk_I
timestamp 1698431365
transform 1 0 12880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_clk_I
timestamp 1698431365
transform 1 0 8848 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_clk_I
timestamp 1698431365
transform 1 0 5040 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_clk_I
timestamp 1698431365
transform -1 0 8288 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_clk_I
timestamp 1698431365
transform 1 0 20160 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_clk_I
timestamp 1698431365
transform 1 0 17472 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_clk_I
timestamp 1698431365
transform 1 0 22512 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_clk_I
timestamp 1698431365
transform 1 0 23408 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_clk_I
timestamp 1698431365
transform 1 0 20944 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_clk_I
timestamp 1698431365
transform 1 0 23296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_clk_I
timestamp 1698431365
transform 1 0 23968 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_clk_I
timestamp 1698431365
transform 1 0 20272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_clk_I
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_clk_I
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_clk_I
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_clk_I
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_clk_I
timestamp 1698431365
transform -1 0 7616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._078__A1
timestamp 1698431365
transform 1 0 28112 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 26880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 18368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 17920 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 16352 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 16800 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 15568 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 14896 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 13552 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 13664 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 14112 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 12208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 27776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 13552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 10752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 9184 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 8736 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 8288 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 7840 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 7504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 6832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 26432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 2464 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 26880 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 28112 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 18816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 25984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 19040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 27328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 1792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 1792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 2464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform 1 0 2240 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 1792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 2128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform 1 0 2464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform 1 0 2464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform 1 0 1792 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform 1 0 2464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform 1 0 2464 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform 1 0 2464 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform 1 0 1792 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform 1 0 1792 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform 1 0 3024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform 1 0 1792 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform 1 0 2240 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform 1 0 1792 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform 1 0 2464 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform 1 0 2464 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform 1 0 4368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform 1 0 2464 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform 1 0 1792 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform 1 0 1792 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform 1 0 1792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform 1 0 1792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform 1 0 4368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform 1 0 2912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform 1 0 27776 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform 1 0 27328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform -1 0 2016 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac._4__I
timestamp 1698431365
transform 1 0 25312 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac._5__A2
timestamp 1698431365
transform 1 0 26208 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 20160 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 21504 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 23632 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 25984 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._4__A2
timestamp 1698431365
transform -1 0 15456 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 18928 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 19376 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 20608 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 21840 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._4__A2
timestamp 1698431365
transform -1 0 15904 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._5__A1
timestamp 1698431365
transform -1 0 13776 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 16128 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 16576 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 16576 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 16576 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 16352 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._4__A2
timestamp 1698431365
transform -1 0 16800 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._5__A1
timestamp 1698431365
transform -1 0 12432 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 13552 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 16352 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 16128 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 16240 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 16352 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref_I
timestamp 1698431365
transform 1 0 16800 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref_I
timestamp 1698431365
transform 1 0 13552 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref_I
timestamp 1698431365
transform 1 0 13776 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref_I
timestamp 1698431365
transform 1 0 12656 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._3__I
timestamp 1698431365
transform 1 0 25312 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A1
timestamp 1698431365
transform -1 0 20048 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A2
timestamp 1698431365
transform -1 0 19600 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 24976 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 22400 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 22624 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 22624 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 19824 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 23968 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref_I
timestamp 1698431365
transform 1 0 24080 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref_I
timestamp 1698431365
transform 1 0 19824 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref_I
timestamp 1698431365
transform 1 0 20832 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref_I
timestamp 1698431365
transform 1 0 20272 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref_I
timestamp 1698431365
transform 1 0 19824 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref_I
timestamp 1698431365
transform 1 0 21840 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref_I
timestamp 1698431365
transform 1 0 19264 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref_I
timestamp 1698431365
transform 1 0 21392 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref_I
timestamp 1698431365
transform 1 0 20720 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref_I
timestamp 1698431365
transform 1 0 22624 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref_I
timestamp 1698431365
transform 1 0 18480 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref_I
timestamp 1698431365
transform 1 0 22624 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.vdac_single.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 26656 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dcdc_EN
timestamp 1698431365
transform 1 0 8064 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_wire4_I
timestamp 1698431365
transform 1 0 5600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0551_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7504 0 1 98784
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0553_
timestamp 1698431365
transform 1 0 9744 0 -1 89376
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0889_
timestamp 1698431365
transform 1 0 11424 0 -1 101920
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0902_
timestamp 1698431365
transform -1 0 23296 0 -1 101920
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk
timestamp 1698431365
transform 1 0 14224 0 1 54880
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_net81
timestamp 1698431365
transform 1 0 13328 0 1 100352
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_temp1.i_precharge_n
timestamp 1698431365
transform 1 0 11424 0 -1 105056
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0551_
timestamp 1698431365
transform -1 0 11872 0 1 95648
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0553_
timestamp 1698431365
transform -1 0 15008 0 -1 86240
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0889_
timestamp 1698431365
transform 1 0 13328 0 1 98784
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0902_
timestamp 1698431365
transform 1 0 17248 0 -1 100352
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 18928 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_net81
timestamp 1698431365
transform -1 0 16800 0 -1 98784
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_temp1.i_precharge_n
timestamp 1698431365
transform -1 0 15680 0 -1 106624
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0551_
timestamp 1698431365
transform 1 0 11424 0 -1 100352
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0553_
timestamp 1698431365
transform 1 0 10864 0 -1 92512
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0889_
timestamp 1698431365
transform 1 0 14000 0 1 101920
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0902_
timestamp 1698431365
transform 1 0 19264 0 -1 105056
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 14112 0 1 76832
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_net81
timestamp 1698431365
transform 1 0 14224 0 1 105056
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_temp1.i_precharge_n
timestamp 1698431365
transform 1 0 15344 0 1 103488
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1698431365
transform 1 0 3584 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1698431365
transform 1 0 3248 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1698431365
transform -1 0 15008 0 -1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1698431365
transform 1 0 7056 0 1 65856
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1698431365
transform -1 0 8848 0 -1 70560
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1698431365
transform 1 0 3584 0 -1 92512
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1698431365
transform 1 0 7504 0 1 97216
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1698431365
transform 1 0 11424 0 -1 78400
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1698431365
transform 1 0 17920 0 -1 86240
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1698431365
transform 1 0 22736 0 1 98784
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1698431365
transform 1 0 22736 0 1 65856
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1698431365
transform 1 0 22736 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1698431365
transform 1 0 14336 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1698431365
transform 1 0 11424 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1698431365
transform -1 0 7504 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  dec1._049_
timestamp 1698431365
transform -1 0 27440 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._050_
timestamp 1698431365
transform 1 0 23744 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  dec1._051_
timestamp 1698431365
transform 1 0 20160 0 -1 83104
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  dec1._052_
timestamp 1698431365
transform 1 0 18704 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._053_
timestamp 1698431365
transform 1 0 19712 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._054_
timestamp 1698431365
transform 1 0 21952 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._055_
timestamp 1698431365
transform 1 0 21168 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  dec1._056_
timestamp 1698431365
transform 1 0 21616 0 -1 84672
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  dec1._057_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._058_
timestamp 1698431365
transform 1 0 21168 0 1 81536
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  dec1._059_
timestamp 1698431365
transform 1 0 21616 0 1 84672
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._060_
timestamp 1698431365
transform 1 0 23632 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._061_
timestamp 1698431365
transform -1 0 20944 0 1 84672
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._062_
timestamp 1698431365
transform 1 0 22960 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  dec1._063_
timestamp 1698431365
transform 1 0 24304 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  dec1._064_
timestamp 1698431365
transform -1 0 20944 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  dec1._065_
timestamp 1698431365
transform -1 0 24080 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  dec1._066_
timestamp 1698431365
transform 1 0 24304 0 1 81536
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  dec1._067_
timestamp 1698431365
transform 1 0 23296 0 -1 84672
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  dec1._068_
timestamp 1698431365
transform 1 0 23856 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  dec1._069_
timestamp 1698431365
transform 1 0 25088 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._070_
timestamp 1698431365
transform 1 0 25424 0 1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._071_
timestamp 1698431365
transform 1 0 24304 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  dec1._072_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 81536
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  dec1._073_
timestamp 1698431365
transform -1 0 28112 0 1 84672
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  dec1._074_
timestamp 1698431365
transform 1 0 25088 0 -1 84672
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  dec1._075_
timestamp 1698431365
transform 1 0 25200 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  dec1._076_
timestamp 1698431365
transform 1 0 25648 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  dec1._077_
timestamp 1698431365
transform 1 0 25872 0 1 84672
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  dec1._078_
timestamp 1698431365
transform -1 0 28336 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._079_
timestamp 1698431365
transform 1 0 19040 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  dec1._080_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24416 0 1 87808
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._081_
timestamp 1698431365
transform 1 0 26096 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._082_
timestamp 1698431365
transform 1 0 26208 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  dec1._083_
timestamp 1698431365
transform -1 0 23184 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  dec1._084_
timestamp 1698431365
transform 1 0 26880 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  dec1._085_
timestamp 1698431365
transform 1 0 26880 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  dec1._086_
timestamp 1698431365
transform 1 0 27104 0 1 81536
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._087_
timestamp 1698431365
transform -1 0 28336 0 -1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  dec1._088_
timestamp 1698431365
transform 1 0 25424 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  dec1._089_
timestamp 1698431365
transform 1 0 27104 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  dec1._090_
timestamp 1698431365
transform 1 0 23744 0 -1 87808
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  dec1._091_
timestamp 1698431365
transform 1 0 24752 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._092_
timestamp 1698431365
transform -1 0 24976 0 1 84672
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._093_
timestamp 1698431365
transform -1 0 24864 0 -1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  dec1._094_
timestamp 1698431365
transform 1 0 25312 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  dec1._095_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28336 0 1 86240
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  dec1._096_
timestamp 1698431365
transform -1 0 25872 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._097_
timestamp 1698431365
transform -1 0 27776 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  dec1._098_
timestamp 1698431365
transform -1 0 27328 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._099_
timestamp 1698431365
transform 1 0 26992 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  dec1._100_
timestamp 1698431365
transform 1 0 26544 0 -1 87808
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._101_
timestamp 1698431365
transform 1 0 26096 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_6
timestamp 1698431365
transform 1 0 2016 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_106 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13216 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_133
timestamp 1698431365
transform 1 0 16240 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_222
timestamp 1698431365
transform 1 0 26208 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_10
timestamp 1698431365
transform 1 0 2464 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_52 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_58
timestamp 1698431365
transform 1 0 7840 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_62
timestamp 1698431365
transform 1 0 8288 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_97
timestamp 1698431365
transform 1 0 12208 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_108
timestamp 1698431365
transform 1 0 13440 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_112
timestamp 1698431365
transform 1 0 13888 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_116
timestamp 1698431365
transform 1 0 14336 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_118
timestamp 1698431365
transform 1 0 14560 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_121
timestamp 1698431365
transform 1 0 14896 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_127
timestamp 1698431365
transform 1 0 15568 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_131
timestamp 1698431365
transform 1 0 16016 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_134
timestamp 1698431365
transform 1 0 16352 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_138
timestamp 1698431365
transform 1 0 16800 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_237
timestamp 1698431365
transform 1 0 27888 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_18
timestamp 1698431365
transform 1 0 3360 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_26
timestamp 1698431365
transform 1 0 4256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_30
timestamp 1698431365
transform 1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_42
timestamp 1698431365
transform 1 0 6048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_46
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_48
timestamp 1698431365
transform 1 0 6720 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_51
timestamp 1698431365
transform 1 0 7056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_111
timestamp 1698431365
transform 1 0 13776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_119
timestamp 1698431365
transform 1 0 14672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_121
timestamp 1698431365
transform 1 0 14896 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_227
timestamp 1698431365
transform 1 0 26768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_235
timestamp 1698431365
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_239
timestamp 1698431365
transform 1 0 28112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_80
timestamp 1698431365
transform 1 0 10304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_86
timestamp 1698431365
transform 1 0 10976 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_95
timestamp 1698431365
transform 1 0 11984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_99 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_131
timestamp 1698431365
transform 1 0 16016 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_165
timestamp 1698431365
transform 1 0 19824 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_226
timestamp 1698431365
transform 1 0 26656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_230
timestamp 1698431365
transform 1 0 27104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_234
timestamp 1698431365
transform 1 0 27552 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_238
timestamp 1698431365
transform 1 0 28000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_240
timestamp 1698431365
transform 1 0 28224 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_8
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_28
timestamp 1698431365
transform 1 0 4480 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_139
timestamp 1698431365
transform 1 0 16912 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_147
timestamp 1698431365
transform 1 0 17808 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_151
timestamp 1698431365
transform 1 0 18256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_153
timestamp 1698431365
transform 1 0 18480 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_156
timestamp 1698431365
transform 1 0 18816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_160
timestamp 1698431365
transform 1 0 19264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_162
timestamp 1698431365
transform 1 0 19488 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_183
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_185
timestamp 1698431365
transform 1 0 22064 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_218
timestamp 1698431365
transform 1 0 25760 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_226
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_230
timestamp 1698431365
transform 1 0 27104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_234
timestamp 1698431365
transform 1 0 27552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_238
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_240
timestamp 1698431365
transform 1 0 28224 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_18
timestamp 1698431365
transform 1 0 3360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_26
timestamp 1698431365
transform 1 0 4256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_30
timestamp 1698431365
transform 1 0 4704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_32
timestamp 1698431365
transform 1 0 4928 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_35
timestamp 1698431365
transform 1 0 5264 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_41
timestamp 1698431365
transform 1 0 5936 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_57
timestamp 1698431365
transform 1 0 7728 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_65
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_152
timestamp 1698431365
transform 1 0 18368 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_238
timestamp 1698431365
transform 1 0 28000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_240
timestamp 1698431365
transform 1 0 28224 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_12
timestamp 1698431365
transform 1 0 2688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_16
timestamp 1698431365
transform 1 0 3136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_20
timestamp 1698431365
transform 1 0 3584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_24
timestamp 1698431365
transform 1 0 4032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_26
timestamp 1698431365
transform 1 0 4256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_33
timestamp 1698431365
transform 1 0 5040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_45
timestamp 1698431365
transform 1 0 6384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_49
timestamp 1698431365
transform 1 0 6832 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_81
timestamp 1698431365
transform 1 0 10416 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_97
timestamp 1698431365
transform 1 0 12208 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_123
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_127
timestamp 1698431365
transform 1 0 15568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_129
timestamp 1698431365
transform 1 0 15792 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_217
timestamp 1698431365
transform 1 0 25648 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_233
timestamp 1698431365
transform 1 0 27440 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_8
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_12
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_39
timestamp 1698431365
transform 1 0 5712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_76
timestamp 1698431365
transform 1 0 9856 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_108
timestamp 1698431365
transform 1 0 13440 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_204
timestamp 1698431365
transform 1 0 24192 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_208
timestamp 1698431365
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_228
timestamp 1698431365
transform 1 0 26880 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_236
timestamp 1698431365
transform 1 0 27776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_240
timestamp 1698431365
transform 1 0 28224 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_63
timestamp 1698431365
transform 1 0 8400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_67
timestamp 1698431365
transform 1 0 8848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_99
timestamp 1698431365
transform 1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_136
timestamp 1698431365
transform 1 0 16576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_140
timestamp 1698431365
transform 1 0 17024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_144
timestamp 1698431365
transform 1 0 17472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_148
timestamp 1698431365
transform 1 0 17920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_152
timestamp 1698431365
transform 1 0 18368 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_154
timestamp 1698431365
transform 1 0 18592 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_157
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_161
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_183
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_218
timestamp 1698431365
transform 1 0 25760 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_234
timestamp 1698431365
transform 1 0 27552 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_238
timestamp 1698431365
transform 1 0 28000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_22
timestamp 1698431365
transform 1 0 3808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_24
timestamp 1698431365
transform 1 0 4032 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_35
timestamp 1698431365
transform 1 0 5264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_39
timestamp 1698431365
transform 1 0 5712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_51
timestamp 1698431365
transform 1 0 7056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_53
timestamp 1698431365
transform 1 0 7280 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_64
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_96
timestamp 1698431365
transform 1 0 12096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_100
timestamp 1698431365
transform 1 0 12544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_112
timestamp 1698431365
transform 1 0 13888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_116
timestamp 1698431365
transform 1 0 14336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_120
timestamp 1698431365
transform 1 0 14784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_124
timestamp 1698431365
transform 1 0 15232 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_134
timestamp 1698431365
transform 1 0 16352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_155
timestamp 1698431365
transform 1 0 18704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_159
timestamp 1698431365
transform 1 0 19152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_163
timestamp 1698431365
transform 1 0 19600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_167
timestamp 1698431365
transform 1 0 20048 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_177
timestamp 1698431365
transform 1 0 21168 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_193
timestamp 1698431365
transform 1 0 22960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_195
timestamp 1698431365
transform 1 0 23184 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_228
timestamp 1698431365
transform 1 0 26880 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_236
timestamp 1698431365
transform 1 0 27776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_240
timestamp 1698431365
transform 1 0 28224 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_68
timestamp 1698431365
transform 1 0 8960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_72
timestamp 1698431365
transform 1 0 9408 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_136
timestamp 1698431365
transform 1 0 16576 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_145
timestamp 1698431365
transform 1 0 17584 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_181
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_183
timestamp 1698431365
transform 1 0 21840 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_186
timestamp 1698431365
transform 1 0 22176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_214
timestamp 1698431365
transform 1 0 25312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_218
timestamp 1698431365
transform 1 0 25760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_222
timestamp 1698431365
transform 1 0 26208 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_238
timestamp 1698431365
transform 1 0 28000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_240
timestamp 1698431365
transform 1 0 28224 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_4
timestamp 1698431365
transform 1 0 1792 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_74
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_77
timestamp 1698431365
transform 1 0 9968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_89
timestamp 1698431365
transform 1 0 11312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_99
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_101
timestamp 1698431365
transform 1 0 12656 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_104
timestamp 1698431365
transform 1 0 12992 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_184
timestamp 1698431365
transform 1 0 21952 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_193
timestamp 1698431365
transform 1 0 22960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_197
timestamp 1698431365
transform 1 0 23408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_201
timestamp 1698431365
transform 1 0 23856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_205
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_238
timestamp 1698431365
transform 1 0 28000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_240
timestamp 1698431365
transform 1 0 28224 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_4
timestamp 1698431365
transform 1 0 1792 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_49
timestamp 1698431365
transform 1 0 6832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_86
timestamp 1698431365
transform 1 0 10976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_90
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_94
timestamp 1698431365
transform 1 0 11872 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_97
timestamp 1698431365
transform 1 0 12208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_161
timestamp 1698431365
transform 1 0 19376 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_206
timestamp 1698431365
transform 1 0 24416 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_233
timestamp 1698431365
transform 1 0 27440 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_20
timestamp 1698431365
transform 1 0 3584 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_55
timestamp 1698431365
transform 1 0 7504 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_59
timestamp 1698431365
transform 1 0 7952 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_62
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_92
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_96
timestamp 1698431365
transform 1 0 12096 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_104
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_108
timestamp 1698431365
transform 1 0 13440 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_118
timestamp 1698431365
transform 1 0 14560 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_126
timestamp 1698431365
transform 1 0 15456 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_148
timestamp 1698431365
transform 1 0 17920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_152
timestamp 1698431365
transform 1 0 18368 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_169
timestamp 1698431365
transform 1 0 20272 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_173
timestamp 1698431365
transform 1 0 20720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_177
timestamp 1698431365
transform 1 0 21168 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_191
timestamp 1698431365
transform 1 0 22736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_195
timestamp 1698431365
transform 1 0 23184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_197
timestamp 1698431365
transform 1 0 23408 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_200
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_204
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_238
timestamp 1698431365
transform 1 0 28000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_240
timestamp 1698431365
transform 1 0 28224 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_57
timestamp 1698431365
transform 1 0 7728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_59
timestamp 1698431365
transform 1 0 7952 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_62
timestamp 1698431365
transform 1 0 8288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_66
timestamp 1698431365
transform 1 0 8736 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_70
timestamp 1698431365
transform 1 0 9184 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_81
timestamp 1698431365
transform 1 0 10416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_83
timestamp 1698431365
transform 1 0 10640 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_86
timestamp 1698431365
transform 1 0 10976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_88
timestamp 1698431365
transform 1 0 11200 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_91
timestamp 1698431365
transform 1 0 11536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_95
timestamp 1698431365
transform 1 0 11984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_99
timestamp 1698431365
transform 1 0 12432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_123
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_158
timestamp 1698431365
transform 1 0 19040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_162
timestamp 1698431365
transform 1 0 19488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_166
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_170
timestamp 1698431365
transform 1 0 20384 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_219
timestamp 1698431365
transform 1 0 25872 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_223
timestamp 1698431365
transform 1 0 26320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_227
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_231
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_6
timestamp 1698431365
transform 1 0 2016 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_15
timestamp 1698431365
transform 1 0 3024 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_20
timestamp 1698431365
transform 1 0 3584 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_24
timestamp 1698431365
transform 1 0 4032 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_56
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_89
timestamp 1698431365
transform 1 0 11312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_122
timestamp 1698431365
transform 1 0 15008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_126
timestamp 1698431365
transform 1 0 15456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_130
timestamp 1698431365
transform 1 0 15904 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_156
timestamp 1698431365
transform 1 0 18816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_160
timestamp 1698431365
transform 1 0 19264 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_164
timestamp 1698431365
transform 1 0 19712 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_166
timestamp 1698431365
transform 1 0 19936 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_196
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_200
timestamp 1698431365
transform 1 0 23744 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_224
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_228
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_232
timestamp 1698431365
transform 1 0 27328 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_240
timestamp 1698431365
transform 1 0 28224 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_4
timestamp 1698431365
transform 1 0 1792 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_17
timestamp 1698431365
transform 1 0 3248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_27
timestamp 1698431365
transform 1 0 4368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_137
timestamp 1698431365
transform 1 0 16688 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1698431365
transform 1 0 22288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_219
timestamp 1698431365
transform 1 0 25872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_223
timestamp 1698431365
transform 1 0 26320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_227
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_231
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_237
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_6
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_17
timestamp 1698431365
transform 1 0 3248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_21
timestamp 1698431365
transform 1 0 3696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_25
timestamp 1698431365
transform 1 0 4144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_29
timestamp 1698431365
transform 1 0 4592 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_37
timestamp 1698431365
transform 1 0 5488 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_40
timestamp 1698431365
transform 1 0 5824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_44
timestamp 1698431365
transform 1 0 6272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_64
timestamp 1698431365
transform 1 0 8512 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_101
timestamp 1698431365
transform 1 0 12656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_103
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_130
timestamp 1698431365
transform 1 0 15904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_134
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_162
timestamp 1698431365
transform 1 0 19488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_166
timestamp 1698431365
transform 1 0 19936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_170
timestamp 1698431365
transform 1 0 20384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_176
timestamp 1698431365
transform 1 0 21056 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_179
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_191
timestamp 1698431365
transform 1 0 22736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_193
timestamp 1698431365
transform 1 0 22960 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_238
timestamp 1698431365
transform 1 0 28000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_240
timestamp 1698431365
transform 1 0 28224 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_19
timestamp 1698431365
transform 1 0 3472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_23
timestamp 1698431365
transform 1 0 3920 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_27
timestamp 1698431365
transform 1 0 4368 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_109
timestamp 1698431365
transform 1 0 13552 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_112
timestamp 1698431365
transform 1 0 13888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_116
timestamp 1698431365
transform 1 0 14336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_120
timestamp 1698431365
transform 1 0 14784 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_150
timestamp 1698431365
transform 1 0 18144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_154
timestamp 1698431365
transform 1 0 18592 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_162
timestamp 1698431365
transform 1 0 19488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_166
timestamp 1698431365
transform 1 0 19936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_168
timestamp 1698431365
transform 1 0 20160 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_227
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_231
timestamp 1698431365
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_235
timestamp 1698431365
transform 1 0 27664 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_31
timestamp 1698431365
transform 1 0 4816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_35
timestamp 1698431365
transform 1 0 5264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_37
timestamp 1698431365
transform 1 0 5488 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_40
timestamp 1698431365
transform 1 0 5824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_52
timestamp 1698431365
transform 1 0 7168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_54
timestamp 1698431365
transform 1 0 7392 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_63
timestamp 1698431365
transform 1 0 8400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_82
timestamp 1698431365
transform 1 0 10528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_86
timestamp 1698431365
transform 1 0 10976 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_90
timestamp 1698431365
transform 1 0 11424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_123
timestamp 1698431365
transform 1 0 15120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_127
timestamp 1698431365
transform 1 0 15568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_131
timestamp 1698431365
transform 1 0 16016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_135
timestamp 1698431365
transform 1 0 16464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_147
timestamp 1698431365
transform 1 0 17808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_151
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_163
timestamp 1698431365
transform 1 0 19600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_167
timestamp 1698431365
transform 1 0 20048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_171
timestamp 1698431365
transform 1 0 20496 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_175
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_184
timestamp 1698431365
transform 1 0 21952 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_188
timestamp 1698431365
transform 1 0 22400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_192
timestamp 1698431365
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_196
timestamp 1698431365
transform 1 0 23296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_200
timestamp 1698431365
transform 1 0 23744 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698431365
transform 1 0 25312 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_10
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_21
timestamp 1698431365
transform 1 0 3696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_23
timestamp 1698431365
transform 1 0 3920 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_66
timestamp 1698431365
transform 1 0 8736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_70
timestamp 1698431365
transform 1 0 9184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_74
timestamp 1698431365
transform 1 0 9632 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_88
timestamp 1698431365
transform 1 0 11200 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_97
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_109
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698431365
transform 1 0 15568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_145
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_16
timestamp 1698431365
transform 1 0 3136 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_19
timestamp 1698431365
transform 1 0 3472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_23
timestamp 1698431365
transform 1 0 3920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_31
timestamp 1698431365
transform 1 0 4816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_62
timestamp 1698431365
transform 1 0 8288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_228
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_232
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_236
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_240
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_41
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_52
timestamp 1698431365
transform 1 0 7168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_62
timestamp 1698431365
transform 1 0 8288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_64
timestamp 1698431365
transform 1 0 8512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_96
timestamp 1698431365
transform 1 0 12096 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_98
timestamp 1698431365
transform 1 0 12320 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_115
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_133
timestamp 1698431365
transform 1 0 16240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_137
timestamp 1698431365
transform 1 0 16688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_139
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_142
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_146
timestamp 1698431365
transform 1 0 17696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_148
timestamp 1698431365
transform 1 0 17920 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_155
timestamp 1698431365
transform 1 0 18704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_159
timestamp 1698431365
transform 1 0 19152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_169
timestamp 1698431365
transform 1 0 20272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_188
timestamp 1698431365
transform 1 0 22400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_192
timestamp 1698431365
transform 1 0 22848 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_222
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_226
timestamp 1698431365
transform 1 0 26656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_230
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_234
timestamp 1698431365
transform 1 0 27552 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_19
timestamp 1698431365
transform 1 0 3472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_21
timestamp 1698431365
transform 1 0 3696 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_30
timestamp 1698431365
transform 1 0 4704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_34
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_38
timestamp 1698431365
transform 1 0 5600 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_46
timestamp 1698431365
transform 1 0 6496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_50
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_54
timestamp 1698431365
transform 1 0 7392 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_76
timestamp 1698431365
transform 1 0 9856 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_79
timestamp 1698431365
transform 1 0 10192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_83
timestamp 1698431365
transform 1 0 10640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_87
timestamp 1698431365
transform 1 0 11088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_89
timestamp 1698431365
transform 1 0 11312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_92
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_125
timestamp 1698431365
transform 1 0 15344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_127
timestamp 1698431365
transform 1 0 15568 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_192
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_196
timestamp 1698431365
transform 1 0 23296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_200
timestamp 1698431365
transform 1 0 23744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_204
timestamp 1698431365
transform 1 0 24192 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_6
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_21
timestamp 1698431365
transform 1 0 3696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_25
timestamp 1698431365
transform 1 0 4144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_29
timestamp 1698431365
transform 1 0 4592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_33
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_41
timestamp 1698431365
transform 1 0 5936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_55
timestamp 1698431365
transform 1 0 7504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_59
timestamp 1698431365
transform 1 0 7952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_63
timestamp 1698431365
transform 1 0 8400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_67
timestamp 1698431365
transform 1 0 8848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_97
timestamp 1698431365
transform 1 0 12208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_117
timestamp 1698431365
transform 1 0 14448 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_187
timestamp 1698431365
transform 1 0 22288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_227
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_235
timestamp 1698431365
transform 1 0 27664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_21
timestamp 1698431365
transform 1 0 3696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_25
timestamp 1698431365
transform 1 0 4144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_29
timestamp 1698431365
transform 1 0 4592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_31
timestamp 1698431365
transform 1 0 4816 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_101
timestamp 1698431365
transform 1 0 12656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_105
timestamp 1698431365
transform 1 0 13104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_109
timestamp 1698431365
transform 1 0 13552 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_113
timestamp 1698431365
transform 1 0 14000 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_120
timestamp 1698431365
transform 1 0 14784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_124
timestamp 1698431365
transform 1 0 15232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_128
timestamp 1698431365
transform 1 0 15680 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698431365
transform 1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_154
timestamp 1698431365
transform 1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_187
timestamp 1698431365
transform 1 0 22288 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_214
timestamp 1698431365
transform 1 0 25312 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_57
timestamp 1698431365
transform 1 0 7728 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_61
timestamp 1698431365
transform 1 0 8176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_65
timestamp 1698431365
transform 1 0 8624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_69
timestamp 1698431365
transform 1 0 9072 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_77
timestamp 1698431365
transform 1 0 9968 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_84
timestamp 1698431365
transform 1 0 10752 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_88
timestamp 1698431365
transform 1 0 11200 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_96
timestamp 1698431365
transform 1 0 12096 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_100
timestamp 1698431365
transform 1 0 12544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_102
timestamp 1698431365
transform 1 0 12768 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_111
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_119
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_125
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_134
timestamp 1698431365
transform 1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_138
timestamp 1698431365
transform 1 0 16800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_142
timestamp 1698431365
transform 1 0 17248 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_146
timestamp 1698431365
transform 1 0 17696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_152
timestamp 1698431365
transform 1 0 18368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_156
timestamp 1698431365
transform 1 0 18816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_160
timestamp 1698431365
transform 1 0 19264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_205
timestamp 1698431365
transform 1 0 24304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_24
timestamp 1698431365
transform 1 0 4032 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_26
timestamp 1698431365
transform 1 0 4256 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_35
timestamp 1698431365
transform 1 0 5264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_39
timestamp 1698431365
transform 1 0 5712 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_45
timestamp 1698431365
transform 1 0 6384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_59
timestamp 1698431365
transform 1 0 7952 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_87
timestamp 1698431365
transform 1 0 11088 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_91
timestamp 1698431365
transform 1 0 11536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_93
timestamp 1698431365
transform 1 0 11760 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_103
timestamp 1698431365
transform 1 0 12880 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_146
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_156
timestamp 1698431365
transform 1 0 18816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_160
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_164
timestamp 1698431365
transform 1 0 19712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_168
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_175
timestamp 1698431365
transform 1 0 20944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_179
timestamp 1698431365
transform 1 0 21392 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_70
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_74
timestamp 1698431365
transform 1 0 9632 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_85
timestamp 1698431365
transform 1 0 10864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_87
timestamp 1698431365
transform 1 0 11088 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698431365
transform 1 0 14224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_125
timestamp 1698431365
transform 1 0 15344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_146
timestamp 1698431365
transform 1 0 17696 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_154
timestamp 1698431365
transform 1 0 18592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_158
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_166
timestamp 1698431365
transform 1 0 19936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_170
timestamp 1698431365
transform 1 0 20384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_193
timestamp 1698431365
transform 1 0 22960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_197
timestamp 1698431365
transform 1 0 23408 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_201
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_204
timestamp 1698431365
transform 1 0 24192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_208
timestamp 1698431365
transform 1 0 24640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_212
timestamp 1698431365
transform 1 0 25088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_216
timestamp 1698431365
transform 1 0 25536 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_218
timestamp 1698431365
transform 1 0 25760 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_229
timestamp 1698431365
transform 1 0 26992 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_233
timestamp 1698431365
transform 1 0 27440 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_237
timestamp 1698431365
transform 1 0 27888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_22
timestamp 1698431365
transform 1 0 3808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_55
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_59
timestamp 1698431365
transform 1 0 7952 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_101
timestamp 1698431365
transform 1 0 12656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_105
timestamp 1698431365
transform 1 0 13104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_109
timestamp 1698431365
transform 1 0 13552 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_113
timestamp 1698431365
transform 1 0 14000 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_117
timestamp 1698431365
transform 1 0 14448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_121
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_125
timestamp 1698431365
transform 1 0 15344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_150
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_183
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_195
timestamp 1698431365
transform 1 0 23184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_199
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_203
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_224
timestamp 1698431365
transform 1 0 26432 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_230
timestamp 1698431365
transform 1 0 27104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_234
timestamp 1698431365
transform 1 0 27552 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_238
timestamp 1698431365
transform 1 0 28000 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_6
timestamp 1698431365
transform 1 0 2016 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_15
timestamp 1698431365
transform 1 0 3024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_17
timestamp 1698431365
transform 1 0 3248 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_47
timestamp 1698431365
transform 1 0 6608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_79
timestamp 1698431365
transform 1 0 10192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_83
timestamp 1698431365
transform 1 0 10640 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_99
timestamp 1698431365
transform 1 0 12432 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698431365
transform 1 0 14000 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_119
timestamp 1698431365
transform 1 0 14672 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_123
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_127
timestamp 1698431365
transform 1 0 15568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_158
timestamp 1698431365
transform 1 0 19040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_162
timestamp 1698431365
transform 1 0 19488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_166
timestamp 1698431365
transform 1 0 19936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_170
timestamp 1698431365
transform 1 0 20384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_179
timestamp 1698431365
transform 1 0 21392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_82
timestamp 1698431365
transform 1 0 10528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_86
timestamp 1698431365
transform 1 0 10976 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_94
timestamp 1698431365
transform 1 0 11872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_98
timestamp 1698431365
transform 1 0 12320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_109
timestamp 1698431365
transform 1 0 13552 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_111
timestamp 1698431365
transform 1 0 13776 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_122
timestamp 1698431365
transform 1 0 15008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_126
timestamp 1698431365
transform 1 0 15456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_130
timestamp 1698431365
transform 1 0 15904 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_158
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_162
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_166
timestamp 1698431365
transform 1 0 19936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_170
timestamp 1698431365
transform 1 0 20384 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_185
timestamp 1698431365
transform 1 0 22064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_195
timestamp 1698431365
transform 1 0 23184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_199
timestamp 1698431365
transform 1 0 23632 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_203
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_224
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_230
timestamp 1698431365
transform 1 0 27104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_234
timestamp 1698431365
transform 1 0 27552 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_238
timestamp 1698431365
transform 1 0 28000 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_16
timestamp 1698431365
transform 1 0 3136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_20
timestamp 1698431365
transform 1 0 3584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_24
timestamp 1698431365
transform 1 0 4032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_55
timestamp 1698431365
transform 1 0 7504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_69
timestamp 1698431365
transform 1 0 9072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_71
timestamp 1698431365
transform 1 0 9296 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_136
timestamp 1698431365
transform 1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_140
timestamp 1698431365
transform 1 0 17024 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_148
timestamp 1698431365
transform 1 0 17920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_152
timestamp 1698431365
transform 1 0 18368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_156
timestamp 1698431365
transform 1 0 18816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_160
timestamp 1698431365
transform 1 0 19264 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_203
timestamp 1698431365
transform 1 0 24080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_205
timestamp 1698431365
transform 1 0 24304 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_208
timestamp 1698431365
transform 1 0 24640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_31
timestamp 1698431365
transform 1 0 4816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_35
timestamp 1698431365
transform 1 0 5264 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_43
timestamp 1698431365
transform 1 0 6160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_49
timestamp 1698431365
transform 1 0 6832 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_65
timestamp 1698431365
transform 1 0 8624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_67
timestamp 1698431365
transform 1 0 8848 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_96
timestamp 1698431365
transform 1 0 12096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_100
timestamp 1698431365
transform 1 0 12544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_104
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_112
timestamp 1698431365
transform 1 0 13888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_116
timestamp 1698431365
transform 1 0 14336 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_126
timestamp 1698431365
transform 1 0 15456 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_130
timestamp 1698431365
transform 1 0 15904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_134
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_154
timestamp 1698431365
transform 1 0 18592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_158
timestamp 1698431365
transform 1 0 19040 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_200
timestamp 1698431365
transform 1 0 23744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_204
timestamp 1698431365
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_234
timestamp 1698431365
transform 1 0 27552 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_238
timestamp 1698431365
transform 1 0 28000 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_240
timestamp 1698431365
transform 1 0 28224 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_43
timestamp 1698431365
transform 1 0 6160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_47
timestamp 1698431365
transform 1 0 6608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_51
timestamp 1698431365
transform 1 0 7056 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_55
timestamp 1698431365
transform 1 0 7504 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_87
timestamp 1698431365
transform 1 0 11088 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_90
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_94
timestamp 1698431365
transform 1 0 11872 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_98
timestamp 1698431365
transform 1 0 12320 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_125
timestamp 1698431365
transform 1 0 15344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_129
timestamp 1698431365
transform 1 0 15792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_133
timestamp 1698431365
transform 1 0 16240 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_227
timestamp 1698431365
transform 1 0 26768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_231
timestamp 1698431365
transform 1 0 27216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_235
timestamp 1698431365
transform 1 0 27664 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_8
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_92
timestamp 1698431365
transform 1 0 11648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_96
timestamp 1698431365
transform 1 0 12096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_100
timestamp 1698431365
transform 1 0 12544 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_130
timestamp 1698431365
transform 1 0 15904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_134
timestamp 1698431365
transform 1 0 16352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_138
timestamp 1698431365
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_158
timestamp 1698431365
transform 1 0 19040 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_162
timestamp 1698431365
transform 1 0 19488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_177
timestamp 1698431365
transform 1 0 21168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_4
timestamp 1698431365
transform 1 0 1792 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_17
timestamp 1698431365
transform 1 0 3248 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_21
timestamp 1698431365
transform 1 0 3696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_25
timestamp 1698431365
transform 1 0 4144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_47
timestamp 1698431365
transform 1 0 6608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_67
timestamp 1698431365
transform 1 0 8848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_88
timestamp 1698431365
transform 1 0 11200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_92
timestamp 1698431365
transform 1 0 11648 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_94
timestamp 1698431365
transform 1 0 11872 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_97
timestamp 1698431365
transform 1 0 12208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_109
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_112
timestamp 1698431365
transform 1 0 13888 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_154
timestamp 1698431365
transform 1 0 18592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_158
timestamp 1698431365
transform 1 0 19040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_162
timestamp 1698431365
transform 1 0 19488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_166
timestamp 1698431365
transform 1 0 19936 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_181
timestamp 1698431365
transform 1 0 21616 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_31
timestamp 1698431365
transform 1 0 4816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_35
timestamp 1698431365
transform 1 0 5264 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_41
timestamp 1698431365
transform 1 0 5936 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_45
timestamp 1698431365
transform 1 0 6384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_65
timestamp 1698431365
transform 1 0 8624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_74
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_77
timestamp 1698431365
transform 1 0 9968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_110
timestamp 1698431365
transform 1 0 13664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_122
timestamp 1698431365
transform 1 0 15008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_124
timestamp 1698431365
transform 1 0 15232 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_132
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_153
timestamp 1698431365
transform 1 0 18480 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_159
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_163
timestamp 1698431365
transform 1 0 19600 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_201
timestamp 1698431365
transform 1 0 23856 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_216
timestamp 1698431365
transform 1 0 25536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_232
timestamp 1698431365
transform 1 0 27328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_236
timestamp 1698431365
transform 1 0 27776 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_238
timestamp 1698431365
transform 1 0 28000 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_15
timestamp 1698431365
transform 1 0 3024 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_20
timestamp 1698431365
transform 1 0 3584 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_22
timestamp 1698431365
transform 1 0 3808 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_39
timestamp 1698431365
transform 1 0 5712 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_71
timestamp 1698431365
transform 1 0 9296 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_81
timestamp 1698431365
transform 1 0 10416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_85
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_157
timestamp 1698431365
transform 1 0 18928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_190
timestamp 1698431365
transform 1 0 22624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_200
timestamp 1698431365
transform 1 0 23744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_206
timestamp 1698431365
transform 1 0 24416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_210
timestamp 1698431365
transform 1 0 24864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_6
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_10
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_13
timestamp 1698431365
transform 1 0 2800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_17
timestamp 1698431365
transform 1 0 3248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_21
timestamp 1698431365
transform 1 0 3696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_25
timestamp 1698431365
transform 1 0 4144 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_57
timestamp 1698431365
transform 1 0 7728 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_65
timestamp 1698431365
transform 1 0 8624 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_80
timestamp 1698431365
transform 1 0 10304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_83
timestamp 1698431365
transform 1 0 10640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_85
timestamp 1698431365
transform 1 0 10864 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_92
timestamp 1698431365
transform 1 0 11648 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_98
timestamp 1698431365
transform 1 0 12320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_131
timestamp 1698431365
transform 1 0 16016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_135
timestamp 1698431365
transform 1 0 16464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_150
timestamp 1698431365
transform 1 0 18144 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_160
timestamp 1698431365
transform 1 0 19264 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_173
timestamp 1698431365
transform 1 0 20720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_177
timestamp 1698431365
transform 1 0 21168 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_218
timestamp 1698431365
transform 1 0 25760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_228
timestamp 1698431365
transform 1 0 26880 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_232
timestamp 1698431365
transform 1 0 27328 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_236
timestamp 1698431365
transform 1 0 27776 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_239
timestamp 1698431365
transform 1 0 28112 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_6
timestamp 1698431365
transform 1 0 2016 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_23
timestamp 1698431365
transform 1 0 3920 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_29
timestamp 1698431365
transform 1 0 4592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_33
timestamp 1698431365
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_66
timestamp 1698431365
transform 1 0 8736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_70
timestamp 1698431365
transform 1 0 9184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_74
timestamp 1698431365
transform 1 0 9632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_76
timestamp 1698431365
transform 1 0 9856 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_90
timestamp 1698431365
transform 1 0 11424 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_100
timestamp 1698431365
transform 1 0 12544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_111
timestamp 1698431365
transform 1 0 13776 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_125
timestamp 1698431365
transform 1 0 15344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_129
timestamp 1698431365
transform 1 0 15792 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_145
timestamp 1698431365
transform 1 0 17584 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_151
timestamp 1698431365
transform 1 0 18256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_155
timestamp 1698431365
transform 1 0 18704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_157
timestamp 1698431365
transform 1 0 18928 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_160
timestamp 1698431365
transform 1 0 19264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_182
timestamp 1698431365
transform 1 0 21728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_184
timestamp 1698431365
transform 1 0 21952 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_194
timestamp 1698431365
transform 1 0 23072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_204
timestamp 1698431365
transform 1 0 24192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_208
timestamp 1698431365
transform 1 0 24640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_31
timestamp 1698431365
transform 1 0 4816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_43
timestamp 1698431365
transform 1 0 6160 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_48
timestamp 1698431365
transform 1 0 6720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_50
timestamp 1698431365
transform 1 0 6944 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_53
timestamp 1698431365
transform 1 0 7280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_89
timestamp 1698431365
transform 1 0 11312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_93
timestamp 1698431365
transform 1 0 11760 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_97
timestamp 1698431365
transform 1 0 12208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_101
timestamp 1698431365
transform 1 0 12656 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_109
timestamp 1698431365
transform 1 0 13552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_113
timestamp 1698431365
transform 1 0 14000 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_121
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_127
timestamp 1698431365
transform 1 0 15568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_131
timestamp 1698431365
transform 1 0 16016 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_146
timestamp 1698431365
transform 1 0 17696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_148
timestamp 1698431365
transform 1 0 17920 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_151
timestamp 1698431365
transform 1 0 18256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_155
timestamp 1698431365
transform 1 0 18704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_159
timestamp 1698431365
transform 1 0 19152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_161
timestamp 1698431365
transform 1 0 19376 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_171
timestamp 1698431365
transform 1 0 20496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_175
timestamp 1698431365
transform 1 0 20944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_179
timestamp 1698431365
transform 1 0 21392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_183
timestamp 1698431365
transform 1 0 21840 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_187
timestamp 1698431365
transform 1 0 22288 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_193
timestamp 1698431365
transform 1 0 22960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_197
timestamp 1698431365
transform 1 0 23408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_201
timestamp 1698431365
transform 1 0 23856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_203
timestamp 1698431365
transform 1 0 24080 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_234
timestamp 1698431365
transform 1 0 27552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_238
timestamp 1698431365
transform 1 0 28000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_240
timestamp 1698431365
transform 1 0 28224 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_8
timestamp 1698431365
transform 1 0 2240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_10
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_21
timestamp 1698431365
transform 1 0 3696 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_29
timestamp 1698431365
transform 1 0 4592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_33
timestamp 1698431365
transform 1 0 5040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_68
timestamp 1698431365
transform 1 0 8960 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_93
timestamp 1698431365
transform 1 0 11760 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_97
timestamp 1698431365
transform 1 0 12208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_111
timestamp 1698431365
transform 1 0 13776 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_123
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_125
timestamp 1698431365
transform 1 0 15344 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_136
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_142
timestamp 1698431365
transform 1 0 17248 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_144
timestamp 1698431365
transform 1 0 17472 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_155
timestamp 1698431365
transform 1 0 18704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_170
timestamp 1698431365
transform 1 0 20384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_181
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_190
timestamp 1698431365
transform 1 0 22624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_194
timestamp 1698431365
transform 1 0 23072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_198
timestamp 1698431365
transform 1 0 23520 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_202
timestamp 1698431365
transform 1 0 23968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_206
timestamp 1698431365
transform 1 0 24416 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_210
timestamp 1698431365
transform 1 0 24864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_214
timestamp 1698431365
transform 1 0 25312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_216
timestamp 1698431365
transform 1 0 25536 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_219
timestamp 1698431365
transform 1 0 25872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_223
timestamp 1698431365
transform 1 0 26320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_227
timestamp 1698431365
transform 1 0 26768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_229
timestamp 1698431365
transform 1 0 26992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_232
timestamp 1698431365
transform 1 0 27328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_234
timestamp 1698431365
transform 1 0 27552 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_237
timestamp 1698431365
transform 1 0 27888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_6
timestamp 1698431365
transform 1 0 2016 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_14
timestamp 1698431365
transform 1 0 2912 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_20
timestamp 1698431365
transform 1 0 3584 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_52
timestamp 1698431365
transform 1 0 7168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_56
timestamp 1698431365
transform 1 0 7616 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_76
timestamp 1698431365
transform 1 0 9856 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_86
timestamp 1698431365
transform 1 0 10976 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_90
timestamp 1698431365
transform 1 0 11424 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_103
timestamp 1698431365
transform 1 0 12880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_105
timestamp 1698431365
transform 1 0 13104 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_135
timestamp 1698431365
transform 1 0 16464 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_171
timestamp 1698431365
transform 1 0 20496 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_202
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_8
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_12
timestamp 1698431365
transform 1 0 2688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_14
timestamp 1698431365
transform 1 0 2912 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_19
timestamp 1698431365
transform 1 0 3472 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_25
timestamp 1698431365
transform 1 0 4144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_57
timestamp 1698431365
transform 1 0 7728 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_59
timestamp 1698431365
transform 1 0 7952 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_73
timestamp 1698431365
transform 1 0 9520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_75
timestamp 1698431365
transform 1 0 9744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_139
timestamp 1698431365
transform 1 0 16912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_143
timestamp 1698431365
transform 1 0 17360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_147
timestamp 1698431365
transform 1 0 17808 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_151
timestamp 1698431365
transform 1 0 18256 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_154
timestamp 1698431365
transform 1 0 18592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_164
timestamp 1698431365
transform 1 0 19712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_168
timestamp 1698431365
transform 1 0 20160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_189
timestamp 1698431365
transform 1 0 22512 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_193
timestamp 1698431365
transform 1 0 22960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_234
timestamp 1698431365
transform 1 0 27552 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_238
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_31
timestamp 1698431365
transform 1 0 4816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_35
timestamp 1698431365
transform 1 0 5264 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_43
timestamp 1698431365
transform 1 0 6160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_47
timestamp 1698431365
transform 1 0 6608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_59
timestamp 1698431365
transform 1 0 7952 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_95
timestamp 1698431365
transform 1 0 11984 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_104
timestamp 1698431365
transform 1 0 12992 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_110
timestamp 1698431365
transform 1 0 13664 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_125
timestamp 1698431365
transform 1 0 15344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_129
timestamp 1698431365
transform 1 0 15792 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_150
timestamp 1698431365
transform 1 0 18144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_163
timestamp 1698431365
transform 1 0 19600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_167
timestamp 1698431365
transform 1 0 20048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_169
timestamp 1698431365
transform 1 0 20272 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_172
timestamp 1698431365
transform 1 0 20608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_176
timestamp 1698431365
transform 1 0 21056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_180
timestamp 1698431365
transform 1 0 21504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_184
timestamp 1698431365
transform 1 0 21952 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_191
timestamp 1698431365
transform 1 0 22736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_195
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_199
timestamp 1698431365
transform 1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_220
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_230
timestamp 1698431365
transform 1 0 27104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_234
timestamp 1698431365
transform 1 0 27552 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_236
timestamp 1698431365
transform 1 0 27776 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_239
timestamp 1698431365
transform 1 0 28112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_16
timestamp 1698431365
transform 1 0 3136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_20
timestamp 1698431365
transform 1 0 3584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_24
timestamp 1698431365
transform 1 0 4032 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_39
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_71
timestamp 1698431365
transform 1 0 9296 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_75
timestamp 1698431365
transform 1 0 9744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_86
timestamp 1698431365
transform 1 0 10976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_90
timestamp 1698431365
transform 1 0 11424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_92
timestamp 1698431365
transform 1 0 11648 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_95
timestamp 1698431365
transform 1 0 11984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_99
timestamp 1698431365
transform 1 0 12432 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_113
timestamp 1698431365
transform 1 0 14000 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_166
timestamp 1698431365
transform 1 0 19936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_170
timestamp 1698431365
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_172
timestamp 1698431365
transform 1 0 20608 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_197
timestamp 1698431365
transform 1 0 23408 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_201
timestamp 1698431365
transform 1 0 23856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_205
timestamp 1698431365
transform 1 0 24304 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_211
timestamp 1698431365
transform 1 0 24976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_215
timestamp 1698431365
transform 1 0 25424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_219
timestamp 1698431365
transform 1 0 25872 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_223
timestamp 1698431365
transform 1 0 26320 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_227
timestamp 1698431365
transform 1 0 26768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_231
timestamp 1698431365
transform 1 0 27216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_235
timestamp 1698431365
transform 1 0 27664 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_6
timestamp 1698431365
transform 1 0 2016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_10
timestamp 1698431365
transform 1 0 2464 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_14
timestamp 1698431365
transform 1 0 2912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_16
timestamp 1698431365
transform 1 0 3136 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_21
timestamp 1698431365
transform 1 0 3696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_25
timestamp 1698431365
transform 1 0 4144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_29
timestamp 1698431365
transform 1 0 4592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_35
timestamp 1698431365
transform 1 0 5264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_39
timestamp 1698431365
transform 1 0 5712 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_55
timestamp 1698431365
transform 1 0 7504 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_63
timestamp 1698431365
transform 1 0 8400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_67
timestamp 1698431365
transform 1 0 8848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_86
timestamp 1698431365
transform 1 0 10976 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_90
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_94
timestamp 1698431365
transform 1 0 11872 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_100
timestamp 1698431365
transform 1 0 12544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_104
timestamp 1698431365
transform 1 0 12992 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_108
timestamp 1698431365
transform 1 0 13440 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_110
timestamp 1698431365
transform 1 0 13664 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_146
timestamp 1698431365
transform 1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_148
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_169
timestamp 1698431365
transform 1 0 20272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1698431365
transform 1 0 24528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_47
timestamp 1698431365
transform 1 0 6608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_51
timestamp 1698431365
transform 1 0 7056 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_54
timestamp 1698431365
transform 1 0 7392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_58
timestamp 1698431365
transform 1 0 7840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_62
timestamp 1698431365
transform 1 0 8288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_66
timestamp 1698431365
transform 1 0 8736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_70
timestamp 1698431365
transform 1 0 9184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_72
timestamp 1698431365
transform 1 0 9408 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_75
timestamp 1698431365
transform 1 0 9744 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_113
timestamp 1698431365
transform 1 0 14000 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_116
timestamp 1698431365
transform 1 0 14336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_128
timestamp 1698431365
transform 1 0 15680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_132
timestamp 1698431365
transform 1 0 16128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_136
timestamp 1698431365
transform 1 0 16576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_138
timestamp 1698431365
transform 1 0 16800 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_141
timestamp 1698431365
transform 1 0 17136 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_145
timestamp 1698431365
transform 1 0 17584 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_148
timestamp 1698431365
transform 1 0 17920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_152
timestamp 1698431365
transform 1 0 18368 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_156
timestamp 1698431365
transform 1 0 18816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_160
timestamp 1698431365
transform 1 0 19264 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_163
timestamp 1698431365
transform 1 0 19600 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_167
timestamp 1698431365
transform 1 0 20048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_181
timestamp 1698431365
transform 1 0 21616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_185
timestamp 1698431365
transform 1 0 22064 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_189
timestamp 1698431365
transform 1 0 22512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_237
timestamp 1698431365
transform 1 0 27888 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_54
timestamp 1698431365
transform 1 0 7392 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_78
timestamp 1698431365
transform 1 0 10080 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_82
timestamp 1698431365
transform 1 0 10528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_102
timestamp 1698431365
transform 1 0 12768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_107
timestamp 1698431365
transform 1 0 13328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_111
timestamp 1698431365
transform 1 0 13776 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_115
timestamp 1698431365
transform 1 0 14224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_119
timestamp 1698431365
transform 1 0 14672 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_125
timestamp 1698431365
transform 1 0 15344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_129
timestamp 1698431365
transform 1 0 15792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_133
timestamp 1698431365
transform 1 0 16240 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_144
timestamp 1698431365
transform 1 0 17472 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_174
timestamp 1698431365
transform 1 0 20832 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_178
timestamp 1698431365
transform 1 0 21280 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_182
timestamp 1698431365
transform 1 0 21728 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_186
timestamp 1698431365
transform 1 0 22176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_190
timestamp 1698431365
transform 1 0 22624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_194
timestamp 1698431365
transform 1 0 23072 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_198
timestamp 1698431365
transform 1 0 23520 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_222
timestamp 1698431365
transform 1 0 26208 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_225
timestamp 1698431365
transform 1 0 26544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_229
timestamp 1698431365
transform 1 0 26992 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_235
timestamp 1698431365
transform 1 0 27664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_4
timestamp 1698431365
transform 1 0 1792 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_7
timestamp 1698431365
transform 1 0 2128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_17
timestamp 1698431365
transform 1 0 3248 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_21
timestamp 1698431365
transform 1 0 3696 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_25
timestamp 1698431365
transform 1 0 4144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_29
timestamp 1698431365
transform 1 0 4592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1698431365
transform 1 0 5040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_39
timestamp 1698431365
transform 1 0 5712 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_46
timestamp 1698431365
transform 1 0 6496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_48
timestamp 1698431365
transform 1 0 6720 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_51
timestamp 1698431365
transform 1 0 7056 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_84
timestamp 1698431365
transform 1 0 10752 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_88
timestamp 1698431365
transform 1 0 11200 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_91
timestamp 1698431365
transform 1 0 11536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_95
timestamp 1698431365
transform 1 0 11984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_99
timestamp 1698431365
transform 1 0 12432 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_115
timestamp 1698431365
transform 1 0 14224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_148
timestamp 1698431365
transform 1 0 17920 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_158
timestamp 1698431365
transform 1 0 19040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_168
timestamp 1698431365
transform 1 0 20160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_181
timestamp 1698431365
transform 1 0 21616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_185
timestamp 1698431365
transform 1 0 22064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_189
timestamp 1698431365
transform 1 0 22512 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_193
timestamp 1698431365
transform 1 0 22960 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_197
timestamp 1698431365
transform 1 0 23408 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_200
timestamp 1698431365
transform 1 0 23744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_204
timestamp 1698431365
transform 1 0 24192 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_210
timestamp 1698431365
transform 1 0 24864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_214
timestamp 1698431365
transform 1 0 25312 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_230
timestamp 1698431365
transform 1 0 27104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_234
timestamp 1698431365
transform 1 0 27552 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_240
timestamp 1698431365
transform 1 0 28224 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_8
timestamp 1698431365
transform 1 0 2240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_19
timestamp 1698431365
transform 1 0 3472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_52
timestamp 1698431365
transform 1 0 7168 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_86
timestamp 1698431365
transform 1 0 10976 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_90
timestamp 1698431365
transform 1 0 11424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_94
timestamp 1698431365
transform 1 0 11872 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_125
timestamp 1698431365
transform 1 0 15344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_137
timestamp 1698431365
transform 1 0 16688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_153
timestamp 1698431365
transform 1 0 18480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_155
timestamp 1698431365
transform 1 0 18704 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_174
timestamp 1698431365
transform 1 0 20832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_191
timestamp 1698431365
transform 1 0 22736 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_195
timestamp 1698431365
transform 1 0 23184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_197
timestamp 1698431365
transform 1 0 23408 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_31
timestamp 1698431365
transform 1 0 4816 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_41
timestamp 1698431365
transform 1 0 5936 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_79
timestamp 1698431365
transform 1 0 10192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_89
timestamp 1698431365
transform 1 0 11312 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_93
timestamp 1698431365
transform 1 0 11760 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_97
timestamp 1698431365
transform 1 0 12208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_159
timestamp 1698431365
transform 1 0 19152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_235
timestamp 1698431365
transform 1 0 27664 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_239
timestamp 1698431365
transform 1 0 28112 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_6
timestamp 1698431365
transform 1 0 2016 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_15
timestamp 1698431365
transform 1 0 3024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_67
timestamp 1698431365
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_87
timestamp 1698431365
transform 1 0 11088 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_117
timestamp 1698431365
transform 1 0 14448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_123
timestamp 1698431365
transform 1 0 15120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_125
timestamp 1698431365
transform 1 0 15344 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_166
timestamp 1698431365
transform 1 0 19936 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_170
timestamp 1698431365
transform 1 0 20384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_174
timestamp 1698431365
transform 1 0 20832 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_176
timestamp 1698431365
transform 1 0 21056 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_179
timestamp 1698431365
transform 1 0 21392 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_183
timestamp 1698431365
transform 1 0 21840 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_187
timestamp 1698431365
transform 1 0 22288 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_191
timestamp 1698431365
transform 1 0 22736 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_195
timestamp 1698431365
transform 1 0 23184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_199
timestamp 1698431365
transform 1 0 23632 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_214
timestamp 1698431365
transform 1 0 25312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_237
timestamp 1698431365
transform 1 0 27888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_8
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_12
timestamp 1698431365
transform 1 0 2688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_16
timestamp 1698431365
transform 1 0 3136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_30
timestamp 1698431365
transform 1 0 4704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_53
timestamp 1698431365
transform 1 0 7280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_55
timestamp 1698431365
transform 1 0 7504 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_72
timestamp 1698431365
transform 1 0 9408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_76
timestamp 1698431365
transform 1 0 9856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_89
timestamp 1698431365
transform 1 0 11312 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_91
timestamp 1698431365
transform 1 0 11536 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_102
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_115
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_117
timestamp 1698431365
transform 1 0 14448 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_127
timestamp 1698431365
transform 1 0 15568 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_173
timestamp 1698431365
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_190
timestamp 1698431365
transform 1 0 22624 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_4
timestamp 1698431365
transform 1 0 1792 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_21
timestamp 1698431365
transform 1 0 3696 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_25
timestamp 1698431365
transform 1 0 4144 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_28
timestamp 1698431365
transform 1 0 4480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_32
timestamp 1698431365
transform 1 0 4928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_36
timestamp 1698431365
transform 1 0 5376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_38
timestamp 1698431365
transform 1 0 5600 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_41
timestamp 1698431365
transform 1 0 5936 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_45
timestamp 1698431365
transform 1 0 6384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_49
timestamp 1698431365
transform 1 0 6832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_53
timestamp 1698431365
transform 1 0 7280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_57
timestamp 1698431365
transform 1 0 7728 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_61
timestamp 1698431365
transform 1 0 8176 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_63
timestamp 1698431365
transform 1 0 8400 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_81
timestamp 1698431365
transform 1 0 10416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_87
timestamp 1698431365
transform 1 0 11088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_91
timestamp 1698431365
transform 1 0 11536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_95
timestamp 1698431365
transform 1 0 11984 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_99
timestamp 1698431365
transform 1 0 12432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_103
timestamp 1698431365
transform 1 0 12880 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_127
timestamp 1698431365
transform 1 0 15568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_146
timestamp 1698431365
transform 1 0 17696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_150
timestamp 1698431365
transform 1 0 18144 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_180
timestamp 1698431365
transform 1 0 21504 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_192
timestamp 1698431365
transform 1 0 22848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_196
timestamp 1698431365
transform 1 0 23296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_200
timestamp 1698431365
transform 1 0 23744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_204
timestamp 1698431365
transform 1 0 24192 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_31
timestamp 1698431365
transform 1 0 4816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_43
timestamp 1698431365
transform 1 0 6160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_55
timestamp 1698431365
transform 1 0 7504 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_64
timestamp 1698431365
transform 1 0 8512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_70
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_74
timestamp 1698431365
transform 1 0 9632 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_78
timestamp 1698431365
transform 1 0 10080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_82
timestamp 1698431365
transform 1 0 10528 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_94
timestamp 1698431365
transform 1 0 11872 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_103
timestamp 1698431365
transform 1 0 12880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_168
timestamp 1698431365
transform 1 0 20160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_172
timestamp 1698431365
transform 1 0 20608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_174
timestamp 1698431365
transform 1 0 20832 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_206
timestamp 1698431365
transform 1 0 24416 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_210
timestamp 1698431365
transform 1 0 24864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_214
timestamp 1698431365
transform 1 0 25312 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_8
timestamp 1698431365
transform 1 0 2240 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_14
timestamp 1698431365
transform 1 0 2912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_18
timestamp 1698431365
transform 1 0 3360 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_22
timestamp 1698431365
transform 1 0 3808 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_26
timestamp 1698431365
transform 1 0 4256 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_65
timestamp 1698431365
transform 1 0 8624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_67
timestamp 1698431365
transform 1 0 8848 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_76
timestamp 1698431365
transform 1 0 9856 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_108
timestamp 1698431365
transform 1 0 13440 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_183
timestamp 1698431365
transform 1 0 21840 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_187
timestamp 1698431365
transform 1 0 22288 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_189
timestamp 1698431365
transform 1 0 22512 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_198
timestamp 1698431365
transform 1 0 23520 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_200
timestamp 1698431365
transform 1 0 23744 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_209
timestamp 1698431365
transform 1 0 24752 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_220
timestamp 1698431365
transform 1 0 25984 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_224
timestamp 1698431365
transform 1 0 26432 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_228
timestamp 1698431365
transform 1 0 26880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_232
timestamp 1698431365
transform 1 0 27328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_236
timestamp 1698431365
transform 1 0 27776 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_238
timestamp 1698431365
transform 1 0 28000 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_8
timestamp 1698431365
transform 1 0 2240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_12
timestamp 1698431365
transform 1 0 2688 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_23
timestamp 1698431365
transform 1 0 3920 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_25
timestamp 1698431365
transform 1 0 4144 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_28
timestamp 1698431365
transform 1 0 4480 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698431365
transform 1 0 4928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_44
timestamp 1698431365
transform 1 0 6272 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_75
timestamp 1698431365
transform 1 0 9744 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_85
timestamp 1698431365
transform 1 0 10864 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_89
timestamp 1698431365
transform 1 0 11312 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_93
timestamp 1698431365
transform 1 0 11760 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_97
timestamp 1698431365
transform 1 0 12208 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_120
timestamp 1698431365
transform 1 0 14784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_122
timestamp 1698431365
transform 1 0 15008 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_160
timestamp 1698431365
transform 1 0 19264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_164
timestamp 1698431365
transform 1 0 19712 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_185
timestamp 1698431365
transform 1 0 22064 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_189
timestamp 1698431365
transform 1 0 22512 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_193
timestamp 1698431365
transform 1 0 22960 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_195
timestamp 1698431365
transform 1 0 23184 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_233
timestamp 1698431365
transform 1 0 27440 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_237
timestamp 1698431365
transform 1 0 27888 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_37
timestamp 1698431365
transform 1 0 5488 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_41
timestamp 1698431365
transform 1 0 5936 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_45
timestamp 1698431365
transform 1 0 6384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_49
timestamp 1698431365
transform 1 0 6832 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_53
timestamp 1698431365
transform 1 0 7280 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_57
timestamp 1698431365
transform 1 0 7728 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_69
timestamp 1698431365
transform 1 0 9072 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_80
timestamp 1698431365
transform 1 0 10304 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_86
timestamp 1698431365
transform 1 0 10976 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_90
timestamp 1698431365
transform 1 0 11424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_92
timestamp 1698431365
transform 1 0 11648 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_95
timestamp 1698431365
transform 1 0 11984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_99
timestamp 1698431365
transform 1 0 12432 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_205
timestamp 1698431365
transform 1 0 24304 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_209
timestamp 1698431365
transform 1 0 24752 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_6
timestamp 1698431365
transform 1 0 2016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_12
timestamp 1698431365
transform 1 0 2688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_16
timestamp 1698431365
transform 1 0 3136 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_28
timestamp 1698431365
transform 1 0 4480 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_43
timestamp 1698431365
transform 1 0 6160 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_47
timestamp 1698431365
transform 1 0 6608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_51
timestamp 1698431365
transform 1 0 7056 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_55
timestamp 1698431365
transform 1 0 7504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_59
timestamp 1698431365
transform 1 0 7952 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_63
timestamp 1698431365
transform 1 0 8400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_67
timestamp 1698431365
transform 1 0 8848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_71
timestamp 1698431365
transform 1 0 9296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_75
timestamp 1698431365
transform 1 0 9744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_79
timestamp 1698431365
transform 1 0 10192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_83
timestamp 1698431365
transform 1 0 10640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_87
timestamp 1698431365
transform 1 0 11088 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_102
timestamp 1698431365
transform 1 0 12768 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_104
timestamp 1698431365
transform 1 0 12992 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_218
timestamp 1698431365
transform 1 0 25760 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_228
timestamp 1698431365
transform 1 0 26880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_232
timestamp 1698431365
transform 1 0 27328 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_236
timestamp 1698431365
transform 1 0 27776 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_240
timestamp 1698431365
transform 1 0 28224 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_8
timestamp 1698431365
transform 1 0 2240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_22
timestamp 1698431365
transform 1 0 3808 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_24
timestamp 1698431365
transform 1 0 4032 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_56
timestamp 1698431365
transform 1 0 7616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_90
timestamp 1698431365
transform 1 0 11424 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_179
timestamp 1698431365
transform 1 0 21392 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_214
timestamp 1698431365
transform 1 0 25312 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_223
timestamp 1698431365
transform 1 0 26320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_227
timestamp 1698431365
transform 1 0 26768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_231
timestamp 1698431365
transform 1 0 27216 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_235
timestamp 1698431365
transform 1 0 27664 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_239
timestamp 1698431365
transform 1 0 28112 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_31
timestamp 1698431365
transform 1 0 4816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_41
timestamp 1698431365
transform 1 0 5936 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_81
timestamp 1698431365
transform 1 0 10416 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_85
timestamp 1698431365
transform 1 0 10864 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_161
timestamp 1698431365
transform 1 0 19376 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_165
timestamp 1698431365
transform 1 0 19824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_169
timestamp 1698431365
transform 1 0 20272 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_173
timestamp 1698431365
transform 1 0 20720 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_203
timestamp 1698431365
transform 1 0 24080 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_207
timestamp 1698431365
transform 1 0 24528 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_238
timestamp 1698431365
transform 1 0 28000 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_240
timestamp 1698431365
transform 1 0 28224 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_14
timestamp 1698431365
transform 1 0 2912 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_18
timestamp 1698431365
transform 1 0 3360 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_27
timestamp 1698431365
transform 1 0 4368 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_31
timestamp 1698431365
transform 1 0 4816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_35
timestamp 1698431365
transform 1 0 5264 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_47
timestamp 1698431365
transform 1 0 6608 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_51
timestamp 1698431365
transform 1 0 7056 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_54
timestamp 1698431365
transform 1 0 7392 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_58
timestamp 1698431365
transform 1 0 7840 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_122
timestamp 1698431365
transform 1 0 15008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_146
timestamp 1698431365
transform 1 0 17696 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_150
timestamp 1698431365
transform 1 0 18144 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_162
timestamp 1698431365
transform 1 0 19488 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_208
timestamp 1698431365
transform 1 0 24640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_216
timestamp 1698431365
transform 1 0 25536 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_220
timestamp 1698431365
transform 1 0 25984 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_229
timestamp 1698431365
transform 1 0 26992 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_233
timestamp 1698431365
transform 1 0 27440 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_237
timestamp 1698431365
transform 1 0 27888 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_6
timestamp 1698431365
transform 1 0 2016 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_15
timestamp 1698431365
transform 1 0 3024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_19
timestamp 1698431365
transform 1 0 3472 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698431365
transform 1 0 4928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_41
timestamp 1698431365
transform 1 0 5936 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_45
timestamp 1698431365
transform 1 0 6384 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_49
timestamp 1698431365
transform 1 0 6832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_100
timestamp 1698431365
transform 1 0 12544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_102
timestamp 1698431365
transform 1 0 12768 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1698431365
transform 1 0 20832 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_195
timestamp 1698431365
transform 1 0 23184 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_199
timestamp 1698431365
transform 1 0 23632 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_203
timestamp 1698431365
transform 1 0 24080 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_207
timestamp 1698431365
transform 1 0 24528 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_211
timestamp 1698431365
transform 1 0 24976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_215
timestamp 1698431365
transform 1 0 25424 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_219
timestamp 1698431365
transform 1 0 25872 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_238
timestamp 1698431365
transform 1 0 28000 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_240
timestamp 1698431365
transform 1 0 28224 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_14
timestamp 1698431365
transform 1 0 2912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_16
timestamp 1698431365
transform 1 0 3136 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_19
timestamp 1698431365
transform 1 0 3472 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_51
timestamp 1698431365
transform 1 0 7056 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_55
timestamp 1698431365
transform 1 0 7504 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_58
timestamp 1698431365
transform 1 0 7840 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_62
timestamp 1698431365
transform 1 0 8288 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_81
timestamp 1698431365
transform 1 0 10416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_83
timestamp 1698431365
transform 1 0 10640 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_86
timestamp 1698431365
transform 1 0 10976 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_179
timestamp 1698431365
transform 1 0 21392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_8
timestamp 1698431365
transform 1 0 2240 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_15
timestamp 1698431365
transform 1 0 3024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_17
timestamp 1698431365
transform 1 0 3248 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_20
timestamp 1698431365
transform 1 0 3584 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_33
timestamp 1698431365
transform 1 0 5040 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_74
timestamp 1698431365
transform 1 0 9632 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_78
timestamp 1698431365
transform 1 0 10080 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_89
timestamp 1698431365
transform 1 0 11312 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_111
timestamp 1698431365
transform 1 0 13776 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_114
timestamp 1698431365
transform 1 0 14112 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_155
timestamp 1698431365
transform 1 0 18704 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_159
timestamp 1698431365
transform 1 0 19152 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_174
timestamp 1698431365
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_188
timestamp 1698431365
transform 1 0 22400 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_206
timestamp 1698431365
transform 1 0 24416 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_210
timestamp 1698431365
transform 1 0 24864 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_214
timestamp 1698431365
transform 1 0 25312 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_216
timestamp 1698431365
transform 1 0 25536 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_233
timestamp 1698431365
transform 1 0 27440 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_237
timestamp 1698431365
transform 1 0 27888 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_8
timestamp 1698431365
transform 1 0 2240 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_22
timestamp 1698431365
transform 1 0 3808 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_26
timestamp 1698431365
transform 1 0 4256 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_29
timestamp 1698431365
transform 1 0 4592 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_33
timestamp 1698431365
transform 1 0 5040 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_37
timestamp 1698431365
transform 1 0 5488 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_41
timestamp 1698431365
transform 1 0 5936 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_45
timestamp 1698431365
transform 1 0 6384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_55
timestamp 1698431365
transform 1 0 7504 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_59
timestamp 1698431365
transform 1 0 7952 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_62
timestamp 1698431365
transform 1 0 8288 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_111
timestamp 1698431365
transform 1 0 13776 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_113
timestamp 1698431365
transform 1 0 14000 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_171
timestamp 1698431365
transform 1 0 20496 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_173
timestamp 1698431365
transform 1 0 20720 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_182
timestamp 1698431365
transform 1 0 21728 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_186
timestamp 1698431365
transform 1 0 22176 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_190
timestamp 1698431365
transform 1 0 22624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_194
timestamp 1698431365
transform 1 0 23072 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_198
timestamp 1698431365
transform 1 0 23520 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_202
timestamp 1698431365
transform 1 0 23968 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_216
timestamp 1698431365
transform 1 0 25536 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_220
timestamp 1698431365
transform 1 0 25984 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_224
timestamp 1698431365
transform 1 0 26432 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_228
timestamp 1698431365
transform 1 0 26880 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_232
timestamp 1698431365
transform 1 0 27328 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_236
timestamp 1698431365
transform 1 0 27776 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_240
timestamp 1698431365
transform 1 0 28224 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_31
timestamp 1698431365
transform 1 0 4816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_43
timestamp 1698431365
transform 1 0 6160 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_49
timestamp 1698431365
transform 1 0 6832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_53
timestamp 1698431365
transform 1 0 7280 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_57
timestamp 1698431365
transform 1 0 7728 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_61
timestamp 1698431365
transform 1 0 8176 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_65
timestamp 1698431365
transform 1 0 8624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_69
timestamp 1698431365
transform 1 0 9072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_73
timestamp 1698431365
transform 1 0 9520 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_77
timestamp 1698431365
transform 1 0 9968 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_81
timestamp 1698431365
transform 1 0 10416 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_85
timestamp 1698431365
transform 1 0 10864 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_89
timestamp 1698431365
transform 1 0 11312 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_93
timestamp 1698431365
transform 1 0 11760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_97
timestamp 1698431365
transform 1 0 12208 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_111
timestamp 1698431365
transform 1 0 13776 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_193
timestamp 1698431365
transform 1 0 22960 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_197
timestamp 1698431365
transform 1 0 23408 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_201
timestamp 1698431365
transform 1 0 23856 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_205
timestamp 1698431365
transform 1 0 24304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_209
timestamp 1698431365
transform 1 0 24752 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_211
timestamp 1698431365
transform 1 0 24976 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_237
timestamp 1698431365
transform 1 0 27888 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_8
timestamp 1698431365
transform 1 0 2240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_12
timestamp 1698431365
transform 1 0 2688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_16
timestamp 1698431365
transform 1 0 3136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_18
timestamp 1698431365
transform 1 0 3360 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_56
timestamp 1698431365
transform 1 0 7616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_58
timestamp 1698431365
transform 1 0 7840 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_69
timestamp 1698431365
transform 1 0 9072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_83
timestamp 1698431365
transform 1 0 10640 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_156
timestamp 1698431365
transform 1 0 18816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_189
timestamp 1698431365
transform 1 0 22512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_193
timestamp 1698431365
transform 1 0 22960 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_203
timestamp 1698431365
transform 1 0 24080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_207
timestamp 1698431365
transform 1 0 24528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_209
timestamp 1698431365
transform 1 0 24752 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_22
timestamp 1698431365
transform 1 0 3808 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_26
timestamp 1698431365
transform 1 0 4256 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_30
timestamp 1698431365
transform 1 0 4704 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_32
timestamp 1698431365
transform 1 0 4928 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_115
timestamp 1698431365
transform 1 0 14224 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_117
timestamp 1698431365
transform 1 0 14448 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_170
timestamp 1698431365
transform 1 0 20384 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_174
timestamp 1698431365
transform 1 0 20832 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_181
timestamp 1698431365
transform 1 0 21616 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_211
timestamp 1698431365
transform 1 0 24976 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_215
timestamp 1698431365
transform 1 0 25424 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_218
timestamp 1698431365
transform 1 0 25760 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_222
timestamp 1698431365
transform 1 0 26208 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_226
timestamp 1698431365
transform 1 0 26656 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_230
timestamp 1698431365
transform 1 0 27104 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_234
timestamp 1698431365
transform 1 0 27552 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_237
timestamp 1698431365
transform 1 0 27888 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_31
timestamp 1698431365
transform 1 0 4816 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_35
timestamp 1698431365
transform 1 0 5264 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_39
timestamp 1698431365
transform 1 0 5712 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_49
timestamp 1698431365
transform 1 0 6832 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_53
timestamp 1698431365
transform 1 0 7280 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_57
timestamp 1698431365
transform 1 0 7728 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_59
timestamp 1698431365
transform 1 0 7952 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_62
timestamp 1698431365
transform 1 0 8288 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_66
timestamp 1698431365
transform 1 0 8736 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_80
timestamp 1698431365
transform 1 0 10304 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_82
timestamp 1698431365
transform 1 0 10528 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_85
timestamp 1698431365
transform 1 0 10864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_89
timestamp 1698431365
transform 1 0 11312 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_101
timestamp 1698431365
transform 1 0 12656 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_103
timestamp 1698431365
transform 1 0 12880 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_106
timestamp 1698431365
transform 1 0 13216 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_110
timestamp 1698431365
transform 1 0 13664 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_114
timestamp 1698431365
transform 1 0 14112 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_120
timestamp 1698431365
transform 1 0 14784 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_179
timestamp 1698431365
transform 1 0 21392 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_183
timestamp 1698431365
transform 1 0 21840 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_187
timestamp 1698431365
transform 1 0 22288 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_207
timestamp 1698431365
transform 1 0 24528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_209
timestamp 1698431365
transform 1 0 24752 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_216
timestamp 1698431365
transform 1 0 25536 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_234
timestamp 1698431365
transform 1 0 27552 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_238
timestamp 1698431365
transform 1 0 28000 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_240
timestamp 1698431365
transform 1 0 28224 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_2
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_6
timestamp 1698431365
transform 1 0 2016 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_26
timestamp 1698431365
transform 1 0 4256 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_30
timestamp 1698431365
transform 1 0 4704 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_45
timestamp 1698431365
transform 1 0 6384 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_61
timestamp 1698431365
transform 1 0 8176 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_69
timestamp 1698431365
transform 1 0 9072 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_72
timestamp 1698431365
transform 1 0 9408 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_76
timestamp 1698431365
transform 1 0 9856 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_80
timestamp 1698431365
transform 1 0 10304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_84
timestamp 1698431365
transform 1 0 10752 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_98
timestamp 1698431365
transform 1 0 12320 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_111
timestamp 1698431365
transform 1 0 13776 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_115
timestamp 1698431365
transform 1 0 14224 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_119
timestamp 1698431365
transform 1 0 14672 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_123
timestamp 1698431365
transform 1 0 15120 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_129
timestamp 1698431365
transform 1 0 15792 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_170
timestamp 1698431365
transform 1 0 20384 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_174
timestamp 1698431365
transform 1 0 20832 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_181
timestamp 1698431365
transform 1 0 21616 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_185
timestamp 1698431365
transform 1 0 22064 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_189
timestamp 1698431365
transform 1 0 22512 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_193
timestamp 1698431365
transform 1 0 22960 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_195
timestamp 1698431365
transform 1 0 23184 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_198
timestamp 1698431365
transform 1 0 23520 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_202
timestamp 1698431365
transform 1 0 23968 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_208
timestamp 1698431365
transform 1 0 24640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_8
timestamp 1698431365
transform 1 0 2240 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_12
timestamp 1698431365
transform 1 0 2688 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_14
timestamp 1698431365
transform 1 0 2912 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_19
timestamp 1698431365
transform 1 0 3472 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_23
timestamp 1698431365
transform 1 0 3920 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_41
timestamp 1698431365
transform 1 0 5936 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_55
timestamp 1698431365
transform 1 0 7504 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_59
timestamp 1698431365
transform 1 0 7952 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_67
timestamp 1698431365
transform 1 0 8848 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_69
timestamp 1698431365
transform 1 0 9072 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_79
timestamp 1698431365
transform 1 0 10192 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_109
timestamp 1698431365
transform 1 0 13552 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_146
timestamp 1698431365
transform 1 0 17696 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_148
timestamp 1698431365
transform 1 0 17920 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_178
timestamp 1698431365
transform 1 0 21280 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_182
timestamp 1698431365
transform 1 0 21728 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_186
timestamp 1698431365
transform 1 0 22176 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_204
timestamp 1698431365
transform 1 0 24192 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_208
timestamp 1698431365
transform 1 0 24640 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_216
timestamp 1698431365
transform 1 0 25536 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_226
timestamp 1698431365
transform 1 0 26656 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_230
timestamp 1698431365
transform 1 0 27104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_234
timestamp 1698431365
transform 1 0 27552 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_238
timestamp 1698431365
transform 1 0 28000 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_31
timestamp 1698431365
transform 1 0 4816 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_66
timestamp 1698431365
transform 1 0 8736 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_70
timestamp 1698431365
transform 1 0 9184 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_78
timestamp 1698431365
transform 1 0 10080 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_80
timestamp 1698431365
transform 1 0 10304 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_83
timestamp 1698431365
transform 1 0 10640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_95
timestamp 1698431365
transform 1 0 11984 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_101
timestamp 1698431365
transform 1 0 12656 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_172
timestamp 1698431365
transform 1 0 20608 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_174
timestamp 1698431365
transform 1 0 20832 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_179
timestamp 1698431365
transform 1 0 21392 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_209
timestamp 1698431365
transform 1 0 24752 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_211
timestamp 1698431365
transform 1 0 24976 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_2
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_4
timestamp 1698431365
transform 1 0 1792 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_23
timestamp 1698431365
transform 1 0 3920 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_60
timestamp 1698431365
transform 1 0 8064 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_64
timestamp 1698431365
transform 1 0 8512 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_74
timestamp 1698431365
transform 1 0 9632 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_85
timestamp 1698431365
transform 1 0 10864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_137
timestamp 1698431365
transform 1 0 16688 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_139
timestamp 1698431365
transform 1 0 16912 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_174
timestamp 1698431365
transform 1 0 20832 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_176
timestamp 1698431365
transform 1 0 21056 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_203
timestamp 1698431365
transform 1 0 24080 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_207
timestamp 1698431365
transform 1 0 24528 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_209
timestamp 1698431365
transform 1 0 24752 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_216
timestamp 1698431365
transform 1 0 25536 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_220
timestamp 1698431365
transform 1 0 25984 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_232
timestamp 1698431365
transform 1 0 27328 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_236
timestamp 1698431365
transform 1 0 27776 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_240
timestamp 1698431365
transform 1 0 28224 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_8
timestamp 1698431365
transform 1 0 2240 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_12
timestamp 1698431365
transform 1 0 2688 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_23
timestamp 1698431365
transform 1 0 3920 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_27
timestamp 1698431365
transform 1 0 4368 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_31
timestamp 1698431365
transform 1 0 4816 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_53
timestamp 1698431365
transform 1 0 7280 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_57
timestamp 1698431365
transform 1 0 7728 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_61
timestamp 1698431365
transform 1 0 8176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_65
timestamp 1698431365
transform 1 0 8624 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_104
timestamp 1698431365
transform 1 0 12992 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_129
timestamp 1698431365
transform 1 0 15792 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_181
timestamp 1698431365
transform 1 0 21616 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_185
timestamp 1698431365
transform 1 0 22064 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_194
timestamp 1698431365
transform 1 0 23072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_198
timestamp 1698431365
transform 1 0 23520 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_200
timestamp 1698431365
transform 1 0 23744 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_210
timestamp 1698431365
transform 1 0 24864 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_214
timestamp 1698431365
transform 1 0 25312 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_12
timestamp 1698431365
transform 1 0 2688 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_16
timestamp 1698431365
transform 1 0 3136 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_22
timestamp 1698431365
transform 1 0 3808 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_38
timestamp 1698431365
transform 1 0 5600 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_46
timestamp 1698431365
transform 1 0 6496 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_49
timestamp 1698431365
transform 1 0 6832 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_53
timestamp 1698431365
transform 1 0 7280 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_64
timestamp 1698431365
transform 1 0 8512 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_68
timestamp 1698431365
transform 1 0 8960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_78
timestamp 1698431365
transform 1 0 10080 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_84
timestamp 1698431365
transform 1 0 10752 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_88
timestamp 1698431365
transform 1 0 11200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_92
timestamp 1698431365
transform 1 0 11648 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_94
timestamp 1698431365
transform 1 0 11872 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_97
timestamp 1698431365
transform 1 0 12208 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_101
timestamp 1698431365
transform 1 0 12656 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_103
timestamp 1698431365
transform 1 0 12880 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_106
timestamp 1698431365
transform 1 0 13216 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_108
timestamp 1698431365
transform 1 0 13440 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_111
timestamp 1698431365
transform 1 0 13776 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_120
timestamp 1698431365
transform 1 0 14784 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_124
timestamp 1698431365
transform 1 0 15232 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_127
timestamp 1698431365
transform 1 0 15568 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_131
timestamp 1698431365
transform 1 0 16016 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_135
timestamp 1698431365
transform 1 0 16464 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_137
timestamp 1698431365
transform 1 0 16688 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_158
timestamp 1698431365
transform 1 0 19040 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_162
timestamp 1698431365
transform 1 0 19488 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_166
timestamp 1698431365
transform 1 0 19936 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_170
timestamp 1698431365
transform 1 0 20384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_174
timestamp 1698431365
transform 1 0 20832 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_176
timestamp 1698431365
transform 1 0 21056 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_206
timestamp 1698431365
transform 1 0 24416 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_31
timestamp 1698431365
transform 1 0 4816 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_45
timestamp 1698431365
transform 1 0 6384 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_84
timestamp 1698431365
transform 1 0 10752 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_86
timestamp 1698431365
transform 1 0 10976 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_95
timestamp 1698431365
transform 1 0 11984 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_104
timestamp 1698431365
transform 1 0 12992 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_111
timestamp 1698431365
transform 1 0 13776 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_115
timestamp 1698431365
transform 1 0 14224 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_119
timestamp 1698431365
transform 1 0 14672 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_139
timestamp 1698431365
transform 1 0 16912 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_143
timestamp 1698431365
transform 1 0 17360 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_145
timestamp 1698431365
transform 1 0 17584 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_148
timestamp 1698431365
transform 1 0 17920 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_150
timestamp 1698431365
transform 1 0 18144 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_161
timestamp 1698431365
transform 1 0 19376 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_165
timestamp 1698431365
transform 1 0 19824 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_169
timestamp 1698431365
transform 1 0 20272 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_173
timestamp 1698431365
transform 1 0 20720 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_227
timestamp 1698431365
transform 1 0 26768 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_231
timestamp 1698431365
transform 1 0 27216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_235
timestamp 1698431365
transform 1 0 27664 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_6
timestamp 1698431365
transform 1 0 2016 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_8
timestamp 1698431365
transform 1 0 2240 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_19
timestamp 1698431365
transform 1 0 3472 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_21
timestamp 1698431365
transform 1 0 3696 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_30
timestamp 1698431365
transform 1 0 4704 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_38
timestamp 1698431365
transform 1 0 5600 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_49
timestamp 1698431365
transform 1 0 6832 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_61
timestamp 1698431365
transform 1 0 8176 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_65
timestamp 1698431365
transform 1 0 8624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_69
timestamp 1698431365
transform 1 0 9072 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_76
timestamp 1698431365
transform 1 0 9856 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_106
timestamp 1698431365
transform 1 0 13216 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_108
timestamp 1698431365
transform 1 0 13440 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_142
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_173
timestamp 1698431365
transform 1 0 20720 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_177
timestamp 1698431365
transform 1 0 21168 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_179
timestamp 1698431365
transform 1 0 21392 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_186
timestamp 1698431365
transform 1 0 22176 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_190
timestamp 1698431365
transform 1 0 22624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_202
timestamp 1698431365
transform 1 0 23968 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_206
timestamp 1698431365
transform 1 0 24416 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_236
timestamp 1698431365
transform 1 0 27776 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_240
timestamp 1698431365
transform 1 0 28224 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_8
timestamp 1698431365
transform 1 0 2240 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_10
timestamp 1698431365
transform 1 0 2464 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_17
timestamp 1698431365
transform 1 0 3248 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_23
timestamp 1698431365
transform 1 0 3920 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_27
timestamp 1698431365
transform 1 0 4368 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_31
timestamp 1698431365
transform 1 0 4816 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_66
timestamp 1698431365
transform 1 0 8736 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_70
timestamp 1698431365
transform 1 0 9184 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_74
timestamp 1698431365
transform 1 0 9632 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_86
timestamp 1698431365
transform 1 0 10976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_90
timestamp 1698431365
transform 1 0 11424 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_98
timestamp 1698431365
transform 1 0 12320 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_100
timestamp 1698431365
transform 1 0 12544 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_103
timestamp 1698431365
transform 1 0 12880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_111
timestamp 1698431365
transform 1 0 13776 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_117
timestamp 1698431365
transform 1 0 14448 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_133
timestamp 1698431365
transform 1 0 16240 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_137
timestamp 1698431365
transform 1 0 16688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_141
timestamp 1698431365
transform 1 0 17136 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_145
timestamp 1698431365
transform 1 0 17584 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_153
timestamp 1698431365
transform 1 0 18480 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_161
timestamp 1698431365
transform 1 0 19376 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_206
timestamp 1698431365
transform 1 0 24416 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_210
timestamp 1698431365
transform 1 0 24864 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_6
timestamp 1698431365
transform 1 0 2016 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_21
timestamp 1698431365
transform 1 0 3696 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_25
timestamp 1698431365
transform 1 0 4144 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_29
timestamp 1698431365
transform 1 0 4592 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_33
timestamp 1698431365
transform 1 0 5040 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_49
timestamp 1698431365
transform 1 0 6832 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_51
timestamp 1698431365
transform 1 0 7056 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_60
timestamp 1698431365
transform 1 0 8064 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_64
timestamp 1698431365
transform 1 0 8512 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_68
timestamp 1698431365
transform 1 0 8960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_101
timestamp 1698431365
transform 1 0 12656 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_115
timestamp 1698431365
transform 1 0 14224 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_124
timestamp 1698431365
transform 1 0 15232 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_128
timestamp 1698431365
transform 1 0 15680 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_132
timestamp 1698431365
transform 1 0 16128 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_136
timestamp 1698431365
transform 1 0 16576 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_153
timestamp 1698431365
transform 1 0 18480 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_157
timestamp 1698431365
transform 1 0 18928 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_163
timestamp 1698431365
transform 1 0 19600 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_167
timestamp 1698431365
transform 1 0 20048 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_177
timestamp 1698431365
transform 1 0 21168 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_181
timestamp 1698431365
transform 1 0 21616 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_185
timestamp 1698431365
transform 1 0 22064 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_189
timestamp 1698431365
transform 1 0 22512 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_200
timestamp 1698431365
transform 1 0 23744 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_204
timestamp 1698431365
transform 1 0 24192 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_208
timestamp 1698431365
transform 1 0 24640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_216
timestamp 1698431365
transform 1 0 25536 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_225
timestamp 1698431365
transform 1 0 26544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_227
timestamp 1698431365
transform 1 0 26768 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_230
timestamp 1698431365
transform 1 0 27104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_234
timestamp 1698431365
transform 1 0 27552 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_238
timestamp 1698431365
transform 1 0 28000 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_240
timestamp 1698431365
transform 1 0 28224 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_31
timestamp 1698431365
transform 1 0 4816 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_47
timestamp 1698431365
transform 1 0 6608 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_101
timestamp 1698431365
transform 1 0 12656 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_136
timestamp 1698431365
transform 1 0 16576 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_140
timestamp 1698431365
transform 1 0 17024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_142
timestamp 1698431365
transform 1 0 17248 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_159
timestamp 1698431365
transform 1 0 19152 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_163
timestamp 1698431365
transform 1 0 19600 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_165
timestamp 1698431365
transform 1 0 19824 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_168
timestamp 1698431365
transform 1 0 20160 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_172
timestamp 1698431365
transform 1 0 20608 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_187
timestamp 1698431365
transform 1 0 22288 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_20
timestamp 1698431365
transform 1 0 3584 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_24
timestamp 1698431365
transform 1 0 4032 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_65
timestamp 1698431365
transform 1 0 8624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_69
timestamp 1698431365
transform 1 0 9072 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_72
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_76
timestamp 1698431365
transform 1 0 9856 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_84
timestamp 1698431365
transform 1 0 10752 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_96
timestamp 1698431365
transform 1 0 12096 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_98
timestamp 1698431365
transform 1 0 12320 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_107
timestamp 1698431365
transform 1 0 13328 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_111
timestamp 1698431365
transform 1 0 13776 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_115
timestamp 1698431365
transform 1 0 14224 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_139
timestamp 1698431365
transform 1 0 16912 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_150
timestamp 1698431365
transform 1 0 18144 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_154
timestamp 1698431365
transform 1 0 18592 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_195
timestamp 1698431365
transform 1 0 23184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_199
timestamp 1698431365
transform 1 0 23632 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_201
timestamp 1698431365
transform 1 0 23856 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_6
timestamp 1698431365
transform 1 0 2016 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_14
timestamp 1698431365
transform 1 0 2912 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_16
timestamp 1698431365
transform 1 0 3136 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_19
timestamp 1698431365
transform 1 0 3472 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_27
timestamp 1698431365
transform 1 0 4368 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_31
timestamp 1698431365
transform 1 0 4816 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_39
timestamp 1698431365
transform 1 0 5712 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_48
timestamp 1698431365
transform 1 0 6720 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_52
timestamp 1698431365
transform 1 0 7168 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_56
timestamp 1698431365
transform 1 0 7616 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_59
timestamp 1698431365
transform 1 0 7952 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_67
timestamp 1698431365
transform 1 0 8848 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_71
timestamp 1698431365
transform 1 0 9296 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_75
timestamp 1698431365
transform 1 0 9744 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_87
timestamp 1698431365
transform 1 0 11088 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_97
timestamp 1698431365
transform 1 0 12208 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_101
timestamp 1698431365
transform 1 0 12656 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_115
timestamp 1698431365
transform 1 0 14224 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_119
timestamp 1698431365
transform 1 0 14672 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_127
timestamp 1698431365
transform 1 0 15568 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_129
timestamp 1698431365
transform 1 0 15792 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_185
timestamp 1698431365
transform 1 0 22064 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_189
timestamp 1698431365
transform 1 0 22512 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_199
timestamp 1698431365
transform 1 0 23632 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_235
timestamp 1698431365
transform 1 0 27664 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_2
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_6
timestamp 1698431365
transform 1 0 2016 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_21
timestamp 1698431365
transform 1 0 3696 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_25
timestamp 1698431365
transform 1 0 4144 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_58
timestamp 1698431365
transform 1 0 7840 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_60
timestamp 1698431365
transform 1 0 8064 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_65
timestamp 1698431365
transform 1 0 8624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_67
timestamp 1698431365
transform 1 0 8848 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_119
timestamp 1698431365
transform 1 0 14672 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_123
timestamp 1698431365
transform 1 0 15120 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_127
timestamp 1698431365
transform 1 0 15568 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_135
timestamp 1698431365
transform 1 0 16464 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_137
timestamp 1698431365
transform 1 0 16688 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_150
timestamp 1698431365
transform 1 0 18144 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_154
timestamp 1698431365
transform 1 0 18592 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_156
timestamp 1698431365
transform 1 0 18816 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_159
timestamp 1698431365
transform 1 0 19152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_163
timestamp 1698431365
transform 1 0 19600 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_167
timestamp 1698431365
transform 1 0 20048 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_171
timestamp 1698431365
transform 1 0 20496 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_175
timestamp 1698431365
transform 1 0 20944 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_179
timestamp 1698431365
transform 1 0 21392 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_181
timestamp 1698431365
transform 1 0 21616 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_31
timestamp 1698431365
transform 1 0 4816 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_37
timestamp 1698431365
transform 1 0 5488 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_53
timestamp 1698431365
transform 1 0 7280 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_57
timestamp 1698431365
transform 1 0 7728 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_64
timestamp 1698431365
transform 1 0 8512 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_74
timestamp 1698431365
transform 1 0 9632 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_78
timestamp 1698431365
transform 1 0 10080 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_80
timestamp 1698431365
transform 1 0 10304 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_83
timestamp 1698431365
transform 1 0 10640 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_91
timestamp 1698431365
transform 1 0 11536 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_95
timestamp 1698431365
transform 1 0 11984 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_103
timestamp 1698431365
transform 1 0 12880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_116
timestamp 1698431365
transform 1 0 14336 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_122
timestamp 1698431365
transform 1 0 15008 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_141
timestamp 1698431365
transform 1 0 17136 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_145
timestamp 1698431365
transform 1 0 17584 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_149
timestamp 1698431365
transform 1 0 18032 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_167
timestamp 1698431365
transform 1 0 20048 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_171
timestamp 1698431365
transform 1 0 20496 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_179
timestamp 1698431365
transform 1 0 21392 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_212
timestamp 1698431365
transform 1 0 25088 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_216
timestamp 1698431365
transform 1 0 25536 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_220
timestamp 1698431365
transform 1 0 25984 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_238
timestamp 1698431365
transform 1 0 28000 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_240
timestamp 1698431365
transform 1 0 28224 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_4
timestamp 1698431365
transform 1 0 1792 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_67
timestamp 1698431365
transform 1 0 8848 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_69
timestamp 1698431365
transform 1 0 9072 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_81
timestamp 1698431365
transform 1 0 10416 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_87
timestamp 1698431365
transform 1 0 11088 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_91
timestamp 1698431365
transform 1 0 11536 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_93
timestamp 1698431365
transform 1 0 11760 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_171
timestamp 1698431365
transform 1 0 20496 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_175
timestamp 1698431365
transform 1 0 20944 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_177
timestamp 1698431365
transform 1 0 21168 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_180
timestamp 1698431365
transform 1 0 21504 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_216
timestamp 1698431365
transform 1 0 25536 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_231
timestamp 1698431365
transform 1 0 27216 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_235
timestamp 1698431365
transform 1 0 27664 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_239
timestamp 1698431365
transform 1 0 28112 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_8
timestamp 1698431365
transform 1 0 2240 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_10
timestamp 1698431365
transform 1 0 2464 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_13
timestamp 1698431365
transform 1 0 2800 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_17
timestamp 1698431365
transform 1 0 3248 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_21
timestamp 1698431365
transform 1 0 3696 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_25
timestamp 1698431365
transform 1 0 4144 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_31
timestamp 1698431365
transform 1 0 4816 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_53
timestamp 1698431365
transform 1 0 7280 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_57
timestamp 1698431365
transform 1 0 7728 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_65
timestamp 1698431365
transform 1 0 8624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_69
timestamp 1698431365
transform 1 0 9072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_79
timestamp 1698431365
transform 1 0 10192 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_83
timestamp 1698431365
transform 1 0 10640 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_87
timestamp 1698431365
transform 1 0 11088 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_90
timestamp 1698431365
transform 1 0 11424 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_98
timestamp 1698431365
transform 1 0 12320 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_101
timestamp 1698431365
transform 1 0 12656 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_154
timestamp 1698431365
transform 1 0 18592 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_158
timestamp 1698431365
transform 1 0 19040 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_177
timestamp 1698431365
transform 1 0 21168 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_207
timestamp 1698431365
transform 1 0 24528 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_211
timestamp 1698431365
transform 1 0 24976 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_6
timestamp 1698431365
transform 1 0 2016 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_21
timestamp 1698431365
transform 1 0 3696 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_54
timestamp 1698431365
transform 1 0 7392 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_58
timestamp 1698431365
transform 1 0 7840 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_88
timestamp 1698431365
transform 1 0 11200 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_97
timestamp 1698431365
transform 1 0 12208 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_101
timestamp 1698431365
transform 1 0 12656 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_105
timestamp 1698431365
transform 1 0 13104 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_118
timestamp 1698431365
transform 1 0 14560 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_122
timestamp 1698431365
transform 1 0 15008 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_137
timestamp 1698431365
transform 1 0 16688 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_139
timestamp 1698431365
transform 1 0 16912 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_193
timestamp 1698431365
transform 1 0 22960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_216
timestamp 1698431365
transform 1 0 25536 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_222
timestamp 1698431365
transform 1 0 26208 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_231
timestamp 1698431365
transform 1 0 27216 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_235
timestamp 1698431365
transform 1 0 27664 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_31
timestamp 1698431365
transform 1 0 4816 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_54
timestamp 1698431365
transform 1 0 7392 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_58
timestamp 1698431365
transform 1 0 7840 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_99
timestamp 1698431365
transform 1 0 12432 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_117
timestamp 1698431365
transform 1 0 14448 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_166
timestamp 1698431365
transform 1 0 19936 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_170
timestamp 1698431365
transform 1 0 20384 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_174
timestamp 1698431365
transform 1 0 20832 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_181
timestamp 1698431365
transform 1 0 21616 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_201
timestamp 1698431365
transform 1 0 23856 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_205
timestamp 1698431365
transform 1 0 24304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_209
timestamp 1698431365
transform 1 0 24752 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_213
timestamp 1698431365
transform 1 0 25200 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_14
timestamp 1698431365
transform 1 0 2912 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_21
timestamp 1698431365
transform 1 0 3696 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_27
timestamp 1698431365
transform 1 0 4368 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_60
timestamp 1698431365
transform 1 0 8064 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_64
timestamp 1698431365
transform 1 0 8512 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_76
timestamp 1698431365
transform 1 0 9856 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_80
timestamp 1698431365
transform 1 0 10304 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_96
timestamp 1698431365
transform 1 0 12096 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_116
timestamp 1698431365
transform 1 0 14336 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_120
timestamp 1698431365
transform 1 0 14784 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_122
timestamp 1698431365
transform 1 0 15008 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_125
timestamp 1698431365
transform 1 0 15344 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_131
timestamp 1698431365
transform 1 0 16016 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_135
timestamp 1698431365
transform 1 0 16464 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_139
timestamp 1698431365
transform 1 0 16912 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_153
timestamp 1698431365
transform 1 0 18480 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_157
timestamp 1698431365
transform 1 0 18928 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_163
timestamp 1698431365
transform 1 0 19600 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_167
timestamp 1698431365
transform 1 0 20048 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_171
timestamp 1698431365
transform 1 0 20496 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_191
timestamp 1698431365
transform 1 0 22736 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_195
timestamp 1698431365
transform 1 0 23184 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_208
timestamp 1698431365
transform 1 0 24640 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_2
timestamp 1698431365
transform 1 0 1568 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_6
timestamp 1698431365
transform 1 0 2016 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_10
timestamp 1698431365
transform 1 0 2464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_16
timestamp 1698431365
transform 1 0 3136 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_22
timestamp 1698431365
transform 1 0 3808 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_26
timestamp 1698431365
transform 1 0 4256 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_30
timestamp 1698431365
transform 1 0 4704 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_33
timestamp 1698431365
transform 1 0 5040 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_41
timestamp 1698431365
transform 1 0 5936 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_45
timestamp 1698431365
transform 1 0 6384 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_47
timestamp 1698431365
transform 1 0 6608 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_50
timestamp 1698431365
transform 1 0 6944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_54
timestamp 1698431365
transform 1 0 7392 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_62
timestamp 1698431365
transform 1 0 8288 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_64
timestamp 1698431365
transform 1 0 8512 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_67
timestamp 1698431365
transform 1 0 8848 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_71
timestamp 1698431365
transform 1 0 9296 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_75
timestamp 1698431365
transform 1 0 9744 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_79
timestamp 1698431365
transform 1 0 10192 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_83
timestamp 1698431365
transform 1 0 10640 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_87
timestamp 1698431365
transform 1 0 11088 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_91
timestamp 1698431365
transform 1 0 11536 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_94
timestamp 1698431365
transform 1 0 11872 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_102
timestamp 1698431365
transform 1 0 12768 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_104
timestamp 1698431365
transform 1 0 12992 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_111
timestamp 1698431365
transform 1 0 13776 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_115
timestamp 1698431365
transform 1 0 14224 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_123
timestamp 1698431365
transform 1 0 15120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_151
timestamp 1698431365
transform 1 0 18256 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_159
timestamp 1698431365
transform 1 0 19152 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_163
timestamp 1698431365
transform 1 0 19600 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_167
timestamp 1698431365
transform 1 0 20048 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_171
timestamp 1698431365
transform 1 0 20496 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_214
timestamp 1698431365
transform 1 0 25312 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_235
timestamp 1698431365
transform 1 0 27664 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_239
timestamp 1698431365
transform 1 0 28112 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_18
timestamp 1698431365
transform 1 0 3360 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_27
timestamp 1698431365
transform 1 0 4368 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_33
timestamp 1698431365
transform 1 0 5040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_53
timestamp 1698431365
transform 1 0 7280 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_57
timestamp 1698431365
transform 1 0 7728 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_81
timestamp 1698431365
transform 1 0 10416 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_95
timestamp 1698431365
transform 1 0 11984 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_97
timestamp 1698431365
transform 1 0 12208 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_100
timestamp 1698431365
transform 1 0 12544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_104
timestamp 1698431365
transform 1 0 12992 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_128
timestamp 1698431365
transform 1 0 15680 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_132
timestamp 1698431365
transform 1 0 16128 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_136
timestamp 1698431365
transform 1 0 16576 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_171
timestamp 1698431365
transform 1 0 20496 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_175
timestamp 1698431365
transform 1 0 20944 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_179
timestamp 1698431365
transform 1 0 21392 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_183
timestamp 1698431365
transform 1 0 21840 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_186
timestamp 1698431365
transform 1 0 22176 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_190
timestamp 1698431365
transform 1 0 22624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_194
timestamp 1698431365
transform 1 0 23072 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_198
timestamp 1698431365
transform 1 0 23520 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_202
timestamp 1698431365
transform 1 0 23968 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_206
timestamp 1698431365
transform 1 0 24416 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_212
timestamp 1698431365
transform 1 0 25088 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_216
timestamp 1698431365
transform 1 0 25536 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_219
timestamp 1698431365
transform 1 0 25872 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_223
timestamp 1698431365
transform 1 0 26320 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_225
timestamp 1698431365
transform 1 0 26544 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_228
timestamp 1698431365
transform 1 0 26880 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_232
timestamp 1698431365
transform 1 0 27328 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_236
timestamp 1698431365
transform 1 0 27776 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_238
timestamp 1698431365
transform 1 0 28000 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_66
timestamp 1698431365
transform 1 0 8736 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_96
timestamp 1698431365
transform 1 0 12096 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_136
timestamp 1698431365
transform 1 0 16576 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_140
timestamp 1698431365
transform 1 0 17024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_144
timestamp 1698431365
transform 1 0 17472 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_155
timestamp 1698431365
transform 1 0 18704 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_161
timestamp 1698431365
transform 1 0 19376 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_172
timestamp 1698431365
transform 1 0 20608 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_174
timestamp 1698431365
transform 1 0 20832 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_181
timestamp 1698431365
transform 1 0 21616 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_185
timestamp 1698431365
transform 1 0 22064 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_189
timestamp 1698431365
transform 1 0 22512 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_219
timestamp 1698431365
transform 1 0 25872 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_221
timestamp 1698431365
transform 1 0 26096 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_230
timestamp 1698431365
transform 1 0 27104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_234
timestamp 1698431365
transform 1 0 27552 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_238
timestamp 1698431365
transform 1 0 28000 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_240
timestamp 1698431365
transform 1 0 28224 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_2
timestamp 1698431365
transform 1 0 1568 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_6
timestamp 1698431365
transform 1 0 2016 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_16
timestamp 1698431365
transform 1 0 3136 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_18
timestamp 1698431365
transform 1 0 3360 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_33
timestamp 1698431365
transform 1 0 5040 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_37
timestamp 1698431365
transform 1 0 5488 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_41
timestamp 1698431365
transform 1 0 5936 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_61
timestamp 1698431365
transform 1 0 8176 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_63
timestamp 1698431365
transform 1 0 8400 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_66
timestamp 1698431365
transform 1 0 8736 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_72
timestamp 1698431365
transform 1 0 9408 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_74
timestamp 1698431365
transform 1 0 9632 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_91
timestamp 1698431365
transform 1 0 11536 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_100
timestamp 1698431365
transform 1 0 12544 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_104
timestamp 1698431365
transform 1 0 12992 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_133
timestamp 1698431365
transform 1 0 16240 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_137
timestamp 1698431365
transform 1 0 16688 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_139
timestamp 1698431365
transform 1 0 16912 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_142
timestamp 1698431365
transform 1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_146
timestamp 1698431365
transform 1 0 17696 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_152
timestamp 1698431365
transform 1 0 18368 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_154
timestamp 1698431365
transform 1 0 18592 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_184
timestamp 1698431365
transform 1 0 21952 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_188
timestamp 1698431365
transform 1 0 22400 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_192
timestamp 1698431365
transform 1 0 22848 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_196
timestamp 1698431365
transform 1 0 23296 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_200
timestamp 1698431365
transform 1 0 23744 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_204
timestamp 1698431365
transform 1 0 24192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_208
timestamp 1698431365
transform 1 0 24640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_212
timestamp 1698431365
transform 1 0 25088 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_216
timestamp 1698431365
transform 1 0 25536 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_218
timestamp 1698431365
transform 1 0 25760 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_235
timestamp 1698431365
transform 1 0 27664 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_2
timestamp 1698431365
transform 1 0 1568 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_6
timestamp 1698431365
transform 1 0 2016 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_15
timestamp 1698431365
transform 1 0 3024 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_17
timestamp 1698431365
transform 1 0 3248 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_26
timestamp 1698431365
transform 1 0 4256 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_28
timestamp 1698431365
transform 1 0 4480 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_31
timestamp 1698431365
transform 1 0 4816 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_66
timestamp 1698431365
transform 1 0 8736 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_72
timestamp 1698431365
transform 1 0 9408 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_107
timestamp 1698431365
transform 1 0 13328 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_112
timestamp 1698431365
transform 1 0 13888 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_164
timestamp 1698431365
transform 1 0 19712 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_168
timestamp 1698431365
transform 1 0 20160 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_177
timestamp 1698431365
transform 1 0 21168 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_181
timestamp 1698431365
transform 1 0 21616 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_197
timestamp 1698431365
transform 1 0 23408 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_201
timestamp 1698431365
transform 1 0 23856 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_203
timestamp 1698431365
transform 1 0 24080 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_22
timestamp 1698431365
transform 1 0 3808 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_26
timestamp 1698431365
transform 1 0 4256 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_30
timestamp 1698431365
transform 1 0 4704 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_33
timestamp 1698431365
transform 1 0 5040 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_37
timestamp 1698431365
transform 1 0 5488 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_43
timestamp 1698431365
transform 1 0 6160 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_47
timestamp 1698431365
transform 1 0 6608 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_49
timestamp 1698431365
transform 1 0 6832 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_52
timestamp 1698431365
transform 1 0 7168 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_56
timestamp 1698431365
transform 1 0 7616 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_158
timestamp 1698431365
transform 1 0 19040 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_162
timestamp 1698431365
transform 1 0 19488 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_166
timestamp 1698431365
transform 1 0 19936 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_170
timestamp 1698431365
transform 1 0 20384 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_174
timestamp 1698431365
transform 1 0 20832 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_178
timestamp 1698431365
transform 1 0 21280 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_180
timestamp 1698431365
transform 1 0 21504 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_31
timestamp 1698431365
transform 1 0 4816 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_47
timestamp 1698431365
transform 1 0 6608 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_51
timestamp 1698431365
transform 1 0 7056 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_55
timestamp 1698431365
transform 1 0 7504 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_57
timestamp 1698431365
transform 1 0 7728 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_60
timestamp 1698431365
transform 1 0 8064 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_90
timestamp 1698431365
transform 1 0 11424 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_107
timestamp 1698431365
transform 1 0 13328 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_173
timestamp 1698431365
transform 1 0 20720 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_183
timestamp 1698431365
transform 1 0 21840 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_187
timestamp 1698431365
transform 1 0 22288 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_194
timestamp 1698431365
transform 1 0 23072 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_198
timestamp 1698431365
transform 1 0 23520 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_202
timestamp 1698431365
transform 1 0 23968 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_206
timestamp 1698431365
transform 1 0 24416 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_210
timestamp 1698431365
transform 1 0 24864 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_214
timestamp 1698431365
transform 1 0 25312 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_218
timestamp 1698431365
transform 1 0 25760 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_222
timestamp 1698431365
transform 1 0 26208 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_226
timestamp 1698431365
transform 1 0 26656 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_230
timestamp 1698431365
transform 1 0 27104 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_234
timestamp 1698431365
transform 1 0 27552 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_238
timestamp 1698431365
transform 1 0 28000 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_99_2
timestamp 1698431365
transform 1 0 1568 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_12
timestamp 1698431365
transform 1 0 2688 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_22
timestamp 1698431365
transform 1 0 3808 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_26
timestamp 1698431365
transform 1 0 4256 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_60
timestamp 1698431365
transform 1 0 8064 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_64
timestamp 1698431365
transform 1 0 8512 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_72
timestamp 1698431365
transform 1 0 9408 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_137
timestamp 1698431365
transform 1 0 16688 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_139
timestamp 1698431365
transform 1 0 16912 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_142
timestamp 1698431365
transform 1 0 17248 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_194
timestamp 1698431365
transform 1 0 23072 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_198
timestamp 1698431365
transform 1 0 23520 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_202
timestamp 1698431365
transform 1 0 23968 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_206
timestamp 1698431365
transform 1 0 24416 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_212
timestamp 1698431365
transform 1 0 25088 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_216
timestamp 1698431365
transform 1 0 25536 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_220
timestamp 1698431365
transform 1 0 25984 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_224
timestamp 1698431365
transform 1 0 26432 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_228
timestamp 1698431365
transform 1 0 26880 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_232
timestamp 1698431365
transform 1 0 27328 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_236
timestamp 1698431365
transform 1 0 27776 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_240
timestamp 1698431365
transform 1 0 28224 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_8
timestamp 1698431365
transform 1 0 2240 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_28
timestamp 1698431365
transform 1 0 4480 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_32
timestamp 1698431365
transform 1 0 4928 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_37
timestamp 1698431365
transform 1 0 5488 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_44
timestamp 1698431365
transform 1 0 6272 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_48
timestamp 1698431365
transform 1 0 6720 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_100_52
timestamp 1698431365
transform 1 0 7168 0 1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_68
timestamp 1698431365
transform 1 0 8960 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_99
timestamp 1698431365
transform 1 0 12432 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_107
timestamp 1698431365
transform 1 0 13328 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_173
timestamp 1698431365
transform 1 0 20720 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_183
timestamp 1698431365
transform 1 0 21840 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_190
timestamp 1698431365
transform 1 0 22624 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_192
timestamp 1698431365
transform 1 0 22848 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_199
timestamp 1698431365
transform 1 0 23632 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_209
timestamp 1698431365
transform 1 0 24752 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_227
timestamp 1698431365
transform 1 0 26768 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_236
timestamp 1698431365
transform 1 0 27776 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_240
timestamp 1698431365
transform 1 0 28224 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_2
timestamp 1698431365
transform 1 0 1568 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_6
timestamp 1698431365
transform 1 0 2016 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_8
timestamp 1698431365
transform 1 0 2240 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_35
timestamp 1698431365
transform 1 0 5264 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_41
timestamp 1698431365
transform 1 0 5936 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_45
timestamp 1698431365
transform 1 0 6384 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_59
timestamp 1698431365
transform 1 0 7952 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_67
timestamp 1698431365
transform 1 0 8848 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_69
timestamp 1698431365
transform 1 0 9072 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_72
timestamp 1698431365
transform 1 0 9408 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_76
timestamp 1698431365
transform 1 0 9856 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_78
timestamp 1698431365
transform 1 0 10080 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_89
timestamp 1698431365
transform 1 0 11312 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_93
timestamp 1698431365
transform 1 0 11760 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_155
timestamp 1698431365
transform 1 0 18704 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_157
timestamp 1698431365
transform 1 0 18928 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_203
timestamp 1698431365
transform 1 0 24080 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_43
timestamp 1698431365
transform 1 0 6160 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_77
timestamp 1698431365
transform 1 0 9968 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_81
timestamp 1698431365
transform 1 0 10416 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_85
timestamp 1698431365
transform 1 0 10864 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_89
timestamp 1698431365
transform 1 0 11312 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_93
timestamp 1698431365
transform 1 0 11760 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_97
timestamp 1698431365
transform 1 0 12208 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_101
timestamp 1698431365
transform 1 0 12656 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_107
timestamp 1698431365
transform 1 0 13328 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_111
timestamp 1698431365
transform 1 0 13776 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_115
timestamp 1698431365
transform 1 0 14224 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_150
timestamp 1698431365
transform 1 0 18144 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_154
timestamp 1698431365
transform 1 0 18592 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_158
timestamp 1698431365
transform 1 0 19040 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_162
timestamp 1698431365
transform 1 0 19488 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_166
timestamp 1698431365
transform 1 0 19936 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_204
timestamp 1698431365
transform 1 0 24192 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_240
timestamp 1698431365
transform 1 0 28224 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_2
timestamp 1698431365
transform 1 0 1568 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_6
timestamp 1698431365
transform 1 0 2016 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_58
timestamp 1698431365
transform 1 0 7840 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_103_62
timestamp 1698431365
transform 1 0 8288 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_72
timestamp 1698431365
transform 1 0 9408 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_78
timestamp 1698431365
transform 1 0 10080 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_82
timestamp 1698431365
transform 1 0 10528 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_94
timestamp 1698431365
transform 1 0 11872 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_96
timestamp 1698431365
transform 1 0 12096 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_123
timestamp 1698431365
transform 1 0 15120 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_125
timestamp 1698431365
transform 1 0 15344 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_139
timestamp 1698431365
transform 1 0 16912 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_142
timestamp 1698431365
transform 1 0 17248 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_146
timestamp 1698431365
transform 1 0 17696 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_150
timestamp 1698431365
transform 1 0 18144 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_152
timestamp 1698431365
transform 1 0 18368 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_155
timestamp 1698431365
transform 1 0 18704 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_159
timestamp 1698431365
transform 1 0 19152 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_163
timestamp 1698431365
transform 1 0 19600 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_236
timestamp 1698431365
transform 1 0 27776 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_240
timestamp 1698431365
transform 1 0 28224 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_8
timestamp 1698431365
transform 1 0 2240 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_12
timestamp 1698431365
transform 1 0 2688 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_15
timestamp 1698431365
transform 1 0 3024 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_19
timestamp 1698431365
transform 1 0 3472 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_23
timestamp 1698431365
transform 1 0 3920 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_27
timestamp 1698431365
transform 1 0 4368 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_31
timestamp 1698431365
transform 1 0 4816 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_51
timestamp 1698431365
transform 1 0 7056 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_55
timestamp 1698431365
transform 1 0 7504 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104_59
timestamp 1698431365
transform 1 0 7952 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_67
timestamp 1698431365
transform 1 0 8848 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_107
timestamp 1698431365
transform 1 0 13328 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_111
timestamp 1698431365
transform 1 0 13776 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_114
timestamp 1698431365
transform 1 0 14112 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_123
timestamp 1698431365
transform 1 0 15120 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_125
timestamp 1698431365
transform 1 0 15344 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_128
timestamp 1698431365
transform 1 0 15680 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_132
timestamp 1698431365
transform 1 0 16128 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_136
timestamp 1698431365
transform 1 0 16576 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_142
timestamp 1698431365
transform 1 0 17248 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_154
timestamp 1698431365
transform 1 0 18592 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_183
timestamp 1698431365
transform 1 0 21840 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_214
timestamp 1698431365
transform 1 0 25312 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_216
timestamp 1698431365
transform 1 0 25536 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_225
timestamp 1698431365
transform 1 0 26544 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_235
timestamp 1698431365
transform 1 0 27664 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_239
timestamp 1698431365
transform 1 0 28112 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_2
timestamp 1698431365
transform 1 0 1568 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_105_12
timestamp 1698431365
transform 1 0 2688 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_28
timestamp 1698431365
transform 1 0 4480 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_32
timestamp 1698431365
transform 1 0 4928 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_34
timestamp 1698431365
transform 1 0 5152 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_37
timestamp 1698431365
transform 1 0 5488 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_105_41
timestamp 1698431365
transform 1 0 5936 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_57
timestamp 1698431365
transform 1 0 7728 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_65
timestamp 1698431365
transform 1 0 8624 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_67
timestamp 1698431365
transform 1 0 8848 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_72
timestamp 1698431365
transform 1 0 9408 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_74
timestamp 1698431365
transform 1 0 9632 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_77
timestamp 1698431365
transform 1 0 9968 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_81
timestamp 1698431365
transform 1 0 10416 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_134
timestamp 1698431365
transform 1 0 16352 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_142
timestamp 1698431365
transform 1 0 17248 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_162
timestamp 1698431365
transform 1 0 19488 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_194
timestamp 1698431365
transform 1 0 23072 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_208
timestamp 1698431365
transform 1 0 24640 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_236
timestamp 1698431365
transform 1 0 27776 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_240
timestamp 1698431365
transform 1 0 28224 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_2
timestamp 1698431365
transform 1 0 1568 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_6
timestamp 1698431365
transform 1 0 2016 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_8
timestamp 1698431365
transform 1 0 2240 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_37
timestamp 1698431365
transform 1 0 5488 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_41
timestamp 1698431365
transform 1 0 5936 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_99
timestamp 1698431365
transform 1 0 12432 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_107
timestamp 1698431365
transform 1 0 13328 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_138
timestamp 1698431365
transform 1 0 16800 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_167
timestamp 1698431365
transform 1 0 20048 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_169
timestamp 1698431365
transform 1 0 20272 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_193
timestamp 1698431365
transform 1 0 22960 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_197
timestamp 1698431365
transform 1 0 23408 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_201
timestamp 1698431365
transform 1 0 23856 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_203
timestamp 1698431365
transform 1 0 24080 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_239
timestamp 1698431365
transform 1 0 28112 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_8
timestamp 1698431365
transform 1 0 2240 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_12
timestamp 1698431365
transform 1 0 2688 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_44
timestamp 1698431365
transform 1 0 6272 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_48
timestamp 1698431365
transform 1 0 6720 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_51
timestamp 1698431365
transform 1 0 7056 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_55
timestamp 1698431365
transform 1 0 7504 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_67
timestamp 1698431365
transform 1 0 8848 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_69
timestamp 1698431365
transform 1 0 9072 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_122
timestamp 1698431365
transform 1 0 15008 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_126
timestamp 1698431365
transform 1 0 15456 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_128
timestamp 1698431365
transform 1 0 15680 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_142
timestamp 1698431365
transform 1 0 17248 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_198
timestamp 1698431365
transform 1 0 23520 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_212
timestamp 1698431365
transform 1 0 25088 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_238
timestamp 1698431365
transform 1 0 28000 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_240
timestamp 1698431365
transform 1 0 28224 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_108_2
timestamp 1698431365
transform 1 0 1568 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_32
timestamp 1698431365
transform 1 0 4928 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_34
timestamp 1698431365
transform 1 0 5152 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_37
timestamp 1698431365
transform 1 0 5488 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_41
timestamp 1698431365
transform 1 0 5936 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_44
timestamp 1698431365
transform 1 0 6272 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_48
timestamp 1698431365
transform 1 0 6720 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_52
timestamp 1698431365
transform 1 0 7168 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_56
timestamp 1698431365
transform 1 0 7616 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_60
timestamp 1698431365
transform 1 0 8064 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_80
timestamp 1698431365
transform 1 0 10304 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_82
timestamp 1698431365
transform 1 0 10528 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_91
timestamp 1698431365
transform 1 0 11536 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_93
timestamp 1698431365
transform 1 0 11760 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_102
timestamp 1698431365
transform 1 0 12768 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_104
timestamp 1698431365
transform 1 0 12992 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_107
timestamp 1698431365
transform 1 0 13328 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_152
timestamp 1698431365
transform 1 0 18368 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_154
timestamp 1698431365
transform 1 0 18592 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_171
timestamp 1698431365
transform 1 0 20496 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_190
timestamp 1698431365
transform 1 0 22624 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_194
timestamp 1698431365
transform 1 0 23072 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_2
timestamp 1698431365
transform 1 0 1568 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_109_6
timestamp 1698431365
transform 1 0 2016 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_22
timestamp 1698431365
transform 1 0 3808 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_26
timestamp 1698431365
transform 1 0 4256 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_126
timestamp 1698431365
transform 1 0 15456 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_139
timestamp 1698431365
transform 1 0 16912 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_142
timestamp 1698431365
transform 1 0 17248 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_154
timestamp 1698431365
transform 1 0 18592 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_158
timestamp 1698431365
transform 1 0 19040 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_160
timestamp 1698431365
transform 1 0 19264 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_163
timestamp 1698431365
transform 1 0 19600 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_167
timestamp 1698431365
transform 1 0 20048 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_171
timestamp 1698431365
transform 1 0 20496 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_175
timestamp 1698431365
transform 1 0 20944 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_179
timestamp 1698431365
transform 1 0 21392 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_109_183
timestamp 1698431365
transform 1 0 21840 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_199
timestamp 1698431365
transform 1 0 23632 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_212
timestamp 1698431365
transform 1 0 25088 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_214
timestamp 1698431365
transform 1 0 25312 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_223
timestamp 1698431365
transform 1 0 26320 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_237
timestamp 1698431365
transform 1 0 27888 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_8
timestamp 1698431365
transform 1 0 2240 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_15
timestamp 1698431365
transform 1 0 3024 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_110_19
timestamp 1698431365
transform 1 0 3472 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_37
timestamp 1698431365
transform 1 0 5488 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_41
timestamp 1698431365
transform 1 0 5936 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_45
timestamp 1698431365
transform 1 0 6384 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_49
timestamp 1698431365
transform 1 0 6832 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_51
timestamp 1698431365
transform 1 0 7056 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_54
timestamp 1698431365
transform 1 0 7392 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_66
timestamp 1698431365
transform 1 0 8736 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_75
timestamp 1698431365
transform 1 0 9744 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_156
timestamp 1698431365
transform 1 0 18816 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_162
timestamp 1698431365
transform 1 0 19488 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_110_177
timestamp 1698431365
transform 1 0 21168 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_185
timestamp 1698431365
transform 1 0 22064 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_110_197
timestamp 1698431365
transform 1 0 23408 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_205
timestamp 1698431365
transform 1 0 24304 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_31
timestamp 1698431365
transform 1 0 4816 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_111_35
timestamp 1698431365
transform 1 0 5264 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_43
timestamp 1698431365
transform 1 0 6160 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_47
timestamp 1698431365
transform 1 0 6608 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_50
timestamp 1698431365
transform 1 0 6944 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_54
timestamp 1698431365
transform 1 0 7392 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_58
timestamp 1698431365
transform 1 0 7840 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_62
timestamp 1698431365
transform 1 0 8288 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_66
timestamp 1698431365
transform 1 0 8736 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_72
timestamp 1698431365
transform 1 0 9408 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_74
timestamp 1698431365
transform 1 0 9632 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_125
timestamp 1698431365
transform 1 0 15344 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_136
timestamp 1698431365
transform 1 0 16576 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_142
timestamp 1698431365
transform 1 0 17248 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_161
timestamp 1698431365
transform 1 0 19376 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_111_165
timestamp 1698431365
transform 1 0 19824 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_173
timestamp 1698431365
transform 1 0 20720 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_177
timestamp 1698431365
transform 1 0 21168 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_209
timestamp 1698431365
transform 1 0 24752 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_220
timestamp 1698431365
transform 1 0 25984 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_112_2
timestamp 1698431365
transform 1 0 1568 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_112_18
timestamp 1698431365
transform 1 0 3360 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_26
timestamp 1698431365
transform 1 0 4256 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_30
timestamp 1698431365
transform 1 0 4704 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_33
timestamp 1698431365
transform 1 0 5040 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_68
timestamp 1698431365
transform 1 0 8960 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_72
timestamp 1698431365
transform 1 0 9408 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_75
timestamp 1698431365
transform 1 0 9744 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_115
timestamp 1698431365
transform 1 0 14224 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_158
timestamp 1698431365
transform 1 0 19040 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_170
timestamp 1698431365
transform 1 0 20384 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_174
timestamp 1698431365
transform 1 0 20832 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_177
timestamp 1698431365
transform 1 0 21168 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_198
timestamp 1698431365
transform 1 0 23520 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_200
timestamp 1698431365
transform 1 0 23744 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_113_2
timestamp 1698431365
transform 1 0 1568 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_113_18
timestamp 1698431365
transform 1 0 3360 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_26
timestamp 1698431365
transform 1 0 4256 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_37
timestamp 1698431365
transform 1 0 5488 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_58
timestamp 1698431365
transform 1 0 7840 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_72
timestamp 1698431365
transform 1 0 9408 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_115
timestamp 1698431365
transform 1 0 14224 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_117
timestamp 1698431365
transform 1 0 14448 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_130
timestamp 1698431365
transform 1 0 15904 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_134
timestamp 1698431365
transform 1 0 16352 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_138
timestamp 1698431365
transform 1 0 16800 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_142
timestamp 1698431365
transform 1 0 17248 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_146
timestamp 1698431365
transform 1 0 17696 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_150
timestamp 1698431365
transform 1 0 18144 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_154
timestamp 1698431365
transform 1 0 18592 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_158
timestamp 1698431365
transform 1 0 19040 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_160
timestamp 1698431365
transform 1 0 19264 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_180
timestamp 1698431365
transform 1 0 21504 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_186
timestamp 1698431365
transform 1 0 22176 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_188
timestamp 1698431365
transform 1 0 22400 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_194
timestamp 1698431365
transform 1 0 23072 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_113_200
timestamp 1698431365
transform 1 0 23744 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_208
timestamp 1698431365
transform 1 0 24640 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_113_212
timestamp 1698431365
transform 1 0 25088 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_220
timestamp 1698431365
transform 1 0 25984 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_224
timestamp 1698431365
transform 1 0 26432 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_31
timestamp 1698431365
transform 1 0 4816 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_55
timestamp 1698431365
transform 1 0 7504 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_86
timestamp 1698431365
transform 1 0 10976 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_92
timestamp 1698431365
transform 1 0 11648 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_143
timestamp 1698431365
transform 1 0 17360 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_145
timestamp 1698431365
transform 1 0 17584 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_114_163
timestamp 1698431365
transform 1 0 19600 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_171
timestamp 1698431365
transform 1 0 20496 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_177
timestamp 1698431365
transform 1 0 21168 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_181
timestamp 1698431365
transform 1 0 21616 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_207
timestamp 1698431365
transform 1 0 24528 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_233
timestamp 1698431365
transform 1 0 27440 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_237
timestamp 1698431365
transform 1 0 27888 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_2
timestamp 1698431365
transform 1 0 1568 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_6
timestamp 1698431365
transform 1 0 2016 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_8
timestamp 1698431365
transform 1 0 2240 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_11
timestamp 1698431365
transform 1 0 2576 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_72
timestamp 1698431365
transform 1 0 9408 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_74
timestamp 1698431365
transform 1 0 9632 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_135
timestamp 1698431365
transform 1 0 16464 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_139
timestamp 1698431365
transform 1 0 16912 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_142
timestamp 1698431365
transform 1 0 17248 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_151
timestamp 1698431365
transform 1 0 18256 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_155
timestamp 1698431365
transform 1 0 18704 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_115_159
timestamp 1698431365
transform 1 0 19152 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_167
timestamp 1698431365
transform 1 0 20048 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_176
timestamp 1698431365
transform 1 0 21056 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_180
timestamp 1698431365
transform 1 0 21504 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_182
timestamp 1698431365
transform 1 0 21728 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_239
timestamp 1698431365
transform 1 0 28112 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_31
timestamp 1698431365
transform 1 0 4816 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_37
timestamp 1698431365
transform 1 0 5488 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_46
timestamp 1698431365
transform 1 0 6496 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_52
timestamp 1698431365
transform 1 0 7168 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_98
timestamp 1698431365
transform 1 0 12320 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_102
timestamp 1698431365
transform 1 0 12768 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_104
timestamp 1698431365
transform 1 0 12992 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_107
timestamp 1698431365
transform 1 0 13328 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_109
timestamp 1698431365
transform 1 0 13552 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_125
timestamp 1698431365
transform 1 0 15344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_156
timestamp 1698431365
transform 1 0 18816 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_160
timestamp 1698431365
transform 1 0 19264 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_172
timestamp 1698431365
transform 1 0 20608 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_174
timestamp 1698431365
transform 1 0 20832 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_194
timestamp 1698431365
transform 1 0 23072 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_205
timestamp 1698431365
transform 1 0 24304 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_213
timestamp 1698431365
transform 1 0 25200 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_232
timestamp 1698431365
transform 1 0 27328 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_240
timestamp 1698431365
transform 1 0 28224 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_117_2
timestamp 1698431365
transform 1 0 1568 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_18
timestamp 1698431365
transform 1 0 3360 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_22
timestamp 1698431365
transform 1 0 3808 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_25
timestamp 1698431365
transform 1 0 4144 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_60
timestamp 1698431365
transform 1 0 8064 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_85
timestamp 1698431365
transform 1 0 10864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_89
timestamp 1698431365
transform 1 0 11312 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_109
timestamp 1698431365
transform 1 0 13552 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_111
timestamp 1698431365
transform 1 0 13776 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_137
timestamp 1698431365
transform 1 0 16688 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_139
timestamp 1698431365
transform 1 0 16912 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_192
timestamp 1698431365
transform 1 0 22848 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_117_196
timestamp 1698431365
transform 1 0 23296 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_204
timestamp 1698431365
transform 1 0 24192 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_208
timestamp 1698431365
transform 1 0 24640 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_117_212
timestamp 1698431365
transform 1 0 25088 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_220
timestamp 1698431365
transform 1 0 25984 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_224
timestamp 1698431365
transform 1 0 26432 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_234
timestamp 1698431365
transform 1 0 27552 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_238
timestamp 1698431365
transform 1 0 28000 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_240
timestamp 1698431365
transform 1 0 28224 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_2
timestamp 1698431365
transform 1 0 1568 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_12
timestamp 1698431365
transform 1 0 2688 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_25
timestamp 1698431365
transform 1 0 4144 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_31
timestamp 1698431365
transform 1 0 4816 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_37
timestamp 1698431365
transform 1 0 5488 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_49
timestamp 1698431365
transform 1 0 6832 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_84
timestamp 1698431365
transform 1 0 10752 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_94
timestamp 1698431365
transform 1 0 11872 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_96
timestamp 1698431365
transform 1 0 12096 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_107
timestamp 1698431365
transform 1 0 13328 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_161
timestamp 1698431365
transform 1 0 19376 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_165
timestamp 1698431365
transform 1 0 19824 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_173
timestamp 1698431365
transform 1 0 20720 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_185
timestamp 1698431365
transform 1 0 22064 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_187
timestamp 1698431365
transform 1 0 22288 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_118_190
timestamp 1698431365
transform 1 0 22624 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_206
timestamp 1698431365
transform 1 0 24416 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_2
timestamp 1698431365
transform 1 0 1568 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_6
timestamp 1698431365
transform 1 0 2016 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_10
timestamp 1698431365
transform 1 0 2464 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_14
timestamp 1698431365
transform 1 0 2912 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_18
timestamp 1698431365
transform 1 0 3360 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_22
timestamp 1698431365
transform 1 0 3808 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_26
timestamp 1698431365
transform 1 0 4256 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_30
timestamp 1698431365
transform 1 0 4704 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_34
timestamp 1698431365
transform 1 0 5152 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_54
timestamp 1698431365
transform 1 0 7392 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_77
timestamp 1698431365
transform 1 0 9968 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_101
timestamp 1698431365
transform 1 0 12656 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_105
timestamp 1698431365
transform 1 0 13104 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_136
timestamp 1698431365
transform 1 0 16576 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_160
timestamp 1698431365
transform 1 0 19264 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_169
timestamp 1698431365
transform 1 0 20272 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_119_173
timestamp 1698431365
transform 1 0 20720 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_119_189
timestamp 1698431365
transform 1 0 22512 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_197
timestamp 1698431365
transform 1 0 23408 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_201
timestamp 1698431365
transform 1 0 23856 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_209
timestamp 1698431365
transform 1 0 24752 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_212
timestamp 1698431365
transform 1 0 25088 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_218
timestamp 1698431365
transform 1 0 25760 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_119_222
timestamp 1698431365
transform 1 0 26208 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_238
timestamp 1698431365
transform 1 0 28000 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_240
timestamp 1698431365
transform 1 0 28224 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_31
timestamp 1698431365
transform 1 0 4816 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_37
timestamp 1698431365
transform 1 0 5488 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_41
timestamp 1698431365
transform 1 0 5936 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_103
timestamp 1698431365
transform 1 0 12880 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_107
timestamp 1698431365
transform 1 0 13328 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_109
timestamp 1698431365
transform 1 0 13552 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_135
timestamp 1698431365
transform 1 0 16464 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_139
timestamp 1698431365
transform 1 0 16912 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_141
timestamp 1698431365
transform 1 0 17136 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_158
timestamp 1698431365
transform 1 0 19040 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_177
timestamp 1698431365
transform 1 0 21168 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_179
timestamp 1698431365
transform 1 0 21392 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_192
timestamp 1698431365
transform 1 0 22848 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_220
timestamp 1698431365
transform 1 0 25984 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_120_224
timestamp 1698431365
transform 1 0 26432 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_240
timestamp 1698431365
transform 1 0 28224 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_2
timestamp 1698431365
transform 1 0 1568 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_19
timestamp 1698431365
transform 1 0 3472 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_121_21
timestamp 1698431365
transform 1 0 3696 0 -1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_121_53
timestamp 1698431365
transform 1 0 7280 0 -1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_72
timestamp 1698431365
transform 1 0 9408 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_103
timestamp 1698431365
transform 1 0 12880 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_130
timestamp 1698431365
transform 1 0 15904 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_160
timestamp 1698431365
transform 1 0 19264 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_164
timestamp 1698431365
transform 1 0 19712 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_181
timestamp 1698431365
transform 1 0 21616 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_121_183
timestamp 1698431365
transform 1 0 21840 0 -1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_122_2
timestamp 1698431365
transform 1 0 1568 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_10
timestamp 1698431365
transform 1 0 2464 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_12
timestamp 1698431365
transform 1 0 2688 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_15
timestamp 1698431365
transform 1 0 3024 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_19
timestamp 1698431365
transform 1 0 3472 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_23
timestamp 1698431365
transform 1 0 3920 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_27
timestamp 1698431365
transform 1 0 4368 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_31
timestamp 1698431365
transform 1 0 4816 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_45
timestamp 1698431365
transform 1 0 6384 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_107
timestamp 1698431365
transform 1 0 13328 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_150
timestamp 1698431365
transform 1 0 18144 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_154
timestamp 1698431365
transform 1 0 18592 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_170
timestamp 1698431365
transform 1 0 20384 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_174
timestamp 1698431365
transform 1 0 20832 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_177
timestamp 1698431365
transform 1 0 21168 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_181
timestamp 1698431365
transform 1 0 21616 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_185
timestamp 1698431365
transform 1 0 22064 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_230
timestamp 1698431365
transform 1 0 27104 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_234
timestamp 1698431365
transform 1 0 27552 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_238
timestamp 1698431365
transform 1 0 28000 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_240
timestamp 1698431365
transform 1 0 28224 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123_2
timestamp 1698431365
transform 1 0 1568 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_6
timestamp 1698431365
transform 1 0 2016 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_123_8
timestamp 1698431365
transform 1 0 2240 0 -1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_11
timestamp 1698431365
transform 1 0 2576 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_20
timestamp 1698431365
transform 1 0 3584 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_123_22
timestamp 1698431365
transform 1 0 3808 0 -1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_25
timestamp 1698431365
transform 1 0 4144 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_29
timestamp 1698431365
transform 1 0 4592 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_68
timestamp 1698431365
transform 1 0 8960 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_123_87
timestamp 1698431365
transform 1 0 11088 0 -1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_138
timestamp 1698431365
transform 1 0 16800 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_123_142
timestamp 1698431365
transform 1 0 17248 0 -1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_161
timestamp 1698431365
transform 1 0 19376 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_123_165
timestamp 1698431365
transform 1 0 19824 0 -1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_181
timestamp 1698431365
transform 1 0 21616 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_185
timestamp 1698431365
transform 1 0 22064 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_189
timestamp 1698431365
transform 1 0 22512 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123_193
timestamp 1698431365
transform 1 0 22960 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_123_209
timestamp 1698431365
transform 1 0 24752 0 -1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_124_31
timestamp 1698431365
transform 1 0 4816 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_124_37
timestamp 1698431365
transform 1 0 5488 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_124_170
timestamp 1698431365
transform 1 0 20384 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_124_174
timestamp 1698431365
transform 1 0 20832 0 1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_124_177
timestamp 1698431365
transform 1 0 21168 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_124_189
timestamp 1698431365
transform 1 0 22512 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_125_2
timestamp 1698431365
transform 1 0 1568 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_125_6
timestamp 1698431365
transform 1 0 2016 0 -1 100352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125_9
timestamp 1698431365
transform 1 0 2352 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_125_21
timestamp 1698431365
transform 1 0 3696 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125_58
timestamp 1698431365
transform 1 0 7840 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125_208
timestamp 1698431365
transform 1 0 24640 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125_220
timestamp 1698431365
transform 1 0 25984 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125_224
timestamp 1698431365
transform 1 0 26432 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_125_228
timestamp 1698431365
transform 1 0 26880 0 -1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_125_236
timestamp 1698431365
transform 1 0 27776 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_125_240
timestamp 1698431365
transform 1 0 28224 0 -1 100352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_126_2
timestamp 1698431365
transform 1 0 1568 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126_8
timestamp 1698431365
transform 1 0 2240 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126_12
timestamp 1698431365
transform 1 0 2688 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_126_24
timestamp 1698431365
transform 1 0 4032 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126_37
timestamp 1698431365
transform 1 0 5488 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126_75
timestamp 1698431365
transform 1 0 9744 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_126_77
timestamp 1698431365
transform 1 0 9968 0 1 100352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_126_157
timestamp 1698431365
transform 1 0 18928 0 1 100352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126_171
timestamp 1698431365
transform 1 0 20496 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_126_235
timestamp 1698431365
transform 1 0 27664 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126_239
timestamp 1698431365
transform 1 0 28112 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127_31
timestamp 1698431365
transform 1 0 4816 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127_35
timestamp 1698431365
transform 1 0 5264 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127_72
timestamp 1698431365
transform 1 0 9408 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_127_74
timestamp 1698431365
transform 1 0 9632 0 -1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127_142
timestamp 1698431365
transform 1 0 17248 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127_212
timestamp 1698431365
transform 1 0 25088 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_127_216
timestamp 1698431365
transform 1 0 25536 0 -1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_127_232
timestamp 1698431365
transform 1 0 27328 0 -1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_127_240
timestamp 1698431365
transform 1 0 28224 0 -1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_128_2
timestamp 1698431365
transform 1 0 1568 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_128_10
timestamp 1698431365
transform 1 0 2464 0 1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_13
timestamp 1698431365
transform 1 0 2800 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_22
timestamp 1698431365
transform 1 0 3808 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_128_24
timestamp 1698431365
transform 1 0 4032 0 1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_27
timestamp 1698431365
transform 1 0 4368 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_31
timestamp 1698431365
transform 1 0 4816 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_128_37
timestamp 1698431365
transform 1 0 5488 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_43
timestamp 1698431365
transform 1 0 6160 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_47
timestamp 1698431365
transform 1 0 6608 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_51
timestamp 1698431365
transform 1 0 7056 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_128_112
timestamp 1698431365
transform 1 0 13888 0 1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_193
timestamp 1698431365
transform 1 0 22960 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_197
timestamp 1698431365
transform 1 0 23408 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_207
timestamp 1698431365
transform 1 0 24528 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_128_211
timestamp 1698431365
transform 1 0 24976 0 1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_128_227
timestamp 1698431365
transform 1 0 26768 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_128_235
timestamp 1698431365
transform 1 0 27664 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_239
timestamp 1698431365
transform 1 0 28112 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129_2
timestamp 1698431365
transform 1 0 1568 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_8
timestamp 1698431365
transform 1 0 2240 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_12
timestamp 1698431365
transform 1 0 2688 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129_29
timestamp 1698431365
transform 1 0 4592 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_129_33
timestamp 1698431365
transform 1 0 5040 0 -1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_36
timestamp 1698431365
transform 1 0 5376 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_40
timestamp 1698431365
transform 1 0 5824 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_44
timestamp 1698431365
transform 1 0 6272 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_137
timestamp 1698431365
transform 1 0 16688 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_129_139
timestamp 1698431365
transform 1 0 16912 0 -1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_207
timestamp 1698431365
transform 1 0 24528 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_129_209
timestamp 1698431365
transform 1 0 24752 0 -1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_212
timestamp 1698431365
transform 1 0 25088 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_129_216
timestamp 1698431365
transform 1 0 25536 0 -1 103488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_129_232
timestamp 1698431365
transform 1 0 27328 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_129_240
timestamp 1698431365
transform 1 0 28224 0 -1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_130_31
timestamp 1698431365
transform 1 0 4816 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_130_37
timestamp 1698431365
transform 1 0 5488 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130_68
timestamp 1698431365
transform 1 0 8960 0 1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130_107
timestamp 1698431365
transform 1 0 13328 0 1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130_124
timestamp 1698431365
transform 1 0 15232 0 1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_130_200
timestamp 1698431365
transform 1 0 23744 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130_204
timestamp 1698431365
transform 1 0 24192 0 1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_130_218
timestamp 1698431365
transform 1 0 25760 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_130_222
timestamp 1698431365
transform 1 0 26208 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_130_230
timestamp 1698431365
transform 1 0 27104 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130_232
timestamp 1698431365
transform 1 0 27328 0 1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_130_237
timestamp 1698431365
transform 1 0 27888 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_131_2
timestamp 1698431365
transform 1 0 1568 0 -1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_10
timestamp 1698431365
transform 1 0 2464 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_131_12
timestamp 1698431365
transform 1 0 2688 0 -1 105056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_15
timestamp 1698431365
transform 1 0 3024 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_28
timestamp 1698431365
transform 1 0 4480 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_32
timestamp 1698431365
transform 1 0 4928 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_36
timestamp 1698431365
transform 1 0 5376 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_40
timestamp 1698431365
transform 1 0 5824 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_53
timestamp 1698431365
transform 1 0 7280 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_131_72
timestamp 1698431365
transform 1 0 9408 0 -1 105056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_142
timestamp 1698431365
transform 1 0 17248 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_131_146
timestamp 1698431365
transform 1 0 17696 0 -1 105056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_239
timestamp 1698431365
transform 1 0 28112 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_31
timestamp 1698431365
transform 1 0 4816 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_70
timestamp 1698431365
transform 1 0 9184 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_95
timestamp 1698431365
transform 1 0 11984 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_173
timestamp 1698431365
transform 1 0 20720 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_183
timestamp 1698431365
transform 1 0 21840 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_191
timestamp 1698431365
transform 1 0 22736 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_220
timestamp 1698431365
transform 1 0 25984 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_224
timestamp 1698431365
transform 1 0 26432 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_132_228
timestamp 1698431365
transform 1 0 26880 0 1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_132_236
timestamp 1698431365
transform 1 0 27776 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_132_240
timestamp 1698431365
transform 1 0 28224 0 1 105056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_133_2
timestamp 1698431365
transform 1 0 1568 0 -1 106624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133_10
timestamp 1698431365
transform 1 0 2464 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_20
timestamp 1698431365
transform 1 0 3584 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133_24
timestamp 1698431365
transform 1 0 4032 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_28
timestamp 1698431365
transform 1 0 4480 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_32
timestamp 1698431365
transform 1 0 4928 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_36
timestamp 1698431365
transform 1 0 5376 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_133_38
timestamp 1698431365
transform 1 0 5600 0 -1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133_47
timestamp 1698431365
transform 1 0 6608 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_133_51
timestamp 1698431365
transform 1 0 7056 0 -1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_54
timestamp 1698431365
transform 1 0 7392 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_58
timestamp 1698431365
transform 1 0 7840 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_62
timestamp 1698431365
transform 1 0 8288 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_66
timestamp 1698431365
transform 1 0 8736 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_72
timestamp 1698431365
transform 1 0 9408 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_133_142
timestamp 1698431365
transform 1 0 17248 0 -1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_166
timestamp 1698431365
transform 1 0 19936 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_133_170
timestamp 1698431365
transform 1 0 20384 0 -1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_193
timestamp 1698431365
transform 1 0 22960 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_207
timestamp 1698431365
transform 1 0 24528 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_133_209
timestamp 1698431365
transform 1 0 24752 0 -1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_212
timestamp 1698431365
transform 1 0 25088 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_216
timestamp 1698431365
transform 1 0 25536 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_134_2
timestamp 1698431365
transform 1 0 1568 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_134_34
timestamp 1698431365
transform 1 0 5152 0 1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_134_37
timestamp 1698431365
transform 1 0 5488 0 1 106624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_53
timestamp 1698431365
transform 1 0 7280 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_57
timestamp 1698431365
transform 1 0 7728 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_134_59
timestamp 1698431365
transform 1 0 7952 0 1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_62
timestamp 1698431365
transform 1 0 8288 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_66
timestamp 1698431365
transform 1 0 8736 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_70
timestamp 1698431365
transform 1 0 9184 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_74
timestamp 1698431365
transform 1 0 9632 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_101
timestamp 1698431365
transform 1 0 12656 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_147
timestamp 1698431365
transform 1 0 17808 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_173
timestamp 1698431365
transform 1 0 20720 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_134_185
timestamp 1698431365
transform 1 0 22064 0 1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_209
timestamp 1698431365
transform 1 0 24752 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134_213
timestamp 1698431365
transform 1 0 25200 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_134_217
timestamp 1698431365
transform 1 0 25648 0 1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_135_2
timestamp 1698431365
transform 1 0 1568 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135_66
timestamp 1698431365
transform 1 0 8736 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_135_103
timestamp 1698431365
transform 1 0 12880 0 -1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_135_148
timestamp 1698431365
transform 1 0 17920 0 -1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135_178
timestamp 1698431365
transform 1 0 21280 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135_182
timestamp 1698431365
transform 1 0 21728 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_135_184
timestamp 1698431365
transform 1 0 21952 0 -1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135_208
timestamp 1698431365
transform 1 0 24640 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_135_212
timestamp 1698431365
transform 1 0 25088 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135_216
timestamp 1698431365
transform 1 0 25536 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_136_2
timestamp 1698431365
transform 1 0 1568 0 1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_34
timestamp 1698431365
transform 1 0 5152 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_136_37
timestamp 1698431365
transform 1 0 5488 0 1 108192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_136_53
timestamp 1698431365
transform 1 0 7280 0 1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_136_61
timestamp 1698431365
transform 1 0 8176 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_65
timestamp 1698431365
transform 1 0 8624 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_136_124
timestamp 1698431365
transform 1 0 15232 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_126
timestamp 1698431365
transform 1 0 15456 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_136_133
timestamp 1698431365
transform 1 0 16240 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_161
timestamp 1698431365
transform 1 0 19376 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_136_181
timestamp 1698431365
transform 1 0 21616 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_185
timestamp 1698431365
transform 1 0 22064 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_136_232
timestamp 1698431365
transform 1 0 27328 0 1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_240
timestamp 1698431365
transform 1 0 28224 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_137_2
timestamp 1698431365
transform 1 0 1568 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_66
timestamp 1698431365
transform 1 0 8736 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_119
timestamp 1698431365
transform 1 0 14672 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_137_123
timestamp 1698431365
transform 1 0 15120 0 -1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_126
timestamp 1698431365
transform 1 0 15456 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_130
timestamp 1698431365
transform 1 0 15904 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_134
timestamp 1698431365
transform 1 0 16352 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_138
timestamp 1698431365
transform 1 0 16800 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_142
timestamp 1698431365
transform 1 0 17248 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_146
timestamp 1698431365
transform 1 0 17696 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_137_148
timestamp 1698431365
transform 1 0 17920 0 -1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_151
timestamp 1698431365
transform 1 0 18256 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_155
timestamp 1698431365
transform 1 0 18704 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_159
timestamp 1698431365
transform 1 0 19152 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_163
timestamp 1698431365
transform 1 0 19600 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_137_167
timestamp 1698431365
transform 1 0 20048 0 -1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_186
timestamp 1698431365
transform 1 0 22176 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_137_190
timestamp 1698431365
transform 1 0 22624 0 -1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_206
timestamp 1698431365
transform 1 0 24416 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_212
timestamp 1698431365
transform 1 0 25088 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_216
timestamp 1698431365
transform 1 0 25536 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138_2
timestamp 1698431365
transform 1 0 1568 0 1 109760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_138_34
timestamp 1698431365
transform 1 0 5152 0 1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_138_37
timestamp 1698431365
transform 1 0 5488 0 1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_138_53
timestamp 1698431365
transform 1 0 7280 0 1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_61
timestamp 1698431365
transform 1 0 8176 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_138_65
timestamp 1698431365
transform 1 0 8624 0 1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138_134
timestamp 1698431365
transform 1 0 16352 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_138_138
timestamp 1698431365
transform 1 0 16800 0 1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_154
timestamp 1698431365
transform 1 0 18592 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138_158
timestamp 1698431365
transform 1 0 19040 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_138_160
timestamp 1698431365
transform 1 0 19264 0 1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138_163
timestamp 1698431365
transform 1 0 19600 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_167
timestamp 1698431365
transform 1 0 20048 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_138_171
timestamp 1698431365
transform 1 0 20496 0 1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_138_174
timestamp 1698431365
transform 1 0 20832 0 1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138_200
timestamp 1698431365
transform 1 0 23744 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_138_204
timestamp 1698431365
transform 1 0 24192 0 1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_212
timestamp 1698431365
transform 1 0 25088 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138_216
timestamp 1698431365
transform 1 0 25536 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_139_2
timestamp 1698431365
transform 1 0 1568 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_139_66
timestamp 1698431365
transform 1 0 8736 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_103
timestamp 1698431365
transform 1 0 12880 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_107
timestamp 1698431365
transform 1 0 13328 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_134
timestamp 1698431365
transform 1 0 16352 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_138
timestamp 1698431365
transform 1 0 16800 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_188
timestamp 1698431365
transform 1 0 22400 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_139_192
timestamp 1698431365
transform 1 0 22848 0 -1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_208
timestamp 1698431365
transform 1 0 24640 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_139_212
timestamp 1698431365
transform 1 0 25088 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_216
timestamp 1698431365
transform 1 0 25536 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_140_2
timestamp 1698431365
transform 1 0 1568 0 1 111328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_140_34
timestamp 1698431365
transform 1 0 5152 0 1 111328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_140_37
timestamp 1698431365
transform 1 0 5488 0 1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_140_45
timestamp 1698431365
transform 1 0 6384 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_140_95
timestamp 1698431365
transform 1 0 11984 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_140_99
timestamp 1698431365
transform 1 0 12432 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_140_103
timestamp 1698431365
transform 1 0 12880 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_140_107
timestamp 1698431365
transform 1 0 13328 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_140_134
timestamp 1698431365
transform 1 0 16352 0 1 111328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_140_158
timestamp 1698431365
transform 1 0 19040 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_140_162
timestamp 1698431365
transform 1 0 19488 0 1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_140_170
timestamp 1698431365
transform 1 0 20384 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_140_174
timestamp 1698431365
transform 1 0 20832 0 1 111328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_140_177
timestamp 1698431365
transform 1 0 21168 0 1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_140_239
timestamp 1698431365
transform 1 0 28112 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_141_2
timestamp 1698431365
transform 1 0 1568 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_141_66
timestamp 1698431365
transform 1 0 8736 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_141_72
timestamp 1698431365
transform 1 0 9408 0 -1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_141_134
timestamp 1698431365
transform 1 0 16352 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_141_138
timestamp 1698431365
transform 1 0 16800 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_141_142
timestamp 1698431365
transform 1 0 17248 0 -1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_141_181
timestamp 1698431365
transform 1 0 21616 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_141_185
timestamp 1698431365
transform 1 0 22064 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_141_212
timestamp 1698431365
transform 1 0 25088 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_141_216
timestamp 1698431365
transform 1 0 25536 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142_2
timestamp 1698431365
transform 1 0 1568 0 1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142_34
timestamp 1698431365
transform 1 0 5152 0 1 112896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_142_37
timestamp 1698431365
transform 1 0 5488 0 1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142_53
timestamp 1698431365
transform 1 0 7280 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142_103
timestamp 1698431365
transform 1 0 12880 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142_107
timestamp 1698431365
transform 1 0 13328 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_142_113
timestamp 1698431365
transform 1 0 14000 0 1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142_129
timestamp 1698431365
transform 1 0 15792 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142_133
timestamp 1698431365
transform 1 0 16240 0 1 112896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_142_136
timestamp 1698431365
transform 1 0 16576 0 1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142_177
timestamp 1698431365
transform 1 0 21168 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142_181
timestamp 1698431365
transform 1 0 21616 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_142_206
timestamp 1698431365
transform 1 0 24416 0 1 112896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142_214
timestamp 1698431365
transform 1 0 25312 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_143_2
timestamp 1698431365
transform 1 0 1568 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_66
timestamp 1698431365
transform 1 0 8736 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_72
timestamp 1698431365
transform 1 0 9408 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_143_99
timestamp 1698431365
transform 1 0 12432 0 -1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_143_107
timestamp 1698431365
transform 1 0 13328 0 -1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_143_131
timestamp 1698431365
transform 1 0 16016 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_135
timestamp 1698431365
transform 1 0 16464 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_143_139
timestamp 1698431365
transform 1 0 16912 0 -1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_143_188
timestamp 1698431365
transform 1 0 22400 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_143_192
timestamp 1698431365
transform 1 0 22848 0 -1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_143_208
timestamp 1698431365
transform 1 0 24640 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_143_212
timestamp 1698431365
transform 1 0 25088 0 -1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_143_228
timestamp 1698431365
transform 1 0 26880 0 -1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_236
timestamp 1698431365
transform 1 0 27776 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_143_240
timestamp 1698431365
transform 1 0 28224 0 -1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_144_2
timestamp 1698431365
transform 1 0 1568 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144_34
timestamp 1698431365
transform 1 0 5152 0 1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_144_37
timestamp 1698431365
transform 1 0 5488 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144_101
timestamp 1698431365
transform 1 0 12656 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_144_107
timestamp 1698431365
transform 1 0 13328 0 1 114464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144_123
timestamp 1698431365
transform 1 0 15120 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144_127
timestamp 1698431365
transform 1 0 15568 0 1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_144_151
timestamp 1698431365
transform 1 0 18256 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_144_155
timestamp 1698431365
transform 1 0 18704 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_144_163
timestamp 1698431365
transform 1 0 19600 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_144_167
timestamp 1698431365
transform 1 0 20048 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144_177
timestamp 1698431365
transform 1 0 21168 0 1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_144_201
timestamp 1698431365
transform 1 0 23856 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_144_205
timestamp 1698431365
transform 1 0 24304 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144_237
timestamp 1698431365
transform 1 0 27888 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_145_6
timestamp 1698431365
transform 1 0 2016 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_72
timestamp 1698431365
transform 1 0 9408 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_145_99
timestamp 1698431365
transform 1 0 12432 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_103
timestamp 1698431365
transform 1 0 12880 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_145_130
timestamp 1698431365
transform 1 0 15904 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_134
timestamp 1698431365
transform 1 0 16352 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_145_138
timestamp 1698431365
transform 1 0 16800 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_145_188
timestamp 1698431365
transform 1 0 22400 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_145_192
timestamp 1698431365
transform 1 0 22848 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_145_208
timestamp 1698431365
transform 1 0 24640 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_145_212
timestamp 1698431365
transform 1 0 25088 0 -1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_145_228
timestamp 1698431365
transform 1 0 26880 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_236
timestamp 1698431365
transform 1 0 27776 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_145_240
timestamp 1698431365
transform 1 0 28224 0 -1 116032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_146_2
timestamp 1698431365
transform 1 0 1568 0 1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_146_34
timestamp 1698431365
transform 1 0 5152 0 1 116032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_146_37
timestamp 1698431365
transform 1 0 5488 0 1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_146_69
timestamp 1698431365
transform 1 0 9072 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_146_77
timestamp 1698431365
transform 1 0 9968 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_146_81
timestamp 1698431365
transform 1 0 10416 0 1 116032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_146_107
timestamp 1698431365
transform 1 0 13328 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_146_134
timestamp 1698431365
transform 1 0 16352 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_146_160
timestamp 1698431365
transform 1 0 19264 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_146_164
timestamp 1698431365
transform 1 0 19712 0 1 116032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_146_167
timestamp 1698431365
transform 1 0 20048 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_146_171
timestamp 1698431365
transform 1 0 20496 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_146_177
timestamp 1698431365
transform 1 0 21168 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_147_2
timestamp 1698431365
transform 1 0 1568 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_147_66
timestamp 1698431365
transform 1 0 8736 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_147_72
timestamp 1698431365
transform 1 0 9408 0 -1 117600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_147_104
timestamp 1698431365
transform 1 0 12992 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_147_108
timestamp 1698431365
transform 1 0 13440 0 -1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147_132
timestamp 1698431365
transform 1 0 16128 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147_136
timestamp 1698431365
transform 1 0 16576 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147_188
timestamp 1698431365
transform 1 0 22400 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_147_192
timestamp 1698431365
transform 1 0 22848 0 -1 117600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_147_212
timestamp 1698431365
transform 1 0 25088 0 -1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_147_219
timestamp 1698431365
transform 1 0 25872 0 -1 117600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_147_235
timestamp 1698431365
transform 1 0 27664 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147_239
timestamp 1698431365
transform 1 0 28112 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_148_6
timestamp 1698431365
transform 1 0 2016 0 1 117600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_148_14
timestamp 1698431365
transform 1 0 2912 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_16
timestamp 1698431365
transform 1 0 3136 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_148_21
timestamp 1698431365
transform 1 0 3696 0 1 117600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_29
timestamp 1698431365
transform 1 0 4592 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_33
timestamp 1698431365
transform 1 0 5040 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_148_40
timestamp 1698431365
transform 1 0 5824 0 1 117600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_48
timestamp 1698431365
transform 1 0 6720 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_148_53
timestamp 1698431365
transform 1 0 7280 0 1 117600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_61
timestamp 1698431365
transform 1 0 8176 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_148_65
timestamp 1698431365
transform 1 0 8624 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_67
timestamp 1698431365
transform 1 0 8848 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_74
timestamp 1698431365
transform 1 0 9632 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_148_78
timestamp 1698431365
transform 1 0 10080 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_80
timestamp 1698431365
transform 1 0 10304 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_148_85
timestamp 1698431365
transform 1 0 10864 0 1 117600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_93
timestamp 1698431365
transform 1 0 11760 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_101
timestamp 1698431365
transform 1 0 12656 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_104
timestamp 1698431365
transform 1 0 12992 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_148_132
timestamp 1698431365
transform 1 0 16128 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_148_138
timestamp 1698431365
transform 1 0 16800 0 1 117600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_146
timestamp 1698431365
transform 1 0 17696 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_148_172
timestamp 1698431365
transform 1 0 20608 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_148_176
timestamp 1698431365
transform 1 0 21056 0 1 117600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_148_192
timestamp 1698431365
transform 1 0 22848 0 1 117600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_200
timestamp 1698431365
transform 1 0 23744 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_148_206
timestamp 1698431365
transform 1 0 24416 0 1 117600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_240
timestamp 1698431365
transform 1 0 28224 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 27216 0 -1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 19152 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 19824 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 17472 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 16800 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 15568 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 14896 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 14896 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 14224 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 12096 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 11424 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 27888 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 11424 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 10080 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 9408 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 9520 0 -1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 8288 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 7616 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 6944 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 6272 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 6272 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input23
timestamp 1698431365
transform -1 0 26208 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 3808 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 3136 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input26
timestamp 1698431365
transform -1 0 25312 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input27
timestamp 1698431365
transform -1 0 23520 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input28
timestamp 1698431365
transform -1 0 22624 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform -1 0 23856 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 21840 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 24192 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 19040 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input33
timestamp 1698431365
transform -1 0 27664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input34
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input45
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 1568 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform 1 0 1568 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform 1 0 1568 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform 1 0 1568 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform 1 0 1568 0 -1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input54
timestamp 1698431365
transform 1 0 1568 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform 1 0 1568 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input56
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input57
timestamp 1698431365
transform 1 0 1568 0 -1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input58
timestamp 1698431365
transform 1 0 1568 0 1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input59
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input66
timestamp 1698431365
transform -1 0 27216 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1698431365
transform -1 0 27888 0 -1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input68
timestamp 1698431365
transform 1 0 2464 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_149 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 28560 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_150
timestamp 1698431365
transform 1 0 1344 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 28560 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_151
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 28560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_152
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_153
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_154
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 28560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_155
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_156
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 28560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_157
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_158
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_159
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_160
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 28560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_161
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_162
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 28560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_163
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_164
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_165
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_166
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_167
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_168
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_169
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_170
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_171
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_172
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_173
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_174
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_175
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_176
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 28560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_177
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_178
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 28560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_179
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_180
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_181
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_182
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 28560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_183
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_184
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 28560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_185
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_186
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 28560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_187
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_188
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 28560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_189
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_190
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 28560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_191
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_192
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 28560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_193
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_194
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 28560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_195
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_196
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 28560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_197
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 28560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_198
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 28560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_199
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_200
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 28560 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_201
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_202
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 28560 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_203
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_204
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 28560 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_205
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 28560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_206
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 28560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_207
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 28560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_208
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 28560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_209
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 28560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_210
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 28560 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_211
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 28560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_212
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 28560 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_213
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 28560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_214
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 28560 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_215
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_216
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 28560 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_217
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 28560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_218
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 28560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_219
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 28560 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_220
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 28560 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_221
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 28560 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_222
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 28560 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_223
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 28560 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_224
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 28560 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_225
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 28560 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_226
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 28560 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_227
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 28560 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_228
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 28560 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_229
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 28560 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_230
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 28560 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_231
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 28560 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_232
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 28560 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_233
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 28560 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_234
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 28560 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_235
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 28560 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_236
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 28560 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_237
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 28560 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_238
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 28560 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_239
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 28560 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_240
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 28560 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_241
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 28560 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_242
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 28560 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Left_243
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Right_94
timestamp 1698431365
transform -1 0 28560 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Left_244
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Right_95
timestamp 1698431365
transform -1 0 28560 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Left_245
timestamp 1698431365
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Right_96
timestamp 1698431365
transform -1 0 28560 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Left_246
timestamp 1698431365
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Right_97
timestamp 1698431365
transform -1 0 28560 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Left_247
timestamp 1698431365
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Right_98
timestamp 1698431365
transform -1 0 28560 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Left_248
timestamp 1698431365
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Right_99
timestamp 1698431365
transform -1 0 28560 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Left_249
timestamp 1698431365
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Right_100
timestamp 1698431365
transform -1 0 28560 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Left_250
timestamp 1698431365
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Right_101
timestamp 1698431365
transform -1 0 28560 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Left_251
timestamp 1698431365
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Right_102
timestamp 1698431365
transform -1 0 28560 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Left_252
timestamp 1698431365
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Right_103
timestamp 1698431365
transform -1 0 28560 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Left_253
timestamp 1698431365
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Right_104
timestamp 1698431365
transform -1 0 28560 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Left_254
timestamp 1698431365
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Right_105
timestamp 1698431365
transform -1 0 28560 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Left_255
timestamp 1698431365
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Right_106
timestamp 1698431365
transform -1 0 28560 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Left_256
timestamp 1698431365
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Right_107
timestamp 1698431365
transform -1 0 28560 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Left_257
timestamp 1698431365
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Right_108
timestamp 1698431365
transform -1 0 28560 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Left_258
timestamp 1698431365
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Right_109
timestamp 1698431365
transform -1 0 28560 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Left_259
timestamp 1698431365
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Right_110
timestamp 1698431365
transform -1 0 28560 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Left_260
timestamp 1698431365
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Right_111
timestamp 1698431365
transform -1 0 28560 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Left_261
timestamp 1698431365
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Right_112
timestamp 1698431365
transform -1 0 28560 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Left_262
timestamp 1698431365
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Right_113
timestamp 1698431365
transform -1 0 28560 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Left_263
timestamp 1698431365
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Right_114
timestamp 1698431365
transform -1 0 28560 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Left_264
timestamp 1698431365
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Right_115
timestamp 1698431365
transform -1 0 28560 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Left_265
timestamp 1698431365
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Right_116
timestamp 1698431365
transform -1 0 28560 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Left_266
timestamp 1698431365
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Right_117
timestamp 1698431365
transform -1 0 28560 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Left_267
timestamp 1698431365
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Right_118
timestamp 1698431365
transform -1 0 28560 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_Left_268
timestamp 1698431365
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_Right_119
timestamp 1698431365
transform -1 0 28560 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_Left_269
timestamp 1698431365
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_Right_120
timestamp 1698431365
transform -1 0 28560 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_Left_270
timestamp 1698431365
transform 1 0 1344 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_Right_121
timestamp 1698431365
transform -1 0 28560 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_Left_271
timestamp 1698431365
transform 1 0 1344 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_Right_122
timestamp 1698431365
transform -1 0 28560 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_123_Left_272
timestamp 1698431365
transform 1 0 1344 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_123_Right_123
timestamp 1698431365
transform -1 0 28560 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_124_Left_273
timestamp 1698431365
transform 1 0 1344 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_124_Right_124
timestamp 1698431365
transform -1 0 28560 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_125_Left_274
timestamp 1698431365
transform 1 0 1344 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_125_Right_125
timestamp 1698431365
transform -1 0 28560 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_126_Left_275
timestamp 1698431365
transform 1 0 1344 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_126_Right_126
timestamp 1698431365
transform -1 0 28560 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_127_Left_276
timestamp 1698431365
transform 1 0 1344 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_127_Right_127
timestamp 1698431365
transform -1 0 28560 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_128_Left_277
timestamp 1698431365
transform 1 0 1344 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_128_Right_128
timestamp 1698431365
transform -1 0 28560 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_129_Left_278
timestamp 1698431365
transform 1 0 1344 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_129_Right_129
timestamp 1698431365
transform -1 0 28560 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_130_Left_279
timestamp 1698431365
transform 1 0 1344 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_130_Right_130
timestamp 1698431365
transform -1 0 28560 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_131_Left_280
timestamp 1698431365
transform 1 0 1344 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_131_Right_131
timestamp 1698431365
transform -1 0 28560 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_132_Left_281
timestamp 1698431365
transform 1 0 1344 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_132_Right_132
timestamp 1698431365
transform -1 0 28560 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_133_Left_282
timestamp 1698431365
transform 1 0 1344 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_133_Right_133
timestamp 1698431365
transform -1 0 28560 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_134_Left_283
timestamp 1698431365
transform 1 0 1344 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_134_Right_134
timestamp 1698431365
transform -1 0 28560 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_135_Left_284
timestamp 1698431365
transform 1 0 1344 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_135_Right_135
timestamp 1698431365
transform -1 0 28560 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_136_Left_285
timestamp 1698431365
transform 1 0 1344 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_136_Right_136
timestamp 1698431365
transform -1 0 28560 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_137_Left_286
timestamp 1698431365
transform 1 0 1344 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_137_Right_137
timestamp 1698431365
transform -1 0 28560 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_138_Left_287
timestamp 1698431365
transform 1 0 1344 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_138_Right_138
timestamp 1698431365
transform -1 0 28560 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_139_Left_288
timestamp 1698431365
transform 1 0 1344 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_139_Right_139
timestamp 1698431365
transform -1 0 28560 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_140_Left_289
timestamp 1698431365
transform 1 0 1344 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_140_Right_140
timestamp 1698431365
transform -1 0 28560 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_141_Left_290
timestamp 1698431365
transform 1 0 1344 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_141_Right_141
timestamp 1698431365
transform -1 0 28560 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_142_Left_291
timestamp 1698431365
transform 1 0 1344 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_142_Right_142
timestamp 1698431365
transform -1 0 28560 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_143_Left_292
timestamp 1698431365
transform 1 0 1344 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_143_Right_143
timestamp 1698431365
transform -1 0 28560 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_144_Left_293
timestamp 1698431365
transform 1 0 1344 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_144_Right_144
timestamp 1698431365
transform -1 0 28560 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_145_Left_294
timestamp 1698431365
transform 1 0 1344 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_145_Right_145
timestamp 1698431365
transform -1 0 28560 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_146_Left_295
timestamp 1698431365
transform 1 0 1344 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_146_Right_146
timestamp 1698431365
transform -1 0 28560 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_147_Left_296
timestamp 1698431365
transform 1 0 1344 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_147_Right_147
timestamp 1698431365
transform -1 0 28560 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_148_Left_297
timestamp 1698431365
transform 1 0 1344 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_148_Right_148
timestamp 1698431365
transform -1 0 28560 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  seg1._26_
timestamp 1698431365
transform 1 0 27440 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  seg1._27_
timestamp 1698431365
transform -1 0 25872 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  seg1._28_
timestamp 1698431365
transform 1 0 25984 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  seg1._29_
timestamp 1698431365
transform 1 0 24976 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  seg1._30_
timestamp 1698431365
transform 1 0 25312 0 1 92512
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  seg1._31_
timestamp 1698431365
transform 1 0 26768 0 1 90944
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._32_
timestamp 1698431365
transform -1 0 25984 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._33_
timestamp 1698431365
transform 1 0 27216 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  seg1._34_
timestamp 1698431365
transform -1 0 27216 0 -1 92512
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  seg1._35_
timestamp 1698431365
transform 1 0 22176 0 -1 89376
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  seg1._36_
timestamp 1698431365
transform -1 0 23520 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._37_
timestamp 1698431365
transform -1 0 23072 0 1 89376
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  seg1._38_
timestamp 1698431365
transform -1 0 27328 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  seg1._39_
timestamp 1698431365
transform -1 0 24752 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._40_
timestamp 1698431365
transform -1 0 24528 0 1 90944
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  seg1._41_
timestamp 1698431365
transform -1 0 23968 0 1 90944
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._42_
timestamp 1698431365
transform -1 0 23072 0 -1 90944
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._43_
timestamp 1698431365
transform -1 0 22176 0 -1 90944
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._44_
timestamp 1698431365
transform 1 0 21616 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  seg1._45_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23184 0 1 90944
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  seg1._46_
timestamp 1698431365
transform 1 0 22736 0 -1 92512
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  seg1._47_
timestamp 1698431365
transform -1 0 23072 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  seg1._48_
timestamp 1698431365
transform -1 0 22848 0 -1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._49_
timestamp 1698431365
transform -1 0 22736 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._50_
timestamp 1698431365
transform 1 0 23184 0 1 92512
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  seg1._51_
timestamp 1698431365
transform 1 0 23744 0 -1 92512
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._52_
timestamp 1698431365
transform -1 0 24304 0 1 92512
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._53_
timestamp 1698431365
transform -1 0 23744 0 -1 90944
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  seg1._54_
timestamp 1698431365
transform -1 0 23408 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._55_
timestamp 1698431365
transform 1 0 21280 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._56_
timestamp 1698431365
transform 1 0 25088 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  seg1._57_
timestamp 1698431365
transform -1 0 26768 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._58_
timestamp 1698431365
transform 1 0 23856 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_298 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_299
timestamp 1698431365
transform 1 0 8960 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_300
timestamp 1698431365
transform 1 0 12768 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_301
timestamp 1698431365
transform 1 0 16576 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_302
timestamp 1698431365
transform 1 0 20384 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_303
timestamp 1698431365
transform 1 0 24192 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_304
timestamp 1698431365
transform 1 0 28000 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_305
timestamp 1698431365
transform 1 0 9184 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_306
timestamp 1698431365
transform 1 0 17024 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_307
timestamp 1698431365
transform 1 0 24864 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_308
timestamp 1698431365
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_309
timestamp 1698431365
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_310
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_311
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_312
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_313
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_314
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_315
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_316
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_317
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_318
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_319
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_320
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_321
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_322
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_323
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_324
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_325
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_326
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_327
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_328
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_329
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_330
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_331
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_332
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_333
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_334
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_335
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_336
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_337
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_338
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_339
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_340
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_341
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_342
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_343
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_344
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_345
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_346
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_347
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_348
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_349
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_350
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_351
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_352
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_353
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_354
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_355
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_356
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_357
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_358
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_359
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_360
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_361
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_362
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_363
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_364
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_365
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_366
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_367
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_368
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_369
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_370
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_371
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_372
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_373
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_374
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_375
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_376
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_377
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_378
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_379
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_380
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_381
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_382
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_383
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_384
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_385
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_386
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_387
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_388
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_389
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_390
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_391
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_392
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_393
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_394
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_395
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_396
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_397
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_398
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_399
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_400
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_401
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_402
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_403
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_404
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_405
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_406
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_407
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_408
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_409
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_410
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_411
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_412
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_413
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_414
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_415
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_416
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_417
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_418
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_422
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_425
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_426
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_427
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_428
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_429
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_430
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_431
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_432
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_433
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_434
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_435
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_436
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_437
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_438
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_439
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_440
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_441
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_442
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_443
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_444
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_445
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_446
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_447
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_448
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_449
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_450
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_451
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_452
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_453
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_454
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_455
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_456
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_457
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_458
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_459
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_460
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_461
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_462
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_463
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_464
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_465
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_466
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_467
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_468
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_469
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_470
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_471
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_472
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_473
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_474
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_475
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_476
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_477
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_478
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_479
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_480
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_481
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_482
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_483
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_484
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_485
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_486
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_487
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_488
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_489
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_490
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_491
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_492
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_493
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_494
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_495
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_496
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_497
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_498
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_499
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_500
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_501
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_502
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_503
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_504
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_505
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_506
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_507
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_508
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_509
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_510
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_511
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_512
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_513
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_514
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_515
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_516
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_517
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_518
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_519
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_520
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_521
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_522
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_523
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_524
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_525
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_526
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_527
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_528
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_529
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_530
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_531
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_532
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_533
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_534
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_535
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_536
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_537
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_538
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_539
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_540
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_541
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_542
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_543
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_544
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_545
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_546
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_547
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_548
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_549
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_550
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_551
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_552
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_553
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_554
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_555
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_556
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_557
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_558
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_559
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_560
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_561
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_562
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_563
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_564
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_565
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_566
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_567
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_568
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_569
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_570
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_571
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_572
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_573
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_574
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_575
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_576
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_577
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_578
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_579
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_580
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_581
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_582
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_583
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_584
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_585
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_586
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_587
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_588
timestamp 1698431365
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_589
timestamp 1698431365
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_590
timestamp 1698431365
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_591
timestamp 1698431365
transform 1 0 13104 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_592
timestamp 1698431365
transform 1 0 20944 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_593
timestamp 1698431365
transform 1 0 9184 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_594
timestamp 1698431365
transform 1 0 17024 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_595
timestamp 1698431365
transform 1 0 24864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_596
timestamp 1698431365
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_597
timestamp 1698431365
transform 1 0 13104 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_598
timestamp 1698431365
transform 1 0 20944 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_599
timestamp 1698431365
transform 1 0 9184 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_600
timestamp 1698431365
transform 1 0 17024 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_601
timestamp 1698431365
transform 1 0 24864 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_602
timestamp 1698431365
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_603
timestamp 1698431365
transform 1 0 13104 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_604
timestamp 1698431365
transform 1 0 20944 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_605
timestamp 1698431365
transform 1 0 9184 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_606
timestamp 1698431365
transform 1 0 17024 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_607
timestamp 1698431365
transform 1 0 24864 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_608
timestamp 1698431365
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_609
timestamp 1698431365
transform 1 0 13104 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_610
timestamp 1698431365
transform 1 0 20944 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_611
timestamp 1698431365
transform 1 0 9184 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_612
timestamp 1698431365
transform 1 0 17024 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_613
timestamp 1698431365
transform 1 0 24864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_614
timestamp 1698431365
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_615
timestamp 1698431365
transform 1 0 13104 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_616
timestamp 1698431365
transform 1 0 20944 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_617
timestamp 1698431365
transform 1 0 9184 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_618
timestamp 1698431365
transform 1 0 17024 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_619
timestamp 1698431365
transform 1 0 24864 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_620
timestamp 1698431365
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_621
timestamp 1698431365
transform 1 0 13104 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_622
timestamp 1698431365
transform 1 0 20944 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_623
timestamp 1698431365
transform 1 0 9184 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_624
timestamp 1698431365
transform 1 0 17024 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_625
timestamp 1698431365
transform 1 0 24864 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_626
timestamp 1698431365
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_627
timestamp 1698431365
transform 1 0 13104 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_628
timestamp 1698431365
transform 1 0 20944 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_629
timestamp 1698431365
transform 1 0 9184 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_630
timestamp 1698431365
transform 1 0 17024 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_631
timestamp 1698431365
transform 1 0 24864 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_632
timestamp 1698431365
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_633
timestamp 1698431365
transform 1 0 13104 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_634
timestamp 1698431365
transform 1 0 20944 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_635
timestamp 1698431365
transform 1 0 9184 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_636
timestamp 1698431365
transform 1 0 17024 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_637
timestamp 1698431365
transform 1 0 24864 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_638
timestamp 1698431365
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_639
timestamp 1698431365
transform 1 0 13104 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_640
timestamp 1698431365
transform 1 0 20944 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_641
timestamp 1698431365
transform 1 0 9184 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_642
timestamp 1698431365
transform 1 0 17024 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_643
timestamp 1698431365
transform 1 0 24864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_644
timestamp 1698431365
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_645
timestamp 1698431365
transform 1 0 13104 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_646
timestamp 1698431365
transform 1 0 20944 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_647
timestamp 1698431365
transform 1 0 9184 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_648
timestamp 1698431365
transform 1 0 17024 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_649
timestamp 1698431365
transform 1 0 24864 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_650
timestamp 1698431365
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_651
timestamp 1698431365
transform 1 0 13104 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_652
timestamp 1698431365
transform 1 0 20944 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_653
timestamp 1698431365
transform 1 0 9184 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_654
timestamp 1698431365
transform 1 0 17024 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_655
timestamp 1698431365
transform 1 0 24864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_656
timestamp 1698431365
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_657
timestamp 1698431365
transform 1 0 13104 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_658
timestamp 1698431365
transform 1 0 20944 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_659
timestamp 1698431365
transform 1 0 9184 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_660
timestamp 1698431365
transform 1 0 17024 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_661
timestamp 1698431365
transform 1 0 24864 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_662
timestamp 1698431365
transform 1 0 5264 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_663
timestamp 1698431365
transform 1 0 13104 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_664
timestamp 1698431365
transform 1 0 20944 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_665
timestamp 1698431365
transform 1 0 9184 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_666
timestamp 1698431365
transform 1 0 17024 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_667
timestamp 1698431365
transform 1 0 24864 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_668
timestamp 1698431365
transform 1 0 5264 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_669
timestamp 1698431365
transform 1 0 13104 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_670
timestamp 1698431365
transform 1 0 20944 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_671
timestamp 1698431365
transform 1 0 9184 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_672
timestamp 1698431365
transform 1 0 17024 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_673
timestamp 1698431365
transform 1 0 24864 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_674
timestamp 1698431365
transform 1 0 5264 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_675
timestamp 1698431365
transform 1 0 13104 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_676
timestamp 1698431365
transform 1 0 20944 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_677
timestamp 1698431365
transform 1 0 9184 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_678
timestamp 1698431365
transform 1 0 17024 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_679
timestamp 1698431365
transform 1 0 24864 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_680
timestamp 1698431365
transform 1 0 5264 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_681
timestamp 1698431365
transform 1 0 13104 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_682
timestamp 1698431365
transform 1 0 20944 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_683
timestamp 1698431365
transform 1 0 9184 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_684
timestamp 1698431365
transform 1 0 17024 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_685
timestamp 1698431365
transform 1 0 24864 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_686
timestamp 1698431365
transform 1 0 5264 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_687
timestamp 1698431365
transform 1 0 13104 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_688
timestamp 1698431365
transform 1 0 20944 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_689
timestamp 1698431365
transform 1 0 9184 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_690
timestamp 1698431365
transform 1 0 17024 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_691
timestamp 1698431365
transform 1 0 24864 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_692
timestamp 1698431365
transform 1 0 5264 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_693
timestamp 1698431365
transform 1 0 13104 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_694
timestamp 1698431365
transform 1 0 20944 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_695
timestamp 1698431365
transform 1 0 9184 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_696
timestamp 1698431365
transform 1 0 17024 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_697
timestamp 1698431365
transform 1 0 24864 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_698
timestamp 1698431365
transform 1 0 5264 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_699
timestamp 1698431365
transform 1 0 13104 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_700
timestamp 1698431365
transform 1 0 20944 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_701
timestamp 1698431365
transform 1 0 9184 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_702
timestamp 1698431365
transform 1 0 17024 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_703
timestamp 1698431365
transform 1 0 24864 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_704
timestamp 1698431365
transform 1 0 5264 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_705
timestamp 1698431365
transform 1 0 13104 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_706
timestamp 1698431365
transform 1 0 20944 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_707
timestamp 1698431365
transform 1 0 9184 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_708
timestamp 1698431365
transform 1 0 17024 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_709
timestamp 1698431365
transform 1 0 24864 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_710
timestamp 1698431365
transform 1 0 5264 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_711
timestamp 1698431365
transform 1 0 13104 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_712
timestamp 1698431365
transform 1 0 20944 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_713
timestamp 1698431365
transform 1 0 9184 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_714
timestamp 1698431365
transform 1 0 17024 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_715
timestamp 1698431365
transform 1 0 24864 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_716
timestamp 1698431365
transform 1 0 5264 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_717
timestamp 1698431365
transform 1 0 13104 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_718
timestamp 1698431365
transform 1 0 20944 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_719
timestamp 1698431365
transform 1 0 9184 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_720
timestamp 1698431365
transform 1 0 17024 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_721
timestamp 1698431365
transform 1 0 24864 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_722
timestamp 1698431365
transform 1 0 5264 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_723
timestamp 1698431365
transform 1 0 13104 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_724
timestamp 1698431365
transform 1 0 20944 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_725
timestamp 1698431365
transform 1 0 9184 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_726
timestamp 1698431365
transform 1 0 17024 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_727
timestamp 1698431365
transform 1 0 24864 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_728
timestamp 1698431365
transform 1 0 5264 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_729
timestamp 1698431365
transform 1 0 13104 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_730
timestamp 1698431365
transform 1 0 20944 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_731
timestamp 1698431365
transform 1 0 9184 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_732
timestamp 1698431365
transform 1 0 17024 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_733
timestamp 1698431365
transform 1 0 24864 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_144_734
timestamp 1698431365
transform 1 0 5264 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_144_735
timestamp 1698431365
transform 1 0 13104 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_144_736
timestamp 1698431365
transform 1 0 20944 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_145_737
timestamp 1698431365
transform 1 0 9184 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_145_738
timestamp 1698431365
transform 1 0 17024 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_145_739
timestamp 1698431365
transform 1 0 24864 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_146_740
timestamp 1698431365
transform 1 0 5264 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_146_741
timestamp 1698431365
transform 1 0 13104 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_146_742
timestamp 1698431365
transform 1 0 20944 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_147_743
timestamp 1698431365
transform 1 0 9184 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_147_744
timestamp 1698431365
transform 1 0 17024 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_147_745
timestamp 1698431365
transform 1 0 24864 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_746
timestamp 1698431365
transform 1 0 5152 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_747
timestamp 1698431365
transform 1 0 8960 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_748
timestamp 1698431365
transform 1 0 12768 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_749
timestamp 1698431365
transform 1 0 16576 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_750
timestamp 1698431365
transform 1 0 20384 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_751
timestamp 1698431365
transform 1 0 24192 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_752
timestamp 1698431365
transform 1 0 28000 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac._4_
timestamp 1698431365
transform -1 0 23184 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac._5_
timestamp 1698431365
transform 1 0 22064 0 1 105056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[0\].vdac_batch._3_
timestamp 1698431365
transform 1 0 18144 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[0\].vdac_batch._4_
timestamp 1698431365
transform 1 0 17808 0 -1 105056
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[0\].vdac_batch._5_
timestamp 1698431365
transform -1 0 20720 0 1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.parallel_cells\[0\].vdac_batch._6_
timestamp 1698431365
transform -1 0 17920 0 -1 108192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[0\].vdac_batch._7_
timestamp 1698431365
transform 1 0 20496 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.parallel_cells\[0\].vdac_batch._8_
timestamp 1698431365
transform 1 0 21168 0 1 105056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17360 0 -1 106624
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 21168 0 1 103488
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[1\].vdac_batch._3_
timestamp 1698431365
transform 1 0 13328 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[1\].vdac_batch._4_
timestamp 1698431365
transform 1 0 13776 0 1 106624
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[1\].vdac_batch._5_
timestamp 1698431365
transform -1 0 18928 0 1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.parallel_cells\[1\].vdac_batch._6_
timestamp 1698431365
transform -1 0 16240 0 1 108192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[1\].vdac_batch._7_
timestamp 1698431365
transform -1 0 19376 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.parallel_cells\[1\].vdac_batch._8_
timestamp 1698431365
transform 1 0 16464 0 1 108192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 15232 0 1 106624
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 18032 0 -1 108192
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform -1 0 17024 0 -1 108192
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_4  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 1 106624
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[2\].vdac_batch._3_
timestamp 1698431365
transform 1 0 9632 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[2\].vdac_batch._4_
timestamp 1698431365
transform -1 0 14448 0 -1 108192
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[2\].vdac_batch._5_
timestamp 1698431365
transform -1 0 13104 0 1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  temp1.dac.parallel_cells\[2\].vdac_batch._6_
timestamp 1698431365
transform -1 0 12656 0 -1 109760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[2\].vdac_batch._7_
timestamp 1698431365
transform -1 0 15232 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  temp1.dac.parallel_cells\[2\].vdac_batch._8_
timestamp 1698431365
transform 1 0 11984 0 1 108192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform -1 0 11984 0 1 108192
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 13776 0 1 109760
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform -1 0 12656 0 1 106624
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform 1 0 13776 0 1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform -1 0 11984 0 -1 108192
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform 1 0 13776 0 -1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform -1 0 11984 0 1 105056
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform 1 0 13776 0 -1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  temp1.dac.parallel_cells\[3\].vdac_batch._3_
timestamp 1698431365
transform -1 0 9408 0 1 108192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[3\].vdac_batch._4_
timestamp 1698431365
transform 1 0 13328 0 1 108192
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[3\].vdac_batch._5_
timestamp 1698431365
transform 1 0 11312 0 1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  temp1.dac.parallel_cells\[3\].vdac_batch._6_
timestamp 1698431365
transform 1 0 11984 0 -1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[3\].vdac_batch._7_
timestamp 1698431365
transform 1 0 13328 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  temp1.dac.parallel_cells\[3\].vdac_batch._8_
timestamp 1698431365
transform 1 0 12656 0 -1 109760
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 9408 0 -1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 13776 0 1 116032
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform -1 0 12432 0 -1 114464
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform 1 0 13328 0 -1 116032
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform -1 0 9408 0 1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform 1 0 13440 0 -1 114464
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform 1 0 9408 0 1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform 1 0 13552 0 1 117600
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1698431365
transform 1 0 8736 0 1 109760
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1698431365
transform 1 0 13552 0 -1 117600
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1698431365
transform 1 0 10304 0 1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1698431365
transform 1 0 10528 0 1 116032
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1698431365
transform -1 0 11984 0 -1 109760
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref
timestamp 1698431365
transform 1 0 11200 0 -1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1698431365
transform 1 0 7728 0 1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1698431365
transform -1 0 12432 0 -1 116032
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  temp1.dac.parallel_cells\[4\].vdac_batch._3_
timestamp 1698431365
transform 1 0 22064 0 -1 106624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[4\].vdac_batch._4_
timestamp 1698431365
transform 1 0 19488 0 1 108192
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[4\].vdac_batch._5_
timestamp 1698431365
transform 1 0 21168 0 1 106624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  temp1.dac.parallel_cells\[4\].vdac_batch._6_
timestamp 1698431365
transform -1 0 22064 0 -1 106624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[4\].vdac_batch._7_
timestamp 1698431365
transform -1 0 21616 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  temp1.dac.parallel_cells\[4\].vdac_batch._8_
timestamp 1698431365
transform -1 0 22176 0 -1 109760
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 25760 0 1 109760
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 19824 0 -1 116032
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform 1 0 22064 0 -1 108192
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform 1 0 19824 0 -1 114464
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform 1 0 25760 0 1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform 1 0 17248 0 -1 114464
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform 1 0 25760 0 -1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform 1 0 21168 0 1 109760
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1698431365
transform 1 0 25760 0 -1 109760
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1698431365
transform 1 0 21280 0 1 114464
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1698431365
transform 1 0 25760 0 1 106624
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1698431365
transform 1 0 17248 0 -1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1698431365
transform 1 0 25760 0 -1 106624
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref
timestamp 1698431365
transform -1 0 20384 0 1 117600
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1698431365
transform 1 0 25760 0 -1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_4  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1698431365
transform 1 0 16576 0 1 116032
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1698431365
transform 1 0 22176 0 1 106624
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1698431365
transform 1 0 17248 0 -1 116032
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1698431365
transform 1 0 22288 0 -1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1698431365
transform 1 0 19040 0 -1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1698431365
transform -1 0 24416 0 1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1698431365
transform 1 0 16464 0 1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1698431365
transform 1 0 22176 0 1 108192
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1698431365
transform 1 0 18368 0 1 112896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1698431365
transform 1 0 25760 0 -1 108192
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1698431365
transform 1 0 17248 0 -1 117600
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1698431365
transform 1 0 25536 0 1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1698431365
transform 1 0 19824 0 -1 117600
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1698431365
transform 1 0 24752 0 1 108192
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1698431365
transform -1 0 18256 0 1 114464
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1698431365
transform 1 0 22960 0 1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1698431365
transform 1 0 19824 0 -1 111328
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.dac.vdac_single._3_
timestamp 1698431365
transform -1 0 27888 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._3__78 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._4__79
timestamp 1698431365
transform -1 0 25536 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._4__80
timestamp 1698431365
transform -1 0 25984 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.vdac_single._4_
timestamp 1698431365
transform -1 0 25760 0 1 103488
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.vdac_single._5_
timestamp 1698431365
transform 1 0 23632 0 -1 106624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.vdac_single._6_
timestamp 1698431365
transform 1 0 24864 0 1 105056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.vdac_single._7_
timestamp 1698431365
transform 1 0 23184 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.vdac_single._8_
timestamp 1698431365
transform -1 0 24528 0 1 101920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 25536 0 -1 105056
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  temp1.dac.vdac_single.einvp_batch\[0\].vref open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 1 105056
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  temp1.dcdc
timestamp 1698431365
transform 1 0 9520 0 -1 105056
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv1_1
timestamp 1698431365
transform 1 0 8736 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv2_2
timestamp 1698431365
transform -1 0 9520 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv2_3
timestamp 1698431365
transform -1 0 16128 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_69
timestamp 1698431365
transform 1 0 13104 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_70
timestamp 1698431365
transform -1 0 12656 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_71
timestamp 1698431365
transform -1 0 10864 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_72
timestamp 1698431365
transform -1 0 9632 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_73
timestamp 1698431365
transform -1 0 7280 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_74
timestamp 1698431365
transform -1 0 5824 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_75
timestamp 1698431365
transform -1 0 3696 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_76
timestamp 1698431365
transform -1 0 2016 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_77
timestamp 1698431365
transform -1 0 2016 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  wire4
timestamp 1698431365
transform 1 0 6720 0 -1 15680
box -86 -86 982 870
<< labels >>
flabel metal2 s 3360 0 3472 400 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 24864 0 24976 400 0 FreeSans 448 90 0 0 i_wb_addr[0]
port 1 nsew signal input
flabel metal2 s 18144 0 18256 400 0 FreeSans 448 90 0 0 i_wb_addr[10]
port 2 nsew signal input
flabel metal2 s 17472 0 17584 400 0 FreeSans 448 90 0 0 i_wb_addr[11]
port 3 nsew signal input
flabel metal2 s 16800 0 16912 400 0 FreeSans 448 90 0 0 i_wb_addr[12]
port 4 nsew signal input
flabel metal2 s 16128 0 16240 400 0 FreeSans 448 90 0 0 i_wb_addr[13]
port 5 nsew signal input
flabel metal2 s 15456 0 15568 400 0 FreeSans 448 90 0 0 i_wb_addr[14]
port 6 nsew signal input
flabel metal2 s 14784 0 14896 400 0 FreeSans 448 90 0 0 i_wb_addr[15]
port 7 nsew signal input
flabel metal2 s 14112 0 14224 400 0 FreeSans 448 90 0 0 i_wb_addr[16]
port 8 nsew signal input
flabel metal2 s 13440 0 13552 400 0 FreeSans 448 90 0 0 i_wb_addr[17]
port 9 nsew signal input
flabel metal2 s 12768 0 12880 400 0 FreeSans 448 90 0 0 i_wb_addr[18]
port 10 nsew signal input
flabel metal2 s 12096 0 12208 400 0 FreeSans 448 90 0 0 i_wb_addr[19]
port 11 nsew signal input
flabel metal2 s 24192 0 24304 400 0 FreeSans 448 90 0 0 i_wb_addr[1]
port 12 nsew signal input
flabel metal2 s 11424 0 11536 400 0 FreeSans 448 90 0 0 i_wb_addr[20]
port 13 nsew signal input
flabel metal2 s 10752 0 10864 400 0 FreeSans 448 90 0 0 i_wb_addr[21]
port 14 nsew signal input
flabel metal2 s 10080 0 10192 400 0 FreeSans 448 90 0 0 i_wb_addr[22]
port 15 nsew signal input
flabel metal2 s 9408 0 9520 400 0 FreeSans 448 90 0 0 i_wb_addr[23]
port 16 nsew signal input
flabel metal2 s 8736 0 8848 400 0 FreeSans 448 90 0 0 i_wb_addr[24]
port 17 nsew signal input
flabel metal2 s 8064 0 8176 400 0 FreeSans 448 90 0 0 i_wb_addr[25]
port 18 nsew signal input
flabel metal2 s 7392 0 7504 400 0 FreeSans 448 90 0 0 i_wb_addr[26]
port 19 nsew signal input
flabel metal2 s 6720 0 6832 400 0 FreeSans 448 90 0 0 i_wb_addr[27]
port 20 nsew signal input
flabel metal2 s 6048 0 6160 400 0 FreeSans 448 90 0 0 i_wb_addr[28]
port 21 nsew signal input
flabel metal2 s 5376 0 5488 400 0 FreeSans 448 90 0 0 i_wb_addr[29]
port 22 nsew signal input
flabel metal2 s 23520 0 23632 400 0 FreeSans 448 90 0 0 i_wb_addr[2]
port 23 nsew signal input
flabel metal2 s 4704 0 4816 400 0 FreeSans 448 90 0 0 i_wb_addr[30]
port 24 nsew signal input
flabel metal2 s 4032 0 4144 400 0 FreeSans 448 90 0 0 i_wb_addr[31]
port 25 nsew signal input
flabel metal2 s 22848 0 22960 400 0 FreeSans 448 90 0 0 i_wb_addr[3]
port 26 nsew signal input
flabel metal2 s 22176 0 22288 400 0 FreeSans 448 90 0 0 i_wb_addr[4]
port 27 nsew signal input
flabel metal2 s 21504 0 21616 400 0 FreeSans 448 90 0 0 i_wb_addr[5]
port 28 nsew signal input
flabel metal2 s 20832 0 20944 400 0 FreeSans 448 90 0 0 i_wb_addr[6]
port 29 nsew signal input
flabel metal2 s 20160 0 20272 400 0 FreeSans 448 90 0 0 i_wb_addr[7]
port 30 nsew signal input
flabel metal2 s 19488 0 19600 400 0 FreeSans 448 90 0 0 i_wb_addr[8]
port 31 nsew signal input
flabel metal2 s 18816 0 18928 400 0 FreeSans 448 90 0 0 i_wb_addr[9]
port 32 nsew signal input
flabel metal2 s 26880 0 26992 400 0 FreeSans 448 90 0 0 i_wb_cyc
port 33 nsew signal input
flabel metal3 s 0 4704 400 4816 0 FreeSans 448 0 0 0 i_wb_data[0]
port 34 nsew signal input
flabel metal3 s 0 31584 400 31696 0 FreeSans 448 0 0 0 i_wb_data[10]
port 35 nsew signal input
flabel metal3 s 0 34272 400 34384 0 FreeSans 448 0 0 0 i_wb_data[11]
port 36 nsew signal input
flabel metal3 s 0 36960 400 37072 0 FreeSans 448 0 0 0 i_wb_data[12]
port 37 nsew signal input
flabel metal3 s 0 39648 400 39760 0 FreeSans 448 0 0 0 i_wb_data[13]
port 38 nsew signal input
flabel metal3 s 0 42336 400 42448 0 FreeSans 448 0 0 0 i_wb_data[14]
port 39 nsew signal input
flabel metal3 s 0 45024 400 45136 0 FreeSans 448 0 0 0 i_wb_data[15]
port 40 nsew signal input
flabel metal3 s 0 47712 400 47824 0 FreeSans 448 0 0 0 i_wb_data[16]
port 41 nsew signal input
flabel metal3 s 0 50400 400 50512 0 FreeSans 448 0 0 0 i_wb_data[17]
port 42 nsew signal input
flabel metal3 s 0 53088 400 53200 0 FreeSans 448 0 0 0 i_wb_data[18]
port 43 nsew signal input
flabel metal3 s 0 55776 400 55888 0 FreeSans 448 0 0 0 i_wb_data[19]
port 44 nsew signal input
flabel metal3 s 0 7392 400 7504 0 FreeSans 448 0 0 0 i_wb_data[1]
port 45 nsew signal input
flabel metal3 s 0 58464 400 58576 0 FreeSans 448 0 0 0 i_wb_data[20]
port 46 nsew signal input
flabel metal3 s 0 61152 400 61264 0 FreeSans 448 0 0 0 i_wb_data[21]
port 47 nsew signal input
flabel metal3 s 0 63840 400 63952 0 FreeSans 448 0 0 0 i_wb_data[22]
port 48 nsew signal input
flabel metal3 s 0 66528 400 66640 0 FreeSans 448 0 0 0 i_wb_data[23]
port 49 nsew signal input
flabel metal3 s 0 69216 400 69328 0 FreeSans 448 0 0 0 i_wb_data[24]
port 50 nsew signal input
flabel metal3 s 0 71904 400 72016 0 FreeSans 448 0 0 0 i_wb_data[25]
port 51 nsew signal input
flabel metal3 s 0 74592 400 74704 0 FreeSans 448 0 0 0 i_wb_data[26]
port 52 nsew signal input
flabel metal3 s 0 77280 400 77392 0 FreeSans 448 0 0 0 i_wb_data[27]
port 53 nsew signal input
flabel metal3 s 0 79968 400 80080 0 FreeSans 448 0 0 0 i_wb_data[28]
port 54 nsew signal input
flabel metal3 s 0 82656 400 82768 0 FreeSans 448 0 0 0 i_wb_data[29]
port 55 nsew signal input
flabel metal3 s 0 10080 400 10192 0 FreeSans 448 0 0 0 i_wb_data[2]
port 56 nsew signal input
flabel metal3 s 0 85344 400 85456 0 FreeSans 448 0 0 0 i_wb_data[30]
port 57 nsew signal input
flabel metal3 s 0 88032 400 88144 0 FreeSans 448 0 0 0 i_wb_data[31]
port 58 nsew signal input
flabel metal3 s 0 12768 400 12880 0 FreeSans 448 0 0 0 i_wb_data[3]
port 59 nsew signal input
flabel metal3 s 0 15456 400 15568 0 FreeSans 448 0 0 0 i_wb_data[4]
port 60 nsew signal input
flabel metal3 s 0 18144 400 18256 0 FreeSans 448 0 0 0 i_wb_data[5]
port 61 nsew signal input
flabel metal3 s 0 20832 400 20944 0 FreeSans 448 0 0 0 i_wb_data[6]
port 62 nsew signal input
flabel metal3 s 0 23520 400 23632 0 FreeSans 448 0 0 0 i_wb_data[7]
port 63 nsew signal input
flabel metal3 s 0 26208 400 26320 0 FreeSans 448 0 0 0 i_wb_data[8]
port 64 nsew signal input
flabel metal3 s 0 28896 400 29008 0 FreeSans 448 0 0 0 i_wb_data[9]
port 65 nsew signal input
flabel metal2 s 26208 0 26320 400 0 FreeSans 448 90 0 0 i_wb_stb
port 66 nsew signal input
flabel metal2 s 25536 0 25648 400 0 FreeSans 448 90 0 0 i_wb_we
port 67 nsew signal input
flabel metal2 s 13888 119600 14000 120000 0 FreeSans 448 90 0 0 io_oeb[0]
port 68 nsew signal tristate
flabel metal2 s 12096 119600 12208 120000 0 FreeSans 448 90 0 0 io_oeb[1]
port 69 nsew signal tristate
flabel metal2 s 10304 119600 10416 120000 0 FreeSans 448 90 0 0 io_oeb[2]
port 70 nsew signal tristate
flabel metal2 s 8512 119600 8624 120000 0 FreeSans 448 90 0 0 io_oeb[3]
port 71 nsew signal tristate
flabel metal2 s 6720 119600 6832 120000 0 FreeSans 448 90 0 0 io_oeb[4]
port 72 nsew signal tristate
flabel metal2 s 4928 119600 5040 120000 0 FreeSans 448 90 0 0 io_oeb[5]
port 73 nsew signal tristate
flabel metal2 s 3136 119600 3248 120000 0 FreeSans 448 90 0 0 io_oeb[6]
port 74 nsew signal tristate
flabel metal2 s 1344 119600 1456 120000 0 FreeSans 448 90 0 0 io_oeb[7]
port 75 nsew signal tristate
flabel metal2 s 28224 119600 28336 120000 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 26432 119600 26544 120000 0 FreeSans 448 90 0 0 io_out[1]
port 77 nsew signal tristate
flabel metal2 s 24640 119600 24752 120000 0 FreeSans 448 90 0 0 io_out[2]
port 78 nsew signal tristate
flabel metal2 s 22848 119600 22960 120000 0 FreeSans 448 90 0 0 io_out[3]
port 79 nsew signal tristate
flabel metal2 s 21056 119600 21168 120000 0 FreeSans 448 90 0 0 io_out[4]
port 80 nsew signal tristate
flabel metal2 s 19264 119600 19376 120000 0 FreeSans 448 90 0 0 io_out[5]
port 81 nsew signal tristate
flabel metal2 s 17472 119600 17584 120000 0 FreeSans 448 90 0 0 io_out[6]
port 82 nsew signal tristate
flabel metal2 s 15680 119600 15792 120000 0 FreeSans 448 90 0 0 io_out[7]
port 83 nsew signal tristate
flabel metal3 s 0 90720 400 90832 0 FreeSans 448 0 0 0 o_wb_ack
port 84 nsew signal tristate
flabel metal3 s 0 93408 400 93520 0 FreeSans 448 0 0 0 o_wb_data[0]
port 85 nsew signal tristate
flabel metal3 s 0 96096 400 96208 0 FreeSans 448 0 0 0 o_wb_data[1]
port 86 nsew signal tristate
flabel metal3 s 0 98784 400 98896 0 FreeSans 448 0 0 0 o_wb_data[2]
port 87 nsew signal tristate
flabel metal3 s 0 101472 400 101584 0 FreeSans 448 0 0 0 o_wb_data[3]
port 88 nsew signal tristate
flabel metal3 s 0 104160 400 104272 0 FreeSans 448 0 0 0 o_wb_data[4]
port 89 nsew signal tristate
flabel metal3 s 0 106848 400 106960 0 FreeSans 448 0 0 0 o_wb_data[5]
port 90 nsew signal tristate
flabel metal3 s 0 109536 400 109648 0 FreeSans 448 0 0 0 o_wb_data[6]
port 91 nsew signal tristate
flabel metal3 s 0 112224 400 112336 0 FreeSans 448 0 0 0 o_wb_data[7]
port 92 nsew signal tristate
flabel metal3 s 0 114912 400 115024 0 FreeSans 448 0 0 0 o_wb_stall
port 93 nsew signal tristate
flabel metal2 s 2688 0 2800 400 0 FreeSans 448 90 0 0 reset
port 94 nsew signal input
flabel metal4 s 4586 1508 4906 118444 0 FreeSans 1280 90 0 0 vdd
port 95 nsew power bidirectional
flabel metal4 s 11390 1508 11710 118444 0 FreeSans 1280 90 0 0 vdd
port 95 nsew power bidirectional
flabel metal4 s 18194 1508 18514 118444 0 FreeSans 1280 90 0 0 vdd
port 95 nsew power bidirectional
flabel metal4 s 24998 1508 25318 118444 0 FreeSans 1280 90 0 0 vdd
port 95 nsew power bidirectional
flabel metal4 s 7988 1508 8308 118444 0 FreeSans 1280 90 0 0 vss
port 96 nsew ground bidirectional
flabel metal4 s 14792 1508 15112 118444 0 FreeSans 1280 90 0 0 vss
port 96 nsew ground bidirectional
flabel metal4 s 21596 1508 21916 118444 0 FreeSans 1280 90 0 0 vss
port 96 nsew ground bidirectional
flabel metal4 s 28400 1508 28720 118444 0 FreeSans 1280 90 0 0 vss
port 96 nsew ground bidirectional
rlabel metal1 14952 118384 14952 118384 0 vdd
rlabel via1 15032 117600 15032 117600 0 vss
rlabel metal2 18984 17304 18984 17304 0 _0000_
rlabel metal2 10472 15400 10472 15400 0 _0001_
rlabel metal2 21336 17304 21336 17304 0 _0002_
rlabel metal2 15848 16352 15848 16352 0 _0003_
rlabel metal2 11928 76888 11928 76888 0 _0004_
rlabel metal3 10024 75768 10024 75768 0 _0005_
rlabel metal2 23576 73584 23576 73584 0 _0006_
rlabel metal3 10360 71960 10360 71960 0 _0007_
rlabel metal2 22792 59640 22792 59640 0 _0008_
rlabel metal2 8456 56504 8456 56504 0 _0009_
rlabel metal2 8232 52472 8232 52472 0 _0010_
rlabel metal2 7448 47824 7448 47824 0 _0011_
rlabel metal2 8568 50204 8568 50204 0 _0012_
rlabel metal2 15848 43120 15848 43120 0 _0013_
rlabel metal2 12152 43848 12152 43848 0 _0014_
rlabel metal2 11256 45920 11256 45920 0 _0015_
rlabel metal2 18536 40712 18536 40712 0 _0016_
rlabel metal2 13608 41496 13608 41496 0 _0017_
rlabel metal2 18088 35280 18088 35280 0 _0018_
rlabel metal2 14728 38976 14728 38976 0 _0019_
rlabel metal2 23016 36120 23016 36120 0 _0020_
rlabel metal3 20384 44072 20384 44072 0 _0021_
rlabel metal2 26040 58072 26040 58072 0 _0022_
rlabel metal2 26040 59640 26040 59640 0 _0023_
rlabel metal2 26152 48328 26152 48328 0 _0024_
rlabel metal2 21448 55664 21448 55664 0 _0025_
rlabel metal2 26488 44352 26488 44352 0 _0026_
rlabel metal2 22680 57064 22680 57064 0 _0027_
rlabel metal2 25480 55496 25480 55496 0 _0028_
rlabel metal2 26040 53256 26040 53256 0 _0029_
rlabel metal2 25704 50232 25704 50232 0 _0030_
rlabel metal2 23912 53256 23912 53256 0 _0031_
rlabel metal2 8568 14168 8568 14168 0 _0032_
rlabel metal2 5992 18760 5992 18760 0 _0033_
rlabel metal2 6552 17304 6552 17304 0 _0034_
rlabel metal2 10024 11760 10024 11760 0 _0035_
rlabel metal2 5208 12320 5208 12320 0 _0036_
rlabel metal2 5320 13888 5320 13888 0 _0037_
rlabel metal2 25368 18872 25368 18872 0 _0038_
rlabel metal2 21000 13944 21000 13944 0 _0039_
rlabel metal2 23408 15288 23408 15288 0 _0040_
rlabel metal2 18200 14168 18200 14168 0 _0041_
rlabel metal2 13832 13048 13832 13048 0 _0042_
rlabel metal2 10640 13944 10640 13944 0 _0043_
rlabel metal2 7896 62776 7896 62776 0 _0044_
rlabel metal2 6328 64344 6328 64344 0 _0045_
rlabel metal2 6104 68208 6104 68208 0 _0046_
rlabel metal2 5992 66416 5992 66416 0 _0047_
rlabel metal2 11312 63224 11312 63224 0 _0048_
rlabel metal2 5376 49896 5376 49896 0 _0049_
rlabel metal2 10360 27440 10360 27440 0 _0050_
rlabel metal3 13944 36512 13944 36512 0 _0051_
rlabel metal2 7336 37688 7336 37688 0 _0052_
rlabel metal2 6888 46256 6888 46256 0 _0053_
rlabel metal2 23128 32144 23128 32144 0 _0054_
rlabel metal2 24024 39256 24024 39256 0 _0055_
rlabel metal2 23912 42392 23912 42392 0 _0056_
rlabel metal2 16296 30800 16296 30800 0 _0057_
rlabel metal2 25704 25144 25704 25144 0 _0058_
rlabel metal2 27384 29008 27384 29008 0 _0059_
rlabel metal2 24640 28728 24640 28728 0 _0060_
rlabel metal2 24136 36848 24136 36848 0 _0061_
rlabel metal2 24248 47096 24248 47096 0 _0062_
rlabel metal2 22232 45528 22232 45528 0 _0063_
rlabel metal2 5264 100072 5264 100072 0 _0064_
rlabel metal2 6328 101136 6328 101136 0 _0065_
rlabel metal2 3752 86184 3752 86184 0 _0066_
rlabel metal3 6608 97720 6608 97720 0 _0067_
rlabel metal2 6216 93296 6216 93296 0 _0068_
rlabel metal2 2520 91504 2520 91504 0 _0069_
rlabel metal2 8008 90216 8008 90216 0 _0070_
rlabel metal2 9744 94584 9744 94584 0 _0071_
rlabel metal2 19880 101080 19880 101080 0 _0072_
rlabel metal2 23464 100408 23464 100408 0 _0073_
rlabel metal2 25368 100408 25368 100408 0 _0074_
rlabel metal2 27384 98224 27384 98224 0 _0075_
rlabel metal2 27328 96936 27328 96936 0 _0076_
rlabel metal2 25760 94584 25760 94584 0 _0077_
rlabel metal2 19768 21896 19768 21896 0 _0078_
rlabel metal2 13048 20216 13048 20216 0 _0079_
rlabel metal2 23352 22120 23352 22120 0 _0080_
rlabel metal2 16744 25872 16744 25872 0 _0081_
rlabel metal2 19152 18424 19152 18424 0 _0082_
rlabel metal2 16520 20440 16520 20440 0 _0083_
rlabel metal3 23408 25368 23408 25368 0 _0084_
rlabel metal2 13608 29008 13608 29008 0 _0085_
rlabel metal2 6888 23576 6888 23576 0 _0086_
rlabel metal2 10304 20552 10304 20552 0 _0087_
rlabel metal2 5880 21224 5880 21224 0 _0088_
rlabel metal2 9800 19936 9800 19936 0 _0089_
rlabel metal2 7896 26208 7896 26208 0 _0090_
rlabel metal2 14280 26712 14280 26712 0 _0091_
rlabel metal2 11424 31080 11424 31080 0 _0092_
rlabel metal2 10808 40040 10808 40040 0 _0093_
rlabel metal2 8456 40824 8456 40824 0 _0094_
rlabel metal2 7224 42896 7224 42896 0 _0095_
rlabel metal2 17696 28504 17696 28504 0 _0096_
rlabel metal3 14504 35560 14504 35560 0 _0097_
rlabel metal2 23464 42392 23464 42392 0 _0098_
rlabel metal2 15680 41272 15680 41272 0 _0099_
rlabel metal2 26712 31416 26712 31416 0 _0100_
rlabel metal3 27216 39368 27216 39368 0 _0101_
rlabel metal2 27048 41384 27048 41384 0 _0102_
rlabel metal2 13720 31808 13720 31808 0 _0103_
rlabel metal2 26712 23408 26712 23408 0 _0104_
rlabel metal2 25984 20104 25984 20104 0 _0105_
rlabel metal2 26712 27608 26712 27608 0 _0106_
rlabel metal2 27328 35784 27328 35784 0 _0107_
rlabel metal2 26712 33880 26712 33880 0 _0108_
rlabel metal2 21336 38668 21336 38668 0 _0109_
rlabel metal2 6888 7784 6888 7784 0 _0110_
rlabel metal2 2520 10528 2520 10528 0 _0111_
rlabel metal2 2968 7896 2968 7896 0 _0112_
rlabel metal2 6664 9464 6664 9464 0 _0113_
rlabel metal2 2576 13048 2576 13048 0 _0114_
rlabel metal2 2464 16744 2464 16744 0 _0115_
rlabel metal2 2464 19320 2464 19320 0 _0116_
rlabel metal2 2520 22008 2520 22008 0 _0117_
rlabel metal2 2520 24472 2520 24472 0 _0118_
rlabel metal2 5208 24864 5208 24864 0 _0119_
rlabel metal2 2520 30408 2520 30408 0 _0120_
rlabel metal2 2520 33544 2520 33544 0 _0121_
rlabel metal3 5264 35784 5264 35784 0 _0122_
rlabel metal2 2520 42392 2520 42392 0 _0123_
rlabel metal2 2520 28168 2520 28168 0 _0124_
rlabel metal2 2632 39704 2632 39704 0 _0125_
rlabel metal2 5880 33712 5880 33712 0 _0126_
rlabel metal2 5152 40264 5152 40264 0 _0127_
rlabel metal2 2520 37576 2520 37576 0 _0128_
rlabel metal2 2576 45752 2576 45752 0 _0129_
rlabel metal2 2520 57960 2520 57960 0 _0130_
rlabel metal2 2520 60536 2520 60536 0 _0131_
rlabel metal2 2464 63224 2464 63224 0 _0132_
rlabel metal2 2520 65912 2520 65912 0 _0133_
rlabel metal2 2576 69272 2576 69272 0 _0134_
rlabel metal2 2520 72184 2520 72184 0 _0135_
rlabel metal2 2520 75320 2520 75320 0 _0136_
rlabel metal2 2520 78456 2520 78456 0 _0137_
rlabel metal2 5320 79016 5320 79016 0 _0138_
rlabel metal2 2464 82040 2464 82040 0 _0139_
rlabel metal2 7224 81592 7224 81592 0 _0140_
rlabel metal3 5264 82824 5264 82824 0 _0141_
rlabel metal2 20328 27216 20328 27216 0 _0142_
rlabel metal3 11424 56952 11424 56952 0 _0143_
rlabel metal3 19264 9912 19264 9912 0 _0144_
rlabel metal2 16856 6888 16856 6888 0 _0145_
rlabel metal2 15512 9856 15512 9856 0 _0146_
rlabel metal2 14280 10416 14280 10416 0 _0147_
rlabel metal2 12824 17976 12824 17976 0 _0148_
rlabel metal2 14392 14896 14392 14896 0 _0149_
rlabel metal2 23464 11704 23464 11704 0 _0150_
rlabel metal2 17080 11760 17080 11760 0 _0151_
rlabel metal3 13776 8344 13776 8344 0 _0152_
rlabel metal2 10472 9968 10472 9968 0 _0153_
rlabel metal2 10360 24136 10360 24136 0 _0154_
rlabel metal2 14280 23296 14280 23296 0 _0155_
rlabel metal2 10472 68208 10472 68208 0 _0156_
rlabel metal2 10360 65072 10360 65072 0 _0157_
rlabel metal2 17864 67480 17864 67480 0 _0158_
rlabel metal2 13608 65968 13608 65968 0 _0159_
rlabel metal3 10024 60984 10024 60984 0 _0160_
rlabel metal2 10696 54152 10696 54152 0 _0161_
rlabel metal2 18648 69608 18648 69608 0 _0162_
rlabel metal2 14280 75320 14280 75320 0 _0163_
rlabel metal2 26096 73416 26096 73416 0 _0164_
rlabel metal2 26096 70392 26096 70392 0 _0165_
rlabel metal2 26040 65072 26040 65072 0 _0166_
rlabel metal2 15176 63280 15176 63280 0 _0167_
rlabel metal2 26264 76888 26264 76888 0 _0168_
rlabel metal2 24472 77560 24472 77560 0 _0169_
rlabel metal2 27384 68768 27384 68768 0 _0170_
rlabel metal2 26600 68264 26600 68264 0 _0171_
rlabel metal2 26600 63336 26600 63336 0 _0172_
rlabel metal3 22288 62216 22288 62216 0 _0173_
rlabel metal2 2520 88480 2520 88480 0 _0174_
rlabel metal2 15680 82040 15680 82040 0 _0175_
rlabel metal2 19656 76048 19656 76048 0 _0176_
rlabel metal2 9128 78456 9128 78456 0 _0177_
rlabel metal2 22456 77448 22456 77448 0 _0178_
rlabel metal2 15624 78456 15624 78456 0 _0179_
rlabel metal2 18200 75208 18200 75208 0 _0180_
rlabel metal2 14448 78568 14448 78568 0 _0181_
rlabel metal2 22232 71680 22232 71680 0 _0182_
rlabel metal2 21952 73528 21952 73528 0 _0183_
rlabel metal2 20832 66920 20832 66920 0 _0184_
rlabel metal2 20776 64512 20776 64512 0 _0185_
rlabel metal2 11256 58800 11256 58800 0 _0186_
rlabel metal2 2968 54880 2968 54880 0 _0187_
rlabel metal2 6888 29680 6888 29680 0 _0188_
rlabel metal3 4648 29512 4648 29512 0 _0189_
rlabel metal2 7056 31640 7056 31640 0 _0190_
rlabel metal2 4872 42000 4872 42000 0 _0191_
rlabel metal2 6440 59640 6440 59640 0 _0192_
rlabel metal2 5320 56224 5320 56224 0 _0193_
rlabel metal3 2856 50456 2856 50456 0 _0194_
rlabel metal2 3080 47824 3080 47824 0 _0195_
rlabel metal2 6440 53368 6440 53368 0 _0196_
rlabel metal2 19544 54824 19544 54824 0 _0197_
rlabel metal2 5096 60984 5096 60984 0 _0198_
rlabel metal2 19264 62888 19264 62888 0 _0199_
rlabel metal2 5152 71736 5152 71736 0 _0200_
rlabel metal2 5824 73192 5824 73192 0 _0201_
rlabel metal2 6440 75320 6440 75320 0 _0202_
rlabel metal2 6440 76888 6440 76888 0 _0203_
rlabel metal2 19992 61208 19992 61208 0 _0204_
rlabel metal3 19656 59304 19656 59304 0 _0205_
rlabel metal3 23016 49672 23016 49672 0 _0206_
rlabel metal2 20832 51464 20832 51464 0 _0207_
rlabel metal2 3864 93296 3864 93296 0 _0208_
rlabel metal2 3864 96432 3864 96432 0 _0209_
rlabel metal2 3864 99400 3864 99400 0 _0210_
rlabel metal2 3808 100856 3808 100856 0 _0211_
rlabel metal2 3808 103208 3808 103208 0 _0212_
rlabel metal2 7112 103544 7112 103544 0 _0213_
rlabel metal2 3304 105896 3304 105896 0 _0214_
rlabel metal3 7056 105560 7056 105560 0 _0215_
rlabel metal2 14448 85176 14448 85176 0 _0216_
rlabel metal2 11816 84672 11816 84672 0 _0217_
rlabel metal2 11256 82992 11256 82992 0 _0218_
rlabel metal2 8232 85708 8232 85708 0 _0219_
rlabel metal2 10752 88312 10752 88312 0 _0220_
rlabel metal2 6888 87976 6888 87976 0 _0221_
rlabel metal2 8680 91000 8680 91000 0 _0222_
rlabel metal2 10136 82264 10136 82264 0 _0223_
rlabel metal2 9240 93464 9240 93464 0 _0224_
rlabel metal2 6664 98616 6664 98616 0 _0225_
rlabel metal2 21896 22960 21896 22960 0 _0226_
rlabel metal2 24696 73640 24696 73640 0 _0227_
rlabel metal2 21560 14560 21560 14560 0 _0228_
rlabel metal3 11312 71848 11312 71848 0 _0229_
rlabel metal3 21728 15176 21728 15176 0 _0230_
rlabel metal2 26992 38136 26992 38136 0 _0231_
rlabel metal3 23296 59192 23296 59192 0 _0232_
rlabel metal2 20216 64288 20216 64288 0 _0233_
rlabel metal3 9240 56168 9240 56168 0 _0234_
rlabel metal3 6384 50008 6384 50008 0 _0235_
rlabel metal2 9800 53368 9800 53368 0 _0236_
rlabel metal2 9128 20944 9128 20944 0 _0237_
rlabel metal2 8904 48160 8904 48160 0 _0238_
rlabel metal2 7448 62188 7448 62188 0 _0239_
rlabel metal2 8904 50512 8904 50512 0 _0240_
rlabel metal2 16072 41384 16072 41384 0 _0241_
rlabel metal3 17752 43512 17752 43512 0 _0242_
rlabel metal2 11816 43120 11816 43120 0 _0243_
rlabel metal2 13664 44296 13664 44296 0 _0244_
rlabel metal2 10696 58296 10696 58296 0 _0245_
rlabel metal3 11984 45752 11984 45752 0 _0246_
rlabel metal2 17864 39144 17864 39144 0 _0247_
rlabel metal3 19208 41272 19208 41272 0 _0248_
rlabel metal3 13776 41048 13776 41048 0 _0249_
rlabel metal2 14168 41160 14168 41160 0 _0250_
rlabel metal2 18200 34832 18200 34832 0 _0251_
rlabel metal2 18592 34888 18592 34888 0 _0252_
rlabel metal2 2072 44800 2072 44800 0 _0253_
rlabel metal3 16464 39480 16464 39480 0 _0254_
rlabel metal3 20272 69160 20272 69160 0 _0255_
rlabel metal2 22008 35672 22008 35672 0 _0256_
rlabel metal2 22568 43344 22568 43344 0 _0257_
rlabel metal2 20440 44800 20440 44800 0 _0258_
rlabel metal2 26264 26684 26264 26684 0 _0259_
rlabel metal3 26712 57624 26712 57624 0 _0260_
rlabel metal2 26936 60144 26936 60144 0 _0261_
rlabel metal2 26488 59864 26488 59864 0 _0262_
rlabel metal2 27720 37128 27720 37128 0 _0263_
rlabel metal2 26936 48216 26936 48216 0 _0264_
rlabel metal2 16968 49224 16968 49224 0 _0265_
rlabel metal2 27272 52696 27272 52696 0 _0266_
rlabel metal2 22120 55272 22120 55272 0 _0267_
rlabel metal2 27048 19712 27048 19712 0 _0268_
rlabel metal3 27048 43512 27048 43512 0 _0269_
rlabel metal2 27552 17752 27552 17752 0 _0270_
rlabel metal3 23716 57736 23716 57736 0 _0271_
rlabel metal2 25592 44520 25592 44520 0 _0272_
rlabel metal3 26544 55160 26544 55160 0 _0273_
rlabel metal2 26040 71344 26040 71344 0 _0274_
rlabel metal3 26600 53704 26600 53704 0 _0275_
rlabel metal3 23856 49000 23856 49000 0 _0276_
rlabel metal2 26152 50148 26152 50148 0 _0277_
rlabel metal2 25144 53312 25144 53312 0 _0278_
rlabel metal3 23744 53816 23744 53816 0 _0279_
rlabel metal2 24024 6552 24024 6552 0 _0280_
rlabel metal2 27048 13104 27048 13104 0 _0281_
rlabel metal2 23240 15400 23240 15400 0 _0282_
rlabel metal2 27888 20552 27888 20552 0 _0283_
rlabel metal2 9016 13888 9016 13888 0 _0284_
rlabel metal3 7336 18984 7336 18984 0 _0285_
rlabel metal2 7112 16968 7112 16968 0 _0286_
rlabel metal2 9688 12264 9688 12264 0 _0287_
rlabel metal3 6664 12824 6664 12824 0 _0288_
rlabel metal3 7056 15288 7056 15288 0 _0289_
rlabel metal3 25984 18424 25984 18424 0 _0290_
rlabel metal2 21896 14560 21896 14560 0 _0291_
rlabel metal2 24584 22512 24584 22512 0 _0292_
rlabel metal2 23800 15456 23800 15456 0 _0293_
rlabel metal2 18872 15148 18872 15148 0 _0294_
rlabel metal2 13496 14056 13496 14056 0 _0295_
rlabel metal3 11816 15848 11816 15848 0 _0296_
rlabel metal3 8792 62440 8792 62440 0 _0297_
rlabel metal2 20776 25760 20776 25760 0 _0298_
rlabel metal2 6664 63840 6664 63840 0 _0299_
rlabel metal2 7448 65576 7448 65576 0 _0300_
rlabel metal2 6440 66584 6440 66584 0 _0301_
rlabel metal2 12376 63056 12376 63056 0 _0302_
rlabel metal2 6552 51016 6552 51016 0 _0303_
rlabel metal2 11032 28000 11032 28000 0 _0304_
rlabel metal3 13328 36344 13328 36344 0 _0305_
rlabel metal2 7896 37352 7896 37352 0 _0306_
rlabel metal2 7616 45864 7616 45864 0 _0307_
rlabel metal2 23576 32424 23576 32424 0 _0308_
rlabel metal2 24360 39536 24360 39536 0 _0309_
rlabel metal2 24248 42504 24248 42504 0 _0310_
rlabel metal2 17864 30016 17864 30016 0 _0311_
rlabel metal2 25368 25032 25368 25032 0 _0312_
rlabel metal3 26096 28616 26096 28616 0 _0313_
rlabel metal2 24248 29736 24248 29736 0 _0314_
rlabel metal3 24976 37240 24976 37240 0 _0315_
rlabel metal3 24976 46648 24976 46648 0 _0316_
rlabel metal2 22680 45528 22680 45528 0 _0317_
rlabel metal2 4480 86856 4480 86856 0 _0318_
rlabel metal2 3864 86464 3864 86464 0 _0319_
rlabel metal3 6440 97608 6440 97608 0 _0320_
rlabel metal2 6328 94024 6328 94024 0 _0321_
rlabel metal2 3416 91840 3416 91840 0 _0322_
rlabel metal2 7000 90832 7000 90832 0 _0323_
rlabel metal2 7280 90552 7280 90552 0 _0324_
rlabel metal2 9128 95144 9128 95144 0 _0325_
rlabel metal2 20272 99176 20272 99176 0 _0326_
rlabel metal2 23576 100800 23576 100800 0 _0327_
rlabel metal2 25200 100184 25200 100184 0 _0328_
rlabel metal2 24024 98168 24024 98168 0 _0329_
rlabel metal3 24864 96040 24864 96040 0 _0330_
rlabel metal3 25816 97496 25816 97496 0 _0331_
rlabel metal3 24416 95816 24416 95816 0 _0332_
rlabel metal2 24584 95648 24584 95648 0 _0333_
rlabel metal3 24808 95256 24808 95256 0 _0334_
rlabel metal2 20664 4536 20664 4536 0 _0335_
rlabel metal2 22456 5544 22456 5544 0 _0336_
rlabel metal2 22456 7168 22456 7168 0 _0337_
rlabel metal3 24808 5880 24808 5880 0 _0338_
rlabel metal3 17472 4200 17472 4200 0 _0339_
rlabel metal2 23016 4760 23016 4760 0 _0340_
rlabel metal3 24808 4312 24808 4312 0 _0341_
rlabel metal2 23240 4704 23240 4704 0 _0342_
rlabel metal2 21784 5544 21784 5544 0 _0343_
rlabel metal2 27440 27944 27440 27944 0 _0344_
rlabel metal3 21840 20552 21840 20552 0 _0345_
rlabel metal2 26936 24192 26936 24192 0 _0346_
rlabel metal2 20216 22848 20216 22848 0 _0347_
rlabel metal2 2968 93072 2968 93072 0 _0348_
rlabel metal2 14056 21056 14056 21056 0 _0349_
rlabel metal3 23744 21784 23744 21784 0 _0350_
rlabel metal3 18200 26040 18200 26040 0 _0351_
rlabel metal3 19824 21000 19824 21000 0 _0352_
rlabel metal2 18312 19376 18312 19376 0 _0353_
rlabel metal2 22792 25312 22792 25312 0 _0354_
rlabel metal3 14560 28616 14560 28616 0 _0355_
rlabel metal2 27048 23128 27048 23128 0 _0356_
rlabel metal2 8344 22960 8344 22960 0 _0357_
rlabel metal2 10024 21448 10024 21448 0 _0358_
rlabel metal2 6888 21168 6888 21168 0 _0359_
rlabel metal3 11368 21000 11368 21000 0 _0360_
rlabel metal2 9632 26488 9632 26488 0 _0361_
rlabel via2 26264 24024 26264 24024 0 _0362_
rlabel metal2 14672 26040 14672 26040 0 _0363_
rlabel metal2 12488 31892 12488 31892 0 _0364_
rlabel metal2 12376 40152 12376 40152 0 _0365_
rlabel metal2 9688 40040 9688 40040 0 _0366_
rlabel metal2 8232 42056 8232 42056 0 _0367_
rlabel metal2 18312 27608 18312 27608 0 _0368_
rlabel metal2 14560 35784 14560 35784 0 _0369_
rlabel metal3 21952 41720 21952 41720 0 _0370_
rlabel metal2 16352 41720 16352 41720 0 _0371_
rlabel metal2 26376 31640 26376 31640 0 _0372_
rlabel metal3 27104 39816 27104 39816 0 _0373_
rlabel metal2 26376 42336 26376 42336 0 _0374_
rlabel metal2 14672 30744 14672 30744 0 _0375_
rlabel metal2 24976 22456 24976 22456 0 _0376_
rlabel metal3 26768 21000 26768 21000 0 _0377_
rlabel metal3 26712 27608 26712 27608 0 _0378_
rlabel metal2 26824 36904 26824 36904 0 _0379_
rlabel metal3 26768 33880 26768 33880 0 _0380_
rlabel metal2 22344 37912 22344 37912 0 _0381_
rlabel metal2 6664 8176 6664 8176 0 _0382_
rlabel metal3 21336 5992 21336 5992 0 _0383_
rlabel metal2 2128 18760 2128 18760 0 _0384_
rlabel metal2 3304 43568 3304 43568 0 _0385_
rlabel metal3 2800 71848 2800 71848 0 _0386_
rlabel metal2 6944 8456 6944 8456 0 _0387_
rlabel metal2 2632 15624 2632 15624 0 _0388_
rlabel metal3 3920 11256 3920 11256 0 _0389_
rlabel metal2 2632 11816 2632 11816 0 _0390_
rlabel metal2 4872 6720 4872 6720 0 _0391_
rlabel metal2 4648 7224 4648 7224 0 _0392_
rlabel metal2 6328 9744 6328 9744 0 _0393_
rlabel metal2 6496 9016 6496 9016 0 _0394_
rlabel metal2 3304 14168 3304 14168 0 _0395_
rlabel metal2 2856 13832 2856 13832 0 _0396_
rlabel metal2 3080 16744 3080 16744 0 _0397_
rlabel metal2 2856 16856 2856 16856 0 _0398_
rlabel metal2 3192 20328 3192 20328 0 _0399_
rlabel metal2 2912 19992 2912 19992 0 _0400_
rlabel metal2 3304 21952 3304 21952 0 _0401_
rlabel metal2 3080 22232 3080 22232 0 _0402_
rlabel metal3 3248 24696 3248 24696 0 _0403_
rlabel metal2 2520 26096 2520 26096 0 _0404_
rlabel metal2 2632 24864 2632 24864 0 _0405_
rlabel metal2 6328 26152 6328 26152 0 _0406_
rlabel metal2 5992 26432 5992 26432 0 _0407_
rlabel metal2 2856 30856 2856 30856 0 _0408_
rlabel metal2 2632 30968 2632 30968 0 _0409_
rlabel metal2 2912 33320 2912 33320 0 _0410_
rlabel metal3 3080 33432 3080 33432 0 _0411_
rlabel metal2 6104 36568 6104 36568 0 _0412_
rlabel metal2 5096 36512 5096 36512 0 _0413_
rlabel metal2 3080 42784 3080 42784 0 _0414_
rlabel metal2 2744 41552 2744 41552 0 _0415_
rlabel metal3 3584 28616 3584 28616 0 _0416_
rlabel metal3 3136 28728 3136 28728 0 _0417_
rlabel metal2 2968 39928 2968 39928 0 _0418_
rlabel metal2 2632 41776 2632 41776 0 _0419_
rlabel metal2 5768 34272 5768 34272 0 _0420_
rlabel metal2 5488 42504 5488 42504 0 _0421_
rlabel metal2 6216 40264 6216 40264 0 _0422_
rlabel metal2 5488 47880 5488 47880 0 _0423_
rlabel metal2 3192 36848 3192 36848 0 _0424_
rlabel metal4 2408 42000 2408 42000 0 _0425_
rlabel metal3 3108 45080 3108 45080 0 _0426_
rlabel metal2 2464 51352 2464 51352 0 _0427_
rlabel metal2 3192 57680 3192 57680 0 _0428_
rlabel metal3 3360 58632 3360 58632 0 _0429_
rlabel metal2 3080 71960 3080 71960 0 _0430_
rlabel metal2 3080 59416 3080 59416 0 _0431_
rlabel metal3 3024 60536 3024 60536 0 _0432_
rlabel metal2 3080 63840 3080 63840 0 _0433_
rlabel metal2 2912 63896 2912 63896 0 _0434_
rlabel metal2 2856 65688 2856 65688 0 _0435_
rlabel metal2 2688 65464 2688 65464 0 _0436_
rlabel metal3 3136 68600 3136 68600 0 _0437_
rlabel metal2 2464 68376 2464 68376 0 _0438_
rlabel metal3 3024 71736 3024 71736 0 _0439_
rlabel metal2 2744 72408 2744 72408 0 _0440_
rlabel metal2 2968 75320 2968 75320 0 _0441_
rlabel metal2 2744 75600 2744 75600 0 _0442_
rlabel metal3 3248 78008 3248 78008 0 _0443_
rlabel metal2 2744 77560 2744 77560 0 _0444_
rlabel metal2 5880 79576 5880 79576 0 _0445_
rlabel metal3 3136 82488 3136 82488 0 _0446_
rlabel metal2 7448 81872 7448 81872 0 _0447_
rlabel metal2 5992 82824 5992 82824 0 _0448_
rlabel metal3 24304 25032 24304 25032 0 _0449_
rlabel metal2 15400 24696 15400 24696 0 _0450_
rlabel metal2 22400 23016 22400 23016 0 _0451_
rlabel metal2 21448 26684 21448 26684 0 _0452_
rlabel metal2 16072 22288 16072 22288 0 _0453_
rlabel metal3 13048 56952 13048 56952 0 _0454_
rlabel metal3 20776 10584 20776 10584 0 _0455_
rlabel metal2 18088 9464 18088 9464 0 _0456_
rlabel metal2 15960 10752 15960 10752 0 _0457_
rlabel metal2 14616 10864 14616 10864 0 _0458_
rlabel metal2 13944 18480 13944 18480 0 _0459_
rlabel metal3 15064 15288 15064 15288 0 _0460_
rlabel metal2 17528 21952 17528 21952 0 _0461_
rlabel metal2 22344 10976 22344 10976 0 _0462_
rlabel metal3 18200 12824 18200 12824 0 _0463_
rlabel metal2 13720 9800 13720 9800 0 _0464_
rlabel metal3 11480 10584 11480 10584 0 _0465_
rlabel metal3 11200 23800 11200 23800 0 _0466_
rlabel metal2 15232 23800 15232 23800 0 _0467_
rlabel metal2 11256 67816 11256 67816 0 _0468_
rlabel metal2 10808 65744 10808 65744 0 _0469_
rlabel metal2 17528 67760 17528 67760 0 _0470_
rlabel metal2 14056 65408 14056 65408 0 _0471_
rlabel metal2 11368 60144 11368 60144 0 _0472_
rlabel metal3 11480 53816 11480 53816 0 _0473_
rlabel metal3 19208 69496 19208 69496 0 _0474_
rlabel metal3 14840 74872 14840 74872 0 _0475_
rlabel metal3 26824 74088 26824 74088 0 _0476_
rlabel metal2 26600 70952 26600 70952 0 _0477_
rlabel metal2 26488 64568 26488 64568 0 _0478_
rlabel metal2 16296 63336 16296 63336 0 _0479_
rlabel metal2 26488 76104 26488 76104 0 _0480_
rlabel metal2 24920 76888 24920 76888 0 _0481_
rlabel metal2 24584 67760 24584 67760 0 _0482_
rlabel metal2 27048 68600 27048 68600 0 _0483_
rlabel metal2 26152 64064 26152 64064 0 _0484_
rlabel metal3 23296 63000 23296 63000 0 _0485_
rlabel metal2 20272 1960 20272 1960 0 _0486_
rlabel metal2 19880 2296 19880 2296 0 _0487_
rlabel metal2 19936 7560 19936 7560 0 _0488_
rlabel metal2 2856 88032 2856 88032 0 _0489_
rlabel metal2 21224 3024 21224 3024 0 _0490_
rlabel metal2 21896 5936 21896 5936 0 _0491_
rlabel metal3 20944 6552 20944 6552 0 _0492_
rlabel metal2 15232 86072 15232 86072 0 _0493_
rlabel metal2 16408 82768 16408 82768 0 _0494_
rlabel metal2 22344 25704 22344 25704 0 _0495_
rlabel metal2 2800 46536 2800 46536 0 _0496_
rlabel metal2 23352 48608 23352 48608 0 _0497_
rlabel metal2 20216 76384 20216 76384 0 _0498_
rlabel metal3 9968 76664 9968 76664 0 _0499_
rlabel metal2 22624 77448 22624 77448 0 _0500_
rlabel metal3 18200 77784 18200 77784 0 _0501_
rlabel metal2 18760 74480 18760 74480 0 _0502_
rlabel metal2 14280 79968 14280 79968 0 _0503_
rlabel metal2 24584 72016 24584 72016 0 _0504_
rlabel metal2 22344 73136 22344 73136 0 _0505_
rlabel metal2 21896 29176 21896 29176 0 _0506_
rlabel metal2 21560 66696 21560 66696 0 _0507_
rlabel metal2 20104 54712 20104 54712 0 _0508_
rlabel metal2 21784 63840 21784 63840 0 _0509_
rlabel metal3 12208 58632 12208 58632 0 _0510_
rlabel metal3 3640 54264 3640 54264 0 _0511_
rlabel metal3 8064 30296 8064 30296 0 _0512_
rlabel metal2 5152 30408 5152 30408 0 _0513_
rlabel metal2 8120 31080 8120 31080 0 _0514_
rlabel metal3 6552 44520 6552 44520 0 _0515_
rlabel metal2 7280 58968 7280 58968 0 _0516_
rlabel metal2 6216 57176 6216 57176 0 _0517_
rlabel metal2 3696 49560 3696 49560 0 _0518_
rlabel metal3 3808 47656 3808 47656 0 _0519_
rlabel metal2 6832 52696 6832 52696 0 _0520_
rlabel metal2 20328 55832 20328 55832 0 _0521_
rlabel metal3 6496 61544 6496 61544 0 _0522_
rlabel metal2 18872 64064 18872 64064 0 _0523_
rlabel metal3 6496 70952 6496 70952 0 _0524_
rlabel metal3 6608 72632 6608 72632 0 _0525_
rlabel metal3 6496 74872 6496 74872 0 _0526_
rlabel metal2 7784 76216 7784 76216 0 _0527_
rlabel metal3 19992 60536 19992 60536 0 _0528_
rlabel metal2 20104 60256 20104 60256 0 _0529_
rlabel metal3 24584 49224 24584 49224 0 _0530_
rlabel metal2 24360 51632 24360 51632 0 _0531_
rlabel metal2 24584 3808 24584 3808 0 _0532_
rlabel metal2 3304 94136 3304 94136 0 _0533_
rlabel metal2 22456 94080 22456 94080 0 _0534_
rlabel metal2 18032 109256 18032 109256 0 _0535_
rlabel metal2 3192 94192 3192 94192 0 _0536_
rlabel metal2 2520 96768 2520 96768 0 _0537_
rlabel metal2 3304 96264 3304 96264 0 _0538_
rlabel metal2 3080 99288 3080 99288 0 _0539_
rlabel metal2 3472 100072 3472 100072 0 _0540_
rlabel metal2 3528 101024 3528 101024 0 _0541_
rlabel metal3 21448 100576 21448 100576 0 _0542_
rlabel metal3 3808 103208 3808 103208 0 _0543_
rlabel metal2 17192 106344 17192 106344 0 _0544_
rlabel metal2 7224 103992 7224 103992 0 _0545_
rlabel metal2 3976 105392 3976 105392 0 _0546_
rlabel metal2 6720 104888 6720 104888 0 _0547_
rlabel metal2 14560 86632 14560 86632 0 _0548_
rlabel metal2 12712 86072 12712 86072 0 _0549_
rlabel metal2 11592 83104 11592 83104 0 _0550_
rlabel metal3 7168 99176 7168 99176 0 _0551_
rlabel metal2 7784 94360 7784 94360 0 _0552_
rlabel metal2 8008 92680 8008 92680 0 _0553_
rlabel metal3 9184 85960 9184 85960 0 _0554_
rlabel metal2 11144 90440 11144 90440 0 _0555_
rlabel metal2 8848 88200 8848 88200 0 _0556_
rlabel metal2 9128 90552 9128 90552 0 _0557_
rlabel metal3 10080 86520 10080 86520 0 _0558_
rlabel metal3 9632 92344 9632 92344 0 _0559_
rlabel metal2 7448 99120 7448 99120 0 _0560_
rlabel metal3 17024 95256 17024 95256 0 _0561_
rlabel metal2 21784 93352 21784 93352 0 _0562_
rlabel metal2 9800 98000 9800 98000 0 _0563_
rlabel metal2 10584 96208 10584 96208 0 _0564_
rlabel metal2 2856 98672 2856 98672 0 _0565_
rlabel via2 6888 95480 6888 95480 0 _0566_
rlabel metal2 6104 94080 6104 94080 0 _0567_
rlabel metal2 17528 95032 17528 95032 0 _0568_
rlabel metal2 18088 95368 18088 95368 0 _0569_
rlabel metal2 24136 100632 24136 100632 0 _0570_
rlabel metal2 24640 98392 24640 98392 0 _0571_
rlabel metal2 23688 96740 23688 96740 0 _0572_
rlabel metal2 7504 100520 7504 100520 0 _0573_
rlabel metal2 22792 96600 22792 96600 0 _0574_
rlabel metal3 22008 95480 22008 95480 0 _0575_
rlabel metal2 11032 98616 11032 98616 0 _0576_
rlabel metal2 11144 101248 11144 101248 0 _0577_
rlabel metal2 8680 102480 8680 102480 0 _0578_
rlabel metal2 8400 102536 8400 102536 0 _0579_
rlabel metal2 16016 45304 16016 45304 0 _0580_
rlabel metal2 17528 44408 17528 44408 0 _0581_
rlabel metal2 16744 87696 16744 87696 0 _0582_
rlabel metal2 22848 47320 22848 47320 0 _0583_
rlabel metal3 21112 86520 21112 86520 0 _0584_
rlabel metal3 17976 85736 17976 85736 0 _0585_
rlabel metal2 20776 71232 20776 71232 0 _0586_
rlabel metal2 24416 48104 24416 48104 0 _0587_
rlabel metal2 15960 48720 15960 48720 0 _0588_
rlabel metal2 11368 49168 11368 49168 0 _0589_
rlabel metal4 16296 63000 16296 63000 0 _0590_
rlabel metal3 15176 48272 15176 48272 0 _0591_
rlabel metal2 15400 48048 15400 48048 0 _0592_
rlabel metal2 20720 47208 20720 47208 0 _0593_
rlabel metal2 23576 46648 23576 46648 0 _0594_
rlabel metal3 22232 44296 22232 44296 0 _0595_
rlabel metal2 5712 53144 5712 53144 0 _0596_
rlabel metal2 20664 49000 20664 49000 0 _0597_
rlabel metal2 27272 50960 27272 50960 0 _0598_
rlabel metal2 13272 69328 13272 69328 0 _0599_
rlabel metal2 6104 54824 6104 54824 0 _0600_
rlabel metal2 20328 53032 20328 53032 0 _0601_
rlabel metal3 26264 52080 26264 52080 0 _0602_
rlabel metal2 16688 66920 16688 66920 0 _0603_
rlabel metal2 12264 70504 12264 70504 0 _0604_
rlabel metal2 27160 53816 27160 53816 0 _0605_
rlabel metal2 26488 54488 26488 54488 0 _0606_
rlabel metal2 16296 46256 16296 46256 0 _0607_
rlabel metal2 20328 10528 20328 10528 0 _0608_
rlabel metal3 16632 45864 16632 45864 0 _0609_
rlabel metal2 19712 10808 19712 10808 0 _0610_
rlabel metal4 20272 15120 20272 15120 0 _0611_
rlabel metal3 17416 23016 17416 23016 0 _0612_
rlabel metal2 21896 47320 21896 47320 0 _0613_
rlabel metal2 21672 47600 21672 47600 0 _0614_
rlabel metal2 21336 49056 21336 49056 0 _0615_
rlabel metal3 19880 70728 19880 70728 0 _0616_
rlabel metal2 23576 65352 23576 65352 0 _0617_
rlabel metal2 23800 71512 23800 71512 0 _0618_
rlabel metal3 21000 71624 21000 71624 0 _0619_
rlabel metal3 23408 26488 23408 26488 0 _0620_
rlabel metal2 15904 17080 15904 17080 0 _0621_
rlabel metal2 23912 22848 23912 22848 0 _0622_
rlabel metal2 15624 50176 15624 50176 0 _0623_
rlabel metal2 16632 44408 16632 44408 0 _0624_
rlabel metal3 20104 42672 20104 42672 0 _0625_
rlabel metal2 20104 42224 20104 42224 0 _0626_
rlabel metal2 13944 48216 13944 48216 0 _0627_
rlabel metal2 18088 33488 18088 33488 0 _0628_
rlabel metal3 20160 41944 20160 41944 0 _0629_
rlabel metal2 18872 42672 18872 42672 0 _0630_
rlabel metal2 23464 47824 23464 47824 0 _0631_
rlabel metal2 19320 42392 19320 42392 0 _0632_
rlabel metal2 19208 42952 19208 42952 0 _0633_
rlabel metal2 12544 70168 12544 70168 0 _0634_
rlabel metal2 11144 48328 11144 48328 0 _0635_
rlabel metal2 13384 69832 13384 69832 0 _0636_
rlabel metal3 12712 69720 12712 69720 0 _0637_
rlabel metal3 13272 71176 13272 71176 0 _0638_
rlabel metal2 13832 70896 13832 70896 0 _0639_
rlabel metal2 14224 70840 14224 70840 0 _0640_
rlabel metal2 14504 71064 14504 71064 0 _0641_
rlabel metal2 14280 71120 14280 71120 0 _0642_
rlabel metal4 9688 65744 9688 65744 0 _0643_
rlabel metal2 13832 60816 13832 60816 0 _0644_
rlabel metal2 9520 71736 9520 71736 0 _0645_
rlabel metal2 15232 57624 15232 57624 0 _0646_
rlabel metal3 10136 70392 10136 70392 0 _0647_
rlabel metal2 9576 71288 9576 71288 0 _0648_
rlabel metal2 17976 71568 17976 71568 0 _0649_
rlabel metal2 11928 28392 11928 28392 0 _0650_
rlabel metal3 10528 33320 10528 33320 0 _0651_
rlabel metal2 10136 45024 10136 45024 0 _0652_
rlabel metal2 9800 44632 9800 44632 0 _0653_
rlabel metal3 10248 33208 10248 33208 0 _0654_
rlabel metal3 11200 47096 11200 47096 0 _0655_
rlabel metal2 12320 41048 12320 41048 0 _0656_
rlabel metal2 9744 30296 9744 30296 0 _0657_
rlabel metal2 16072 43680 16072 43680 0 _0658_
rlabel metal2 15400 45864 15400 45864 0 _0659_
rlabel metal3 11592 33320 11592 33320 0 _0660_
rlabel metal2 17528 71176 17528 71176 0 _0661_
rlabel metal3 18312 71512 18312 71512 0 _0662_
rlabel metal2 19712 84280 19712 84280 0 _0663_
rlabel metal2 21560 83832 21560 83832 0 _0664_
rlabel metal2 18592 73192 18592 73192 0 _0665_
rlabel metal2 19768 52528 19768 52528 0 _0666_
rlabel metal2 19992 52192 19992 52192 0 _0667_
rlabel metal4 18984 19628 18984 19628 0 _0668_
rlabel metal2 23016 51856 23016 51856 0 _0669_
rlabel metal2 21560 46704 21560 46704 0 _0670_
rlabel metal3 21504 52136 21504 52136 0 _0671_
rlabel metal3 20328 72296 20328 72296 0 _0672_
rlabel metal2 23240 72296 23240 72296 0 _0673_
rlabel metal2 19264 22680 19264 22680 0 _0674_
rlabel metal3 16380 41944 16380 41944 0 _0675_
rlabel metal2 17920 34664 17920 34664 0 _0676_
rlabel metal2 18200 42448 18200 42448 0 _0677_
rlabel metal3 18256 41944 18256 41944 0 _0678_
rlabel metal2 13160 57008 13160 57008 0 _0679_
rlabel metal3 13496 72296 13496 72296 0 _0680_
rlabel metal2 2632 81984 2632 81984 0 _0681_
rlabel metal2 13944 72688 13944 72688 0 _0682_
rlabel metal1 12992 74648 12992 74648 0 _0683_
rlabel metal3 14392 73416 14392 73416 0 _0684_
rlabel metal2 13720 72800 13720 72800 0 _0685_
rlabel metal2 8456 71456 8456 71456 0 _0686_
rlabel metal2 8512 71960 8512 71960 0 _0687_
rlabel metal2 8904 72240 8904 72240 0 _0688_
rlabel metal2 14280 73024 14280 73024 0 _0689_
rlabel metal2 10136 34608 10136 34608 0 _0690_
rlabel metal2 10808 34888 10808 34888 0 _0691_
rlabel metal2 10920 31360 10920 31360 0 _0692_
rlabel metal3 11872 34888 11872 34888 0 _0693_
rlabel metal2 15960 73248 15960 73248 0 _0694_
rlabel metal2 17304 72800 17304 72800 0 _0695_
rlabel metal2 18984 79072 18984 79072 0 _0696_
rlabel metal2 19096 79128 19096 79128 0 _0697_
rlabel metal2 20552 71960 20552 71960 0 _0698_
rlabel metal2 18424 51632 18424 51632 0 _0699_
rlabel metal2 27496 52472 27496 52472 0 _0700_
rlabel metal3 18368 10808 18368 10808 0 _0701_
rlabel metal2 19320 24304 19320 24304 0 _0702_
rlabel metal3 18704 24136 18704 24136 0 _0703_
rlabel metal3 18928 24920 18928 24920 0 _0704_
rlabel metal2 19432 51688 19432 51688 0 _0705_
rlabel metal2 19712 67032 19712 67032 0 _0706_
rlabel metal2 23016 27888 23016 27888 0 _0707_
rlabel metal2 20104 34552 20104 34552 0 _0708_
rlabel metal2 20216 32928 20216 32928 0 _0709_
rlabel metal2 19656 34608 19656 34608 0 _0710_
rlabel metal2 19992 65800 19992 65800 0 _0711_
rlabel metal2 16744 67984 16744 67984 0 _0712_
rlabel metal2 9800 80976 9800 80976 0 _0713_
rlabel metal2 17304 71120 17304 71120 0 _0714_
rlabel metal3 20216 71736 20216 71736 0 _0715_
rlabel metal2 25592 72856 25592 72856 0 _0716_
rlabel metal2 16352 71624 16352 71624 0 _0717_
rlabel metal2 8344 70000 8344 70000 0 _0718_
rlabel metal2 10248 73248 10248 73248 0 _0719_
rlabel metal3 16184 71568 16184 71568 0 _0720_
rlabel metal2 17864 70056 17864 70056 0 _0721_
rlabel metal3 10808 37240 10808 37240 0 _0722_
rlabel metal2 8680 36960 8680 36960 0 _0723_
rlabel metal2 9968 31864 9968 31864 0 _0724_
rlabel metal2 10528 37240 10528 37240 0 _0725_
rlabel metal3 19208 66024 19208 66024 0 _0726_
rlabel metal2 18760 67592 18760 67592 0 _0727_
rlabel metal2 19152 72744 19152 72744 0 _0728_
rlabel metal2 21336 78904 21336 78904 0 _0729_
rlabel metal2 17472 69944 17472 69944 0 _0730_
rlabel metal3 20664 53760 20664 53760 0 _0731_
rlabel metal2 20552 53536 20552 53536 0 _0732_
rlabel metal4 20384 20970 20384 20970 0 _0733_
rlabel metal2 13496 24136 13496 24136 0 _0734_
rlabel metal2 12824 23576 12824 23576 0 _0735_
rlabel metal2 20104 53648 20104 53648 0 _0736_
rlabel metal2 19432 63560 19432 63560 0 _0737_
rlabel metal3 20776 65352 20776 65352 0 _0738_
rlabel metal2 19096 38080 19096 38080 0 _0739_
rlabel metal2 18872 39592 18872 39592 0 _0740_
rlabel metal2 18760 34020 18760 34020 0 _0741_
rlabel metal3 19152 38808 19152 38808 0 _0742_
rlabel metal2 17696 56168 17696 56168 0 _0743_
rlabel metal2 15904 67144 15904 67144 0 _0744_
rlabel metal2 6776 82880 6776 82880 0 _0745_
rlabel metal2 16184 70056 16184 70056 0 _0746_
rlabel metal2 15120 71176 15120 71176 0 _0747_
rlabel metal2 15848 70336 15848 70336 0 _0748_
rlabel metal2 15792 69384 15792 69384 0 _0749_
rlabel metal2 8456 68992 8456 68992 0 _0750_
rlabel metal2 8680 71064 8680 71064 0 _0751_
rlabel metal3 12320 69272 12320 69272 0 _0752_
rlabel metal2 16520 68432 16520 68432 0 _0753_
rlabel metal2 10360 42336 10360 42336 0 _0754_
rlabel metal2 10024 43624 10024 43624 0 _0755_
rlabel metal2 10752 42840 10752 42840 0 _0756_
rlabel metal2 10808 43792 10808 43792 0 _0757_
rlabel metal2 16968 65128 16968 65128 0 _0758_
rlabel metal3 17920 65464 17920 65464 0 _0759_
rlabel metal2 17864 66640 17864 66640 0 _0760_
rlabel metal2 21672 80864 21672 80864 0 _0761_
rlabel metal2 19432 72464 19432 72464 0 _0762_
rlabel metal2 19096 31472 19096 31472 0 _0763_
rlabel metal2 20552 30408 20552 30408 0 _0764_
rlabel metal2 21224 41328 21224 41328 0 _0765_
rlabel metal2 15512 31136 15512 31136 0 _0766_
rlabel metal2 16072 31360 16072 31360 0 _0767_
rlabel metal2 19880 31192 19880 31192 0 _0768_
rlabel metal3 22008 33096 22008 33096 0 _0769_
rlabel metal3 21336 33376 21336 33376 0 _0770_
rlabel metal2 21504 30968 21504 30968 0 _0771_
rlabel metal2 20328 25592 20328 25592 0 _0772_
rlabel metal2 20440 29176 20440 29176 0 _0773_
rlabel metal2 20664 25368 20664 25368 0 _0774_
rlabel metal2 10584 29568 10584 29568 0 _0775_
rlabel metal2 21112 30240 21112 30240 0 _0776_
rlabel metal2 21000 25256 21000 25256 0 _0777_
rlabel metal3 20552 24920 20552 24920 0 _0778_
rlabel metal3 20496 33320 20496 33320 0 _0779_
rlabel metal2 22568 31360 22568 31360 0 _0780_
rlabel metal2 22008 71232 22008 71232 0 _0781_
rlabel metal2 14168 61880 14168 61880 0 _0782_
rlabel metal2 9968 58968 9968 58968 0 _0783_
rlabel metal3 15344 61544 15344 61544 0 _0784_
rlabel metal2 17416 60144 17416 60144 0 _0785_
rlabel metal2 17136 78008 17136 78008 0 _0786_
rlabel metal2 14392 60480 14392 60480 0 _0787_
rlabel metal2 13888 59976 13888 59976 0 _0788_
rlabel metal2 17360 60760 17360 60760 0 _0789_
rlabel metal2 16968 60200 16968 60200 0 _0790_
rlabel metal2 14168 25760 14168 25760 0 _0791_
rlabel metal2 14224 45192 14224 45192 0 _0792_
rlabel metal2 15288 44744 15288 44744 0 _0793_
rlabel metal2 15512 45920 15512 45920 0 _0794_
rlabel metal3 18592 62104 18592 62104 0 _0795_
rlabel metal3 15288 61152 15288 61152 0 _0796_
rlabel metal3 13552 62328 13552 62328 0 _0797_
rlabel metal2 14728 61656 14728 61656 0 _0798_
rlabel metal2 22624 65128 22624 65128 0 _0799_
rlabel metal2 19488 73416 19488 73416 0 _0800_
rlabel metal3 20160 86632 20160 86632 0 _0801_
rlabel metal2 20776 83608 20776 83608 0 _0802_
rlabel metal3 13328 56056 13328 56056 0 _0803_
rlabel metal2 14056 45416 14056 45416 0 _0804_
rlabel metal2 8456 44856 8456 44856 0 _0805_
rlabel metal2 14784 56056 14784 56056 0 _0806_
rlabel metal3 17976 56112 17976 56112 0 _0807_
rlabel metal2 11928 56448 11928 56448 0 _0808_
rlabel metal2 23464 56000 23464 56000 0 _0809_
rlabel metal2 15848 24360 15848 24360 0 _0810_
rlabel metal3 16576 24136 16576 24136 0 _0811_
rlabel metal2 15680 24920 15680 24920 0 _0812_
rlabel metal2 16632 24416 16632 24416 0 _0813_
rlabel metal2 16968 25032 16968 25032 0 _0814_
rlabel metal3 18648 56056 18648 56056 0 _0815_
rlabel metal2 10472 55944 10472 55944 0 _0816_
rlabel metal3 15512 56000 15512 56000 0 _0817_
rlabel metal2 15736 35112 15736 35112 0 _0818_
rlabel metal2 15960 33936 15960 33936 0 _0819_
rlabel metal2 15960 35168 15960 35168 0 _0820_
rlabel metal3 17696 53480 17696 53480 0 _0821_
rlabel metal2 15680 56168 15680 56168 0 _0822_
rlabel metal2 12712 51800 12712 51800 0 _0823_
rlabel metal2 14112 40936 14112 40936 0 _0824_
rlabel metal2 13608 27496 13608 27496 0 _0825_
rlabel metal2 15624 36120 15624 36120 0 _0826_
rlabel metal2 22904 37520 22904 37520 0 _0827_
rlabel metal3 15400 37464 15400 37464 0 _0828_
rlabel metal3 17304 55944 17304 55944 0 _0829_
rlabel metal2 17808 56280 17808 56280 0 _0830_
rlabel metal2 18032 83496 18032 83496 0 _0831_
rlabel metal2 18424 83552 18424 83552 0 _0832_
rlabel metal2 13496 82936 13496 82936 0 _0833_
rlabel metal2 16520 93184 16520 93184 0 _0834_
rlabel metal2 15624 90104 15624 90104 0 _0835_
rlabel metal3 12824 93688 12824 93688 0 _0836_
rlabel metal2 12040 95648 12040 95648 0 _0837_
rlabel metal2 15736 91056 15736 91056 0 _0838_
rlabel metal2 13384 90776 13384 90776 0 _0839_
rlabel metal2 14168 94976 14168 94976 0 _0840_
rlabel metal2 14280 91504 14280 91504 0 _0841_
rlabel metal2 17976 90048 17976 90048 0 _0842_
rlabel metal2 19208 93968 19208 93968 0 _0843_
rlabel metal2 18200 94416 18200 94416 0 _0844_
rlabel metal2 16408 89264 16408 89264 0 _0845_
rlabel metal2 18424 95144 18424 95144 0 _0846_
rlabel metal2 17864 80472 17864 80472 0 _0847_
rlabel metal2 18312 88256 18312 88256 0 _0848_
rlabel metal3 20776 92232 20776 92232 0 _0849_
rlabel metal2 18984 91504 18984 91504 0 _0850_
rlabel metal2 18088 92232 18088 92232 0 _0851_
rlabel metal2 18312 94528 18312 94528 0 _0852_
rlabel metal2 18704 92792 18704 92792 0 _0853_
rlabel metal3 16016 94360 16016 94360 0 _0854_
rlabel metal2 16800 92792 16800 92792 0 _0855_
rlabel metal3 17080 94024 17080 94024 0 _0856_
rlabel metal2 13776 94472 13776 94472 0 _0857_
rlabel metal2 14056 94752 14056 94752 0 _0858_
rlabel metal2 12376 95200 12376 95200 0 _0859_
rlabel metal2 11032 94192 11032 94192 0 _0860_
rlabel metal2 20216 84448 20216 84448 0 _0861_
rlabel metal2 20048 86856 20048 86856 0 _0862_
rlabel metal2 20440 90496 20440 90496 0 _0863_
rlabel metal2 20104 92904 20104 92904 0 _0864_
rlabel metal2 14280 97328 14280 97328 0 _0865_
rlabel metal2 15624 95872 15624 95872 0 _0866_
rlabel metal2 14728 95312 14728 95312 0 _0867_
rlabel metal3 14168 93240 14168 93240 0 _0868_
rlabel metal2 12376 91392 12376 91392 0 _0869_
rlabel metal2 15848 96320 15848 96320 0 _0870_
rlabel metal2 12824 94192 12824 94192 0 _0871_
rlabel metal2 8568 99736 8568 99736 0 _0872_
rlabel metal2 15176 95648 15176 95648 0 _0873_
rlabel metal3 11032 94472 11032 94472 0 _0874_
rlabel metal3 11480 96152 11480 96152 0 _0875_
rlabel metal2 10248 95424 10248 95424 0 _0876_
rlabel metal3 25032 117208 25032 117208 0 _0877_
rlabel metal2 18088 80752 18088 80752 0 _0878_
rlabel metal2 18984 86184 18984 86184 0 _0879_
rlabel metal2 19208 88872 19208 88872 0 _0880_
rlabel metal2 19208 93128 19208 93128 0 _0881_
rlabel metal3 18592 97496 18592 97496 0 _0882_
rlabel metal2 18200 96264 18200 96264 0 _0883_
rlabel metal2 15288 93968 15288 93968 0 _0884_
rlabel metal3 8792 96768 8792 96768 0 _0885_
rlabel metal2 15176 88200 15176 88200 0 _0886_
rlabel metal2 8568 97132 8568 97132 0 _0887_
rlabel metal2 9688 103264 9688 103264 0 _0888_
rlabel metal2 12264 101808 12264 101808 0 _0889_
rlabel metal2 10248 103488 10248 103488 0 _0890_
rlabel metal2 19768 79296 19768 79296 0 _0891_
rlabel metal2 19992 79576 19992 79576 0 _0892_
rlabel metal2 21448 93576 21448 93576 0 _0893_
rlabel metal2 21672 93464 21672 93464 0 _0894_
rlabel metal3 19264 98392 19264 98392 0 _0895_
rlabel metal2 18536 97328 18536 97328 0 _0896_
rlabel metal2 19992 100800 19992 100800 0 _0897_
rlabel metal3 16464 90552 16464 90552 0 _0898_
rlabel metal3 14728 102200 14728 102200 0 _0899_
rlabel metal2 21672 102312 21672 102312 0 _0900_
rlabel metal2 22456 102872 22456 102872 0 _0901_
rlabel metal2 22232 101808 22232 101808 0 _0902_
rlabel metal2 22568 103040 22568 103040 0 _0903_
rlabel metal2 19320 80640 19320 80640 0 _0904_
rlabel metal2 20160 81704 20160 81704 0 _0905_
rlabel metal2 20440 92568 20440 92568 0 _0906_
rlabel metal2 19992 94528 19992 94528 0 _0907_
rlabel metal2 19544 96712 19544 96712 0 _0908_
rlabel metal2 16856 96880 16856 96880 0 _0909_
rlabel metal2 17752 100408 17752 100408 0 _0910_
rlabel metal2 17080 93660 17080 93660 0 _0911_
rlabel metal2 18760 99736 18760 99736 0 _0912_
rlabel metal3 16968 106008 16968 106008 0 _0913_
rlabel metal2 16856 107128 16856 107128 0 _0914_
rlabel metal3 20328 88312 20328 88312 0 _0915_
rlabel metal2 19768 87584 19768 87584 0 _0916_
rlabel metal2 17416 92176 17416 92176 0 _0917_
rlabel metal2 16968 94528 16968 94528 0 _0918_
rlabel metal2 17696 94360 17696 94360 0 _0919_
rlabel metal2 16072 93968 16072 93968 0 _0920_
rlabel metal2 15176 94024 15176 94024 0 _0921_
rlabel metal2 15624 93800 15624 93800 0 _0922_
rlabel metal2 16296 94416 16296 94416 0 _0923_
rlabel metal2 13160 104160 13160 104160 0 _0924_
rlabel metal2 8960 102984 8960 102984 0 _0925_
rlabel metal2 17584 88312 17584 88312 0 _0926_
rlabel metal2 17752 95592 17752 95592 0 _0927_
rlabel metal2 18648 95536 18648 95536 0 _0928_
rlabel metal2 17752 95928 17752 95928 0 _0929_
rlabel metal2 16744 98336 16744 98336 0 _0930_
rlabel metal2 15176 98448 15176 98448 0 _0931_
rlabel metal2 12488 104832 12488 104832 0 _0932_
rlabel metal2 15960 87864 15960 87864 0 _0933_
rlabel metal3 15512 90944 15512 90944 0 _0934_
rlabel metal2 14336 93912 14336 93912 0 _0935_
rlabel metal2 13888 102312 13888 102312 0 _0936_
rlabel metal2 13608 104944 13608 104944 0 _0937_
rlabel metal2 8120 102984 8120 102984 0 _0938_
rlabel metal2 7672 103376 7672 103376 0 _0939_
rlabel metal2 19880 22848 19880 22848 0 _0940_
rlabel metal2 25480 5600 25480 5600 0 _0941_
rlabel metal3 18704 1848 18704 1848 0 _0942_
rlabel metal2 18648 2296 18648 2296 0 _0943_
rlabel metal3 22624 3304 22624 3304 0 _0944_
rlabel metal2 24304 5992 24304 5992 0 _0945_
rlabel metal2 22120 7952 22120 7952 0 _0946_
rlabel metal2 11312 2632 11312 2632 0 _0947_
rlabel metal2 11704 2856 11704 2856 0 _0948_
rlabel metal2 12152 2968 12152 2968 0 _0949_
rlabel metal2 5992 2968 5992 2968 0 _0950_
rlabel metal2 6328 2968 6328 2968 0 _0951_
rlabel metal2 11032 3584 11032 3584 0 _0952_
rlabel metal2 20328 3640 20328 3640 0 _0953_
rlabel metal3 24416 2968 24416 2968 0 _0954_
rlabel metal2 17528 3080 17528 3080 0 _0955_
rlabel metal2 20776 2464 20776 2464 0 _0956_
rlabel metal3 20888 3640 20888 3640 0 _0957_
rlabel metal2 23912 5768 23912 5768 0 _0958_
rlabel metal2 22680 8680 22680 8680 0 _0959_
rlabel metal2 27048 52472 27048 52472 0 _0960_
rlabel metal2 25256 17584 25256 17584 0 _0961_
rlabel metal2 28168 54656 28168 54656 0 _0962_
rlabel metal2 22792 21728 22792 21728 0 _0963_
rlabel metal2 22064 69496 22064 69496 0 _0964_
rlabel metal3 2912 92232 2912 92232 0 _0965_
rlabel metal2 19544 16968 19544 16968 0 _0966_
rlabel metal2 12488 20944 12488 20944 0 _0967_
rlabel metal2 11312 17640 11312 17640 0 _0968_
rlabel metal2 21952 22456 21952 22456 0 _0969_
rlabel metal2 21672 16968 21672 16968 0 _0970_
rlabel metal2 15456 16856 15456 16856 0 _0971_
rlabel metal2 16856 17752 16856 17752 0 _0972_
rlabel metal2 17920 65240 17920 65240 0 _0973_
rlabel metal2 12432 75768 12432 75768 0 _0974_
rlabel metal2 15400 20216 15400 20216 0 _0975_
rlabel metal3 17024 64456 17024 64456 0 _0976_
rlabel metal2 27272 60872 27272 60872 0 _0977_
rlabel metal2 11368 75208 11368 75208 0 _0978_
rlabel metal2 16352 87192 16352 87192 0 cal_ena
rlabel metal2 9520 23800 9520 23800 0 cal_lut\[100\]
rlabel metal2 7504 33992 7504 33992 0 cal_lut\[101\]
rlabel metal2 6104 16072 6104 16072 0 cal_lut\[102\]
rlabel metal2 23128 18984 23128 18984 0 cal_lut\[103\]
rlabel metal2 23184 15624 23184 15624 0 cal_lut\[104\]
rlabel metal2 24360 16016 24360 16016 0 cal_lut\[105\]
rlabel metal2 19936 16968 19936 16968 0 cal_lut\[106\]
rlabel metal2 13608 15792 13608 15792 0 cal_lut\[107\]
rlabel metal2 12488 16072 12488 16072 0 cal_lut\[108\]
rlabel metal2 9632 63224 9632 63224 0 cal_lut\[109\]
rlabel via2 22904 64792 22904 64792 0 cal_lut\[10\]
rlabel metal2 8512 64792 8512 64792 0 cal_lut\[110\]
rlabel metal2 7560 68488 7560 68488 0 cal_lut\[111\]
rlabel metal2 8288 67256 8288 67256 0 cal_lut\[112\]
rlabel metal3 12992 63112 12992 63112 0 cal_lut\[113\]
rlabel metal2 7448 50036 7448 50036 0 cal_lut\[114\]
rlabel metal2 12488 27608 12488 27608 0 cal_lut\[115\]
rlabel metal2 12152 36008 12152 36008 0 cal_lut\[116\]
rlabel metal3 8792 38136 8792 38136 0 cal_lut\[117\]
rlabel metal3 8120 45864 8120 45864 0 cal_lut\[118\]
rlabel metal2 23688 32760 23688 32760 0 cal_lut\[119\]
rlabel metal2 13384 59024 13384 59024 0 cal_lut\[11\]
rlabel metal2 23016 39760 23016 39760 0 cal_lut\[120\]
rlabel metal2 20664 41888 20664 41888 0 cal_lut\[121\]
rlabel metal2 17696 29624 17696 29624 0 cal_lut\[122\]
rlabel metal3 24528 26264 24528 26264 0 cal_lut\[123\]
rlabel metal2 19096 32368 19096 32368 0 cal_lut\[124\]
rlabel metal2 21784 29456 21784 29456 0 cal_lut\[125\]
rlabel metal2 25480 36960 25480 36960 0 cal_lut\[126\]
rlabel metal2 25480 47040 25480 47040 0 cal_lut\[127\]
rlabel metal3 22288 46648 22288 46648 0 cal_lut\[128\]
rlabel metal2 17640 24416 17640 24416 0 cal_lut\[129\]
rlabel metal3 8400 56056 8400 56056 0 cal_lut\[12\]
rlabel metal2 11928 21672 11928 21672 0 cal_lut\[130\]
rlabel metal3 17752 24584 17752 24584 0 cal_lut\[131\]
rlabel metal2 12152 22624 12152 22624 0 cal_lut\[132\]
rlabel metal3 4200 13608 4200 13608 0 cal_lut\[133\]
rlabel metal3 4088 18424 4088 18424 0 cal_lut\[134\]
rlabel metal2 3304 23128 3304 23128 0 cal_lut\[135\]
rlabel metal2 3864 24080 3864 24080 0 cal_lut\[136\]
rlabel metal3 15400 30240 15400 30240 0 cal_lut\[137\]
rlabel metal2 6608 28056 6608 28056 0 cal_lut\[138\]
rlabel metal2 4648 31416 4648 31416 0 cal_lut\[139\]
rlabel metal2 9016 29680 9016 29680 0 cal_lut\[13\]
rlabel metal2 4648 34440 4648 34440 0 cal_lut\[140\]
rlabel metal3 8736 37128 8736 37128 0 cal_lut\[141\]
rlabel metal2 4648 42728 4648 42728 0 cal_lut\[142\]
rlabel metal2 4312 29064 4312 29064 0 cal_lut\[143\]
rlabel metal2 15344 36456 15344 36456 0 cal_lut\[144\]
rlabel metal2 8624 33432 8624 33432 0 cal_lut\[145\]
rlabel metal2 7280 40264 7280 40264 0 cal_lut\[146\]
rlabel metal2 3304 36624 3304 36624 0 cal_lut\[147\]
rlabel metal2 4648 45584 4648 45584 0 cal_lut\[148\]
rlabel metal3 5544 34328 5544 34328 0 cal_lut\[149\]
rlabel metal3 7728 30184 7728 30184 0 cal_lut\[14\]
rlabel metal2 3304 59584 3304 59584 0 cal_lut\[150\]
rlabel metal3 4200 63224 4200 63224 0 cal_lut\[151\]
rlabel metal2 5544 54488 5544 54488 0 cal_lut\[152\]
rlabel metal2 4760 51912 4760 51912 0 cal_lut\[153\]
rlabel metal2 3528 71400 3528 71400 0 cal_lut\[154\]
rlabel metal3 7560 45080 7560 45080 0 cal_lut\[155\]
rlabel metal2 11368 48384 11368 48384 0 cal_lut\[156\]
rlabel metal2 7448 79520 7448 79520 0 cal_lut\[157\]
rlabel metal2 4816 82040 4816 82040 0 cal_lut\[158\]
rlabel metal2 9688 82096 9688 82096 0 cal_lut\[159\]
rlabel metal2 9128 31416 9128 31416 0 cal_lut\[15\]
rlabel metal2 7000 82992 7000 82992 0 cal_lut\[160\]
rlabel metal2 20776 22288 20776 22288 0 cal_lut\[161\]
rlabel metal2 16520 22680 16520 22680 0 cal_lut\[162\]
rlabel metal2 28000 18424 28000 18424 0 cal_lut\[163\]
rlabel metal2 18536 26768 18536 26768 0 cal_lut\[164\]
rlabel metal2 20048 20776 20048 20776 0 cal_lut\[165\]
rlabel metal2 18704 20888 18704 20888 0 cal_lut\[166\]
rlabel metal2 21672 25928 21672 25928 0 cal_lut\[167\]
rlabel metal2 15176 29344 15176 29344 0 cal_lut\[168\]
rlabel metal2 8568 23184 8568 23184 0 cal_lut\[169\]
rlabel metal2 7000 42168 7000 42168 0 cal_lut\[16\]
rlabel metal2 10472 22456 10472 22456 0 cal_lut\[170\]
rlabel metal3 9184 21672 9184 21672 0 cal_lut\[171\]
rlabel metal2 13272 21784 13272 21784 0 cal_lut\[172\]
rlabel metal2 9968 26264 9968 26264 0 cal_lut\[173\]
rlabel metal2 16408 27496 16408 27496 0 cal_lut\[174\]
rlabel metal2 12600 31920 12600 31920 0 cal_lut\[175\]
rlabel metal2 12544 37688 12544 37688 0 cal_lut\[176\]
rlabel metal2 10024 40376 10024 40376 0 cal_lut\[177\]
rlabel via2 9688 42952 9688 42952 0 cal_lut\[178\]
rlabel metal2 18928 29400 18928 29400 0 cal_lut\[179\]
rlabel metal2 8568 59752 8568 59752 0 cal_lut\[17\]
rlabel metal2 16240 35560 16240 35560 0 cal_lut\[180\]
rlabel metal2 21336 42672 21336 42672 0 cal_lut\[181\]
rlabel metal2 18760 42392 18760 42392 0 cal_lut\[182\]
rlabel metal2 25256 31920 25256 31920 0 cal_lut\[183\]
rlabel metal2 25256 38808 25256 38808 0 cal_lut\[184\]
rlabel metal3 21448 43792 21448 43792 0 cal_lut\[185\]
rlabel metal2 15176 34608 15176 34608 0 cal_lut\[186\]
rlabel metal2 25256 23128 25256 23128 0 cal_lut\[187\]
rlabel metal3 27664 20776 27664 20776 0 cal_lut\[188\]
rlabel metal2 27160 27608 27160 27608 0 cal_lut\[189\]
rlabel metal3 7056 55944 7056 55944 0 cal_lut\[18\]
rlabel metal2 18984 37128 18984 37128 0 cal_lut\[190\]
rlabel metal2 27160 33768 27160 33768 0 cal_lut\[191\]
rlabel metal3 23128 38024 23128 38024 0 cal_lut\[192\]
rlabel metal2 4648 50736 4648 50736 0 cal_lut\[19\]
rlabel metal3 21224 76328 21224 76328 0 cal_lut\[1\]
rlabel metal2 4648 48048 4648 48048 0 cal_lut\[20\]
rlabel metal2 8568 52752 8568 52752 0 cal_lut\[21\]
rlabel metal3 17080 47768 17080 47768 0 cal_lut\[22\]
rlabel metal2 7112 61488 7112 61488 0 cal_lut\[23\]
rlabel metal2 17640 63560 17640 63560 0 cal_lut\[24\]
rlabel metal2 7112 70672 7112 70672 0 cal_lut\[25\]
rlabel metal2 7896 72968 7896 72968 0 cal_lut\[26\]
rlabel metal2 8568 75600 8568 75600 0 cal_lut\[27\]
rlabel metal2 8232 76440 8232 76440 0 cal_lut\[28\]
rlabel metal2 17864 61432 17864 61432 0 cal_lut\[29\]
rlabel metal2 11256 77784 11256 77784 0 cal_lut\[2\]
rlabel metal2 18200 59528 18200 59528 0 cal_lut\[30\]
rlabel metal2 24696 49336 24696 49336 0 cal_lut\[31\]
rlabel metal3 23856 51352 23856 51352 0 cal_lut\[32\]
rlabel metal2 19768 19656 19768 19656 0 cal_lut\[33\]
rlabel metal3 12152 17640 12152 17640 0 cal_lut\[34\]
rlabel metal2 21896 19656 21896 19656 0 cal_lut\[35\]
rlabel metal2 17136 17640 17136 17640 0 cal_lut\[36\]
rlabel metal2 12600 76496 12600 76496 0 cal_lut\[37\]
rlabel metal3 11984 74872 11984 74872 0 cal_lut\[38\]
rlabel metal2 24472 73248 24472 73248 0 cal_lut\[39\]
rlabel metal2 23240 77952 23240 77952 0 cal_lut\[3\]
rlabel metal2 11704 72016 11704 72016 0 cal_lut\[40\]
rlabel metal2 23688 59752 23688 59752 0 cal_lut\[41\]
rlabel metal2 9688 56784 9688 56784 0 cal_lut\[42\]
rlabel metal2 10976 50008 10976 50008 0 cal_lut\[43\]
rlabel metal2 9576 47488 9576 47488 0 cal_lut\[44\]
rlabel metal2 10024 50680 10024 50680 0 cal_lut\[45\]
rlabel metal2 17976 43232 17976 43232 0 cal_lut\[46\]
rlabel metal2 14280 43848 14280 43848 0 cal_lut\[47\]
rlabel metal3 17976 44912 17976 44912 0 cal_lut\[48\]
rlabel metal2 19656 40600 19656 40600 0 cal_lut\[49\]
rlabel metal2 18536 78120 18536 78120 0 cal_lut\[4\]
rlabel metal2 18312 42560 18312 42560 0 cal_lut\[50\]
rlabel metal3 19768 35560 19768 35560 0 cal_lut\[51\]
rlabel metal3 18144 38696 18144 38696 0 cal_lut\[52\]
rlabel metal2 20832 35560 20832 35560 0 cal_lut\[53\]
rlabel metal2 18424 45080 18424 45080 0 cal_lut\[54\]
rlabel metal2 27048 57344 27048 57344 0 cal_lut\[55\]
rlabel metal2 26376 58744 26376 58744 0 cal_lut\[56\]
rlabel metal1 27720 51128 27720 51128 0 cal_lut\[57\]
rlabel metal2 22456 54880 22456 54880 0 cal_lut\[58\]
rlabel metal2 25256 44912 25256 44912 0 cal_lut\[59\]
rlabel metal1 19824 74312 19824 74312 0 cal_lut\[5\]
rlabel metal2 24024 56896 24024 56896 0 cal_lut\[60\]
rlabel metal3 27776 55272 27776 55272 0 cal_lut\[61\]
rlabel metal2 26824 52472 26824 52472 0 cal_lut\[62\]
rlabel via2 27832 51352 27832 51352 0 cal_lut\[63\]
rlabel metal3 23128 53592 23128 53592 0 cal_lut\[64\]
rlabel metal2 21784 26488 21784 26488 0 cal_lut\[65\]
rlabel metal2 12936 56728 12936 56728 0 cal_lut\[66\]
rlabel metal2 20888 10472 20888 10472 0 cal_lut\[67\]
rlabel metal2 18200 9296 18200 9296 0 cal_lut\[68\]
rlabel metal3 16744 10584 16744 10584 0 cal_lut\[69\]
rlabel metal2 16632 81200 16632 81200 0 cal_lut\[6\]
rlabel metal2 15848 10584 15848 10584 0 cal_lut\[70\]
rlabel metal2 14056 18368 14056 18368 0 cal_lut\[71\]
rlabel metal2 15344 15512 15344 15512 0 cal_lut\[72\]
rlabel metal3 20664 11480 20664 11480 0 cal_lut\[73\]
rlabel metal2 19544 12096 19544 12096 0 cal_lut\[74\]
rlabel metal2 16464 8344 16464 8344 0 cal_lut\[75\]
rlabel metal2 11928 11088 11928 11088 0 cal_lut\[76\]
rlabel metal2 12488 24920 12488 24920 0 cal_lut\[77\]
rlabel metal2 16408 23072 16408 23072 0 cal_lut\[78\]
rlabel metal2 12488 68152 12488 68152 0 cal_lut\[79\]
rlabel metal2 24192 71736 24192 71736 0 cal_lut\[7\]
rlabel metal3 12096 67032 12096 67032 0 cal_lut\[80\]
rlabel metal2 16072 68264 16072 68264 0 cal_lut\[81\]
rlabel metal2 15288 66304 15288 66304 0 cal_lut\[82\]
rlabel metal2 11704 60088 11704 60088 0 cal_lut\[83\]
rlabel metal2 12488 54936 12488 54936 0 cal_lut\[84\]
rlabel metal2 19544 69832 19544 69832 0 cal_lut\[85\]
rlabel metal3 15792 75096 15792 75096 0 cal_lut\[86\]
rlabel metal3 27664 73976 27664 73976 0 cal_lut\[87\]
rlabel metal2 27048 71008 27048 71008 0 cal_lut\[88\]
rlabel metal2 24304 61544 24304 61544 0 cal_lut\[89\]
rlabel metal2 22568 73752 22568 73752 0 cal_lut\[8\]
rlabel metal2 16856 63280 16856 63280 0 cal_lut\[90\]
rlabel metal3 24584 73528 24584 73528 0 cal_lut\[91\]
rlabel metal2 27160 75992 27160 75992 0 cal_lut\[92\]
rlabel metal2 24472 67816 24472 67816 0 cal_lut\[93\]
rlabel metal2 25256 66864 25256 66864 0 cal_lut\[94\]
rlabel metal2 25368 62216 25368 62216 0 cal_lut\[95\]
rlabel metal3 23912 62216 23912 62216 0 cal_lut\[96\]
rlabel metal3 9016 23464 9016 23464 0 cal_lut\[97\]
rlabel metal3 8176 19208 8176 19208 0 cal_lut\[98\]
rlabel metal2 8568 17920 8568 17920 0 cal_lut\[99\]
rlabel metal3 22400 67816 22400 67816 0 cal_lut\[9\]
rlabel metal3 4760 15176 4760 15176 0 clk
rlabel metal2 11816 99624 11816 99624 0 clknet_0__0551_
rlabel metal2 13384 88424 13384 88424 0 clknet_0__0553_
rlabel metal2 14280 100296 14280 100296 0 clknet_0__0889_
rlabel metal2 19432 103152 19432 103152 0 clknet_0__0902_
rlabel metal2 17304 33824 17304 33824 0 clknet_0_clk
rlabel metal3 15512 100688 15512 100688 0 clknet_0_net81
rlabel metal2 15512 104216 15512 104216 0 clknet_0_temp1.i_precharge_n
rlabel metal3 6104 96152 6104 96152 0 clknet_1_0__leaf__0551_
rlabel metal2 10808 86184 10808 86184 0 clknet_1_0__leaf__0553_
rlabel metal2 11032 101192 11032 101192 0 clknet_1_0__leaf__0889_
rlabel metal2 21280 102088 21280 102088 0 clknet_1_0__leaf__0902_
rlabel metal3 20832 16072 20832 16072 0 clknet_1_0__leaf_clk
rlabel metal2 9352 103040 9352 103040 0 clknet_1_0__leaf_net81
rlabel metal2 11256 105392 11256 105392 0 clknet_1_0__leaf_temp1.i_precharge_n
rlabel metal2 7112 99456 7112 99456 0 clknet_1_1__leaf__0551_
rlabel metal3 12488 90776 12488 90776 0 clknet_1_1__leaf__0553_
rlabel metal2 16856 103152 16856 103152 0 clknet_1_1__leaf__0889_
rlabel metal2 22232 103824 22232 103824 0 clknet_1_1__leaf__0902_
rlabel metal2 19432 87192 19432 87192 0 clknet_1_1__leaf_clk
rlabel metal2 15960 105896 15960 105896 0 clknet_1_1__leaf_net81
rlabel metal3 14336 103768 14336 103768 0 clknet_1_1__leaf_temp1.i_precharge_n
rlabel metal2 1848 18032 1848 18032 0 clknet_leaf_0_clk
rlabel metal2 28112 59416 28112 59416 0 clknet_leaf_10_clk
rlabel metal2 27720 52416 27720 52416 0 clknet_leaf_11_clk
rlabel metal2 28168 30800 28168 30800 0 clknet_leaf_12_clk
rlabel metal2 28168 23408 28168 23408 0 clknet_leaf_13_clk
rlabel metal3 18312 21560 18312 21560 0 clknet_leaf_14_clk
rlabel metal3 16800 16184 16800 16184 0 clknet_leaf_15_clk
rlabel metal3 17752 30184 17752 30184 0 clknet_leaf_16_clk
rlabel metal2 15736 14112 15736 14112 0 clknet_leaf_17_clk
rlabel metal2 9688 24976 9688 24976 0 clknet_leaf_18_clk
rlabel metal2 2240 10696 2240 10696 0 clknet_leaf_19_clk
rlabel metal2 1848 47040 1848 47040 0 clknet_leaf_1_clk
rlabel metal2 13608 39256 13608 39256 0 clknet_leaf_2_clk
rlabel metal3 8680 72632 8680 72632 0 clknet_leaf_3_clk
rlabel metal2 1736 66304 1736 66304 0 clknet_leaf_4_clk
rlabel metal2 1848 91672 1848 91672 0 clknet_leaf_5_clk
rlabel metal3 10808 93912 10808 93912 0 clknet_leaf_6_clk
rlabel metal2 13496 66696 13496 66696 0 clknet_leaf_7_clk
rlabel metal2 21448 72688 21448 72688 0 clknet_leaf_8_clk
rlabel metal2 27384 100352 27384 100352 0 clknet_leaf_9_clk
rlabel metal2 11816 103264 11816 103264 0 ctr\[0\]
rlabel metal2 21952 96264 21952 96264 0 ctr\[10\]
rlabel metal2 22176 96264 22176 96264 0 ctr\[11\]
rlabel metal2 22344 95984 22344 95984 0 ctr\[12\]
rlabel metal2 8792 101136 8792 101136 0 ctr\[1\]
rlabel metal2 19656 95256 19656 95256 0 ctr\[2\]
rlabel metal4 10920 93240 10920 93240 0 ctr\[3\]
rlabel metal2 18816 88984 18816 88984 0 ctr\[4\]
rlabel metal2 4648 91112 4648 91112 0 ctr\[5\]
rlabel metal2 19376 92680 19376 92680 0 ctr\[6\]
rlabel metal2 16296 95424 16296 95424 0 ctr\[7\]
rlabel metal2 21672 95872 21672 95872 0 ctr\[8\]
rlabel metal2 21336 96880 21336 96880 0 ctr\[9\]
rlabel metal2 9352 85120 9352 85120 0 dbg3\[0\]
rlabel metal2 12936 88256 12936 88256 0 dbg3\[1\]
rlabel metal2 9016 87360 9016 87360 0 dbg3\[2\]
rlabel metal2 10808 90608 10808 90608 0 dbg3\[3\]
rlabel metal2 12264 80808 12264 80808 0 dbg3\[4\]
rlabel metal2 16184 93072 16184 93072 0 dbg3\[5\]
rlabel metal2 27160 89712 27160 89712 0 dec1._000_
rlabel metal3 25928 85568 25928 85568 0 dec1._001_
rlabel metal2 21112 83048 21112 83048 0 dec1._002_
rlabel metal3 20832 83608 20832 83608 0 dec1._003_
rlabel metal2 19992 83216 19992 83216 0 dec1._004_
rlabel metal2 23464 83048 23464 83048 0 dec1._005_
rlabel metal2 21784 84392 21784 84392 0 dec1._006_
rlabel metal2 24248 83328 24248 83328 0 dec1._007_
rlabel metal3 25424 86632 25424 86632 0 dec1._008_
rlabel metal2 22008 82600 22008 82600 0 dec1._009_
rlabel metal2 22792 84448 22792 84448 0 dec1._010_
rlabel metal3 25424 82824 25424 82824 0 dec1._011_
rlabel metal2 23464 81816 23464 81816 0 dec1._012_
rlabel metal2 24472 80416 24472 80416 0 dec1._013_
rlabel metal3 25424 82712 25424 82712 0 dec1._014_
rlabel metal3 22288 81256 22288 81256 0 dec1._015_
rlabel metal2 23800 81704 23800 81704 0 dec1._016_
rlabel metal2 26264 82040 26264 82040 0 dec1._017_
rlabel metal3 25032 84280 25032 84280 0 dec1._018_
rlabel metal3 24696 81032 24696 81032 0 dec1._019_
rlabel metal2 26600 81984 26600 81984 0 dec1._020_
rlabel metal2 26152 83776 26152 83776 0 dec1._021_
rlabel metal3 25032 80920 25032 80920 0 dec1._022_
rlabel metal2 24808 84504 24808 84504 0 dec1._023_
rlabel metal2 27272 84952 27272 84952 0 dec1._024_
rlabel metal2 27160 85848 27160 85848 0 dec1._025_
rlabel metal2 25704 80136 25704 80136 0 dec1._026_
rlabel metal2 26320 85064 26320 85064 0 dec1._027_
rlabel metal3 26152 87416 26152 87416 0 dec1._028_
rlabel metal2 27160 88144 27160 88144 0 dec1._029_
rlabel metal3 21952 88200 21952 88200 0 dec1._030_
rlabel metal2 26600 80640 26600 80640 0 dec1._031_
rlabel metal2 26488 80752 26488 80752 0 dec1._032_
rlabel metal2 22960 81368 22960 81368 0 dec1._033_
rlabel metal2 27160 82208 27160 82208 0 dec1._034_
rlabel metal2 27944 86156 27944 86156 0 dec1._035_
rlabel metal2 28168 81424 28168 81424 0 dec1._036_
rlabel metal2 27272 88256 27272 88256 0 dec1._037_
rlabel metal2 26152 88704 26152 88704 0 dec1._038_
rlabel metal2 27832 86352 27832 86352 0 dec1._039_
rlabel metal2 24696 88592 24696 88592 0 dec1._040_
rlabel metal3 25088 85848 25088 85848 0 dec1._041_
rlabel metal3 25480 85736 25480 85736 0 dec1._042_
rlabel metal2 25032 86352 25032 86352 0 dec1._043_
rlabel metal3 25928 87192 25928 87192 0 dec1._044_
rlabel metal2 27104 84056 27104 84056 0 dec1._045_
rlabel metal2 26656 84392 26656 84392 0 dec1._046_
rlabel metal2 27496 85848 27496 85848 0 dec1._047_
rlabel metal2 26376 87808 26376 87808 0 dec1._048_
rlabel metal3 18872 88088 18872 88088 0 dec1.i_bin\[0\]
rlabel metal2 24472 86688 24472 86688 0 dec1.i_bin\[1\]
rlabel metal3 20888 79800 20888 79800 0 dec1.i_bin\[2\]
rlabel metal3 23016 80136 23016 80136 0 dec1.i_bin\[3\]
rlabel metal2 20328 83048 20328 83048 0 dec1.i_bin\[4\]
rlabel metal3 20888 81928 20888 81928 0 dec1.i_bin\[5\]
rlabel metal2 22568 82320 22568 82320 0 dec1.i_bin\[6\]
rlabel metal2 28168 91504 28168 91504 0 dec1.i_ones
rlabel metal2 26936 94024 26936 94024 0 dec1.i_tens
rlabel metal2 24360 88592 24360 88592 0 dec1.o_dec\[0\]
rlabel metal3 27020 91112 27020 91112 0 dec1.o_dec\[1\]
rlabel metal2 26208 92904 26208 92904 0 dec1.o_dec\[2\]
rlabel metal2 26376 89768 26376 89768 0 dec1.o_dec\[3\]
rlabel metal2 16632 85120 16632 85120 0 en_dbg\[0\]
rlabel metal2 15512 94472 15512 94472 0 en_dbg\[1\]
rlabel metal2 12376 83160 12376 83160 0 en_dbg\[2\]
rlabel metal2 27048 2240 27048 2240 0 i_wb_addr[0]
rlabel metal2 18312 4144 18312 4144 0 i_wb_addr[10]
rlabel metal3 19544 1848 19544 1848 0 i_wb_addr[11]
rlabel metal2 17640 2296 17640 2296 0 i_wb_addr[12]
rlabel metal3 16576 1848 16576 1848 0 i_wb_addr[13]
rlabel metal2 15624 1848 15624 1848 0 i_wb_addr[14]
rlabel metal2 15064 1792 15064 1792 0 i_wb_addr[15]
rlabel metal3 14112 1960 14112 1960 0 i_wb_addr[16]
rlabel metal2 13944 1736 13944 1736 0 i_wb_addr[17]
rlabel metal2 12376 2072 12376 2072 0 i_wb_addr[18]
rlabel metal2 11760 1960 11760 1960 0 i_wb_addr[19]
rlabel metal2 27608 2016 27608 2016 0 i_wb_addr[1]
rlabel metal2 11256 2184 11256 2184 0 i_wb_addr[20]
rlabel metal2 10360 2016 10360 2016 0 i_wb_addr[21]
rlabel metal2 9744 1960 9744 1960 0 i_wb_addr[22]
rlabel metal2 9688 2464 9688 2464 0 i_wb_addr[23]
rlabel metal2 8232 2296 8232 2296 0 i_wb_addr[24]
rlabel metal2 7896 1680 7896 1680 0 i_wb_addr[25]
rlabel metal2 7224 2632 7224 2632 0 i_wb_addr[26]
rlabel metal2 6552 2632 6552 2632 0 i_wb_addr[27]
rlabel metal2 6104 2632 6104 2632 0 i_wb_addr[28]
rlabel metal2 4760 1904 4760 1904 0 i_wb_addr[29]
rlabel metal2 25816 1960 25816 1960 0 i_wb_addr[2]
rlabel metal2 4088 1792 4088 1792 0 i_wb_addr[30]
rlabel metal3 3640 1848 3640 1848 0 i_wb_addr[31]
rlabel metal2 24976 1960 24976 1960 0 i_wb_addr[3]
rlabel metal2 22232 406 22232 406 0 i_wb_addr[4]
rlabel metal2 22456 2296 22456 2296 0 i_wb_addr[5]
rlabel metal2 20776 1848 20776 1848 0 i_wb_addr[6]
rlabel metal2 20328 1736 20328 1736 0 i_wb_addr[7]
rlabel metal3 25032 4872 25032 4872 0 i_wb_addr[8]
rlabel metal2 18816 1512 18816 1512 0 i_wb_addr[9]
rlabel metal2 27496 2464 27496 2464 0 i_wb_cyc
rlabel metal2 1736 4928 1736 4928 0 i_wb_data[0]
rlabel metal3 1022 31640 1022 31640 0 i_wb_data[10]
rlabel metal2 1736 34552 1736 34552 0 i_wb_data[11]
rlabel metal2 1736 36736 1736 36736 0 i_wb_data[12]
rlabel via2 1736 39704 1736 39704 0 i_wb_data[13]
rlabel metal2 1736 41272 1736 41272 0 i_wb_data[14]
rlabel metal2 1736 45192 1736 45192 0 i_wb_data[15]
rlabel metal3 2184 47320 2184 47320 0 i_wb_data[16]
rlabel metal2 1736 48664 1736 48664 0 i_wb_data[17]
rlabel metal2 1904 49112 1904 49112 0 i_wb_data[18]
rlabel metal2 1736 55944 1736 55944 0 i_wb_data[19]
rlabel metal3 1022 7448 1022 7448 0 i_wb_data[1]
rlabel metal2 1736 58856 1736 58856 0 i_wb_data[20]
rlabel metal2 1736 61320 1736 61320 0 i_wb_data[21]
rlabel metal3 1078 63896 1078 63896 0 i_wb_data[22]
rlabel metal2 1736 66808 1736 66808 0 i_wb_data[23]
rlabel metal2 1848 70112 1848 70112 0 i_wb_data[24]
rlabel metal2 1736 72632 1736 72632 0 i_wb_data[25]
rlabel metal2 1736 74760 1736 74760 0 i_wb_data[26]
rlabel metal2 1736 77672 1736 77672 0 i_wb_data[27]
rlabel metal2 1736 80080 1736 80080 0 i_wb_data[28]
rlabel metal2 1736 83048 1736 83048 0 i_wb_data[29]
rlabel metal2 2744 11144 2744 11144 0 i_wb_data[2]
rlabel metal3 1022 85400 1022 85400 0 i_wb_data[30]
rlabel metal3 1022 88088 1022 88088 0 i_wb_data[31]
rlabel metal2 1736 10248 1736 10248 0 i_wb_data[3]
rlabel metal3 1078 15512 1078 15512 0 i_wb_data[4]
rlabel metal2 1736 18312 1736 18312 0 i_wb_data[5]
rlabel metal3 1078 20888 1078 20888 0 i_wb_data[6]
rlabel metal2 1736 22624 1736 22624 0 i_wb_data[7]
rlabel metal3 1022 26264 1022 26264 0 i_wb_data[8]
rlabel metal2 1736 29008 1736 29008 0 i_wb_data[9]
rlabel metal2 26936 2464 26936 2464 0 i_wb_stb
rlabel metal2 27608 3136 27608 3136 0 i_wb_we
rlabel metal2 28280 116942 28280 116942 0 io_out[0]
rlabel metal2 25704 118552 25704 118552 0 io_out[1]
rlabel metal2 24024 119672 24024 119672 0 io_out[2]
rlabel metal3 23520 114408 23520 114408 0 io_out[3]
rlabel metal2 21112 113834 21112 113834 0 io_out[4]
rlabel metal2 19320 116942 19320 116942 0 io_out[5]
rlabel metal2 17584 116984 17584 116984 0 io_out[6]
rlabel metal2 15624 116984 15624 116984 0 io_out[7]
rlabel metal2 26712 2800 26712 2800 0 net1
rlabel metal2 12600 2184 12600 2184 0 net10
rlabel metal2 11928 2296 11928 2296 0 net11
rlabel metal2 24360 2296 24360 2296 0 net12
rlabel metal3 10920 1960 10920 1960 0 net13
rlabel metal2 10584 1904 10584 1904 0 net14
rlabel metal2 9912 2184 9912 2184 0 net15
rlabel metal3 10304 2744 10304 2744 0 net16
rlabel metal3 9240 3528 9240 3528 0 net17
rlabel metal2 8120 2408 8120 2408 0 net18
rlabel metal2 7448 2352 7448 2352 0 net19
rlabel metal2 19600 2856 19600 2856 0 net2
rlabel metal2 6888 1848 6888 1848 0 net20
rlabel metal2 5712 1848 5712 1848 0 net21
rlabel metal3 5376 3416 5376 3416 0 net22
rlabel metal2 25368 2520 25368 2520 0 net23
rlabel metal2 4312 2296 4312 2296 0 net24
rlabel metal2 3640 2016 3640 2016 0 net25
rlabel metal2 24752 2072 24752 2072 0 net26
rlabel metal2 22904 2408 22904 2408 0 net27
rlabel metal2 21840 2856 21840 2856 0 net28
rlabel metal3 22176 3416 22176 3416 0 net29
rlabel metal2 19320 2296 19320 2296 0 net3
rlabel metal2 21224 4872 21224 4872 0 net30
rlabel metal2 23688 2352 23688 2352 0 net31
rlabel metal2 18032 2856 18032 2856 0 net32
rlabel metal2 26152 3192 26152 3192 0 net33
rlabel metal2 2072 5656 2072 5656 0 net34
rlabel metal2 2072 31696 2072 31696 0 net35
rlabel metal2 2800 34888 2800 34888 0 net36
rlabel metal3 2716 36232 2716 36232 0 net37
rlabel metal2 2856 40656 2856 40656 0 net38
rlabel metal2 2128 41160 2128 41160 0 net39
rlabel metal2 17920 1848 17920 1848 0 net4
rlabel metal2 2856 44184 2856 44184 0 net40
rlabel metal2 5096 47040 5096 47040 0 net41
rlabel metal2 5656 49504 5656 49504 0 net42
rlabel metal2 2520 52528 2520 52528 0 net43
rlabel metal2 2464 53704 2464 53704 0 net44
rlabel metal2 2072 8960 2072 8960 0 net45
rlabel metal2 2072 58856 2072 58856 0 net46
rlabel metal2 3304 61152 3304 61152 0 net47
rlabel metal3 2464 64456 2464 64456 0 net48
rlabel metal2 2912 67032 2912 67032 0 net49
rlabel metal2 17304 2604 17304 2604 0 net5
rlabel metal2 2408 70392 2408 70392 0 net50
rlabel metal2 2968 73304 2968 73304 0 net51
rlabel metal2 2072 74928 2072 74928 0 net52
rlabel metal3 2408 77112 2408 77112 0 net53
rlabel metal3 17864 80024 17864 80024 0 net54
rlabel metal2 3304 81144 3304 81144 0 net55
rlabel metal2 4536 10976 4536 10976 0 net56
rlabel metal2 22120 80416 22120 80416 0 net57
rlabel metal2 2072 87752 2072 87752 0 net58
rlabel metal2 2072 11816 2072 11816 0 net59
rlabel metal2 16072 2352 16072 2352 0 net6
rlabel metal2 2184 15848 2184 15848 0 net60
rlabel metal2 2968 17584 2968 17584 0 net61
rlabel metal3 2408 20776 2408 20776 0 net62
rlabel metal3 2632 23352 2632 23352 0 net63
rlabel metal2 2744 25424 2744 25424 0 net64
rlabel metal2 2184 28672 2184 28672 0 net65
rlabel metal2 25368 2688 25368 2688 0 net66
rlabel metal3 25088 2856 25088 2856 0 net67
rlabel metal2 2968 2296 2968 2296 0 net68
rlabel metal2 13384 118328 13384 118328 0 net69
rlabel metal2 15288 1848 15288 1848 0 net7
rlabel metal2 12264 117880 12264 117880 0 net70
rlabel metal2 10472 117880 10472 117880 0 net71
rlabel metal2 9352 118328 9352 118328 0 net72
rlabel metal2 6888 117880 6888 117880 0 net73
rlabel metal2 5544 118328 5544 118328 0 net74
rlabel metal2 3304 117880 3304 117880 0 net75
rlabel metal2 1736 118272 1736 118272 0 net76
rlabel metal3 1022 114968 1022 114968 0 net77
rlabel metal2 26936 103824 26936 103824 0 net78
rlabel metal2 25088 104776 25088 104776 0 net79
rlabel metal2 14392 2184 14392 2184 0 net8
rlabel metal2 24696 104608 24696 104608 0 net80
rlabel metal2 9072 105224 9072 105224 0 net81
rlabel metal2 6552 99456 6552 99456 0 net82
rlabel metal2 15848 105168 15848 105168 0 net83
rlabel metal3 9072 15400 9072 15400 0 net84
rlabel metal2 13720 2016 13720 2016 0 net9
rlabel metal3 1022 90776 1022 90776 0 o_wb_ack
rlabel metal2 1736 93240 1736 93240 0 o_wb_data[0]
rlabel metal3 1022 96152 1022 96152 0 o_wb_data[1]
rlabel metal2 1736 99064 1736 99064 0 o_wb_data[2]
rlabel metal2 1736 101528 1736 101528 0 o_wb_data[3]
rlabel metal2 1736 103656 1736 103656 0 o_wb_data[4]
rlabel metal2 5880 104608 5880 104608 0 o_wb_data[5]
rlabel metal2 1736 107576 1736 107576 0 o_wb_data[6]
rlabel metal3 2142 112280 2142 112280 0 o_wb_data[7]
rlabel metal2 2744 1134 2744 1134 0 reset
rlabel metal2 27160 92624 27160 92624 0 seg1._00_
rlabel metal2 25816 91728 25816 91728 0 seg1._01_
rlabel metal2 26488 92400 26488 92400 0 seg1._02_
rlabel metal2 22008 89488 22008 89488 0 seg1._03_
rlabel metal2 26208 92120 26208 92120 0 seg1._04_
rlabel metal2 27440 91560 27440 91560 0 seg1._05_
rlabel metal2 27160 92120 27160 92120 0 seg1._06_
rlabel metal2 27272 91896 27272 91896 0 seg1._07_
rlabel metal3 22792 89544 22792 89544 0 seg1._08_
rlabel metal2 22904 89880 22904 89880 0 seg1._09_
rlabel metal2 22120 89432 22120 89432 0 seg1._10_
rlabel metal3 27048 92176 27048 92176 0 seg1._11_
rlabel metal3 22176 91336 22176 91336 0 seg1._12_
rlabel metal2 22568 91672 22568 91672 0 seg1._13_
rlabel metal2 22904 90776 22904 90776 0 seg1._14_
rlabel metal2 22288 90552 22288 90552 0 seg1._15_
rlabel metal2 22232 92120 22232 92120 0 seg1._16_
rlabel metal2 23464 91952 23464 91952 0 seg1._17_
rlabel metal2 22400 93128 22400 93128 0 seg1._18_
rlabel metal2 22456 92568 22456 92568 0 seg1._19_
rlabel metal2 24024 92848 24024 92848 0 seg1._20_
rlabel metal2 24136 92624 24136 92624 0 seg1._21_
rlabel metal2 23464 89824 23464 89824 0 seg1._22_
rlabel metal2 22680 88704 22680 88704 0 seg1._23_
rlabel metal3 24696 88984 24696 88984 0 seg1._24_
rlabel metal2 24584 90496 24584 90496 0 seg1._25_
rlabel metal2 19208 91616 19208 91616 0 seg1.o_segments\[0\]
rlabel metal2 21672 90440 21672 90440 0 seg1.o_segments\[1\]
rlabel metal3 20944 89656 20944 89656 0 seg1.o_segments\[2\]
rlabel metal2 21896 94584 21896 94584 0 seg1.o_segments\[3\]
rlabel metal2 20664 92456 20664 92456 0 seg1.o_segments\[4\]
rlabel metal2 20776 88536 20776 88536 0 seg1.o_segments\[5\]
rlabel metal2 17976 89040 17976 89040 0 seg1.o_segments\[6\]
rlabel metal3 22960 106120 22960 106120 0 temp1.dac._0_
rlabel metal2 22904 104384 22904 104384 0 temp1.dac._1_
rlabel metal2 18312 103264 18312 103264 0 temp1.dac.i_data\[0\]
rlabel metal2 15736 96824 15736 96824 0 temp1.dac.i_data\[1\]
rlabel metal2 9800 107072 9800 107072 0 temp1.dac.i_data\[2\]
rlabel metal3 11480 108472 11480 108472 0 temp1.dac.i_data\[3\]
rlabel metal2 19992 109228 19992 109228 0 temp1.dac.i_data\[4\]
rlabel metal3 20300 109256 20300 109256 0 temp1.dac.i_data\[5\]
rlabel metal3 15624 109256 15624 109256 0 temp1.dac.i_enable
rlabel metal2 20776 103992 20776 103992 0 temp1.dac.parallel_cells\[0\].vdac_batch._0_
rlabel metal2 20328 105112 20328 105112 0 temp1.dac.parallel_cells\[0\].vdac_batch._1_
rlabel metal2 19992 106344 19992 106344 0 temp1.dac.parallel_cells\[0\].vdac_batch._2_
rlabel metal2 17472 107912 17472 107912 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal2 21448 104552 21448 104552 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal2 18200 106232 18200 106232 0 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel metal3 24472 114632 24472 114632 0 temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
rlabel metal2 16968 108472 16968 108472 0 temp1.dac.parallel_cells\[1\].vdac_batch._0_
rlabel metal2 16632 108360 16632 108360 0 temp1.dac.parallel_cells\[1\].vdac_batch._1_
rlabel metal3 17136 108472 17136 108472 0 temp1.dac.parallel_cells\[1\].vdac_batch._2_
rlabel metal2 15736 107688 15736 107688 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal2 18088 107800 18088 107800 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal2 16072 107408 16072 107408 0 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal3 13776 108584 13776 108584 0 temp1.dac.parallel_cells\[2\].vdac_batch._0_
rlabel metal2 12824 108248 12824 108248 0 temp1.dac.parallel_cells\[2\].vdac_batch._1_
rlabel metal2 12376 109648 12376 109648 0 temp1.dac.parallel_cells\[2\].vdac_batch._2_
rlabel metal3 12152 107016 12152 107016 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal2 13944 110096 13944 110096 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel metal2 10808 108192 10808 108192 0 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal2 13608 109648 13608 109648 0 temp1.dac.parallel_cells\[3\].vdac_batch._0_
rlabel metal2 14280 109816 14280 109816 0 temp1.dac.parallel_cells\[3\].vdac_batch._1_
rlabel metal2 12040 110656 12040 110656 0 temp1.dac.parallel_cells\[3\].vdac_batch._2_
rlabel metal2 8008 113232 8008 113232 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal2 13440 115640 13440 115640 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal2 8344 112112 8344 112112 0 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal2 21336 109088 21336 109088 0 temp1.dac.parallel_cells\[4\].vdac_batch._0_
rlabel metal2 20608 109480 20608 109480 0 temp1.dac.parallel_cells\[4\].vdac_batch._1_
rlabel metal2 21952 106344 21952 106344 0 temp1.dac.parallel_cells\[4\].vdac_batch._2_
rlabel metal2 25928 109760 25928 109760 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal2 21448 114576 21448 114576 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal2 26712 109760 26712 109760 0 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal2 24024 102256 24024 102256 0 temp1.dac.vdac_single._0_
rlabel metal2 24472 103992 24472 103992 0 temp1.dac.vdac_single._1_
rlabel metal2 24976 105448 24976 105448 0 temp1.dac.vdac_single._2_
rlabel metal2 25368 104944 25368 104944 0 temp1.dac.vdac_single.en_pupd
rlabel metal2 24304 102424 24304 102424 0 temp1.dac.vdac_single.en_vref
rlabel metal2 26712 104384 26712 104384 0 temp1.dac.vdac_single.npu_pd
rlabel metal2 10472 105056 10472 105056 0 temp1.dcdel_capnode_notouch_
rlabel metal2 9016 104720 9016 104720 0 temp1.i_precharge_n
rlabel metal2 8792 98336 8792 98336 0 temp_delay_last
<< properties >>
string FIXED_BBOX 0 0 30000 120000
<< end >>
